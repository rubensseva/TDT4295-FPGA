module VideoBuffer(
  input         clock,
  input         reset,
  input  [3:0]  io_pixelVal_in_0,
  input  [3:0]  io_pixelVal_in_1,
  input  [3:0]  io_pixelVal_in_2,
  input  [3:0]  io_pixelVal_in_3,
  input  [3:0]  io_pixelVal_in_4,
  input  [3:0]  io_pixelVal_in_5,
  input  [3:0]  io_pixelVal_in_6,
  input  [3:0]  io_pixelVal_in_7,
  input         io_valid_in,
  input  [10:0] io_rowIndex,
  input  [10:0] io_colIndex,
  output [3:0]  io_pixelVal_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [17:0] _T = io_rowIndex * 11'h40; // @[VideoBuffer.scala 29:46]
  wire [17:0] _GEN_30722 = {{7'd0}, io_colIndex}; // @[VideoBuffer.scala 29:61]
  wire [17:0] _T_2 = _T + _GEN_30722; // @[VideoBuffer.scala 29:61]
  reg [31:0] pixelIndex; // @[VideoBuffer.scala 31:33]
  wire [31:0] _T_26 = pixelIndex + 32'h7; // @[VideoBuffer.scala 35:42]
  wire [31:0] _T_23 = pixelIndex + 32'h6; // @[VideoBuffer.scala 35:42]
  wire [31:0] _T_20 = pixelIndex + 32'h5; // @[VideoBuffer.scala 35:42]
  wire [31:0] _T_17 = pixelIndex + 32'h4; // @[VideoBuffer.scala 35:42]
  wire [31:0] _T_14 = pixelIndex + 32'h3; // @[VideoBuffer.scala 35:42]
  wire [31:0] _T_11 = pixelIndex + 32'h2; // @[VideoBuffer.scala 35:42]
  wire [31:0] _T_8 = pixelIndex + 32'h1; // @[VideoBuffer.scala 35:42]
  wire [32:0] _T_4 = {{1'd0}, pixelIndex}; // @[VideoBuffer.scala 35:42]
  wire [3:0] _GEN_3072 = 12'h0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6144 = 12'h0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3072; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9216 = 12'h0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6144; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12288 = 12'h0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9216; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15360 = 12'h0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12288; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18432 = 12'h0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15360; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21504 = 12'h0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18432; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24576 = 12'h0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21504; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_0 = io_valid_in ? _GEN_24576 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3073 = 12'h1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6145 = 12'h1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3073; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9217 = 12'h1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6145; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12289 = 12'h1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9217; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15361 = 12'h1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12289; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18433 = 12'h1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15361; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21505 = 12'h1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18433; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24577 = 12'h1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21505; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1 = io_valid_in ? _GEN_24577 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1 = 12'h1 == _T_2[11:0] ? image_1 : image_0; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3074 = 12'h2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6146 = 12'h2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3074; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9218 = 12'h2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6146; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12290 = 12'h2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9218; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15362 = 12'h2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12290; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18434 = 12'h2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15362; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21506 = 12'h2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18434; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24578 = 12'h2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21506; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2 = io_valid_in ? _GEN_24578 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2 = 12'h2 == _T_2[11:0] ? image_2 : _GEN_1; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3075 = 12'h3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6147 = 12'h3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3075; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9219 = 12'h3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6147; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12291 = 12'h3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9219; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15363 = 12'h3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12291; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18435 = 12'h3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15363; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21507 = 12'h3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18435; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24579 = 12'h3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21507; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3 = io_valid_in ? _GEN_24579 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3 = 12'h3 == _T_2[11:0] ? image_3 : _GEN_2; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3076 = 12'h4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6148 = 12'h4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3076; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9220 = 12'h4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6148; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12292 = 12'h4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9220; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15364 = 12'h4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12292; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18436 = 12'h4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15364; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21508 = 12'h4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18436; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24580 = 12'h4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21508; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_4 = io_valid_in ? _GEN_24580 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_4 = 12'h4 == _T_2[11:0] ? image_4 : _GEN_3; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3077 = 12'h5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6149 = 12'h5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3077; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9221 = 12'h5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6149; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12293 = 12'h5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9221; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15365 = 12'h5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12293; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18437 = 12'h5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15365; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21509 = 12'h5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18437; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24581 = 12'h5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21509; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_5 = io_valid_in ? _GEN_24581 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_5 = 12'h5 == _T_2[11:0] ? image_5 : _GEN_4; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3078 = 12'h6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6150 = 12'h6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3078; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9222 = 12'h6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6150; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12294 = 12'h6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9222; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15366 = 12'h6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12294; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18438 = 12'h6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15366; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21510 = 12'h6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18438; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24582 = 12'h6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21510; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_6 = io_valid_in ? _GEN_24582 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_6 = 12'h6 == _T_2[11:0] ? image_6 : _GEN_5; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3079 = 12'h7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6151 = 12'h7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3079; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9223 = 12'h7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6151; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12295 = 12'h7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9223; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15367 = 12'h7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12295; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18439 = 12'h7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15367; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21511 = 12'h7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18439; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24583 = 12'h7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21511; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_7 = io_valid_in ? _GEN_24583 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_7 = 12'h7 == _T_2[11:0] ? image_7 : _GEN_6; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3080 = 12'h8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6152 = 12'h8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3080; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9224 = 12'h8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6152; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12296 = 12'h8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9224; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15368 = 12'h8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12296; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18440 = 12'h8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15368; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21512 = 12'h8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18440; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24584 = 12'h8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21512; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_8 = io_valid_in ? _GEN_24584 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_8 = 12'h8 == _T_2[11:0] ? image_8 : _GEN_7; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3081 = 12'h9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6153 = 12'h9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3081; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9225 = 12'h9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6153; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12297 = 12'h9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9225; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15369 = 12'h9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12297; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18441 = 12'h9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15369; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21513 = 12'h9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18441; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24585 = 12'h9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21513; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_9 = io_valid_in ? _GEN_24585 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_9 = 12'h9 == _T_2[11:0] ? image_9 : _GEN_8; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3082 = 12'ha == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6154 = 12'ha == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3082; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9226 = 12'ha == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6154; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12298 = 12'ha == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9226; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15370 = 12'ha == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12298; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18442 = 12'ha == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15370; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21514 = 12'ha == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18442; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24586 = 12'ha == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21514; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_10 = io_valid_in ? _GEN_24586 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_10 = 12'ha == _T_2[11:0] ? image_10 : _GEN_9; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3083 = 12'hb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6155 = 12'hb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3083; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9227 = 12'hb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6155; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12299 = 12'hb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9227; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15371 = 12'hb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12299; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18443 = 12'hb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15371; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21515 = 12'hb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18443; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24587 = 12'hb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21515; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_11 = io_valid_in ? _GEN_24587 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_11 = 12'hb == _T_2[11:0] ? image_11 : _GEN_10; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3084 = 12'hc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6156 = 12'hc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3084; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9228 = 12'hc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6156; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12300 = 12'hc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9228; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15372 = 12'hc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12300; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18444 = 12'hc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15372; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21516 = 12'hc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18444; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24588 = 12'hc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21516; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_12 = io_valid_in ? _GEN_24588 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_12 = 12'hc == _T_2[11:0] ? image_12 : _GEN_11; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3085 = 12'hd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6157 = 12'hd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3085; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9229 = 12'hd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6157; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12301 = 12'hd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9229; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15373 = 12'hd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12301; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18445 = 12'hd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15373; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21517 = 12'hd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18445; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24589 = 12'hd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21517; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_13 = io_valid_in ? _GEN_24589 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_13 = 12'hd == _T_2[11:0] ? image_13 : _GEN_12; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3086 = 12'he == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6158 = 12'he == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3086; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9230 = 12'he == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6158; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12302 = 12'he == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9230; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15374 = 12'he == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12302; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18446 = 12'he == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15374; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21518 = 12'he == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18446; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24590 = 12'he == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21518; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_14 = io_valid_in ? _GEN_24590 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_14 = 12'he == _T_2[11:0] ? image_14 : _GEN_13; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3087 = 12'hf == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6159 = 12'hf == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3087; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9231 = 12'hf == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6159; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12303 = 12'hf == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9231; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15375 = 12'hf == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12303; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18447 = 12'hf == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15375; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21519 = 12'hf == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18447; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24591 = 12'hf == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21519; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_15 = io_valid_in ? _GEN_24591 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_15 = 12'hf == _T_2[11:0] ? image_15 : _GEN_14; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3088 = 12'h10 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6160 = 12'h10 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3088; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9232 = 12'h10 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6160; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12304 = 12'h10 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9232; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15376 = 12'h10 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12304; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18448 = 12'h10 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15376; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21520 = 12'h10 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18448; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24592 = 12'h10 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21520; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_16 = io_valid_in ? _GEN_24592 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_16 = 12'h10 == _T_2[11:0] ? image_16 : _GEN_15; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3089 = 12'h11 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6161 = 12'h11 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3089; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9233 = 12'h11 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6161; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12305 = 12'h11 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9233; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15377 = 12'h11 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12305; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18449 = 12'h11 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15377; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21521 = 12'h11 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18449; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24593 = 12'h11 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21521; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_17 = io_valid_in ? _GEN_24593 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_17 = 12'h11 == _T_2[11:0] ? image_17 : _GEN_16; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3090 = 12'h12 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6162 = 12'h12 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3090; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9234 = 12'h12 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6162; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12306 = 12'h12 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9234; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15378 = 12'h12 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12306; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18450 = 12'h12 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15378; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21522 = 12'h12 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18450; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24594 = 12'h12 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21522; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_18 = io_valid_in ? _GEN_24594 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_18 = 12'h12 == _T_2[11:0] ? image_18 : _GEN_17; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3091 = 12'h13 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6163 = 12'h13 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3091; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9235 = 12'h13 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6163; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12307 = 12'h13 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9235; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15379 = 12'h13 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12307; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18451 = 12'h13 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15379; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21523 = 12'h13 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18451; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24595 = 12'h13 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21523; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_19 = io_valid_in ? _GEN_24595 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_19 = 12'h13 == _T_2[11:0] ? image_19 : _GEN_18; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3092 = 12'h14 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6164 = 12'h14 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3092; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9236 = 12'h14 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6164; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12308 = 12'h14 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9236; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15380 = 12'h14 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12308; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18452 = 12'h14 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15380; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21524 = 12'h14 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18452; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24596 = 12'h14 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21524; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_20 = io_valid_in ? _GEN_24596 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_20 = 12'h14 == _T_2[11:0] ? image_20 : _GEN_19; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3093 = 12'h15 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6165 = 12'h15 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3093; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9237 = 12'h15 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6165; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12309 = 12'h15 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9237; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15381 = 12'h15 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12309; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18453 = 12'h15 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15381; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21525 = 12'h15 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18453; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24597 = 12'h15 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21525; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_21 = io_valid_in ? _GEN_24597 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_21 = 12'h15 == _T_2[11:0] ? image_21 : _GEN_20; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3094 = 12'h16 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6166 = 12'h16 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3094; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9238 = 12'h16 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6166; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12310 = 12'h16 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9238; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15382 = 12'h16 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12310; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18454 = 12'h16 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15382; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21526 = 12'h16 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18454; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24598 = 12'h16 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21526; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_22 = io_valid_in ? _GEN_24598 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_22 = 12'h16 == _T_2[11:0] ? image_22 : _GEN_21; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3095 = 12'h17 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6167 = 12'h17 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3095; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9239 = 12'h17 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6167; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12311 = 12'h17 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9239; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15383 = 12'h17 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12311; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18455 = 12'h17 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15383; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21527 = 12'h17 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18455; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24599 = 12'h17 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21527; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_23 = io_valid_in ? _GEN_24599 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_23 = 12'h17 == _T_2[11:0] ? image_23 : _GEN_22; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3096 = 12'h18 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6168 = 12'h18 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3096; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9240 = 12'h18 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6168; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12312 = 12'h18 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9240; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15384 = 12'h18 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12312; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18456 = 12'h18 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15384; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21528 = 12'h18 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18456; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24600 = 12'h18 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21528; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_24 = io_valid_in ? _GEN_24600 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_24 = 12'h18 == _T_2[11:0] ? image_24 : _GEN_23; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3097 = 12'h19 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6169 = 12'h19 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3097; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9241 = 12'h19 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6169; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12313 = 12'h19 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9241; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15385 = 12'h19 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12313; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18457 = 12'h19 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15385; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21529 = 12'h19 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18457; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24601 = 12'h19 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21529; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_25 = io_valid_in ? _GEN_24601 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_25 = 12'h19 == _T_2[11:0] ? image_25 : _GEN_24; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3098 = 12'h1a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6170 = 12'h1a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3098; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9242 = 12'h1a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6170; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12314 = 12'h1a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9242; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15386 = 12'h1a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12314; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18458 = 12'h1a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15386; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21530 = 12'h1a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18458; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24602 = 12'h1a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21530; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_26 = io_valid_in ? _GEN_24602 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_26 = 12'h1a == _T_2[11:0] ? image_26 : _GEN_25; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3099 = 12'h1b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6171 = 12'h1b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3099; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9243 = 12'h1b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6171; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12315 = 12'h1b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9243; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15387 = 12'h1b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12315; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18459 = 12'h1b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15387; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21531 = 12'h1b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18459; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24603 = 12'h1b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21531; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_27 = io_valid_in ? _GEN_24603 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_27 = 12'h1b == _T_2[11:0] ? image_27 : _GEN_26; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3100 = 12'h1c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6172 = 12'h1c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3100; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9244 = 12'h1c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6172; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12316 = 12'h1c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9244; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15388 = 12'h1c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12316; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18460 = 12'h1c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15388; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21532 = 12'h1c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18460; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24604 = 12'h1c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21532; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_28 = io_valid_in ? _GEN_24604 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_28 = 12'h1c == _T_2[11:0] ? image_28 : _GEN_27; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3101 = 12'h1d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6173 = 12'h1d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3101; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9245 = 12'h1d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6173; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12317 = 12'h1d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9245; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15389 = 12'h1d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12317; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18461 = 12'h1d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15389; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21533 = 12'h1d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18461; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24605 = 12'h1d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21533; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_29 = io_valid_in ? _GEN_24605 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_29 = 12'h1d == _T_2[11:0] ? image_29 : _GEN_28; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3102 = 12'h1e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6174 = 12'h1e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3102; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9246 = 12'h1e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6174; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12318 = 12'h1e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9246; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15390 = 12'h1e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12318; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18462 = 12'h1e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15390; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21534 = 12'h1e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18462; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24606 = 12'h1e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21534; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_30 = io_valid_in ? _GEN_24606 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_30 = 12'h1e == _T_2[11:0] ? image_30 : _GEN_29; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3103 = 12'h1f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6175 = 12'h1f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3103; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9247 = 12'h1f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6175; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12319 = 12'h1f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9247; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15391 = 12'h1f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12319; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18463 = 12'h1f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15391; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21535 = 12'h1f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18463; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24607 = 12'h1f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21535; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_31 = io_valid_in ? _GEN_24607 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_31 = 12'h1f == _T_2[11:0] ? image_31 : _GEN_30; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3104 = 12'h20 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6176 = 12'h20 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3104; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9248 = 12'h20 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6176; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12320 = 12'h20 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9248; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15392 = 12'h20 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12320; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18464 = 12'h20 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15392; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21536 = 12'h20 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18464; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24608 = 12'h20 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21536; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_32 = io_valid_in ? _GEN_24608 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_32 = 12'h20 == _T_2[11:0] ? image_32 : _GEN_31; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3105 = 12'h21 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6177 = 12'h21 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3105; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9249 = 12'h21 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6177; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12321 = 12'h21 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9249; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15393 = 12'h21 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12321; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18465 = 12'h21 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15393; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21537 = 12'h21 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18465; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24609 = 12'h21 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21537; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_33 = io_valid_in ? _GEN_24609 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_33 = 12'h21 == _T_2[11:0] ? image_33 : _GEN_32; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3106 = 12'h22 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6178 = 12'h22 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3106; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9250 = 12'h22 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6178; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12322 = 12'h22 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9250; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15394 = 12'h22 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12322; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18466 = 12'h22 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15394; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21538 = 12'h22 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18466; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24610 = 12'h22 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21538; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_34 = io_valid_in ? _GEN_24610 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_34 = 12'h22 == _T_2[11:0] ? image_34 : _GEN_33; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3107 = 12'h23 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6179 = 12'h23 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3107; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9251 = 12'h23 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6179; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12323 = 12'h23 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9251; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15395 = 12'h23 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12323; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18467 = 12'h23 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15395; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21539 = 12'h23 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18467; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24611 = 12'h23 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21539; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_35 = io_valid_in ? _GEN_24611 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_35 = 12'h23 == _T_2[11:0] ? image_35 : _GEN_34; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3108 = 12'h24 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6180 = 12'h24 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3108; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9252 = 12'h24 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6180; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12324 = 12'h24 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9252; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15396 = 12'h24 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12324; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18468 = 12'h24 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15396; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21540 = 12'h24 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18468; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24612 = 12'h24 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21540; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_36 = io_valid_in ? _GEN_24612 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_36 = 12'h24 == _T_2[11:0] ? image_36 : _GEN_35; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3109 = 12'h25 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6181 = 12'h25 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3109; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9253 = 12'h25 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6181; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12325 = 12'h25 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9253; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15397 = 12'h25 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12325; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18469 = 12'h25 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15397; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21541 = 12'h25 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18469; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24613 = 12'h25 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21541; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_37 = io_valid_in ? _GEN_24613 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_37 = 12'h25 == _T_2[11:0] ? image_37 : _GEN_36; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3110 = 12'h26 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6182 = 12'h26 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3110; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9254 = 12'h26 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6182; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12326 = 12'h26 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9254; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15398 = 12'h26 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12326; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18470 = 12'h26 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15398; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21542 = 12'h26 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18470; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24614 = 12'h26 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21542; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_38 = io_valid_in ? _GEN_24614 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_38 = 12'h26 == _T_2[11:0] ? image_38 : _GEN_37; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3111 = 12'h27 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6183 = 12'h27 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3111; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9255 = 12'h27 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6183; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12327 = 12'h27 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9255; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15399 = 12'h27 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12327; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18471 = 12'h27 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15399; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21543 = 12'h27 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18471; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24615 = 12'h27 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21543; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_39 = io_valid_in ? _GEN_24615 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_39 = 12'h27 == _T_2[11:0] ? image_39 : _GEN_38; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3112 = 12'h28 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6184 = 12'h28 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3112; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9256 = 12'h28 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6184; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12328 = 12'h28 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9256; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15400 = 12'h28 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12328; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18472 = 12'h28 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15400; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21544 = 12'h28 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18472; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24616 = 12'h28 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21544; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_40 = io_valid_in ? _GEN_24616 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_40 = 12'h28 == _T_2[11:0] ? image_40 : _GEN_39; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3113 = 12'h29 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6185 = 12'h29 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3113; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9257 = 12'h29 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6185; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12329 = 12'h29 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9257; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15401 = 12'h29 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12329; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18473 = 12'h29 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15401; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21545 = 12'h29 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18473; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24617 = 12'h29 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21545; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_41 = io_valid_in ? _GEN_24617 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_41 = 12'h29 == _T_2[11:0] ? image_41 : _GEN_40; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3114 = 12'h2a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6186 = 12'h2a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3114; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9258 = 12'h2a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6186; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12330 = 12'h2a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9258; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15402 = 12'h2a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12330; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18474 = 12'h2a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15402; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21546 = 12'h2a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18474; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24618 = 12'h2a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21546; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_42 = io_valid_in ? _GEN_24618 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_42 = 12'h2a == _T_2[11:0] ? image_42 : _GEN_41; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3115 = 12'h2b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6187 = 12'h2b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3115; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9259 = 12'h2b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6187; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12331 = 12'h2b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9259; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15403 = 12'h2b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12331; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18475 = 12'h2b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15403; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21547 = 12'h2b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18475; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24619 = 12'h2b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21547; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_43 = io_valid_in ? _GEN_24619 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_43 = 12'h2b == _T_2[11:0] ? image_43 : _GEN_42; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3116 = 12'h2c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6188 = 12'h2c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3116; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9260 = 12'h2c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6188; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12332 = 12'h2c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9260; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15404 = 12'h2c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12332; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18476 = 12'h2c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15404; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21548 = 12'h2c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18476; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24620 = 12'h2c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21548; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_44 = io_valid_in ? _GEN_24620 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_44 = 12'h2c == _T_2[11:0] ? image_44 : _GEN_43; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3117 = 12'h2d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6189 = 12'h2d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3117; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9261 = 12'h2d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6189; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12333 = 12'h2d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9261; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15405 = 12'h2d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12333; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18477 = 12'h2d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15405; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21549 = 12'h2d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18477; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24621 = 12'h2d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21549; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_45 = io_valid_in ? _GEN_24621 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_45 = 12'h2d == _T_2[11:0] ? image_45 : _GEN_44; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3118 = 12'h2e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6190 = 12'h2e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3118; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9262 = 12'h2e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6190; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12334 = 12'h2e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9262; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15406 = 12'h2e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12334; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18478 = 12'h2e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15406; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21550 = 12'h2e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18478; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24622 = 12'h2e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21550; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_46 = io_valid_in ? _GEN_24622 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_46 = 12'h2e == _T_2[11:0] ? image_46 : _GEN_45; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3119 = 12'h2f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6191 = 12'h2f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3119; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9263 = 12'h2f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6191; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12335 = 12'h2f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9263; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15407 = 12'h2f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12335; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18479 = 12'h2f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15407; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21551 = 12'h2f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18479; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24623 = 12'h2f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21551; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_47 = io_valid_in ? _GEN_24623 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_47 = 12'h2f == _T_2[11:0] ? image_47 : _GEN_46; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3120 = 12'h30 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6192 = 12'h30 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3120; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9264 = 12'h30 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6192; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12336 = 12'h30 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9264; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15408 = 12'h30 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12336; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18480 = 12'h30 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15408; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21552 = 12'h30 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18480; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24624 = 12'h30 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21552; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_48 = io_valid_in ? _GEN_24624 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_48 = 12'h30 == _T_2[11:0] ? image_48 : _GEN_47; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3121 = 12'h31 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6193 = 12'h31 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3121; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9265 = 12'h31 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6193; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12337 = 12'h31 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9265; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15409 = 12'h31 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12337; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18481 = 12'h31 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15409; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21553 = 12'h31 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18481; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24625 = 12'h31 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21553; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_49 = io_valid_in ? _GEN_24625 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_49 = 12'h31 == _T_2[11:0] ? image_49 : _GEN_48; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3122 = 12'h32 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6194 = 12'h32 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3122; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9266 = 12'h32 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6194; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12338 = 12'h32 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9266; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15410 = 12'h32 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12338; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18482 = 12'h32 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15410; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21554 = 12'h32 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18482; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24626 = 12'h32 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21554; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_50 = io_valid_in ? _GEN_24626 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_50 = 12'h32 == _T_2[11:0] ? image_50 : _GEN_49; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3123 = 12'h33 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6195 = 12'h33 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3123; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9267 = 12'h33 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6195; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12339 = 12'h33 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9267; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15411 = 12'h33 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12339; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18483 = 12'h33 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15411; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21555 = 12'h33 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18483; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24627 = 12'h33 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21555; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_51 = io_valid_in ? _GEN_24627 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_51 = 12'h33 == _T_2[11:0] ? image_51 : _GEN_50; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3124 = 12'h34 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6196 = 12'h34 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3124; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9268 = 12'h34 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6196; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12340 = 12'h34 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9268; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15412 = 12'h34 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12340; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18484 = 12'h34 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15412; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21556 = 12'h34 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18484; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24628 = 12'h34 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21556; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_52 = io_valid_in ? _GEN_24628 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_52 = 12'h34 == _T_2[11:0] ? image_52 : _GEN_51; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3125 = 12'h35 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6197 = 12'h35 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3125; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9269 = 12'h35 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6197; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12341 = 12'h35 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9269; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15413 = 12'h35 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12341; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18485 = 12'h35 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15413; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21557 = 12'h35 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18485; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24629 = 12'h35 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21557; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_53 = io_valid_in ? _GEN_24629 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_53 = 12'h35 == _T_2[11:0] ? image_53 : _GEN_52; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3126 = 12'h36 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6198 = 12'h36 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3126; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9270 = 12'h36 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6198; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12342 = 12'h36 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9270; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15414 = 12'h36 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12342; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18486 = 12'h36 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15414; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21558 = 12'h36 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18486; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24630 = 12'h36 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21558; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_54 = io_valid_in ? _GEN_24630 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_54 = 12'h36 == _T_2[11:0] ? image_54 : _GEN_53; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3127 = 12'h37 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6199 = 12'h37 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3127; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9271 = 12'h37 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6199; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12343 = 12'h37 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9271; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15415 = 12'h37 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12343; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18487 = 12'h37 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15415; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21559 = 12'h37 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18487; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24631 = 12'h37 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21559; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_55 = io_valid_in ? _GEN_24631 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_55 = 12'h37 == _T_2[11:0] ? image_55 : _GEN_54; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3128 = 12'h38 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6200 = 12'h38 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3128; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9272 = 12'h38 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6200; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12344 = 12'h38 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9272; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15416 = 12'h38 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12344; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18488 = 12'h38 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15416; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21560 = 12'h38 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18488; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24632 = 12'h38 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21560; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_56 = io_valid_in ? _GEN_24632 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_56 = 12'h38 == _T_2[11:0] ? image_56 : _GEN_55; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3129 = 12'h39 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6201 = 12'h39 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3129; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9273 = 12'h39 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6201; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12345 = 12'h39 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9273; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15417 = 12'h39 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12345; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18489 = 12'h39 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15417; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21561 = 12'h39 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18489; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24633 = 12'h39 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21561; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_57 = io_valid_in ? _GEN_24633 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_57 = 12'h39 == _T_2[11:0] ? image_57 : _GEN_56; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3130 = 12'h3a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6202 = 12'h3a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3130; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9274 = 12'h3a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6202; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12346 = 12'h3a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9274; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15418 = 12'h3a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12346; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18490 = 12'h3a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15418; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21562 = 12'h3a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18490; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24634 = 12'h3a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21562; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_58 = io_valid_in ? _GEN_24634 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_58 = 12'h3a == _T_2[11:0] ? image_58 : _GEN_57; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3131 = 12'h3b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6203 = 12'h3b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3131; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9275 = 12'h3b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6203; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12347 = 12'h3b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9275; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15419 = 12'h3b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12347; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18491 = 12'h3b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15419; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21563 = 12'h3b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18491; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24635 = 12'h3b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21563; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_59 = io_valid_in ? _GEN_24635 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_59 = 12'h3b == _T_2[11:0] ? image_59 : _GEN_58; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3132 = 12'h3c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6204 = 12'h3c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3132; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9276 = 12'h3c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6204; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12348 = 12'h3c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9276; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15420 = 12'h3c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12348; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18492 = 12'h3c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15420; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21564 = 12'h3c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18492; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24636 = 12'h3c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21564; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_60 = io_valid_in ? _GEN_24636 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_60 = 12'h3c == _T_2[11:0] ? image_60 : _GEN_59; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3133 = 12'h3d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6205 = 12'h3d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3133; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9277 = 12'h3d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6205; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12349 = 12'h3d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9277; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15421 = 12'h3d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12349; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18493 = 12'h3d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15421; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21565 = 12'h3d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18493; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24637 = 12'h3d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21565; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_61 = io_valid_in ? _GEN_24637 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_61 = 12'h3d == _T_2[11:0] ? image_61 : _GEN_60; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3134 = 12'h3e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6206 = 12'h3e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3134; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9278 = 12'h3e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6206; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12350 = 12'h3e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9278; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15422 = 12'h3e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12350; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18494 = 12'h3e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15422; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21566 = 12'h3e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18494; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24638 = 12'h3e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21566; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_62 = io_valid_in ? _GEN_24638 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_62 = 12'h3e == _T_2[11:0] ? image_62 : _GEN_61; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3135 = 12'h3f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6207 = 12'h3f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3135; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9279 = 12'h3f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6207; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12351 = 12'h3f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9279; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15423 = 12'h3f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12351; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18495 = 12'h3f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15423; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21567 = 12'h3f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18495; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24639 = 12'h3f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21567; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_63 = io_valid_in ? _GEN_24639 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_63 = 12'h3f == _T_2[11:0] ? image_63 : _GEN_62; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3136 = 12'h40 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6208 = 12'h40 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3136; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9280 = 12'h40 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6208; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12352 = 12'h40 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9280; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15424 = 12'h40 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12352; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18496 = 12'h40 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15424; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21568 = 12'h40 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18496; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24640 = 12'h40 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21568; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_64 = io_valid_in ? _GEN_24640 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_64 = 12'h40 == _T_2[11:0] ? image_64 : _GEN_63; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3137 = 12'h41 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6209 = 12'h41 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3137; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9281 = 12'h41 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6209; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12353 = 12'h41 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9281; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15425 = 12'h41 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12353; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18497 = 12'h41 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15425; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21569 = 12'h41 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18497; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24641 = 12'h41 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21569; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_65 = io_valid_in ? _GEN_24641 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_65 = 12'h41 == _T_2[11:0] ? image_65 : _GEN_64; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3138 = 12'h42 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6210 = 12'h42 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3138; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9282 = 12'h42 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6210; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12354 = 12'h42 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9282; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15426 = 12'h42 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12354; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18498 = 12'h42 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15426; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21570 = 12'h42 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18498; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24642 = 12'h42 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21570; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_66 = io_valid_in ? _GEN_24642 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_66 = 12'h42 == _T_2[11:0] ? image_66 : _GEN_65; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3139 = 12'h43 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6211 = 12'h43 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3139; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9283 = 12'h43 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6211; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12355 = 12'h43 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9283; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15427 = 12'h43 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12355; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18499 = 12'h43 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15427; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21571 = 12'h43 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18499; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24643 = 12'h43 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21571; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_67 = io_valid_in ? _GEN_24643 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_67 = 12'h43 == _T_2[11:0] ? image_67 : _GEN_66; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3140 = 12'h44 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6212 = 12'h44 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3140; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9284 = 12'h44 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6212; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12356 = 12'h44 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9284; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15428 = 12'h44 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12356; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18500 = 12'h44 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15428; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21572 = 12'h44 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18500; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24644 = 12'h44 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21572; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_68 = io_valid_in ? _GEN_24644 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_68 = 12'h44 == _T_2[11:0] ? image_68 : _GEN_67; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3141 = 12'h45 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6213 = 12'h45 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3141; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9285 = 12'h45 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6213; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12357 = 12'h45 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9285; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15429 = 12'h45 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12357; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18501 = 12'h45 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15429; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21573 = 12'h45 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18501; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24645 = 12'h45 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21573; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_69 = io_valid_in ? _GEN_24645 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_69 = 12'h45 == _T_2[11:0] ? image_69 : _GEN_68; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3142 = 12'h46 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6214 = 12'h46 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3142; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9286 = 12'h46 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6214; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12358 = 12'h46 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9286; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15430 = 12'h46 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12358; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18502 = 12'h46 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15430; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21574 = 12'h46 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18502; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24646 = 12'h46 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21574; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_70 = io_valid_in ? _GEN_24646 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_70 = 12'h46 == _T_2[11:0] ? image_70 : _GEN_69; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3143 = 12'h47 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6215 = 12'h47 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3143; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9287 = 12'h47 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6215; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12359 = 12'h47 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9287; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15431 = 12'h47 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12359; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18503 = 12'h47 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15431; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21575 = 12'h47 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18503; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24647 = 12'h47 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21575; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_71 = io_valid_in ? _GEN_24647 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_71 = 12'h47 == _T_2[11:0] ? image_71 : _GEN_70; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3144 = 12'h48 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6216 = 12'h48 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3144; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9288 = 12'h48 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6216; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12360 = 12'h48 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9288; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15432 = 12'h48 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12360; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18504 = 12'h48 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15432; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21576 = 12'h48 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18504; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24648 = 12'h48 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21576; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_72 = io_valid_in ? _GEN_24648 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_72 = 12'h48 == _T_2[11:0] ? image_72 : _GEN_71; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3145 = 12'h49 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6217 = 12'h49 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3145; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9289 = 12'h49 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6217; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12361 = 12'h49 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9289; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15433 = 12'h49 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12361; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18505 = 12'h49 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15433; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21577 = 12'h49 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18505; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24649 = 12'h49 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21577; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_73 = io_valid_in ? _GEN_24649 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_73 = 12'h49 == _T_2[11:0] ? image_73 : _GEN_72; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3146 = 12'h4a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6218 = 12'h4a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3146; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9290 = 12'h4a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6218; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12362 = 12'h4a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9290; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15434 = 12'h4a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12362; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18506 = 12'h4a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15434; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21578 = 12'h4a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18506; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24650 = 12'h4a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21578; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_74 = io_valid_in ? _GEN_24650 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_74 = 12'h4a == _T_2[11:0] ? image_74 : _GEN_73; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3147 = 12'h4b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6219 = 12'h4b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3147; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9291 = 12'h4b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6219; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12363 = 12'h4b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9291; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15435 = 12'h4b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12363; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18507 = 12'h4b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15435; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21579 = 12'h4b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18507; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24651 = 12'h4b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21579; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_75 = io_valid_in ? _GEN_24651 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_75 = 12'h4b == _T_2[11:0] ? image_75 : _GEN_74; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3148 = 12'h4c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6220 = 12'h4c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3148; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9292 = 12'h4c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6220; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12364 = 12'h4c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9292; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15436 = 12'h4c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12364; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18508 = 12'h4c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15436; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21580 = 12'h4c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18508; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24652 = 12'h4c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21580; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_76 = io_valid_in ? _GEN_24652 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_76 = 12'h4c == _T_2[11:0] ? image_76 : _GEN_75; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3149 = 12'h4d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6221 = 12'h4d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3149; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9293 = 12'h4d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6221; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12365 = 12'h4d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9293; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15437 = 12'h4d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12365; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18509 = 12'h4d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15437; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21581 = 12'h4d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18509; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24653 = 12'h4d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21581; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_77 = io_valid_in ? _GEN_24653 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_77 = 12'h4d == _T_2[11:0] ? image_77 : _GEN_76; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3150 = 12'h4e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6222 = 12'h4e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3150; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9294 = 12'h4e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6222; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12366 = 12'h4e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9294; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15438 = 12'h4e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12366; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18510 = 12'h4e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15438; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21582 = 12'h4e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18510; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24654 = 12'h4e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21582; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_78 = io_valid_in ? _GEN_24654 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_78 = 12'h4e == _T_2[11:0] ? image_78 : _GEN_77; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3151 = 12'h4f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6223 = 12'h4f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3151; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9295 = 12'h4f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6223; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12367 = 12'h4f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9295; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15439 = 12'h4f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12367; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18511 = 12'h4f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15439; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21583 = 12'h4f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18511; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24655 = 12'h4f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21583; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_79 = io_valid_in ? _GEN_24655 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_79 = 12'h4f == _T_2[11:0] ? image_79 : _GEN_78; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3152 = 12'h50 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6224 = 12'h50 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3152; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9296 = 12'h50 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6224; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12368 = 12'h50 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9296; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15440 = 12'h50 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12368; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18512 = 12'h50 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15440; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21584 = 12'h50 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18512; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24656 = 12'h50 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21584; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_80 = io_valid_in ? _GEN_24656 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_80 = 12'h50 == _T_2[11:0] ? image_80 : _GEN_79; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3153 = 12'h51 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6225 = 12'h51 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3153; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9297 = 12'h51 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6225; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12369 = 12'h51 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9297; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15441 = 12'h51 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12369; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18513 = 12'h51 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15441; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21585 = 12'h51 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18513; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24657 = 12'h51 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21585; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_81 = io_valid_in ? _GEN_24657 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_81 = 12'h51 == _T_2[11:0] ? image_81 : _GEN_80; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3154 = 12'h52 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6226 = 12'h52 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3154; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9298 = 12'h52 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6226; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12370 = 12'h52 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9298; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15442 = 12'h52 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12370; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18514 = 12'h52 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15442; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21586 = 12'h52 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18514; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24658 = 12'h52 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21586; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_82 = io_valid_in ? _GEN_24658 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_82 = 12'h52 == _T_2[11:0] ? image_82 : _GEN_81; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3155 = 12'h53 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6227 = 12'h53 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3155; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9299 = 12'h53 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6227; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12371 = 12'h53 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9299; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15443 = 12'h53 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12371; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18515 = 12'h53 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15443; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21587 = 12'h53 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18515; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24659 = 12'h53 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21587; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_83 = io_valid_in ? _GEN_24659 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_83 = 12'h53 == _T_2[11:0] ? image_83 : _GEN_82; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3156 = 12'h54 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6228 = 12'h54 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3156; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9300 = 12'h54 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6228; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12372 = 12'h54 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9300; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15444 = 12'h54 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12372; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18516 = 12'h54 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15444; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21588 = 12'h54 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18516; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24660 = 12'h54 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21588; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_84 = io_valid_in ? _GEN_24660 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_84 = 12'h54 == _T_2[11:0] ? image_84 : _GEN_83; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3157 = 12'h55 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6229 = 12'h55 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3157; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9301 = 12'h55 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6229; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12373 = 12'h55 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9301; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15445 = 12'h55 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12373; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18517 = 12'h55 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15445; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21589 = 12'h55 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18517; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24661 = 12'h55 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21589; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_85 = io_valid_in ? _GEN_24661 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_85 = 12'h55 == _T_2[11:0] ? image_85 : _GEN_84; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3158 = 12'h56 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6230 = 12'h56 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3158; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9302 = 12'h56 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6230; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12374 = 12'h56 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9302; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15446 = 12'h56 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12374; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18518 = 12'h56 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15446; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21590 = 12'h56 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18518; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24662 = 12'h56 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21590; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_86 = io_valid_in ? _GEN_24662 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_86 = 12'h56 == _T_2[11:0] ? image_86 : _GEN_85; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3159 = 12'h57 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6231 = 12'h57 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3159; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9303 = 12'h57 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6231; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12375 = 12'h57 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9303; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15447 = 12'h57 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12375; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18519 = 12'h57 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15447; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21591 = 12'h57 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18519; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24663 = 12'h57 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21591; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_87 = io_valid_in ? _GEN_24663 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_87 = 12'h57 == _T_2[11:0] ? image_87 : _GEN_86; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3160 = 12'h58 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6232 = 12'h58 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3160; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9304 = 12'h58 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6232; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12376 = 12'h58 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9304; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15448 = 12'h58 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12376; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18520 = 12'h58 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15448; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21592 = 12'h58 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18520; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24664 = 12'h58 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21592; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_88 = io_valid_in ? _GEN_24664 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_88 = 12'h58 == _T_2[11:0] ? image_88 : _GEN_87; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3161 = 12'h59 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6233 = 12'h59 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3161; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9305 = 12'h59 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6233; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12377 = 12'h59 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9305; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15449 = 12'h59 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12377; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18521 = 12'h59 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15449; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21593 = 12'h59 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18521; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24665 = 12'h59 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21593; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_89 = io_valid_in ? _GEN_24665 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_89 = 12'h59 == _T_2[11:0] ? image_89 : _GEN_88; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3162 = 12'h5a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6234 = 12'h5a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3162; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9306 = 12'h5a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6234; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12378 = 12'h5a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9306; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15450 = 12'h5a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12378; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18522 = 12'h5a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15450; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21594 = 12'h5a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18522; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24666 = 12'h5a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21594; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_90 = io_valid_in ? _GEN_24666 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_90 = 12'h5a == _T_2[11:0] ? image_90 : _GEN_89; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3163 = 12'h5b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6235 = 12'h5b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3163; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9307 = 12'h5b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6235; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12379 = 12'h5b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9307; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15451 = 12'h5b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12379; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18523 = 12'h5b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15451; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21595 = 12'h5b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18523; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24667 = 12'h5b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21595; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_91 = io_valid_in ? _GEN_24667 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_91 = 12'h5b == _T_2[11:0] ? image_91 : _GEN_90; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3164 = 12'h5c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6236 = 12'h5c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3164; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9308 = 12'h5c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6236; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12380 = 12'h5c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9308; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15452 = 12'h5c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12380; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18524 = 12'h5c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15452; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21596 = 12'h5c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18524; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24668 = 12'h5c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21596; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_92 = io_valid_in ? _GEN_24668 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_92 = 12'h5c == _T_2[11:0] ? image_92 : _GEN_91; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3165 = 12'h5d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6237 = 12'h5d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3165; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9309 = 12'h5d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6237; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12381 = 12'h5d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9309; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15453 = 12'h5d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12381; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18525 = 12'h5d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15453; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21597 = 12'h5d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18525; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24669 = 12'h5d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21597; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_93 = io_valid_in ? _GEN_24669 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_93 = 12'h5d == _T_2[11:0] ? image_93 : _GEN_92; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3166 = 12'h5e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6238 = 12'h5e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3166; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9310 = 12'h5e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6238; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12382 = 12'h5e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9310; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15454 = 12'h5e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12382; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18526 = 12'h5e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15454; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21598 = 12'h5e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18526; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24670 = 12'h5e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21598; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_94 = io_valid_in ? _GEN_24670 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_94 = 12'h5e == _T_2[11:0] ? image_94 : _GEN_93; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3167 = 12'h5f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6239 = 12'h5f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3167; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9311 = 12'h5f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6239; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12383 = 12'h5f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9311; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15455 = 12'h5f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12383; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18527 = 12'h5f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15455; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21599 = 12'h5f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18527; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24671 = 12'h5f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21599; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_95 = io_valid_in ? _GEN_24671 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_95 = 12'h5f == _T_2[11:0] ? image_95 : _GEN_94; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3168 = 12'h60 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6240 = 12'h60 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3168; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9312 = 12'h60 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6240; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12384 = 12'h60 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9312; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15456 = 12'h60 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12384; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18528 = 12'h60 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15456; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21600 = 12'h60 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18528; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24672 = 12'h60 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21600; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_96 = io_valid_in ? _GEN_24672 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_96 = 12'h60 == _T_2[11:0] ? image_96 : _GEN_95; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3169 = 12'h61 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6241 = 12'h61 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3169; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9313 = 12'h61 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6241; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12385 = 12'h61 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9313; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15457 = 12'h61 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12385; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18529 = 12'h61 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15457; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21601 = 12'h61 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18529; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24673 = 12'h61 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21601; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_97 = io_valid_in ? _GEN_24673 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_97 = 12'h61 == _T_2[11:0] ? image_97 : _GEN_96; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3170 = 12'h62 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6242 = 12'h62 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3170; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9314 = 12'h62 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6242; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12386 = 12'h62 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9314; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15458 = 12'h62 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12386; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18530 = 12'h62 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15458; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21602 = 12'h62 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18530; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24674 = 12'h62 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21602; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_98 = io_valid_in ? _GEN_24674 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_98 = 12'h62 == _T_2[11:0] ? image_98 : _GEN_97; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3171 = 12'h63 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6243 = 12'h63 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3171; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9315 = 12'h63 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6243; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12387 = 12'h63 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9315; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15459 = 12'h63 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12387; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18531 = 12'h63 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15459; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21603 = 12'h63 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18531; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24675 = 12'h63 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21603; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_99 = io_valid_in ? _GEN_24675 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_99 = 12'h63 == _T_2[11:0] ? image_99 : _GEN_98; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3172 = 12'h64 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6244 = 12'h64 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3172; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9316 = 12'h64 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6244; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12388 = 12'h64 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9316; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15460 = 12'h64 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12388; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18532 = 12'h64 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15460; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21604 = 12'h64 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18532; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24676 = 12'h64 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21604; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_100 = io_valid_in ? _GEN_24676 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_100 = 12'h64 == _T_2[11:0] ? image_100 : _GEN_99; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3173 = 12'h65 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6245 = 12'h65 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3173; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9317 = 12'h65 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6245; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12389 = 12'h65 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9317; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15461 = 12'h65 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12389; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18533 = 12'h65 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15461; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21605 = 12'h65 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18533; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24677 = 12'h65 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21605; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_101 = io_valid_in ? _GEN_24677 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_101 = 12'h65 == _T_2[11:0] ? image_101 : _GEN_100; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3174 = 12'h66 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6246 = 12'h66 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3174; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9318 = 12'h66 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6246; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12390 = 12'h66 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9318; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15462 = 12'h66 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12390; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18534 = 12'h66 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15462; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21606 = 12'h66 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18534; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24678 = 12'h66 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21606; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_102 = io_valid_in ? _GEN_24678 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_102 = 12'h66 == _T_2[11:0] ? image_102 : _GEN_101; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3175 = 12'h67 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6247 = 12'h67 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3175; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9319 = 12'h67 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6247; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12391 = 12'h67 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9319; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15463 = 12'h67 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12391; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18535 = 12'h67 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15463; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21607 = 12'h67 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18535; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24679 = 12'h67 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21607; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_103 = io_valid_in ? _GEN_24679 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_103 = 12'h67 == _T_2[11:0] ? image_103 : _GEN_102; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3176 = 12'h68 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6248 = 12'h68 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3176; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9320 = 12'h68 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6248; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12392 = 12'h68 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9320; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15464 = 12'h68 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12392; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18536 = 12'h68 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15464; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21608 = 12'h68 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18536; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24680 = 12'h68 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21608; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_104 = io_valid_in ? _GEN_24680 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_104 = 12'h68 == _T_2[11:0] ? image_104 : _GEN_103; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3177 = 12'h69 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6249 = 12'h69 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3177; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9321 = 12'h69 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6249; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12393 = 12'h69 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9321; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15465 = 12'h69 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12393; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18537 = 12'h69 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15465; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21609 = 12'h69 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18537; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24681 = 12'h69 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21609; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_105 = io_valid_in ? _GEN_24681 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_105 = 12'h69 == _T_2[11:0] ? image_105 : _GEN_104; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3178 = 12'h6a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6250 = 12'h6a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3178; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9322 = 12'h6a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6250; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12394 = 12'h6a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9322; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15466 = 12'h6a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12394; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18538 = 12'h6a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15466; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21610 = 12'h6a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18538; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24682 = 12'h6a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21610; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_106 = io_valid_in ? _GEN_24682 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_106 = 12'h6a == _T_2[11:0] ? image_106 : _GEN_105; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3179 = 12'h6b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6251 = 12'h6b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3179; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9323 = 12'h6b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6251; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12395 = 12'h6b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9323; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15467 = 12'h6b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12395; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18539 = 12'h6b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15467; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21611 = 12'h6b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18539; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24683 = 12'h6b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21611; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_107 = io_valid_in ? _GEN_24683 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_107 = 12'h6b == _T_2[11:0] ? image_107 : _GEN_106; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3180 = 12'h6c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6252 = 12'h6c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3180; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9324 = 12'h6c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6252; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12396 = 12'h6c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9324; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15468 = 12'h6c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12396; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18540 = 12'h6c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15468; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21612 = 12'h6c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18540; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24684 = 12'h6c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21612; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_108 = io_valid_in ? _GEN_24684 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_108 = 12'h6c == _T_2[11:0] ? image_108 : _GEN_107; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3181 = 12'h6d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6253 = 12'h6d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3181; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9325 = 12'h6d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6253; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12397 = 12'h6d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9325; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15469 = 12'h6d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12397; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18541 = 12'h6d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15469; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21613 = 12'h6d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18541; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24685 = 12'h6d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21613; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_109 = io_valid_in ? _GEN_24685 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_109 = 12'h6d == _T_2[11:0] ? image_109 : _GEN_108; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3182 = 12'h6e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6254 = 12'h6e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3182; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9326 = 12'h6e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6254; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12398 = 12'h6e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9326; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15470 = 12'h6e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12398; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18542 = 12'h6e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15470; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21614 = 12'h6e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18542; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24686 = 12'h6e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21614; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_110 = io_valid_in ? _GEN_24686 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_110 = 12'h6e == _T_2[11:0] ? image_110 : _GEN_109; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3183 = 12'h6f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6255 = 12'h6f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3183; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9327 = 12'h6f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6255; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12399 = 12'h6f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9327; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15471 = 12'h6f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12399; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18543 = 12'h6f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15471; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21615 = 12'h6f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18543; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24687 = 12'h6f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21615; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_111 = io_valid_in ? _GEN_24687 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_111 = 12'h6f == _T_2[11:0] ? image_111 : _GEN_110; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3184 = 12'h70 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6256 = 12'h70 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3184; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9328 = 12'h70 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6256; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12400 = 12'h70 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9328; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15472 = 12'h70 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12400; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18544 = 12'h70 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15472; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21616 = 12'h70 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18544; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24688 = 12'h70 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21616; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_112 = io_valid_in ? _GEN_24688 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_112 = 12'h70 == _T_2[11:0] ? image_112 : _GEN_111; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3185 = 12'h71 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6257 = 12'h71 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3185; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9329 = 12'h71 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6257; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12401 = 12'h71 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9329; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15473 = 12'h71 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12401; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18545 = 12'h71 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15473; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21617 = 12'h71 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18545; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24689 = 12'h71 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21617; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_113 = io_valid_in ? _GEN_24689 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_113 = 12'h71 == _T_2[11:0] ? image_113 : _GEN_112; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3186 = 12'h72 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6258 = 12'h72 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3186; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9330 = 12'h72 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6258; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12402 = 12'h72 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9330; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15474 = 12'h72 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12402; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18546 = 12'h72 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15474; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21618 = 12'h72 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18546; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24690 = 12'h72 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21618; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_114 = io_valid_in ? _GEN_24690 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_114 = 12'h72 == _T_2[11:0] ? image_114 : _GEN_113; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3187 = 12'h73 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6259 = 12'h73 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3187; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9331 = 12'h73 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6259; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12403 = 12'h73 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9331; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15475 = 12'h73 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12403; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18547 = 12'h73 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15475; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21619 = 12'h73 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18547; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24691 = 12'h73 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21619; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_115 = io_valid_in ? _GEN_24691 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_115 = 12'h73 == _T_2[11:0] ? image_115 : _GEN_114; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3188 = 12'h74 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6260 = 12'h74 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3188; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9332 = 12'h74 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6260; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12404 = 12'h74 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9332; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15476 = 12'h74 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12404; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18548 = 12'h74 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15476; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21620 = 12'h74 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18548; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24692 = 12'h74 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21620; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_116 = io_valid_in ? _GEN_24692 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_116 = 12'h74 == _T_2[11:0] ? image_116 : _GEN_115; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3189 = 12'h75 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6261 = 12'h75 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3189; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9333 = 12'h75 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6261; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12405 = 12'h75 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9333; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15477 = 12'h75 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12405; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18549 = 12'h75 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15477; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21621 = 12'h75 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18549; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24693 = 12'h75 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21621; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_117 = io_valid_in ? _GEN_24693 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_117 = 12'h75 == _T_2[11:0] ? image_117 : _GEN_116; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3190 = 12'h76 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6262 = 12'h76 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3190; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9334 = 12'h76 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6262; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12406 = 12'h76 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9334; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15478 = 12'h76 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12406; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18550 = 12'h76 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15478; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21622 = 12'h76 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18550; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24694 = 12'h76 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21622; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_118 = io_valid_in ? _GEN_24694 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_118 = 12'h76 == _T_2[11:0] ? image_118 : _GEN_117; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3191 = 12'h77 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6263 = 12'h77 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3191; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9335 = 12'h77 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6263; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12407 = 12'h77 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9335; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15479 = 12'h77 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12407; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18551 = 12'h77 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15479; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21623 = 12'h77 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18551; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24695 = 12'h77 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21623; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_119 = io_valid_in ? _GEN_24695 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_119 = 12'h77 == _T_2[11:0] ? image_119 : _GEN_118; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3192 = 12'h78 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6264 = 12'h78 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3192; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9336 = 12'h78 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6264; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12408 = 12'h78 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9336; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15480 = 12'h78 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12408; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18552 = 12'h78 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15480; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21624 = 12'h78 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18552; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24696 = 12'h78 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21624; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_120 = io_valid_in ? _GEN_24696 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_120 = 12'h78 == _T_2[11:0] ? image_120 : _GEN_119; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3193 = 12'h79 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6265 = 12'h79 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3193; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9337 = 12'h79 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6265; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12409 = 12'h79 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9337; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15481 = 12'h79 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12409; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18553 = 12'h79 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15481; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21625 = 12'h79 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18553; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24697 = 12'h79 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21625; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_121 = io_valid_in ? _GEN_24697 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_121 = 12'h79 == _T_2[11:0] ? image_121 : _GEN_120; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3194 = 12'h7a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6266 = 12'h7a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3194; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9338 = 12'h7a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6266; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12410 = 12'h7a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9338; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15482 = 12'h7a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12410; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18554 = 12'h7a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15482; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21626 = 12'h7a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18554; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24698 = 12'h7a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21626; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_122 = io_valid_in ? _GEN_24698 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_122 = 12'h7a == _T_2[11:0] ? image_122 : _GEN_121; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3195 = 12'h7b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6267 = 12'h7b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3195; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9339 = 12'h7b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6267; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12411 = 12'h7b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9339; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15483 = 12'h7b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12411; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18555 = 12'h7b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15483; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21627 = 12'h7b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18555; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24699 = 12'h7b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21627; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_123 = io_valid_in ? _GEN_24699 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_123 = 12'h7b == _T_2[11:0] ? image_123 : _GEN_122; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3196 = 12'h7c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6268 = 12'h7c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3196; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9340 = 12'h7c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6268; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12412 = 12'h7c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9340; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15484 = 12'h7c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12412; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18556 = 12'h7c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15484; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21628 = 12'h7c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18556; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24700 = 12'h7c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21628; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_124 = io_valid_in ? _GEN_24700 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_124 = 12'h7c == _T_2[11:0] ? image_124 : _GEN_123; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3197 = 12'h7d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6269 = 12'h7d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3197; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9341 = 12'h7d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6269; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12413 = 12'h7d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9341; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15485 = 12'h7d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12413; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18557 = 12'h7d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15485; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21629 = 12'h7d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18557; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24701 = 12'h7d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21629; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_125 = io_valid_in ? _GEN_24701 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_125 = 12'h7d == _T_2[11:0] ? image_125 : _GEN_124; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3198 = 12'h7e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6270 = 12'h7e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3198; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9342 = 12'h7e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6270; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12414 = 12'h7e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9342; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15486 = 12'h7e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12414; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18558 = 12'h7e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15486; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21630 = 12'h7e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18558; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24702 = 12'h7e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21630; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_126 = io_valid_in ? _GEN_24702 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_126 = 12'h7e == _T_2[11:0] ? image_126 : _GEN_125; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3199 = 12'h7f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6271 = 12'h7f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3199; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9343 = 12'h7f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6271; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12415 = 12'h7f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9343; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15487 = 12'h7f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12415; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18559 = 12'h7f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15487; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21631 = 12'h7f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18559; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24703 = 12'h7f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21631; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_127 = io_valid_in ? _GEN_24703 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_127 = 12'h7f == _T_2[11:0] ? image_127 : _GEN_126; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3200 = 12'h80 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6272 = 12'h80 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3200; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9344 = 12'h80 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6272; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12416 = 12'h80 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9344; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15488 = 12'h80 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12416; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18560 = 12'h80 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15488; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21632 = 12'h80 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18560; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24704 = 12'h80 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21632; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_128 = io_valid_in ? _GEN_24704 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_128 = 12'h80 == _T_2[11:0] ? image_128 : _GEN_127; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3201 = 12'h81 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6273 = 12'h81 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3201; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9345 = 12'h81 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6273; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12417 = 12'h81 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9345; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15489 = 12'h81 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12417; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18561 = 12'h81 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15489; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21633 = 12'h81 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18561; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24705 = 12'h81 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21633; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_129 = io_valid_in ? _GEN_24705 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_129 = 12'h81 == _T_2[11:0] ? image_129 : _GEN_128; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3202 = 12'h82 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6274 = 12'h82 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3202; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9346 = 12'h82 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6274; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12418 = 12'h82 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9346; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15490 = 12'h82 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12418; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18562 = 12'h82 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15490; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21634 = 12'h82 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18562; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24706 = 12'h82 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21634; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_130 = io_valid_in ? _GEN_24706 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_130 = 12'h82 == _T_2[11:0] ? image_130 : _GEN_129; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3203 = 12'h83 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6275 = 12'h83 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3203; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9347 = 12'h83 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6275; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12419 = 12'h83 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9347; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15491 = 12'h83 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12419; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18563 = 12'h83 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15491; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21635 = 12'h83 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18563; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24707 = 12'h83 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21635; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_131 = io_valid_in ? _GEN_24707 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_131 = 12'h83 == _T_2[11:0] ? image_131 : _GEN_130; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3204 = 12'h84 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6276 = 12'h84 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3204; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9348 = 12'h84 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6276; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12420 = 12'h84 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9348; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15492 = 12'h84 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12420; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18564 = 12'h84 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15492; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21636 = 12'h84 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18564; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24708 = 12'h84 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21636; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_132 = io_valid_in ? _GEN_24708 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_132 = 12'h84 == _T_2[11:0] ? image_132 : _GEN_131; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3205 = 12'h85 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6277 = 12'h85 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3205; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9349 = 12'h85 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6277; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12421 = 12'h85 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9349; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15493 = 12'h85 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12421; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18565 = 12'h85 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15493; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21637 = 12'h85 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18565; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24709 = 12'h85 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21637; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_133 = io_valid_in ? _GEN_24709 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_133 = 12'h85 == _T_2[11:0] ? image_133 : _GEN_132; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3206 = 12'h86 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6278 = 12'h86 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3206; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9350 = 12'h86 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6278; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12422 = 12'h86 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9350; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15494 = 12'h86 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12422; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18566 = 12'h86 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15494; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21638 = 12'h86 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18566; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24710 = 12'h86 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21638; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_134 = io_valid_in ? _GEN_24710 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_134 = 12'h86 == _T_2[11:0] ? image_134 : _GEN_133; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3207 = 12'h87 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6279 = 12'h87 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3207; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9351 = 12'h87 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6279; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12423 = 12'h87 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9351; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15495 = 12'h87 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12423; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18567 = 12'h87 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15495; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21639 = 12'h87 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18567; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24711 = 12'h87 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21639; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_135 = io_valid_in ? _GEN_24711 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_135 = 12'h87 == _T_2[11:0] ? image_135 : _GEN_134; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3208 = 12'h88 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6280 = 12'h88 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3208; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9352 = 12'h88 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6280; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12424 = 12'h88 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9352; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15496 = 12'h88 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12424; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18568 = 12'h88 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15496; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21640 = 12'h88 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18568; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24712 = 12'h88 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21640; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_136 = io_valid_in ? _GEN_24712 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_136 = 12'h88 == _T_2[11:0] ? image_136 : _GEN_135; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3209 = 12'h89 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6281 = 12'h89 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3209; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9353 = 12'h89 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6281; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12425 = 12'h89 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9353; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15497 = 12'h89 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12425; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18569 = 12'h89 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15497; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21641 = 12'h89 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18569; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24713 = 12'h89 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21641; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_137 = io_valid_in ? _GEN_24713 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_137 = 12'h89 == _T_2[11:0] ? image_137 : _GEN_136; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3210 = 12'h8a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6282 = 12'h8a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3210; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9354 = 12'h8a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6282; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12426 = 12'h8a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9354; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15498 = 12'h8a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12426; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18570 = 12'h8a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15498; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21642 = 12'h8a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18570; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24714 = 12'h8a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21642; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_138 = io_valid_in ? _GEN_24714 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_138 = 12'h8a == _T_2[11:0] ? image_138 : _GEN_137; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3211 = 12'h8b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6283 = 12'h8b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3211; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9355 = 12'h8b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6283; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12427 = 12'h8b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9355; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15499 = 12'h8b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12427; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18571 = 12'h8b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15499; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21643 = 12'h8b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18571; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24715 = 12'h8b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21643; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_139 = io_valid_in ? _GEN_24715 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_139 = 12'h8b == _T_2[11:0] ? image_139 : _GEN_138; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3212 = 12'h8c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6284 = 12'h8c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3212; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9356 = 12'h8c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6284; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12428 = 12'h8c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9356; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15500 = 12'h8c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12428; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18572 = 12'h8c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15500; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21644 = 12'h8c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18572; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24716 = 12'h8c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21644; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_140 = io_valid_in ? _GEN_24716 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_140 = 12'h8c == _T_2[11:0] ? image_140 : _GEN_139; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3213 = 12'h8d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6285 = 12'h8d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3213; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9357 = 12'h8d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6285; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12429 = 12'h8d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9357; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15501 = 12'h8d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12429; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18573 = 12'h8d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15501; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21645 = 12'h8d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18573; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24717 = 12'h8d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21645; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_141 = io_valid_in ? _GEN_24717 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_141 = 12'h8d == _T_2[11:0] ? image_141 : _GEN_140; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3214 = 12'h8e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6286 = 12'h8e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3214; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9358 = 12'h8e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6286; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12430 = 12'h8e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9358; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15502 = 12'h8e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12430; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18574 = 12'h8e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15502; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21646 = 12'h8e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18574; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24718 = 12'h8e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21646; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_142 = io_valid_in ? _GEN_24718 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_142 = 12'h8e == _T_2[11:0] ? image_142 : _GEN_141; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3215 = 12'h8f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6287 = 12'h8f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3215; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9359 = 12'h8f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6287; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12431 = 12'h8f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9359; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15503 = 12'h8f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12431; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18575 = 12'h8f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15503; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21647 = 12'h8f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18575; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24719 = 12'h8f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21647; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_143 = io_valid_in ? _GEN_24719 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_143 = 12'h8f == _T_2[11:0] ? image_143 : _GEN_142; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3216 = 12'h90 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6288 = 12'h90 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3216; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9360 = 12'h90 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6288; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12432 = 12'h90 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9360; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15504 = 12'h90 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12432; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18576 = 12'h90 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15504; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21648 = 12'h90 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18576; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24720 = 12'h90 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21648; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_144 = io_valid_in ? _GEN_24720 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_144 = 12'h90 == _T_2[11:0] ? image_144 : _GEN_143; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3217 = 12'h91 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6289 = 12'h91 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3217; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9361 = 12'h91 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6289; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12433 = 12'h91 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9361; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15505 = 12'h91 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12433; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18577 = 12'h91 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15505; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21649 = 12'h91 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18577; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24721 = 12'h91 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21649; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_145 = io_valid_in ? _GEN_24721 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_145 = 12'h91 == _T_2[11:0] ? image_145 : _GEN_144; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3218 = 12'h92 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6290 = 12'h92 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3218; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9362 = 12'h92 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6290; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12434 = 12'h92 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9362; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15506 = 12'h92 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12434; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18578 = 12'h92 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15506; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21650 = 12'h92 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18578; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24722 = 12'h92 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21650; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_146 = io_valid_in ? _GEN_24722 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_146 = 12'h92 == _T_2[11:0] ? image_146 : _GEN_145; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3219 = 12'h93 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6291 = 12'h93 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3219; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9363 = 12'h93 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6291; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12435 = 12'h93 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9363; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15507 = 12'h93 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12435; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18579 = 12'h93 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15507; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21651 = 12'h93 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18579; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24723 = 12'h93 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21651; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_147 = io_valid_in ? _GEN_24723 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_147 = 12'h93 == _T_2[11:0] ? image_147 : _GEN_146; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3220 = 12'h94 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6292 = 12'h94 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3220; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9364 = 12'h94 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6292; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12436 = 12'h94 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9364; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15508 = 12'h94 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12436; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18580 = 12'h94 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15508; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21652 = 12'h94 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18580; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24724 = 12'h94 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21652; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_148 = io_valid_in ? _GEN_24724 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_148 = 12'h94 == _T_2[11:0] ? image_148 : _GEN_147; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3221 = 12'h95 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6293 = 12'h95 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3221; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9365 = 12'h95 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6293; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12437 = 12'h95 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9365; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15509 = 12'h95 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12437; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18581 = 12'h95 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15509; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21653 = 12'h95 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18581; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24725 = 12'h95 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21653; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_149 = io_valid_in ? _GEN_24725 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_149 = 12'h95 == _T_2[11:0] ? image_149 : _GEN_148; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3222 = 12'h96 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6294 = 12'h96 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3222; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9366 = 12'h96 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6294; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12438 = 12'h96 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9366; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15510 = 12'h96 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12438; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18582 = 12'h96 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15510; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21654 = 12'h96 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18582; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24726 = 12'h96 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21654; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_150 = io_valid_in ? _GEN_24726 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_150 = 12'h96 == _T_2[11:0] ? image_150 : _GEN_149; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3223 = 12'h97 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6295 = 12'h97 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3223; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9367 = 12'h97 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6295; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12439 = 12'h97 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9367; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15511 = 12'h97 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12439; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18583 = 12'h97 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15511; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21655 = 12'h97 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18583; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24727 = 12'h97 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21655; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_151 = io_valid_in ? _GEN_24727 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_151 = 12'h97 == _T_2[11:0] ? image_151 : _GEN_150; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3224 = 12'h98 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6296 = 12'h98 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3224; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9368 = 12'h98 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6296; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12440 = 12'h98 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9368; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15512 = 12'h98 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12440; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18584 = 12'h98 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15512; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21656 = 12'h98 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18584; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24728 = 12'h98 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21656; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_152 = io_valid_in ? _GEN_24728 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_152 = 12'h98 == _T_2[11:0] ? image_152 : _GEN_151; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3225 = 12'h99 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6297 = 12'h99 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3225; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9369 = 12'h99 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6297; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12441 = 12'h99 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9369; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15513 = 12'h99 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12441; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18585 = 12'h99 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15513; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21657 = 12'h99 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18585; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24729 = 12'h99 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21657; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_153 = io_valid_in ? _GEN_24729 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_153 = 12'h99 == _T_2[11:0] ? image_153 : _GEN_152; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3226 = 12'h9a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6298 = 12'h9a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3226; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9370 = 12'h9a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6298; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12442 = 12'h9a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9370; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15514 = 12'h9a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12442; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18586 = 12'h9a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15514; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21658 = 12'h9a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18586; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24730 = 12'h9a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21658; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_154 = io_valid_in ? _GEN_24730 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_154 = 12'h9a == _T_2[11:0] ? image_154 : _GEN_153; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3227 = 12'h9b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6299 = 12'h9b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3227; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9371 = 12'h9b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6299; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12443 = 12'h9b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9371; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15515 = 12'h9b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12443; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18587 = 12'h9b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15515; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21659 = 12'h9b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18587; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24731 = 12'h9b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21659; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_155 = io_valid_in ? _GEN_24731 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_155 = 12'h9b == _T_2[11:0] ? image_155 : _GEN_154; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3228 = 12'h9c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6300 = 12'h9c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3228; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9372 = 12'h9c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6300; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12444 = 12'h9c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9372; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15516 = 12'h9c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12444; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18588 = 12'h9c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15516; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21660 = 12'h9c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18588; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24732 = 12'h9c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21660; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_156 = io_valid_in ? _GEN_24732 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_156 = 12'h9c == _T_2[11:0] ? image_156 : _GEN_155; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3229 = 12'h9d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6301 = 12'h9d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3229; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9373 = 12'h9d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6301; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12445 = 12'h9d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9373; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15517 = 12'h9d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12445; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18589 = 12'h9d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15517; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21661 = 12'h9d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18589; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24733 = 12'h9d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21661; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_157 = io_valid_in ? _GEN_24733 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_157 = 12'h9d == _T_2[11:0] ? image_157 : _GEN_156; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3230 = 12'h9e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6302 = 12'h9e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3230; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9374 = 12'h9e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6302; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12446 = 12'h9e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9374; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15518 = 12'h9e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12446; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18590 = 12'h9e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15518; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21662 = 12'h9e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18590; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24734 = 12'h9e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21662; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_158 = io_valid_in ? _GEN_24734 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_158 = 12'h9e == _T_2[11:0] ? image_158 : _GEN_157; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3231 = 12'h9f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6303 = 12'h9f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3231; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9375 = 12'h9f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6303; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12447 = 12'h9f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9375; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15519 = 12'h9f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12447; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18591 = 12'h9f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15519; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21663 = 12'h9f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18591; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24735 = 12'h9f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21663; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_159 = io_valid_in ? _GEN_24735 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_159 = 12'h9f == _T_2[11:0] ? image_159 : _GEN_158; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3232 = 12'ha0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6304 = 12'ha0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3232; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9376 = 12'ha0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6304; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12448 = 12'ha0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9376; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15520 = 12'ha0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12448; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18592 = 12'ha0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15520; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21664 = 12'ha0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18592; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24736 = 12'ha0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21664; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_160 = io_valid_in ? _GEN_24736 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_160 = 12'ha0 == _T_2[11:0] ? image_160 : _GEN_159; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3233 = 12'ha1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6305 = 12'ha1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3233; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9377 = 12'ha1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6305; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12449 = 12'ha1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9377; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15521 = 12'ha1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12449; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18593 = 12'ha1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15521; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21665 = 12'ha1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18593; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24737 = 12'ha1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21665; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_161 = io_valid_in ? _GEN_24737 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_161 = 12'ha1 == _T_2[11:0] ? image_161 : _GEN_160; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3234 = 12'ha2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6306 = 12'ha2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3234; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9378 = 12'ha2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6306; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12450 = 12'ha2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9378; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15522 = 12'ha2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12450; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18594 = 12'ha2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15522; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21666 = 12'ha2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18594; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24738 = 12'ha2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21666; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_162 = io_valid_in ? _GEN_24738 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_162 = 12'ha2 == _T_2[11:0] ? image_162 : _GEN_161; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3235 = 12'ha3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6307 = 12'ha3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3235; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9379 = 12'ha3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6307; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12451 = 12'ha3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9379; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15523 = 12'ha3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12451; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18595 = 12'ha3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15523; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21667 = 12'ha3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18595; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24739 = 12'ha3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21667; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_163 = io_valid_in ? _GEN_24739 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_163 = 12'ha3 == _T_2[11:0] ? image_163 : _GEN_162; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3236 = 12'ha4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6308 = 12'ha4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3236; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9380 = 12'ha4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6308; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12452 = 12'ha4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9380; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15524 = 12'ha4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12452; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18596 = 12'ha4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15524; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21668 = 12'ha4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18596; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24740 = 12'ha4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21668; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_164 = io_valid_in ? _GEN_24740 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_164 = 12'ha4 == _T_2[11:0] ? image_164 : _GEN_163; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3237 = 12'ha5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6309 = 12'ha5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3237; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9381 = 12'ha5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6309; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12453 = 12'ha5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9381; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15525 = 12'ha5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12453; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18597 = 12'ha5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15525; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21669 = 12'ha5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18597; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24741 = 12'ha5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21669; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_165 = io_valid_in ? _GEN_24741 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_165 = 12'ha5 == _T_2[11:0] ? image_165 : _GEN_164; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3238 = 12'ha6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6310 = 12'ha6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3238; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9382 = 12'ha6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6310; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12454 = 12'ha6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9382; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15526 = 12'ha6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12454; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18598 = 12'ha6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15526; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21670 = 12'ha6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18598; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24742 = 12'ha6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21670; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_166 = io_valid_in ? _GEN_24742 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_166 = 12'ha6 == _T_2[11:0] ? image_166 : _GEN_165; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3239 = 12'ha7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6311 = 12'ha7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3239; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9383 = 12'ha7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6311; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12455 = 12'ha7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9383; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15527 = 12'ha7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12455; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18599 = 12'ha7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15527; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21671 = 12'ha7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18599; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24743 = 12'ha7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21671; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_167 = io_valid_in ? _GEN_24743 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_167 = 12'ha7 == _T_2[11:0] ? image_167 : _GEN_166; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3240 = 12'ha8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6312 = 12'ha8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3240; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9384 = 12'ha8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6312; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12456 = 12'ha8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9384; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15528 = 12'ha8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12456; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18600 = 12'ha8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15528; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21672 = 12'ha8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18600; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24744 = 12'ha8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21672; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_168 = io_valid_in ? _GEN_24744 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_168 = 12'ha8 == _T_2[11:0] ? image_168 : _GEN_167; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3241 = 12'ha9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6313 = 12'ha9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3241; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9385 = 12'ha9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6313; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12457 = 12'ha9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9385; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15529 = 12'ha9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12457; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18601 = 12'ha9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15529; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21673 = 12'ha9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18601; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24745 = 12'ha9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21673; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_169 = io_valid_in ? _GEN_24745 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_169 = 12'ha9 == _T_2[11:0] ? image_169 : _GEN_168; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3242 = 12'haa == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6314 = 12'haa == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3242; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9386 = 12'haa == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6314; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12458 = 12'haa == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9386; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15530 = 12'haa == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12458; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18602 = 12'haa == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15530; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21674 = 12'haa == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18602; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24746 = 12'haa == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21674; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_170 = io_valid_in ? _GEN_24746 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_170 = 12'haa == _T_2[11:0] ? image_170 : _GEN_169; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3243 = 12'hab == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6315 = 12'hab == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3243; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9387 = 12'hab == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6315; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12459 = 12'hab == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9387; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15531 = 12'hab == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12459; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18603 = 12'hab == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15531; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21675 = 12'hab == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18603; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24747 = 12'hab == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21675; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_171 = io_valid_in ? _GEN_24747 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_171 = 12'hab == _T_2[11:0] ? image_171 : _GEN_170; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3244 = 12'hac == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6316 = 12'hac == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3244; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9388 = 12'hac == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6316; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12460 = 12'hac == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9388; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15532 = 12'hac == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12460; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18604 = 12'hac == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15532; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21676 = 12'hac == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18604; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24748 = 12'hac == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21676; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_172 = io_valid_in ? _GEN_24748 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_172 = 12'hac == _T_2[11:0] ? image_172 : _GEN_171; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3245 = 12'had == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6317 = 12'had == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3245; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9389 = 12'had == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6317; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12461 = 12'had == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9389; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15533 = 12'had == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12461; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18605 = 12'had == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15533; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21677 = 12'had == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18605; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24749 = 12'had == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21677; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_173 = io_valid_in ? _GEN_24749 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_173 = 12'had == _T_2[11:0] ? image_173 : _GEN_172; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3246 = 12'hae == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6318 = 12'hae == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3246; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9390 = 12'hae == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6318; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12462 = 12'hae == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9390; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15534 = 12'hae == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12462; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18606 = 12'hae == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15534; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21678 = 12'hae == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18606; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24750 = 12'hae == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21678; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_174 = io_valid_in ? _GEN_24750 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_174 = 12'hae == _T_2[11:0] ? image_174 : _GEN_173; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3247 = 12'haf == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6319 = 12'haf == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3247; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9391 = 12'haf == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6319; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12463 = 12'haf == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9391; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15535 = 12'haf == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12463; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18607 = 12'haf == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15535; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21679 = 12'haf == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18607; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24751 = 12'haf == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21679; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_175 = io_valid_in ? _GEN_24751 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_175 = 12'haf == _T_2[11:0] ? image_175 : _GEN_174; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3248 = 12'hb0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6320 = 12'hb0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3248; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9392 = 12'hb0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6320; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12464 = 12'hb0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9392; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15536 = 12'hb0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12464; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18608 = 12'hb0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15536; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21680 = 12'hb0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18608; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24752 = 12'hb0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21680; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_176 = io_valid_in ? _GEN_24752 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_176 = 12'hb0 == _T_2[11:0] ? image_176 : _GEN_175; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3249 = 12'hb1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6321 = 12'hb1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3249; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9393 = 12'hb1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6321; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12465 = 12'hb1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9393; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15537 = 12'hb1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12465; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18609 = 12'hb1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15537; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21681 = 12'hb1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18609; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24753 = 12'hb1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21681; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_177 = io_valid_in ? _GEN_24753 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_177 = 12'hb1 == _T_2[11:0] ? image_177 : _GEN_176; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3250 = 12'hb2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6322 = 12'hb2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3250; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9394 = 12'hb2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6322; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12466 = 12'hb2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9394; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15538 = 12'hb2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12466; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18610 = 12'hb2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15538; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21682 = 12'hb2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18610; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24754 = 12'hb2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21682; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_178 = io_valid_in ? _GEN_24754 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_178 = 12'hb2 == _T_2[11:0] ? image_178 : _GEN_177; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3251 = 12'hb3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6323 = 12'hb3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3251; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9395 = 12'hb3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6323; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12467 = 12'hb3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9395; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15539 = 12'hb3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12467; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18611 = 12'hb3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15539; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21683 = 12'hb3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18611; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24755 = 12'hb3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21683; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_179 = io_valid_in ? _GEN_24755 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_179 = 12'hb3 == _T_2[11:0] ? image_179 : _GEN_178; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3252 = 12'hb4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6324 = 12'hb4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3252; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9396 = 12'hb4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6324; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12468 = 12'hb4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9396; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15540 = 12'hb4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12468; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18612 = 12'hb4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15540; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21684 = 12'hb4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18612; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24756 = 12'hb4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21684; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_180 = io_valid_in ? _GEN_24756 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_180 = 12'hb4 == _T_2[11:0] ? image_180 : _GEN_179; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3253 = 12'hb5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6325 = 12'hb5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3253; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9397 = 12'hb5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6325; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12469 = 12'hb5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9397; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15541 = 12'hb5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12469; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18613 = 12'hb5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15541; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21685 = 12'hb5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18613; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24757 = 12'hb5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21685; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_181 = io_valid_in ? _GEN_24757 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_181 = 12'hb5 == _T_2[11:0] ? image_181 : _GEN_180; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3254 = 12'hb6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6326 = 12'hb6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3254; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9398 = 12'hb6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6326; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12470 = 12'hb6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9398; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15542 = 12'hb6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12470; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18614 = 12'hb6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15542; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21686 = 12'hb6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18614; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24758 = 12'hb6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21686; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_182 = io_valid_in ? _GEN_24758 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_182 = 12'hb6 == _T_2[11:0] ? image_182 : _GEN_181; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3255 = 12'hb7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6327 = 12'hb7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3255; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9399 = 12'hb7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6327; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12471 = 12'hb7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9399; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15543 = 12'hb7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12471; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18615 = 12'hb7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15543; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21687 = 12'hb7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18615; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24759 = 12'hb7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21687; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_183 = io_valid_in ? _GEN_24759 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_183 = 12'hb7 == _T_2[11:0] ? image_183 : _GEN_182; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3256 = 12'hb8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6328 = 12'hb8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3256; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9400 = 12'hb8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6328; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12472 = 12'hb8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9400; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15544 = 12'hb8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12472; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18616 = 12'hb8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15544; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21688 = 12'hb8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18616; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24760 = 12'hb8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21688; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_184 = io_valid_in ? _GEN_24760 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_184 = 12'hb8 == _T_2[11:0] ? image_184 : _GEN_183; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3257 = 12'hb9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6329 = 12'hb9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3257; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9401 = 12'hb9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6329; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12473 = 12'hb9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9401; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15545 = 12'hb9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12473; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18617 = 12'hb9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15545; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21689 = 12'hb9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18617; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24761 = 12'hb9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21689; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_185 = io_valid_in ? _GEN_24761 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_185 = 12'hb9 == _T_2[11:0] ? image_185 : _GEN_184; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3258 = 12'hba == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6330 = 12'hba == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3258; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9402 = 12'hba == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6330; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12474 = 12'hba == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9402; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15546 = 12'hba == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12474; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18618 = 12'hba == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15546; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21690 = 12'hba == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18618; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24762 = 12'hba == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21690; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_186 = io_valid_in ? _GEN_24762 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_186 = 12'hba == _T_2[11:0] ? image_186 : _GEN_185; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3259 = 12'hbb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6331 = 12'hbb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3259; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9403 = 12'hbb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6331; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12475 = 12'hbb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9403; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15547 = 12'hbb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12475; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18619 = 12'hbb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15547; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21691 = 12'hbb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18619; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24763 = 12'hbb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21691; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_187 = io_valid_in ? _GEN_24763 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_187 = 12'hbb == _T_2[11:0] ? image_187 : _GEN_186; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3260 = 12'hbc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6332 = 12'hbc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3260; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9404 = 12'hbc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6332; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12476 = 12'hbc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9404; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15548 = 12'hbc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12476; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18620 = 12'hbc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15548; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21692 = 12'hbc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18620; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24764 = 12'hbc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21692; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_188 = io_valid_in ? _GEN_24764 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_188 = 12'hbc == _T_2[11:0] ? image_188 : _GEN_187; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3261 = 12'hbd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6333 = 12'hbd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3261; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9405 = 12'hbd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6333; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12477 = 12'hbd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9405; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15549 = 12'hbd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12477; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18621 = 12'hbd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15549; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21693 = 12'hbd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18621; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24765 = 12'hbd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21693; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_189 = io_valid_in ? _GEN_24765 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_189 = 12'hbd == _T_2[11:0] ? image_189 : _GEN_188; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3262 = 12'hbe == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6334 = 12'hbe == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3262; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9406 = 12'hbe == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6334; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12478 = 12'hbe == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9406; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15550 = 12'hbe == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12478; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18622 = 12'hbe == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15550; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21694 = 12'hbe == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18622; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24766 = 12'hbe == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21694; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_190 = io_valid_in ? _GEN_24766 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_190 = 12'hbe == _T_2[11:0] ? image_190 : _GEN_189; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3263 = 12'hbf == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6335 = 12'hbf == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3263; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9407 = 12'hbf == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6335; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12479 = 12'hbf == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9407; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15551 = 12'hbf == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12479; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18623 = 12'hbf == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15551; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21695 = 12'hbf == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18623; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24767 = 12'hbf == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21695; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_191 = io_valid_in ? _GEN_24767 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_191 = 12'hbf == _T_2[11:0] ? image_191 : _GEN_190; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3264 = 12'hc0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6336 = 12'hc0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3264; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9408 = 12'hc0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6336; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12480 = 12'hc0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9408; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15552 = 12'hc0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12480; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18624 = 12'hc0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15552; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21696 = 12'hc0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18624; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24768 = 12'hc0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21696; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_192 = io_valid_in ? _GEN_24768 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_192 = 12'hc0 == _T_2[11:0] ? image_192 : _GEN_191; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3265 = 12'hc1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6337 = 12'hc1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3265; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9409 = 12'hc1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6337; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12481 = 12'hc1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9409; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15553 = 12'hc1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12481; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18625 = 12'hc1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15553; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21697 = 12'hc1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18625; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24769 = 12'hc1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21697; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_193 = io_valid_in ? _GEN_24769 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_193 = 12'hc1 == _T_2[11:0] ? image_193 : _GEN_192; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3266 = 12'hc2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6338 = 12'hc2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3266; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9410 = 12'hc2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6338; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12482 = 12'hc2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9410; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15554 = 12'hc2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12482; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18626 = 12'hc2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15554; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21698 = 12'hc2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18626; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24770 = 12'hc2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21698; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_194 = io_valid_in ? _GEN_24770 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_194 = 12'hc2 == _T_2[11:0] ? image_194 : _GEN_193; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3267 = 12'hc3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6339 = 12'hc3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3267; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9411 = 12'hc3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6339; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12483 = 12'hc3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9411; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15555 = 12'hc3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12483; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18627 = 12'hc3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15555; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21699 = 12'hc3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18627; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24771 = 12'hc3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21699; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_195 = io_valid_in ? _GEN_24771 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_195 = 12'hc3 == _T_2[11:0] ? image_195 : _GEN_194; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3268 = 12'hc4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6340 = 12'hc4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3268; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9412 = 12'hc4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6340; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12484 = 12'hc4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9412; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15556 = 12'hc4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12484; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18628 = 12'hc4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15556; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21700 = 12'hc4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18628; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24772 = 12'hc4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21700; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_196 = io_valid_in ? _GEN_24772 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_196 = 12'hc4 == _T_2[11:0] ? image_196 : _GEN_195; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3269 = 12'hc5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6341 = 12'hc5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3269; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9413 = 12'hc5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6341; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12485 = 12'hc5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9413; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15557 = 12'hc5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12485; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18629 = 12'hc5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15557; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21701 = 12'hc5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18629; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24773 = 12'hc5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21701; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_197 = io_valid_in ? _GEN_24773 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_197 = 12'hc5 == _T_2[11:0] ? image_197 : _GEN_196; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3270 = 12'hc6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6342 = 12'hc6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3270; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9414 = 12'hc6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6342; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12486 = 12'hc6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9414; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15558 = 12'hc6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12486; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18630 = 12'hc6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15558; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21702 = 12'hc6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18630; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24774 = 12'hc6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21702; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_198 = io_valid_in ? _GEN_24774 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_198 = 12'hc6 == _T_2[11:0] ? image_198 : _GEN_197; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3271 = 12'hc7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6343 = 12'hc7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3271; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9415 = 12'hc7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6343; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12487 = 12'hc7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9415; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15559 = 12'hc7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12487; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18631 = 12'hc7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15559; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21703 = 12'hc7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18631; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24775 = 12'hc7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21703; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_199 = io_valid_in ? _GEN_24775 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_199 = 12'hc7 == _T_2[11:0] ? image_199 : _GEN_198; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3272 = 12'hc8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6344 = 12'hc8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3272; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9416 = 12'hc8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6344; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12488 = 12'hc8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9416; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15560 = 12'hc8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12488; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18632 = 12'hc8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15560; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21704 = 12'hc8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18632; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24776 = 12'hc8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21704; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_200 = io_valid_in ? _GEN_24776 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_200 = 12'hc8 == _T_2[11:0] ? image_200 : _GEN_199; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3273 = 12'hc9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6345 = 12'hc9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3273; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9417 = 12'hc9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6345; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12489 = 12'hc9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9417; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15561 = 12'hc9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12489; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18633 = 12'hc9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15561; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21705 = 12'hc9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18633; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24777 = 12'hc9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21705; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_201 = io_valid_in ? _GEN_24777 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_201 = 12'hc9 == _T_2[11:0] ? image_201 : _GEN_200; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3274 = 12'hca == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6346 = 12'hca == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3274; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9418 = 12'hca == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6346; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12490 = 12'hca == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9418; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15562 = 12'hca == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12490; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18634 = 12'hca == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15562; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21706 = 12'hca == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18634; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24778 = 12'hca == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21706; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_202 = io_valid_in ? _GEN_24778 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_202 = 12'hca == _T_2[11:0] ? image_202 : _GEN_201; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3275 = 12'hcb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6347 = 12'hcb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3275; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9419 = 12'hcb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6347; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12491 = 12'hcb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9419; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15563 = 12'hcb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12491; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18635 = 12'hcb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15563; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21707 = 12'hcb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18635; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24779 = 12'hcb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21707; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_203 = io_valid_in ? _GEN_24779 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_203 = 12'hcb == _T_2[11:0] ? image_203 : _GEN_202; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3276 = 12'hcc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6348 = 12'hcc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3276; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9420 = 12'hcc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6348; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12492 = 12'hcc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9420; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15564 = 12'hcc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12492; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18636 = 12'hcc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15564; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21708 = 12'hcc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18636; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24780 = 12'hcc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21708; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_204 = io_valid_in ? _GEN_24780 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_204 = 12'hcc == _T_2[11:0] ? image_204 : _GEN_203; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3277 = 12'hcd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6349 = 12'hcd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3277; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9421 = 12'hcd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6349; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12493 = 12'hcd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9421; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15565 = 12'hcd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12493; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18637 = 12'hcd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15565; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21709 = 12'hcd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18637; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24781 = 12'hcd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21709; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_205 = io_valid_in ? _GEN_24781 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_205 = 12'hcd == _T_2[11:0] ? image_205 : _GEN_204; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3278 = 12'hce == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6350 = 12'hce == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3278; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9422 = 12'hce == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6350; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12494 = 12'hce == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9422; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15566 = 12'hce == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12494; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18638 = 12'hce == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15566; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21710 = 12'hce == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18638; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24782 = 12'hce == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21710; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_206 = io_valid_in ? _GEN_24782 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_206 = 12'hce == _T_2[11:0] ? image_206 : _GEN_205; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3279 = 12'hcf == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6351 = 12'hcf == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3279; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9423 = 12'hcf == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6351; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12495 = 12'hcf == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9423; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15567 = 12'hcf == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12495; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18639 = 12'hcf == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15567; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21711 = 12'hcf == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18639; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24783 = 12'hcf == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21711; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_207 = io_valid_in ? _GEN_24783 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_207 = 12'hcf == _T_2[11:0] ? image_207 : _GEN_206; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3280 = 12'hd0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6352 = 12'hd0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3280; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9424 = 12'hd0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6352; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12496 = 12'hd0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9424; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15568 = 12'hd0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12496; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18640 = 12'hd0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15568; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21712 = 12'hd0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18640; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24784 = 12'hd0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21712; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_208 = io_valid_in ? _GEN_24784 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_208 = 12'hd0 == _T_2[11:0] ? image_208 : _GEN_207; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3281 = 12'hd1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6353 = 12'hd1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3281; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9425 = 12'hd1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6353; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12497 = 12'hd1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9425; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15569 = 12'hd1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12497; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18641 = 12'hd1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15569; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21713 = 12'hd1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18641; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24785 = 12'hd1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21713; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_209 = io_valid_in ? _GEN_24785 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_209 = 12'hd1 == _T_2[11:0] ? image_209 : _GEN_208; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3282 = 12'hd2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6354 = 12'hd2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3282; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9426 = 12'hd2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6354; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12498 = 12'hd2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9426; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15570 = 12'hd2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12498; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18642 = 12'hd2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15570; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21714 = 12'hd2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18642; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24786 = 12'hd2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21714; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_210 = io_valid_in ? _GEN_24786 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_210 = 12'hd2 == _T_2[11:0] ? image_210 : _GEN_209; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3283 = 12'hd3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6355 = 12'hd3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3283; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9427 = 12'hd3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6355; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12499 = 12'hd3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9427; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15571 = 12'hd3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12499; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18643 = 12'hd3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15571; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21715 = 12'hd3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18643; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24787 = 12'hd3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21715; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_211 = io_valid_in ? _GEN_24787 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_211 = 12'hd3 == _T_2[11:0] ? image_211 : _GEN_210; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3284 = 12'hd4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6356 = 12'hd4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3284; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9428 = 12'hd4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6356; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12500 = 12'hd4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9428; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15572 = 12'hd4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12500; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18644 = 12'hd4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15572; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21716 = 12'hd4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18644; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24788 = 12'hd4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21716; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_212 = io_valid_in ? _GEN_24788 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_212 = 12'hd4 == _T_2[11:0] ? image_212 : _GEN_211; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3285 = 12'hd5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6357 = 12'hd5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3285; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9429 = 12'hd5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6357; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12501 = 12'hd5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9429; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15573 = 12'hd5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12501; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18645 = 12'hd5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15573; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21717 = 12'hd5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18645; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24789 = 12'hd5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21717; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_213 = io_valid_in ? _GEN_24789 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_213 = 12'hd5 == _T_2[11:0] ? image_213 : _GEN_212; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3286 = 12'hd6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6358 = 12'hd6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3286; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9430 = 12'hd6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6358; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12502 = 12'hd6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9430; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15574 = 12'hd6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12502; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18646 = 12'hd6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15574; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21718 = 12'hd6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18646; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24790 = 12'hd6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21718; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_214 = io_valid_in ? _GEN_24790 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_214 = 12'hd6 == _T_2[11:0] ? image_214 : _GEN_213; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3287 = 12'hd7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6359 = 12'hd7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3287; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9431 = 12'hd7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6359; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12503 = 12'hd7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9431; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15575 = 12'hd7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12503; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18647 = 12'hd7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15575; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21719 = 12'hd7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18647; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24791 = 12'hd7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21719; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_215 = io_valid_in ? _GEN_24791 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_215 = 12'hd7 == _T_2[11:0] ? image_215 : _GEN_214; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3288 = 12'hd8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6360 = 12'hd8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3288; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9432 = 12'hd8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6360; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12504 = 12'hd8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9432; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15576 = 12'hd8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12504; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18648 = 12'hd8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15576; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21720 = 12'hd8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18648; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24792 = 12'hd8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21720; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_216 = io_valid_in ? _GEN_24792 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_216 = 12'hd8 == _T_2[11:0] ? image_216 : _GEN_215; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3289 = 12'hd9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6361 = 12'hd9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3289; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9433 = 12'hd9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6361; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12505 = 12'hd9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9433; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15577 = 12'hd9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12505; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18649 = 12'hd9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15577; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21721 = 12'hd9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18649; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24793 = 12'hd9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21721; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_217 = io_valid_in ? _GEN_24793 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_217 = 12'hd9 == _T_2[11:0] ? image_217 : _GEN_216; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3290 = 12'hda == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6362 = 12'hda == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3290; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9434 = 12'hda == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6362; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12506 = 12'hda == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9434; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15578 = 12'hda == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12506; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18650 = 12'hda == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15578; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21722 = 12'hda == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18650; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24794 = 12'hda == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21722; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_218 = io_valid_in ? _GEN_24794 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_218 = 12'hda == _T_2[11:0] ? image_218 : _GEN_217; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3291 = 12'hdb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6363 = 12'hdb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3291; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9435 = 12'hdb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6363; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12507 = 12'hdb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9435; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15579 = 12'hdb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12507; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18651 = 12'hdb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15579; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21723 = 12'hdb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18651; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24795 = 12'hdb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21723; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_219 = io_valid_in ? _GEN_24795 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_219 = 12'hdb == _T_2[11:0] ? image_219 : _GEN_218; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3292 = 12'hdc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6364 = 12'hdc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3292; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9436 = 12'hdc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6364; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12508 = 12'hdc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9436; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15580 = 12'hdc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12508; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18652 = 12'hdc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15580; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21724 = 12'hdc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18652; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24796 = 12'hdc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21724; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_220 = io_valid_in ? _GEN_24796 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_220 = 12'hdc == _T_2[11:0] ? image_220 : _GEN_219; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3293 = 12'hdd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6365 = 12'hdd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3293; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9437 = 12'hdd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6365; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12509 = 12'hdd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9437; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15581 = 12'hdd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12509; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18653 = 12'hdd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15581; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21725 = 12'hdd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18653; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24797 = 12'hdd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21725; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_221 = io_valid_in ? _GEN_24797 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_221 = 12'hdd == _T_2[11:0] ? image_221 : _GEN_220; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3294 = 12'hde == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6366 = 12'hde == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3294; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9438 = 12'hde == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6366; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12510 = 12'hde == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9438; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15582 = 12'hde == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12510; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18654 = 12'hde == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15582; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21726 = 12'hde == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18654; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24798 = 12'hde == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21726; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_222 = io_valid_in ? _GEN_24798 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_222 = 12'hde == _T_2[11:0] ? image_222 : _GEN_221; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3295 = 12'hdf == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6367 = 12'hdf == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3295; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9439 = 12'hdf == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6367; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12511 = 12'hdf == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9439; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15583 = 12'hdf == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12511; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18655 = 12'hdf == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15583; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21727 = 12'hdf == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18655; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24799 = 12'hdf == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21727; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_223 = io_valid_in ? _GEN_24799 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_223 = 12'hdf == _T_2[11:0] ? image_223 : _GEN_222; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3296 = 12'he0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6368 = 12'he0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3296; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9440 = 12'he0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6368; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12512 = 12'he0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9440; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15584 = 12'he0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12512; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18656 = 12'he0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15584; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21728 = 12'he0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18656; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24800 = 12'he0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21728; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_224 = io_valid_in ? _GEN_24800 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_224 = 12'he0 == _T_2[11:0] ? image_224 : _GEN_223; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3297 = 12'he1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6369 = 12'he1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3297; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9441 = 12'he1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6369; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12513 = 12'he1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9441; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15585 = 12'he1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12513; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18657 = 12'he1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15585; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21729 = 12'he1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18657; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24801 = 12'he1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21729; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_225 = io_valid_in ? _GEN_24801 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_225 = 12'he1 == _T_2[11:0] ? image_225 : _GEN_224; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3298 = 12'he2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6370 = 12'he2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3298; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9442 = 12'he2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6370; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12514 = 12'he2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9442; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15586 = 12'he2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12514; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18658 = 12'he2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15586; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21730 = 12'he2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18658; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24802 = 12'he2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21730; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_226 = io_valid_in ? _GEN_24802 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_226 = 12'he2 == _T_2[11:0] ? image_226 : _GEN_225; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3299 = 12'he3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6371 = 12'he3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3299; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9443 = 12'he3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6371; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12515 = 12'he3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9443; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15587 = 12'he3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12515; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18659 = 12'he3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15587; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21731 = 12'he3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18659; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24803 = 12'he3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21731; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_227 = io_valid_in ? _GEN_24803 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_227 = 12'he3 == _T_2[11:0] ? image_227 : _GEN_226; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3300 = 12'he4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6372 = 12'he4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3300; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9444 = 12'he4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6372; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12516 = 12'he4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9444; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15588 = 12'he4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12516; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18660 = 12'he4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15588; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21732 = 12'he4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18660; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24804 = 12'he4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21732; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_228 = io_valid_in ? _GEN_24804 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_228 = 12'he4 == _T_2[11:0] ? image_228 : _GEN_227; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3301 = 12'he5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6373 = 12'he5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3301; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9445 = 12'he5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6373; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12517 = 12'he5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9445; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15589 = 12'he5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12517; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18661 = 12'he5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15589; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21733 = 12'he5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18661; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24805 = 12'he5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21733; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_229 = io_valid_in ? _GEN_24805 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_229 = 12'he5 == _T_2[11:0] ? image_229 : _GEN_228; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3302 = 12'he6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6374 = 12'he6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3302; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9446 = 12'he6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6374; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12518 = 12'he6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9446; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15590 = 12'he6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12518; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18662 = 12'he6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15590; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21734 = 12'he6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18662; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24806 = 12'he6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21734; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_230 = io_valid_in ? _GEN_24806 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_230 = 12'he6 == _T_2[11:0] ? image_230 : _GEN_229; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3303 = 12'he7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6375 = 12'he7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3303; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9447 = 12'he7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6375; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12519 = 12'he7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9447; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15591 = 12'he7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12519; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18663 = 12'he7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15591; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21735 = 12'he7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18663; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24807 = 12'he7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21735; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_231 = io_valid_in ? _GEN_24807 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_231 = 12'he7 == _T_2[11:0] ? image_231 : _GEN_230; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3304 = 12'he8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6376 = 12'he8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3304; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9448 = 12'he8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6376; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12520 = 12'he8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9448; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15592 = 12'he8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12520; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18664 = 12'he8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15592; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21736 = 12'he8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18664; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24808 = 12'he8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21736; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_232 = io_valid_in ? _GEN_24808 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_232 = 12'he8 == _T_2[11:0] ? image_232 : _GEN_231; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3305 = 12'he9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6377 = 12'he9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3305; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9449 = 12'he9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6377; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12521 = 12'he9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9449; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15593 = 12'he9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12521; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18665 = 12'he9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15593; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21737 = 12'he9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18665; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24809 = 12'he9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21737; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_233 = io_valid_in ? _GEN_24809 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_233 = 12'he9 == _T_2[11:0] ? image_233 : _GEN_232; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3306 = 12'hea == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6378 = 12'hea == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3306; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9450 = 12'hea == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6378; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12522 = 12'hea == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9450; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15594 = 12'hea == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12522; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18666 = 12'hea == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15594; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21738 = 12'hea == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18666; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24810 = 12'hea == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21738; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_234 = io_valid_in ? _GEN_24810 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_234 = 12'hea == _T_2[11:0] ? image_234 : _GEN_233; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3307 = 12'heb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6379 = 12'heb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3307; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9451 = 12'heb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6379; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12523 = 12'heb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9451; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15595 = 12'heb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12523; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18667 = 12'heb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15595; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21739 = 12'heb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18667; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24811 = 12'heb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21739; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_235 = io_valid_in ? _GEN_24811 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_235 = 12'heb == _T_2[11:0] ? image_235 : _GEN_234; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3308 = 12'hec == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6380 = 12'hec == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3308; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9452 = 12'hec == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6380; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12524 = 12'hec == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9452; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15596 = 12'hec == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12524; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18668 = 12'hec == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15596; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21740 = 12'hec == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18668; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24812 = 12'hec == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21740; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_236 = io_valid_in ? _GEN_24812 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_236 = 12'hec == _T_2[11:0] ? image_236 : _GEN_235; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3309 = 12'hed == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6381 = 12'hed == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3309; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9453 = 12'hed == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6381; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12525 = 12'hed == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9453; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15597 = 12'hed == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12525; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18669 = 12'hed == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15597; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21741 = 12'hed == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18669; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24813 = 12'hed == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21741; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_237 = io_valid_in ? _GEN_24813 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_237 = 12'hed == _T_2[11:0] ? image_237 : _GEN_236; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3310 = 12'hee == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6382 = 12'hee == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3310; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9454 = 12'hee == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6382; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12526 = 12'hee == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9454; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15598 = 12'hee == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12526; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18670 = 12'hee == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15598; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21742 = 12'hee == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18670; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24814 = 12'hee == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21742; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_238 = io_valid_in ? _GEN_24814 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_238 = 12'hee == _T_2[11:0] ? image_238 : _GEN_237; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3311 = 12'hef == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6383 = 12'hef == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3311; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9455 = 12'hef == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6383; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12527 = 12'hef == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9455; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15599 = 12'hef == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12527; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18671 = 12'hef == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15599; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21743 = 12'hef == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18671; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24815 = 12'hef == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21743; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_239 = io_valid_in ? _GEN_24815 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_239 = 12'hef == _T_2[11:0] ? image_239 : _GEN_238; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3312 = 12'hf0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6384 = 12'hf0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3312; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9456 = 12'hf0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6384; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12528 = 12'hf0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9456; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15600 = 12'hf0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12528; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18672 = 12'hf0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15600; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21744 = 12'hf0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18672; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24816 = 12'hf0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21744; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_240 = io_valid_in ? _GEN_24816 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_240 = 12'hf0 == _T_2[11:0] ? image_240 : _GEN_239; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3313 = 12'hf1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6385 = 12'hf1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3313; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9457 = 12'hf1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6385; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12529 = 12'hf1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9457; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15601 = 12'hf1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12529; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18673 = 12'hf1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15601; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21745 = 12'hf1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18673; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24817 = 12'hf1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21745; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_241 = io_valid_in ? _GEN_24817 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_241 = 12'hf1 == _T_2[11:0] ? image_241 : _GEN_240; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3314 = 12'hf2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6386 = 12'hf2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3314; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9458 = 12'hf2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6386; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12530 = 12'hf2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9458; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15602 = 12'hf2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12530; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18674 = 12'hf2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15602; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21746 = 12'hf2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18674; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24818 = 12'hf2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21746; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_242 = io_valid_in ? _GEN_24818 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_242 = 12'hf2 == _T_2[11:0] ? image_242 : _GEN_241; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3315 = 12'hf3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6387 = 12'hf3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3315; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9459 = 12'hf3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6387; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12531 = 12'hf3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9459; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15603 = 12'hf3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12531; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18675 = 12'hf3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15603; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21747 = 12'hf3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18675; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24819 = 12'hf3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21747; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_243 = io_valid_in ? _GEN_24819 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_243 = 12'hf3 == _T_2[11:0] ? image_243 : _GEN_242; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3316 = 12'hf4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6388 = 12'hf4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3316; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9460 = 12'hf4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6388; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12532 = 12'hf4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9460; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15604 = 12'hf4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12532; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18676 = 12'hf4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15604; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21748 = 12'hf4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18676; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24820 = 12'hf4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21748; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_244 = io_valid_in ? _GEN_24820 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_244 = 12'hf4 == _T_2[11:0] ? image_244 : _GEN_243; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3317 = 12'hf5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6389 = 12'hf5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3317; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9461 = 12'hf5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6389; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12533 = 12'hf5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9461; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15605 = 12'hf5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12533; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18677 = 12'hf5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15605; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21749 = 12'hf5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18677; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24821 = 12'hf5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21749; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_245 = io_valid_in ? _GEN_24821 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_245 = 12'hf5 == _T_2[11:0] ? image_245 : _GEN_244; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3318 = 12'hf6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6390 = 12'hf6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3318; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9462 = 12'hf6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6390; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12534 = 12'hf6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9462; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15606 = 12'hf6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12534; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18678 = 12'hf6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15606; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21750 = 12'hf6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18678; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24822 = 12'hf6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21750; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_246 = io_valid_in ? _GEN_24822 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_246 = 12'hf6 == _T_2[11:0] ? image_246 : _GEN_245; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3319 = 12'hf7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6391 = 12'hf7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3319; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9463 = 12'hf7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6391; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12535 = 12'hf7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9463; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15607 = 12'hf7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12535; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18679 = 12'hf7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15607; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21751 = 12'hf7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18679; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24823 = 12'hf7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21751; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_247 = io_valid_in ? _GEN_24823 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_247 = 12'hf7 == _T_2[11:0] ? image_247 : _GEN_246; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3320 = 12'hf8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6392 = 12'hf8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3320; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9464 = 12'hf8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6392; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12536 = 12'hf8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9464; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15608 = 12'hf8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12536; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18680 = 12'hf8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15608; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21752 = 12'hf8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18680; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24824 = 12'hf8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21752; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_248 = io_valid_in ? _GEN_24824 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_248 = 12'hf8 == _T_2[11:0] ? image_248 : _GEN_247; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3321 = 12'hf9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6393 = 12'hf9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3321; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9465 = 12'hf9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6393; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12537 = 12'hf9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9465; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15609 = 12'hf9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12537; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18681 = 12'hf9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15609; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21753 = 12'hf9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18681; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24825 = 12'hf9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21753; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_249 = io_valid_in ? _GEN_24825 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_249 = 12'hf9 == _T_2[11:0] ? image_249 : _GEN_248; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3322 = 12'hfa == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6394 = 12'hfa == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3322; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9466 = 12'hfa == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6394; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12538 = 12'hfa == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9466; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15610 = 12'hfa == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12538; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18682 = 12'hfa == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15610; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21754 = 12'hfa == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18682; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24826 = 12'hfa == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21754; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_250 = io_valid_in ? _GEN_24826 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_250 = 12'hfa == _T_2[11:0] ? image_250 : _GEN_249; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3323 = 12'hfb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6395 = 12'hfb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3323; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9467 = 12'hfb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6395; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12539 = 12'hfb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9467; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15611 = 12'hfb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12539; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18683 = 12'hfb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15611; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21755 = 12'hfb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18683; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24827 = 12'hfb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21755; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_251 = io_valid_in ? _GEN_24827 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_251 = 12'hfb == _T_2[11:0] ? image_251 : _GEN_250; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3324 = 12'hfc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6396 = 12'hfc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3324; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9468 = 12'hfc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6396; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12540 = 12'hfc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9468; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15612 = 12'hfc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12540; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18684 = 12'hfc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15612; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21756 = 12'hfc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18684; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24828 = 12'hfc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21756; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_252 = io_valid_in ? _GEN_24828 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_252 = 12'hfc == _T_2[11:0] ? image_252 : _GEN_251; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3325 = 12'hfd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6397 = 12'hfd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3325; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9469 = 12'hfd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6397; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12541 = 12'hfd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9469; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15613 = 12'hfd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12541; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18685 = 12'hfd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15613; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21757 = 12'hfd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18685; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24829 = 12'hfd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21757; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_253 = io_valid_in ? _GEN_24829 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_253 = 12'hfd == _T_2[11:0] ? image_253 : _GEN_252; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3326 = 12'hfe == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6398 = 12'hfe == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3326; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9470 = 12'hfe == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6398; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12542 = 12'hfe == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9470; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15614 = 12'hfe == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12542; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18686 = 12'hfe == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15614; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21758 = 12'hfe == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18686; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24830 = 12'hfe == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21758; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_254 = io_valid_in ? _GEN_24830 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_254 = 12'hfe == _T_2[11:0] ? image_254 : _GEN_253; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3327 = 12'hff == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6399 = 12'hff == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3327; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9471 = 12'hff == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6399; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12543 = 12'hff == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9471; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15615 = 12'hff == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12543; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18687 = 12'hff == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15615; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21759 = 12'hff == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18687; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24831 = 12'hff == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21759; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_255 = io_valid_in ? _GEN_24831 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_255 = 12'hff == _T_2[11:0] ? image_255 : _GEN_254; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3328 = 12'h100 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6400 = 12'h100 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3328; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9472 = 12'h100 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6400; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12544 = 12'h100 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9472; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15616 = 12'h100 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12544; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18688 = 12'h100 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15616; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21760 = 12'h100 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18688; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24832 = 12'h100 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21760; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_256 = io_valid_in ? _GEN_24832 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_256 = 12'h100 == _T_2[11:0] ? image_256 : _GEN_255; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3329 = 12'h101 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6401 = 12'h101 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3329; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9473 = 12'h101 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6401; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12545 = 12'h101 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9473; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15617 = 12'h101 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12545; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18689 = 12'h101 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15617; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21761 = 12'h101 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18689; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24833 = 12'h101 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21761; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_257 = io_valid_in ? _GEN_24833 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_257 = 12'h101 == _T_2[11:0] ? image_257 : _GEN_256; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3330 = 12'h102 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6402 = 12'h102 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3330; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9474 = 12'h102 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6402; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12546 = 12'h102 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9474; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15618 = 12'h102 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12546; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18690 = 12'h102 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15618; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21762 = 12'h102 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18690; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24834 = 12'h102 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21762; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_258 = io_valid_in ? _GEN_24834 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_258 = 12'h102 == _T_2[11:0] ? image_258 : _GEN_257; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3331 = 12'h103 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6403 = 12'h103 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3331; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9475 = 12'h103 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6403; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12547 = 12'h103 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9475; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15619 = 12'h103 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12547; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18691 = 12'h103 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15619; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21763 = 12'h103 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18691; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24835 = 12'h103 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21763; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_259 = io_valid_in ? _GEN_24835 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_259 = 12'h103 == _T_2[11:0] ? image_259 : _GEN_258; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3332 = 12'h104 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6404 = 12'h104 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3332; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9476 = 12'h104 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6404; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12548 = 12'h104 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9476; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15620 = 12'h104 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12548; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18692 = 12'h104 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15620; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21764 = 12'h104 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18692; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24836 = 12'h104 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21764; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_260 = io_valid_in ? _GEN_24836 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_260 = 12'h104 == _T_2[11:0] ? image_260 : _GEN_259; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3333 = 12'h105 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6405 = 12'h105 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3333; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9477 = 12'h105 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6405; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12549 = 12'h105 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9477; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15621 = 12'h105 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12549; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18693 = 12'h105 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15621; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21765 = 12'h105 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18693; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24837 = 12'h105 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21765; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_261 = io_valid_in ? _GEN_24837 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_261 = 12'h105 == _T_2[11:0] ? image_261 : _GEN_260; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3334 = 12'h106 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6406 = 12'h106 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3334; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9478 = 12'h106 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6406; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12550 = 12'h106 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9478; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15622 = 12'h106 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12550; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18694 = 12'h106 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15622; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21766 = 12'h106 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18694; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24838 = 12'h106 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21766; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_262 = io_valid_in ? _GEN_24838 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_262 = 12'h106 == _T_2[11:0] ? image_262 : _GEN_261; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3335 = 12'h107 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6407 = 12'h107 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3335; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9479 = 12'h107 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6407; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12551 = 12'h107 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9479; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15623 = 12'h107 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12551; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18695 = 12'h107 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15623; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21767 = 12'h107 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18695; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24839 = 12'h107 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21767; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_263 = io_valid_in ? _GEN_24839 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_263 = 12'h107 == _T_2[11:0] ? image_263 : _GEN_262; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3336 = 12'h108 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6408 = 12'h108 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3336; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9480 = 12'h108 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6408; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12552 = 12'h108 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9480; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15624 = 12'h108 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12552; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18696 = 12'h108 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15624; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21768 = 12'h108 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18696; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24840 = 12'h108 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21768; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_264 = io_valid_in ? _GEN_24840 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_264 = 12'h108 == _T_2[11:0] ? image_264 : _GEN_263; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3337 = 12'h109 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6409 = 12'h109 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3337; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9481 = 12'h109 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6409; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12553 = 12'h109 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9481; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15625 = 12'h109 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12553; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18697 = 12'h109 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15625; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21769 = 12'h109 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18697; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24841 = 12'h109 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21769; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_265 = io_valid_in ? _GEN_24841 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_265 = 12'h109 == _T_2[11:0] ? image_265 : _GEN_264; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3338 = 12'h10a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6410 = 12'h10a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3338; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9482 = 12'h10a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6410; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12554 = 12'h10a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9482; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15626 = 12'h10a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12554; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18698 = 12'h10a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15626; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21770 = 12'h10a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18698; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24842 = 12'h10a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21770; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_266 = io_valid_in ? _GEN_24842 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_266 = 12'h10a == _T_2[11:0] ? image_266 : _GEN_265; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3339 = 12'h10b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6411 = 12'h10b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3339; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9483 = 12'h10b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6411; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12555 = 12'h10b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9483; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15627 = 12'h10b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12555; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18699 = 12'h10b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15627; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21771 = 12'h10b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18699; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24843 = 12'h10b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21771; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_267 = io_valid_in ? _GEN_24843 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_267 = 12'h10b == _T_2[11:0] ? image_267 : _GEN_266; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3340 = 12'h10c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6412 = 12'h10c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3340; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9484 = 12'h10c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6412; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12556 = 12'h10c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9484; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15628 = 12'h10c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12556; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18700 = 12'h10c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15628; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21772 = 12'h10c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18700; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24844 = 12'h10c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21772; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_268 = io_valid_in ? _GEN_24844 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_268 = 12'h10c == _T_2[11:0] ? image_268 : _GEN_267; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3341 = 12'h10d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6413 = 12'h10d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3341; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9485 = 12'h10d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6413; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12557 = 12'h10d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9485; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15629 = 12'h10d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12557; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18701 = 12'h10d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15629; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21773 = 12'h10d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18701; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24845 = 12'h10d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21773; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_269 = io_valid_in ? _GEN_24845 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_269 = 12'h10d == _T_2[11:0] ? image_269 : _GEN_268; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3342 = 12'h10e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6414 = 12'h10e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3342; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9486 = 12'h10e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6414; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12558 = 12'h10e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9486; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15630 = 12'h10e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12558; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18702 = 12'h10e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15630; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21774 = 12'h10e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18702; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24846 = 12'h10e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21774; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_270 = io_valid_in ? _GEN_24846 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_270 = 12'h10e == _T_2[11:0] ? image_270 : _GEN_269; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3343 = 12'h10f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6415 = 12'h10f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3343; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9487 = 12'h10f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6415; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12559 = 12'h10f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9487; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15631 = 12'h10f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12559; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18703 = 12'h10f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15631; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21775 = 12'h10f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18703; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24847 = 12'h10f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21775; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_271 = io_valid_in ? _GEN_24847 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_271 = 12'h10f == _T_2[11:0] ? image_271 : _GEN_270; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3344 = 12'h110 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6416 = 12'h110 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3344; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9488 = 12'h110 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6416; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12560 = 12'h110 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9488; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15632 = 12'h110 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12560; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18704 = 12'h110 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15632; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21776 = 12'h110 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18704; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24848 = 12'h110 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21776; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_272 = io_valid_in ? _GEN_24848 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_272 = 12'h110 == _T_2[11:0] ? image_272 : _GEN_271; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3345 = 12'h111 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6417 = 12'h111 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3345; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9489 = 12'h111 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6417; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12561 = 12'h111 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9489; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15633 = 12'h111 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12561; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18705 = 12'h111 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15633; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21777 = 12'h111 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18705; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24849 = 12'h111 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21777; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_273 = io_valid_in ? _GEN_24849 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_273 = 12'h111 == _T_2[11:0] ? image_273 : _GEN_272; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3346 = 12'h112 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6418 = 12'h112 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3346; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9490 = 12'h112 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6418; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12562 = 12'h112 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9490; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15634 = 12'h112 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12562; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18706 = 12'h112 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15634; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21778 = 12'h112 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18706; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24850 = 12'h112 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21778; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_274 = io_valid_in ? _GEN_24850 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_274 = 12'h112 == _T_2[11:0] ? image_274 : _GEN_273; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3347 = 12'h113 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6419 = 12'h113 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3347; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9491 = 12'h113 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6419; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12563 = 12'h113 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9491; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15635 = 12'h113 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12563; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18707 = 12'h113 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15635; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21779 = 12'h113 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18707; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24851 = 12'h113 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21779; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_275 = io_valid_in ? _GEN_24851 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_275 = 12'h113 == _T_2[11:0] ? image_275 : _GEN_274; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3348 = 12'h114 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6420 = 12'h114 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3348; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9492 = 12'h114 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6420; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12564 = 12'h114 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9492; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15636 = 12'h114 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12564; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18708 = 12'h114 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15636; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21780 = 12'h114 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18708; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24852 = 12'h114 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21780; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_276 = io_valid_in ? _GEN_24852 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_276 = 12'h114 == _T_2[11:0] ? image_276 : _GEN_275; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3349 = 12'h115 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6421 = 12'h115 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3349; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9493 = 12'h115 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6421; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12565 = 12'h115 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9493; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15637 = 12'h115 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12565; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18709 = 12'h115 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15637; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21781 = 12'h115 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18709; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24853 = 12'h115 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21781; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_277 = io_valid_in ? _GEN_24853 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_277 = 12'h115 == _T_2[11:0] ? image_277 : _GEN_276; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3350 = 12'h116 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6422 = 12'h116 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3350; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9494 = 12'h116 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6422; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12566 = 12'h116 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9494; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15638 = 12'h116 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12566; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18710 = 12'h116 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15638; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21782 = 12'h116 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18710; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24854 = 12'h116 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21782; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_278 = io_valid_in ? _GEN_24854 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_278 = 12'h116 == _T_2[11:0] ? image_278 : _GEN_277; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3351 = 12'h117 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6423 = 12'h117 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3351; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9495 = 12'h117 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6423; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12567 = 12'h117 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9495; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15639 = 12'h117 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12567; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18711 = 12'h117 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15639; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21783 = 12'h117 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18711; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24855 = 12'h117 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21783; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_279 = io_valid_in ? _GEN_24855 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_279 = 12'h117 == _T_2[11:0] ? image_279 : _GEN_278; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3352 = 12'h118 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6424 = 12'h118 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3352; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9496 = 12'h118 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6424; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12568 = 12'h118 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9496; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15640 = 12'h118 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12568; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18712 = 12'h118 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15640; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21784 = 12'h118 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18712; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24856 = 12'h118 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21784; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_280 = io_valid_in ? _GEN_24856 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_280 = 12'h118 == _T_2[11:0] ? image_280 : _GEN_279; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3353 = 12'h119 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6425 = 12'h119 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3353; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9497 = 12'h119 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6425; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12569 = 12'h119 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9497; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15641 = 12'h119 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12569; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18713 = 12'h119 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15641; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21785 = 12'h119 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18713; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24857 = 12'h119 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21785; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_281 = io_valid_in ? _GEN_24857 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_281 = 12'h119 == _T_2[11:0] ? image_281 : _GEN_280; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3354 = 12'h11a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6426 = 12'h11a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3354; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9498 = 12'h11a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6426; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12570 = 12'h11a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9498; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15642 = 12'h11a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12570; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18714 = 12'h11a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15642; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21786 = 12'h11a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18714; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24858 = 12'h11a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21786; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_282 = io_valid_in ? _GEN_24858 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_282 = 12'h11a == _T_2[11:0] ? image_282 : _GEN_281; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3355 = 12'h11b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6427 = 12'h11b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3355; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9499 = 12'h11b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6427; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12571 = 12'h11b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9499; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15643 = 12'h11b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12571; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18715 = 12'h11b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15643; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21787 = 12'h11b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18715; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24859 = 12'h11b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21787; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_283 = io_valid_in ? _GEN_24859 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_283 = 12'h11b == _T_2[11:0] ? image_283 : _GEN_282; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3356 = 12'h11c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6428 = 12'h11c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3356; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9500 = 12'h11c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6428; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12572 = 12'h11c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9500; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15644 = 12'h11c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12572; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18716 = 12'h11c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15644; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21788 = 12'h11c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18716; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24860 = 12'h11c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21788; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_284 = io_valid_in ? _GEN_24860 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_284 = 12'h11c == _T_2[11:0] ? image_284 : _GEN_283; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3357 = 12'h11d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6429 = 12'h11d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3357; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9501 = 12'h11d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6429; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12573 = 12'h11d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9501; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15645 = 12'h11d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12573; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18717 = 12'h11d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15645; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21789 = 12'h11d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18717; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24861 = 12'h11d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21789; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_285 = io_valid_in ? _GEN_24861 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_285 = 12'h11d == _T_2[11:0] ? image_285 : _GEN_284; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3358 = 12'h11e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6430 = 12'h11e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3358; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9502 = 12'h11e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6430; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12574 = 12'h11e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9502; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15646 = 12'h11e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12574; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18718 = 12'h11e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15646; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21790 = 12'h11e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18718; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24862 = 12'h11e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21790; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_286 = io_valid_in ? _GEN_24862 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_286 = 12'h11e == _T_2[11:0] ? image_286 : _GEN_285; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3359 = 12'h11f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6431 = 12'h11f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3359; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9503 = 12'h11f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6431; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12575 = 12'h11f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9503; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15647 = 12'h11f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12575; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18719 = 12'h11f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15647; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21791 = 12'h11f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18719; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24863 = 12'h11f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21791; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_287 = io_valid_in ? _GEN_24863 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_287 = 12'h11f == _T_2[11:0] ? image_287 : _GEN_286; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3360 = 12'h120 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6432 = 12'h120 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3360; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9504 = 12'h120 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6432; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12576 = 12'h120 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9504; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15648 = 12'h120 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12576; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18720 = 12'h120 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15648; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21792 = 12'h120 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18720; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24864 = 12'h120 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21792; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_288 = io_valid_in ? _GEN_24864 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_288 = 12'h120 == _T_2[11:0] ? image_288 : _GEN_287; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3361 = 12'h121 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6433 = 12'h121 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3361; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9505 = 12'h121 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6433; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12577 = 12'h121 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9505; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15649 = 12'h121 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12577; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18721 = 12'h121 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15649; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21793 = 12'h121 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18721; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24865 = 12'h121 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21793; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_289 = io_valid_in ? _GEN_24865 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_289 = 12'h121 == _T_2[11:0] ? image_289 : _GEN_288; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3362 = 12'h122 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6434 = 12'h122 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3362; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9506 = 12'h122 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6434; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12578 = 12'h122 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9506; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15650 = 12'h122 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12578; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18722 = 12'h122 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15650; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21794 = 12'h122 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18722; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24866 = 12'h122 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21794; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_290 = io_valid_in ? _GEN_24866 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_290 = 12'h122 == _T_2[11:0] ? image_290 : _GEN_289; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3363 = 12'h123 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6435 = 12'h123 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3363; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9507 = 12'h123 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6435; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12579 = 12'h123 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9507; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15651 = 12'h123 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12579; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18723 = 12'h123 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15651; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21795 = 12'h123 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18723; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24867 = 12'h123 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21795; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_291 = io_valid_in ? _GEN_24867 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_291 = 12'h123 == _T_2[11:0] ? image_291 : _GEN_290; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3364 = 12'h124 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6436 = 12'h124 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3364; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9508 = 12'h124 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6436; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12580 = 12'h124 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9508; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15652 = 12'h124 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12580; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18724 = 12'h124 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15652; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21796 = 12'h124 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18724; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24868 = 12'h124 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21796; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_292 = io_valid_in ? _GEN_24868 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_292 = 12'h124 == _T_2[11:0] ? image_292 : _GEN_291; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3365 = 12'h125 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6437 = 12'h125 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3365; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9509 = 12'h125 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6437; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12581 = 12'h125 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9509; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15653 = 12'h125 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12581; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18725 = 12'h125 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15653; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21797 = 12'h125 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18725; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24869 = 12'h125 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21797; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_293 = io_valid_in ? _GEN_24869 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_293 = 12'h125 == _T_2[11:0] ? image_293 : _GEN_292; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3366 = 12'h126 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6438 = 12'h126 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3366; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9510 = 12'h126 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6438; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12582 = 12'h126 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9510; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15654 = 12'h126 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12582; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18726 = 12'h126 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15654; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21798 = 12'h126 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18726; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24870 = 12'h126 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21798; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_294 = io_valid_in ? _GEN_24870 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_294 = 12'h126 == _T_2[11:0] ? image_294 : _GEN_293; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3367 = 12'h127 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6439 = 12'h127 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3367; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9511 = 12'h127 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6439; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12583 = 12'h127 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9511; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15655 = 12'h127 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12583; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18727 = 12'h127 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15655; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21799 = 12'h127 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18727; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24871 = 12'h127 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21799; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_295 = io_valid_in ? _GEN_24871 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_295 = 12'h127 == _T_2[11:0] ? image_295 : _GEN_294; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3368 = 12'h128 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6440 = 12'h128 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3368; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9512 = 12'h128 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6440; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12584 = 12'h128 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9512; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15656 = 12'h128 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12584; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18728 = 12'h128 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15656; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21800 = 12'h128 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18728; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24872 = 12'h128 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21800; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_296 = io_valid_in ? _GEN_24872 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_296 = 12'h128 == _T_2[11:0] ? image_296 : _GEN_295; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3369 = 12'h129 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6441 = 12'h129 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3369; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9513 = 12'h129 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6441; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12585 = 12'h129 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9513; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15657 = 12'h129 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12585; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18729 = 12'h129 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15657; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21801 = 12'h129 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18729; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24873 = 12'h129 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21801; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_297 = io_valid_in ? _GEN_24873 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_297 = 12'h129 == _T_2[11:0] ? image_297 : _GEN_296; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3370 = 12'h12a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6442 = 12'h12a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3370; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9514 = 12'h12a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6442; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12586 = 12'h12a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9514; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15658 = 12'h12a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12586; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18730 = 12'h12a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15658; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21802 = 12'h12a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18730; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24874 = 12'h12a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21802; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_298 = io_valid_in ? _GEN_24874 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_298 = 12'h12a == _T_2[11:0] ? image_298 : _GEN_297; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3371 = 12'h12b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6443 = 12'h12b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3371; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9515 = 12'h12b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6443; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12587 = 12'h12b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9515; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15659 = 12'h12b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12587; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18731 = 12'h12b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15659; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21803 = 12'h12b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18731; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24875 = 12'h12b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21803; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_299 = io_valid_in ? _GEN_24875 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_299 = 12'h12b == _T_2[11:0] ? image_299 : _GEN_298; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3372 = 12'h12c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6444 = 12'h12c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3372; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9516 = 12'h12c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6444; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12588 = 12'h12c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9516; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15660 = 12'h12c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12588; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18732 = 12'h12c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15660; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21804 = 12'h12c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18732; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24876 = 12'h12c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21804; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_300 = io_valid_in ? _GEN_24876 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_300 = 12'h12c == _T_2[11:0] ? image_300 : _GEN_299; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3373 = 12'h12d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6445 = 12'h12d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3373; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9517 = 12'h12d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6445; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12589 = 12'h12d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9517; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15661 = 12'h12d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12589; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18733 = 12'h12d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15661; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21805 = 12'h12d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18733; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24877 = 12'h12d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21805; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_301 = io_valid_in ? _GEN_24877 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_301 = 12'h12d == _T_2[11:0] ? image_301 : _GEN_300; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3374 = 12'h12e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6446 = 12'h12e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3374; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9518 = 12'h12e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6446; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12590 = 12'h12e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9518; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15662 = 12'h12e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12590; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18734 = 12'h12e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15662; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21806 = 12'h12e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18734; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24878 = 12'h12e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21806; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_302 = io_valid_in ? _GEN_24878 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_302 = 12'h12e == _T_2[11:0] ? image_302 : _GEN_301; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3375 = 12'h12f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6447 = 12'h12f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3375; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9519 = 12'h12f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6447; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12591 = 12'h12f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9519; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15663 = 12'h12f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12591; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18735 = 12'h12f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15663; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21807 = 12'h12f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18735; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24879 = 12'h12f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21807; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_303 = io_valid_in ? _GEN_24879 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_303 = 12'h12f == _T_2[11:0] ? image_303 : _GEN_302; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3376 = 12'h130 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6448 = 12'h130 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3376; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9520 = 12'h130 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6448; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12592 = 12'h130 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9520; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15664 = 12'h130 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12592; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18736 = 12'h130 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15664; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21808 = 12'h130 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18736; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24880 = 12'h130 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21808; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_304 = io_valid_in ? _GEN_24880 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_304 = 12'h130 == _T_2[11:0] ? image_304 : _GEN_303; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3377 = 12'h131 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6449 = 12'h131 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3377; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9521 = 12'h131 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6449; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12593 = 12'h131 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9521; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15665 = 12'h131 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12593; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18737 = 12'h131 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15665; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21809 = 12'h131 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18737; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24881 = 12'h131 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21809; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_305 = io_valid_in ? _GEN_24881 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_305 = 12'h131 == _T_2[11:0] ? image_305 : _GEN_304; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3378 = 12'h132 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6450 = 12'h132 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3378; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9522 = 12'h132 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6450; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12594 = 12'h132 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9522; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15666 = 12'h132 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12594; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18738 = 12'h132 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15666; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21810 = 12'h132 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18738; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24882 = 12'h132 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21810; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_306 = io_valid_in ? _GEN_24882 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_306 = 12'h132 == _T_2[11:0] ? image_306 : _GEN_305; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3379 = 12'h133 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6451 = 12'h133 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3379; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9523 = 12'h133 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6451; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12595 = 12'h133 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9523; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15667 = 12'h133 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12595; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18739 = 12'h133 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15667; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21811 = 12'h133 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18739; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24883 = 12'h133 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21811; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_307 = io_valid_in ? _GEN_24883 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_307 = 12'h133 == _T_2[11:0] ? image_307 : _GEN_306; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3380 = 12'h134 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6452 = 12'h134 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3380; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9524 = 12'h134 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6452; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12596 = 12'h134 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9524; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15668 = 12'h134 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12596; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18740 = 12'h134 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15668; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21812 = 12'h134 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18740; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24884 = 12'h134 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21812; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_308 = io_valid_in ? _GEN_24884 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_308 = 12'h134 == _T_2[11:0] ? image_308 : _GEN_307; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3381 = 12'h135 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6453 = 12'h135 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3381; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9525 = 12'h135 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6453; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12597 = 12'h135 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9525; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15669 = 12'h135 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12597; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18741 = 12'h135 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15669; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21813 = 12'h135 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18741; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24885 = 12'h135 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21813; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_309 = io_valid_in ? _GEN_24885 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_309 = 12'h135 == _T_2[11:0] ? image_309 : _GEN_308; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3382 = 12'h136 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6454 = 12'h136 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3382; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9526 = 12'h136 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6454; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12598 = 12'h136 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9526; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15670 = 12'h136 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12598; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18742 = 12'h136 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15670; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21814 = 12'h136 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18742; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24886 = 12'h136 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21814; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_310 = io_valid_in ? _GEN_24886 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_310 = 12'h136 == _T_2[11:0] ? image_310 : _GEN_309; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3383 = 12'h137 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6455 = 12'h137 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3383; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9527 = 12'h137 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6455; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12599 = 12'h137 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9527; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15671 = 12'h137 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12599; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18743 = 12'h137 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15671; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21815 = 12'h137 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18743; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24887 = 12'h137 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21815; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_311 = io_valid_in ? _GEN_24887 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_311 = 12'h137 == _T_2[11:0] ? image_311 : _GEN_310; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3384 = 12'h138 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6456 = 12'h138 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3384; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9528 = 12'h138 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6456; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12600 = 12'h138 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9528; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15672 = 12'h138 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12600; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18744 = 12'h138 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15672; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21816 = 12'h138 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18744; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24888 = 12'h138 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21816; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_312 = io_valid_in ? _GEN_24888 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_312 = 12'h138 == _T_2[11:0] ? image_312 : _GEN_311; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3385 = 12'h139 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6457 = 12'h139 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3385; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9529 = 12'h139 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6457; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12601 = 12'h139 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9529; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15673 = 12'h139 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12601; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18745 = 12'h139 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15673; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21817 = 12'h139 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18745; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24889 = 12'h139 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21817; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_313 = io_valid_in ? _GEN_24889 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_313 = 12'h139 == _T_2[11:0] ? image_313 : _GEN_312; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3386 = 12'h13a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6458 = 12'h13a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3386; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9530 = 12'h13a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6458; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12602 = 12'h13a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9530; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15674 = 12'h13a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12602; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18746 = 12'h13a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15674; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21818 = 12'h13a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18746; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24890 = 12'h13a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21818; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_314 = io_valid_in ? _GEN_24890 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_314 = 12'h13a == _T_2[11:0] ? image_314 : _GEN_313; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3387 = 12'h13b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6459 = 12'h13b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3387; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9531 = 12'h13b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6459; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12603 = 12'h13b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9531; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15675 = 12'h13b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12603; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18747 = 12'h13b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15675; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21819 = 12'h13b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18747; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24891 = 12'h13b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21819; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_315 = io_valid_in ? _GEN_24891 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_315 = 12'h13b == _T_2[11:0] ? image_315 : _GEN_314; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3388 = 12'h13c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6460 = 12'h13c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3388; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9532 = 12'h13c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6460; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12604 = 12'h13c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9532; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15676 = 12'h13c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12604; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18748 = 12'h13c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15676; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21820 = 12'h13c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18748; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24892 = 12'h13c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21820; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_316 = io_valid_in ? _GEN_24892 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_316 = 12'h13c == _T_2[11:0] ? image_316 : _GEN_315; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3389 = 12'h13d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6461 = 12'h13d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3389; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9533 = 12'h13d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6461; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12605 = 12'h13d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9533; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15677 = 12'h13d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12605; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18749 = 12'h13d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15677; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21821 = 12'h13d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18749; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24893 = 12'h13d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21821; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_317 = io_valid_in ? _GEN_24893 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_317 = 12'h13d == _T_2[11:0] ? image_317 : _GEN_316; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3390 = 12'h13e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6462 = 12'h13e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3390; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9534 = 12'h13e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6462; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12606 = 12'h13e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9534; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15678 = 12'h13e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12606; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18750 = 12'h13e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15678; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21822 = 12'h13e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18750; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24894 = 12'h13e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21822; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_318 = io_valid_in ? _GEN_24894 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_318 = 12'h13e == _T_2[11:0] ? image_318 : _GEN_317; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3391 = 12'h13f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6463 = 12'h13f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3391; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9535 = 12'h13f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6463; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12607 = 12'h13f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9535; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15679 = 12'h13f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12607; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18751 = 12'h13f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15679; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21823 = 12'h13f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18751; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24895 = 12'h13f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21823; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_319 = io_valid_in ? _GEN_24895 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_319 = 12'h13f == _T_2[11:0] ? image_319 : _GEN_318; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3392 = 12'h140 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6464 = 12'h140 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3392; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9536 = 12'h140 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6464; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12608 = 12'h140 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9536; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15680 = 12'h140 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12608; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18752 = 12'h140 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15680; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21824 = 12'h140 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18752; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24896 = 12'h140 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21824; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_320 = io_valid_in ? _GEN_24896 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_320 = 12'h140 == _T_2[11:0] ? image_320 : _GEN_319; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3393 = 12'h141 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6465 = 12'h141 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3393; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9537 = 12'h141 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6465; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12609 = 12'h141 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9537; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15681 = 12'h141 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12609; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18753 = 12'h141 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15681; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21825 = 12'h141 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18753; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24897 = 12'h141 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21825; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_321 = io_valid_in ? _GEN_24897 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_321 = 12'h141 == _T_2[11:0] ? image_321 : _GEN_320; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3394 = 12'h142 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6466 = 12'h142 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3394; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9538 = 12'h142 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6466; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12610 = 12'h142 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9538; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15682 = 12'h142 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12610; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18754 = 12'h142 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15682; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21826 = 12'h142 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18754; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24898 = 12'h142 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21826; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_322 = io_valid_in ? _GEN_24898 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_322 = 12'h142 == _T_2[11:0] ? image_322 : _GEN_321; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3395 = 12'h143 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6467 = 12'h143 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3395; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9539 = 12'h143 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6467; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12611 = 12'h143 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9539; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15683 = 12'h143 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12611; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18755 = 12'h143 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15683; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21827 = 12'h143 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18755; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24899 = 12'h143 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21827; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_323 = io_valid_in ? _GEN_24899 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_323 = 12'h143 == _T_2[11:0] ? image_323 : _GEN_322; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3396 = 12'h144 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6468 = 12'h144 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3396; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9540 = 12'h144 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6468; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12612 = 12'h144 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9540; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15684 = 12'h144 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12612; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18756 = 12'h144 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15684; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21828 = 12'h144 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18756; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24900 = 12'h144 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21828; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_324 = io_valid_in ? _GEN_24900 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_324 = 12'h144 == _T_2[11:0] ? image_324 : _GEN_323; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3397 = 12'h145 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6469 = 12'h145 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3397; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9541 = 12'h145 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6469; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12613 = 12'h145 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9541; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15685 = 12'h145 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12613; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18757 = 12'h145 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15685; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21829 = 12'h145 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18757; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24901 = 12'h145 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21829; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_325 = io_valid_in ? _GEN_24901 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_325 = 12'h145 == _T_2[11:0] ? image_325 : _GEN_324; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3398 = 12'h146 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6470 = 12'h146 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3398; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9542 = 12'h146 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6470; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12614 = 12'h146 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9542; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15686 = 12'h146 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12614; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18758 = 12'h146 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15686; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21830 = 12'h146 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18758; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24902 = 12'h146 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21830; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_326 = io_valid_in ? _GEN_24902 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_326 = 12'h146 == _T_2[11:0] ? image_326 : _GEN_325; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3399 = 12'h147 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6471 = 12'h147 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3399; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9543 = 12'h147 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6471; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12615 = 12'h147 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9543; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15687 = 12'h147 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12615; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18759 = 12'h147 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15687; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21831 = 12'h147 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18759; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24903 = 12'h147 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21831; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_327 = io_valid_in ? _GEN_24903 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_327 = 12'h147 == _T_2[11:0] ? image_327 : _GEN_326; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3400 = 12'h148 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6472 = 12'h148 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3400; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9544 = 12'h148 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6472; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12616 = 12'h148 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9544; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15688 = 12'h148 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12616; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18760 = 12'h148 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15688; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21832 = 12'h148 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18760; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24904 = 12'h148 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21832; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_328 = io_valid_in ? _GEN_24904 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_328 = 12'h148 == _T_2[11:0] ? image_328 : _GEN_327; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3401 = 12'h149 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6473 = 12'h149 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3401; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9545 = 12'h149 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6473; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12617 = 12'h149 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9545; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15689 = 12'h149 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12617; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18761 = 12'h149 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15689; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21833 = 12'h149 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18761; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24905 = 12'h149 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21833; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_329 = io_valid_in ? _GEN_24905 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_329 = 12'h149 == _T_2[11:0] ? image_329 : _GEN_328; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3402 = 12'h14a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6474 = 12'h14a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3402; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9546 = 12'h14a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6474; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12618 = 12'h14a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9546; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15690 = 12'h14a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12618; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18762 = 12'h14a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15690; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21834 = 12'h14a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18762; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24906 = 12'h14a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21834; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_330 = io_valid_in ? _GEN_24906 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_330 = 12'h14a == _T_2[11:0] ? image_330 : _GEN_329; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3403 = 12'h14b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6475 = 12'h14b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3403; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9547 = 12'h14b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6475; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12619 = 12'h14b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9547; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15691 = 12'h14b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12619; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18763 = 12'h14b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15691; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21835 = 12'h14b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18763; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24907 = 12'h14b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21835; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_331 = io_valid_in ? _GEN_24907 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_331 = 12'h14b == _T_2[11:0] ? image_331 : _GEN_330; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3404 = 12'h14c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6476 = 12'h14c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3404; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9548 = 12'h14c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6476; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12620 = 12'h14c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9548; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15692 = 12'h14c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12620; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18764 = 12'h14c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15692; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21836 = 12'h14c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18764; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24908 = 12'h14c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21836; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_332 = io_valid_in ? _GEN_24908 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_332 = 12'h14c == _T_2[11:0] ? image_332 : _GEN_331; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3405 = 12'h14d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6477 = 12'h14d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3405; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9549 = 12'h14d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6477; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12621 = 12'h14d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9549; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15693 = 12'h14d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12621; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18765 = 12'h14d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15693; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21837 = 12'h14d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18765; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24909 = 12'h14d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21837; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_333 = io_valid_in ? _GEN_24909 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_333 = 12'h14d == _T_2[11:0] ? image_333 : _GEN_332; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3406 = 12'h14e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6478 = 12'h14e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3406; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9550 = 12'h14e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6478; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12622 = 12'h14e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9550; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15694 = 12'h14e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12622; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18766 = 12'h14e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15694; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21838 = 12'h14e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18766; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24910 = 12'h14e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21838; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_334 = io_valid_in ? _GEN_24910 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_334 = 12'h14e == _T_2[11:0] ? image_334 : _GEN_333; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3407 = 12'h14f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6479 = 12'h14f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3407; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9551 = 12'h14f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6479; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12623 = 12'h14f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9551; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15695 = 12'h14f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12623; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18767 = 12'h14f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15695; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21839 = 12'h14f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18767; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24911 = 12'h14f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21839; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_335 = io_valid_in ? _GEN_24911 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_335 = 12'h14f == _T_2[11:0] ? image_335 : _GEN_334; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3408 = 12'h150 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6480 = 12'h150 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3408; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9552 = 12'h150 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6480; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12624 = 12'h150 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9552; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15696 = 12'h150 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12624; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18768 = 12'h150 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15696; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21840 = 12'h150 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18768; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24912 = 12'h150 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21840; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_336 = io_valid_in ? _GEN_24912 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_336 = 12'h150 == _T_2[11:0] ? image_336 : _GEN_335; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3409 = 12'h151 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6481 = 12'h151 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3409; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9553 = 12'h151 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6481; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12625 = 12'h151 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9553; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15697 = 12'h151 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12625; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18769 = 12'h151 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15697; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21841 = 12'h151 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18769; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24913 = 12'h151 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21841; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_337 = io_valid_in ? _GEN_24913 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_337 = 12'h151 == _T_2[11:0] ? image_337 : _GEN_336; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3410 = 12'h152 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6482 = 12'h152 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3410; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9554 = 12'h152 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6482; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12626 = 12'h152 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9554; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15698 = 12'h152 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12626; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18770 = 12'h152 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15698; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21842 = 12'h152 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18770; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24914 = 12'h152 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21842; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_338 = io_valid_in ? _GEN_24914 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_338 = 12'h152 == _T_2[11:0] ? image_338 : _GEN_337; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3411 = 12'h153 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6483 = 12'h153 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3411; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9555 = 12'h153 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6483; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12627 = 12'h153 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9555; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15699 = 12'h153 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12627; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18771 = 12'h153 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15699; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21843 = 12'h153 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18771; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24915 = 12'h153 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21843; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_339 = io_valid_in ? _GEN_24915 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_339 = 12'h153 == _T_2[11:0] ? image_339 : _GEN_338; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3412 = 12'h154 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6484 = 12'h154 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3412; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9556 = 12'h154 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6484; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12628 = 12'h154 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9556; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15700 = 12'h154 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12628; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18772 = 12'h154 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15700; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21844 = 12'h154 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18772; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24916 = 12'h154 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21844; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_340 = io_valid_in ? _GEN_24916 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_340 = 12'h154 == _T_2[11:0] ? image_340 : _GEN_339; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3413 = 12'h155 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6485 = 12'h155 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3413; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9557 = 12'h155 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6485; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12629 = 12'h155 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9557; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15701 = 12'h155 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12629; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18773 = 12'h155 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15701; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21845 = 12'h155 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18773; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24917 = 12'h155 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21845; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_341 = io_valid_in ? _GEN_24917 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_341 = 12'h155 == _T_2[11:0] ? image_341 : _GEN_340; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3414 = 12'h156 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6486 = 12'h156 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3414; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9558 = 12'h156 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6486; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12630 = 12'h156 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9558; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15702 = 12'h156 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12630; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18774 = 12'h156 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15702; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21846 = 12'h156 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18774; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24918 = 12'h156 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21846; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_342 = io_valid_in ? _GEN_24918 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_342 = 12'h156 == _T_2[11:0] ? image_342 : _GEN_341; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3415 = 12'h157 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6487 = 12'h157 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3415; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9559 = 12'h157 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6487; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12631 = 12'h157 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9559; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15703 = 12'h157 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12631; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18775 = 12'h157 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15703; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21847 = 12'h157 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18775; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24919 = 12'h157 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21847; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_343 = io_valid_in ? _GEN_24919 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_343 = 12'h157 == _T_2[11:0] ? image_343 : _GEN_342; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3416 = 12'h158 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6488 = 12'h158 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3416; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9560 = 12'h158 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6488; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12632 = 12'h158 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9560; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15704 = 12'h158 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12632; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18776 = 12'h158 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15704; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21848 = 12'h158 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18776; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24920 = 12'h158 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21848; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_344 = io_valid_in ? _GEN_24920 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_344 = 12'h158 == _T_2[11:0] ? image_344 : _GEN_343; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3417 = 12'h159 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6489 = 12'h159 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3417; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9561 = 12'h159 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6489; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12633 = 12'h159 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9561; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15705 = 12'h159 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12633; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18777 = 12'h159 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15705; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21849 = 12'h159 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18777; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24921 = 12'h159 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21849; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_345 = io_valid_in ? _GEN_24921 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_345 = 12'h159 == _T_2[11:0] ? image_345 : _GEN_344; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3418 = 12'h15a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6490 = 12'h15a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3418; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9562 = 12'h15a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6490; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12634 = 12'h15a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9562; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15706 = 12'h15a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12634; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18778 = 12'h15a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15706; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21850 = 12'h15a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18778; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24922 = 12'h15a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21850; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_346 = io_valid_in ? _GEN_24922 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_346 = 12'h15a == _T_2[11:0] ? image_346 : _GEN_345; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3419 = 12'h15b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6491 = 12'h15b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3419; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9563 = 12'h15b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6491; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12635 = 12'h15b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9563; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15707 = 12'h15b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12635; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18779 = 12'h15b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15707; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21851 = 12'h15b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18779; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24923 = 12'h15b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21851; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_347 = io_valid_in ? _GEN_24923 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_347 = 12'h15b == _T_2[11:0] ? image_347 : _GEN_346; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3420 = 12'h15c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6492 = 12'h15c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3420; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9564 = 12'h15c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6492; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12636 = 12'h15c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9564; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15708 = 12'h15c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12636; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18780 = 12'h15c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15708; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21852 = 12'h15c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18780; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24924 = 12'h15c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21852; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_348 = io_valid_in ? _GEN_24924 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_348 = 12'h15c == _T_2[11:0] ? image_348 : _GEN_347; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3421 = 12'h15d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6493 = 12'h15d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3421; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9565 = 12'h15d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6493; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12637 = 12'h15d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9565; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15709 = 12'h15d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12637; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18781 = 12'h15d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15709; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21853 = 12'h15d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18781; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24925 = 12'h15d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21853; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_349 = io_valid_in ? _GEN_24925 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_349 = 12'h15d == _T_2[11:0] ? image_349 : _GEN_348; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3422 = 12'h15e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6494 = 12'h15e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3422; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9566 = 12'h15e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6494; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12638 = 12'h15e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9566; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15710 = 12'h15e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12638; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18782 = 12'h15e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15710; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21854 = 12'h15e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18782; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24926 = 12'h15e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21854; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_350 = io_valid_in ? _GEN_24926 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_350 = 12'h15e == _T_2[11:0] ? image_350 : _GEN_349; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3423 = 12'h15f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6495 = 12'h15f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3423; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9567 = 12'h15f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6495; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12639 = 12'h15f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9567; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15711 = 12'h15f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12639; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18783 = 12'h15f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15711; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21855 = 12'h15f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18783; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24927 = 12'h15f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21855; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_351 = io_valid_in ? _GEN_24927 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_351 = 12'h15f == _T_2[11:0] ? image_351 : _GEN_350; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3424 = 12'h160 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6496 = 12'h160 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3424; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9568 = 12'h160 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6496; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12640 = 12'h160 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9568; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15712 = 12'h160 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12640; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18784 = 12'h160 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15712; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21856 = 12'h160 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18784; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24928 = 12'h160 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21856; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_352 = io_valid_in ? _GEN_24928 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_352 = 12'h160 == _T_2[11:0] ? image_352 : _GEN_351; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3425 = 12'h161 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6497 = 12'h161 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3425; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9569 = 12'h161 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6497; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12641 = 12'h161 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9569; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15713 = 12'h161 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12641; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18785 = 12'h161 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15713; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21857 = 12'h161 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18785; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24929 = 12'h161 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21857; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_353 = io_valid_in ? _GEN_24929 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_353 = 12'h161 == _T_2[11:0] ? image_353 : _GEN_352; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3426 = 12'h162 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6498 = 12'h162 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3426; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9570 = 12'h162 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6498; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12642 = 12'h162 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9570; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15714 = 12'h162 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12642; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18786 = 12'h162 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15714; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21858 = 12'h162 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18786; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24930 = 12'h162 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21858; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_354 = io_valid_in ? _GEN_24930 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_354 = 12'h162 == _T_2[11:0] ? image_354 : _GEN_353; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3427 = 12'h163 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6499 = 12'h163 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3427; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9571 = 12'h163 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6499; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12643 = 12'h163 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9571; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15715 = 12'h163 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12643; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18787 = 12'h163 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15715; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21859 = 12'h163 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18787; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24931 = 12'h163 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21859; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_355 = io_valid_in ? _GEN_24931 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_355 = 12'h163 == _T_2[11:0] ? image_355 : _GEN_354; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3428 = 12'h164 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6500 = 12'h164 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3428; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9572 = 12'h164 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6500; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12644 = 12'h164 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9572; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15716 = 12'h164 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12644; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18788 = 12'h164 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15716; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21860 = 12'h164 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18788; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24932 = 12'h164 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21860; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_356 = io_valid_in ? _GEN_24932 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_356 = 12'h164 == _T_2[11:0] ? image_356 : _GEN_355; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3429 = 12'h165 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6501 = 12'h165 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3429; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9573 = 12'h165 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6501; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12645 = 12'h165 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9573; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15717 = 12'h165 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12645; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18789 = 12'h165 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15717; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21861 = 12'h165 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18789; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24933 = 12'h165 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21861; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_357 = io_valid_in ? _GEN_24933 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_357 = 12'h165 == _T_2[11:0] ? image_357 : _GEN_356; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3430 = 12'h166 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6502 = 12'h166 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3430; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9574 = 12'h166 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6502; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12646 = 12'h166 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9574; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15718 = 12'h166 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12646; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18790 = 12'h166 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15718; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21862 = 12'h166 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18790; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24934 = 12'h166 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21862; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_358 = io_valid_in ? _GEN_24934 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_358 = 12'h166 == _T_2[11:0] ? image_358 : _GEN_357; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3431 = 12'h167 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6503 = 12'h167 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3431; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9575 = 12'h167 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6503; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12647 = 12'h167 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9575; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15719 = 12'h167 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12647; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18791 = 12'h167 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15719; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21863 = 12'h167 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18791; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24935 = 12'h167 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21863; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_359 = io_valid_in ? _GEN_24935 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_359 = 12'h167 == _T_2[11:0] ? image_359 : _GEN_358; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3432 = 12'h168 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6504 = 12'h168 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3432; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9576 = 12'h168 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6504; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12648 = 12'h168 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9576; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15720 = 12'h168 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12648; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18792 = 12'h168 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15720; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21864 = 12'h168 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18792; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24936 = 12'h168 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21864; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_360 = io_valid_in ? _GEN_24936 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_360 = 12'h168 == _T_2[11:0] ? image_360 : _GEN_359; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3433 = 12'h169 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6505 = 12'h169 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3433; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9577 = 12'h169 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6505; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12649 = 12'h169 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9577; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15721 = 12'h169 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12649; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18793 = 12'h169 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15721; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21865 = 12'h169 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18793; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24937 = 12'h169 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21865; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_361 = io_valid_in ? _GEN_24937 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_361 = 12'h169 == _T_2[11:0] ? image_361 : _GEN_360; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3434 = 12'h16a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6506 = 12'h16a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3434; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9578 = 12'h16a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6506; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12650 = 12'h16a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9578; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15722 = 12'h16a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12650; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18794 = 12'h16a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15722; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21866 = 12'h16a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18794; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24938 = 12'h16a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21866; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_362 = io_valid_in ? _GEN_24938 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_362 = 12'h16a == _T_2[11:0] ? image_362 : _GEN_361; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3435 = 12'h16b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6507 = 12'h16b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3435; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9579 = 12'h16b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6507; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12651 = 12'h16b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9579; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15723 = 12'h16b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12651; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18795 = 12'h16b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15723; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21867 = 12'h16b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18795; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24939 = 12'h16b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21867; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_363 = io_valid_in ? _GEN_24939 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_363 = 12'h16b == _T_2[11:0] ? image_363 : _GEN_362; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3436 = 12'h16c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6508 = 12'h16c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3436; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9580 = 12'h16c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6508; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12652 = 12'h16c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9580; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15724 = 12'h16c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12652; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18796 = 12'h16c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15724; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21868 = 12'h16c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18796; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24940 = 12'h16c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21868; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_364 = io_valid_in ? _GEN_24940 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_364 = 12'h16c == _T_2[11:0] ? image_364 : _GEN_363; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3437 = 12'h16d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6509 = 12'h16d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3437; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9581 = 12'h16d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6509; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12653 = 12'h16d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9581; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15725 = 12'h16d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12653; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18797 = 12'h16d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15725; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21869 = 12'h16d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18797; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24941 = 12'h16d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21869; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_365 = io_valid_in ? _GEN_24941 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_365 = 12'h16d == _T_2[11:0] ? image_365 : _GEN_364; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3438 = 12'h16e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6510 = 12'h16e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3438; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9582 = 12'h16e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6510; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12654 = 12'h16e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9582; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15726 = 12'h16e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12654; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18798 = 12'h16e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15726; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21870 = 12'h16e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18798; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24942 = 12'h16e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21870; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_366 = io_valid_in ? _GEN_24942 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_366 = 12'h16e == _T_2[11:0] ? image_366 : _GEN_365; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3439 = 12'h16f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6511 = 12'h16f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3439; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9583 = 12'h16f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6511; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12655 = 12'h16f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9583; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15727 = 12'h16f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12655; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18799 = 12'h16f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15727; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21871 = 12'h16f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18799; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24943 = 12'h16f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21871; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_367 = io_valid_in ? _GEN_24943 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_367 = 12'h16f == _T_2[11:0] ? image_367 : _GEN_366; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3440 = 12'h170 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6512 = 12'h170 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3440; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9584 = 12'h170 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6512; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12656 = 12'h170 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9584; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15728 = 12'h170 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12656; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18800 = 12'h170 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15728; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21872 = 12'h170 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18800; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24944 = 12'h170 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21872; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_368 = io_valid_in ? _GEN_24944 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_368 = 12'h170 == _T_2[11:0] ? image_368 : _GEN_367; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3441 = 12'h171 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6513 = 12'h171 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3441; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9585 = 12'h171 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6513; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12657 = 12'h171 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9585; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15729 = 12'h171 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12657; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18801 = 12'h171 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15729; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21873 = 12'h171 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18801; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24945 = 12'h171 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21873; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_369 = io_valid_in ? _GEN_24945 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_369 = 12'h171 == _T_2[11:0] ? image_369 : _GEN_368; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3442 = 12'h172 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6514 = 12'h172 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3442; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9586 = 12'h172 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6514; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12658 = 12'h172 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9586; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15730 = 12'h172 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12658; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18802 = 12'h172 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15730; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21874 = 12'h172 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18802; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24946 = 12'h172 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21874; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_370 = io_valid_in ? _GEN_24946 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_370 = 12'h172 == _T_2[11:0] ? image_370 : _GEN_369; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3443 = 12'h173 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6515 = 12'h173 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3443; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9587 = 12'h173 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6515; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12659 = 12'h173 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9587; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15731 = 12'h173 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12659; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18803 = 12'h173 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15731; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21875 = 12'h173 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18803; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24947 = 12'h173 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21875; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_371 = io_valid_in ? _GEN_24947 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_371 = 12'h173 == _T_2[11:0] ? image_371 : _GEN_370; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3444 = 12'h174 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6516 = 12'h174 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3444; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9588 = 12'h174 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6516; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12660 = 12'h174 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9588; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15732 = 12'h174 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12660; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18804 = 12'h174 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15732; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21876 = 12'h174 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18804; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24948 = 12'h174 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21876; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_372 = io_valid_in ? _GEN_24948 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_372 = 12'h174 == _T_2[11:0] ? image_372 : _GEN_371; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3445 = 12'h175 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6517 = 12'h175 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3445; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9589 = 12'h175 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6517; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12661 = 12'h175 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9589; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15733 = 12'h175 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12661; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18805 = 12'h175 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15733; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21877 = 12'h175 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18805; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24949 = 12'h175 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21877; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_373 = io_valid_in ? _GEN_24949 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_373 = 12'h175 == _T_2[11:0] ? image_373 : _GEN_372; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3446 = 12'h176 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6518 = 12'h176 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3446; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9590 = 12'h176 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6518; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12662 = 12'h176 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9590; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15734 = 12'h176 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12662; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18806 = 12'h176 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15734; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21878 = 12'h176 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18806; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24950 = 12'h176 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21878; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_374 = io_valid_in ? _GEN_24950 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_374 = 12'h176 == _T_2[11:0] ? image_374 : _GEN_373; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3447 = 12'h177 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6519 = 12'h177 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3447; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9591 = 12'h177 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6519; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12663 = 12'h177 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9591; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15735 = 12'h177 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12663; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18807 = 12'h177 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15735; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21879 = 12'h177 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18807; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24951 = 12'h177 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21879; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_375 = io_valid_in ? _GEN_24951 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_375 = 12'h177 == _T_2[11:0] ? image_375 : _GEN_374; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3448 = 12'h178 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6520 = 12'h178 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3448; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9592 = 12'h178 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6520; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12664 = 12'h178 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9592; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15736 = 12'h178 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12664; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18808 = 12'h178 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15736; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21880 = 12'h178 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18808; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24952 = 12'h178 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21880; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_376 = io_valid_in ? _GEN_24952 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_376 = 12'h178 == _T_2[11:0] ? image_376 : _GEN_375; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3449 = 12'h179 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6521 = 12'h179 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3449; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9593 = 12'h179 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6521; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12665 = 12'h179 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9593; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15737 = 12'h179 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12665; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18809 = 12'h179 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15737; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21881 = 12'h179 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18809; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24953 = 12'h179 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21881; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_377 = io_valid_in ? _GEN_24953 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_377 = 12'h179 == _T_2[11:0] ? image_377 : _GEN_376; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3450 = 12'h17a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6522 = 12'h17a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3450; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9594 = 12'h17a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6522; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12666 = 12'h17a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9594; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15738 = 12'h17a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12666; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18810 = 12'h17a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15738; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21882 = 12'h17a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18810; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24954 = 12'h17a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21882; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_378 = io_valid_in ? _GEN_24954 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_378 = 12'h17a == _T_2[11:0] ? image_378 : _GEN_377; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3451 = 12'h17b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6523 = 12'h17b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3451; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9595 = 12'h17b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6523; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12667 = 12'h17b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9595; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15739 = 12'h17b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12667; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18811 = 12'h17b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15739; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21883 = 12'h17b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18811; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24955 = 12'h17b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21883; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_379 = io_valid_in ? _GEN_24955 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_379 = 12'h17b == _T_2[11:0] ? image_379 : _GEN_378; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3452 = 12'h17c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6524 = 12'h17c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3452; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9596 = 12'h17c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6524; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12668 = 12'h17c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9596; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15740 = 12'h17c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12668; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18812 = 12'h17c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15740; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21884 = 12'h17c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18812; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24956 = 12'h17c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21884; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_380 = io_valid_in ? _GEN_24956 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_380 = 12'h17c == _T_2[11:0] ? image_380 : _GEN_379; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3453 = 12'h17d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6525 = 12'h17d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3453; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9597 = 12'h17d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6525; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12669 = 12'h17d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9597; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15741 = 12'h17d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12669; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18813 = 12'h17d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15741; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21885 = 12'h17d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18813; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24957 = 12'h17d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21885; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_381 = io_valid_in ? _GEN_24957 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_381 = 12'h17d == _T_2[11:0] ? image_381 : _GEN_380; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3454 = 12'h17e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6526 = 12'h17e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3454; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9598 = 12'h17e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6526; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12670 = 12'h17e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9598; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15742 = 12'h17e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12670; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18814 = 12'h17e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15742; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21886 = 12'h17e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18814; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24958 = 12'h17e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21886; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_382 = io_valid_in ? _GEN_24958 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_382 = 12'h17e == _T_2[11:0] ? image_382 : _GEN_381; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3455 = 12'h17f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6527 = 12'h17f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3455; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9599 = 12'h17f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6527; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12671 = 12'h17f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9599; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15743 = 12'h17f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12671; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18815 = 12'h17f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15743; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21887 = 12'h17f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18815; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24959 = 12'h17f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21887; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_383 = io_valid_in ? _GEN_24959 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_383 = 12'h17f == _T_2[11:0] ? image_383 : _GEN_382; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3456 = 12'h180 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6528 = 12'h180 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3456; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9600 = 12'h180 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6528; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12672 = 12'h180 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9600; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15744 = 12'h180 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12672; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18816 = 12'h180 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15744; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21888 = 12'h180 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18816; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24960 = 12'h180 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21888; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_384 = io_valid_in ? _GEN_24960 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_384 = 12'h180 == _T_2[11:0] ? image_384 : _GEN_383; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3457 = 12'h181 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6529 = 12'h181 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3457; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9601 = 12'h181 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6529; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12673 = 12'h181 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9601; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15745 = 12'h181 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12673; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18817 = 12'h181 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15745; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21889 = 12'h181 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18817; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24961 = 12'h181 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21889; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_385 = io_valid_in ? _GEN_24961 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_385 = 12'h181 == _T_2[11:0] ? image_385 : _GEN_384; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3458 = 12'h182 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6530 = 12'h182 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3458; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9602 = 12'h182 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6530; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12674 = 12'h182 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9602; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15746 = 12'h182 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12674; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18818 = 12'h182 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15746; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21890 = 12'h182 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18818; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24962 = 12'h182 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21890; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_386 = io_valid_in ? _GEN_24962 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_386 = 12'h182 == _T_2[11:0] ? image_386 : _GEN_385; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3459 = 12'h183 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6531 = 12'h183 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3459; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9603 = 12'h183 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6531; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12675 = 12'h183 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9603; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15747 = 12'h183 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12675; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18819 = 12'h183 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15747; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21891 = 12'h183 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18819; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24963 = 12'h183 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21891; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_387 = io_valid_in ? _GEN_24963 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_387 = 12'h183 == _T_2[11:0] ? image_387 : _GEN_386; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3460 = 12'h184 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6532 = 12'h184 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3460; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9604 = 12'h184 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6532; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12676 = 12'h184 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9604; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15748 = 12'h184 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12676; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18820 = 12'h184 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15748; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21892 = 12'h184 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18820; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24964 = 12'h184 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21892; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_388 = io_valid_in ? _GEN_24964 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_388 = 12'h184 == _T_2[11:0] ? image_388 : _GEN_387; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3461 = 12'h185 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6533 = 12'h185 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3461; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9605 = 12'h185 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6533; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12677 = 12'h185 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9605; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15749 = 12'h185 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12677; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18821 = 12'h185 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15749; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21893 = 12'h185 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18821; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24965 = 12'h185 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21893; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_389 = io_valid_in ? _GEN_24965 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_389 = 12'h185 == _T_2[11:0] ? image_389 : _GEN_388; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3462 = 12'h186 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6534 = 12'h186 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3462; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9606 = 12'h186 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6534; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12678 = 12'h186 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9606; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15750 = 12'h186 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12678; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18822 = 12'h186 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15750; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21894 = 12'h186 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18822; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24966 = 12'h186 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21894; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_390 = io_valid_in ? _GEN_24966 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_390 = 12'h186 == _T_2[11:0] ? image_390 : _GEN_389; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3463 = 12'h187 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6535 = 12'h187 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3463; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9607 = 12'h187 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6535; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12679 = 12'h187 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9607; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15751 = 12'h187 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12679; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18823 = 12'h187 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15751; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21895 = 12'h187 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18823; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24967 = 12'h187 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21895; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_391 = io_valid_in ? _GEN_24967 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_391 = 12'h187 == _T_2[11:0] ? image_391 : _GEN_390; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3464 = 12'h188 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6536 = 12'h188 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3464; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9608 = 12'h188 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6536; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12680 = 12'h188 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9608; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15752 = 12'h188 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12680; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18824 = 12'h188 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15752; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21896 = 12'h188 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18824; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24968 = 12'h188 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21896; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_392 = io_valid_in ? _GEN_24968 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_392 = 12'h188 == _T_2[11:0] ? image_392 : _GEN_391; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3465 = 12'h189 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6537 = 12'h189 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3465; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9609 = 12'h189 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6537; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12681 = 12'h189 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9609; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15753 = 12'h189 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12681; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18825 = 12'h189 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15753; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21897 = 12'h189 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18825; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24969 = 12'h189 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21897; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_393 = io_valid_in ? _GEN_24969 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_393 = 12'h189 == _T_2[11:0] ? image_393 : _GEN_392; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3466 = 12'h18a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6538 = 12'h18a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3466; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9610 = 12'h18a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6538; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12682 = 12'h18a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9610; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15754 = 12'h18a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12682; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18826 = 12'h18a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15754; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21898 = 12'h18a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18826; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24970 = 12'h18a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21898; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_394 = io_valid_in ? _GEN_24970 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_394 = 12'h18a == _T_2[11:0] ? image_394 : _GEN_393; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3467 = 12'h18b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6539 = 12'h18b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3467; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9611 = 12'h18b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6539; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12683 = 12'h18b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9611; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15755 = 12'h18b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12683; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18827 = 12'h18b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15755; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21899 = 12'h18b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18827; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24971 = 12'h18b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21899; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_395 = io_valid_in ? _GEN_24971 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_395 = 12'h18b == _T_2[11:0] ? image_395 : _GEN_394; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3468 = 12'h18c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6540 = 12'h18c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3468; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9612 = 12'h18c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6540; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12684 = 12'h18c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9612; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15756 = 12'h18c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12684; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18828 = 12'h18c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15756; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21900 = 12'h18c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18828; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24972 = 12'h18c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21900; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_396 = io_valid_in ? _GEN_24972 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_396 = 12'h18c == _T_2[11:0] ? image_396 : _GEN_395; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3469 = 12'h18d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6541 = 12'h18d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3469; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9613 = 12'h18d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6541; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12685 = 12'h18d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9613; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15757 = 12'h18d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12685; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18829 = 12'h18d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15757; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21901 = 12'h18d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18829; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24973 = 12'h18d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21901; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_397 = io_valid_in ? _GEN_24973 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_397 = 12'h18d == _T_2[11:0] ? image_397 : _GEN_396; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3470 = 12'h18e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6542 = 12'h18e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3470; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9614 = 12'h18e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6542; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12686 = 12'h18e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9614; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15758 = 12'h18e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12686; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18830 = 12'h18e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15758; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21902 = 12'h18e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18830; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24974 = 12'h18e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21902; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_398 = io_valid_in ? _GEN_24974 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_398 = 12'h18e == _T_2[11:0] ? image_398 : _GEN_397; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3471 = 12'h18f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6543 = 12'h18f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3471; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9615 = 12'h18f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6543; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12687 = 12'h18f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9615; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15759 = 12'h18f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12687; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18831 = 12'h18f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15759; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21903 = 12'h18f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18831; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24975 = 12'h18f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21903; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_399 = io_valid_in ? _GEN_24975 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_399 = 12'h18f == _T_2[11:0] ? image_399 : _GEN_398; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3472 = 12'h190 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6544 = 12'h190 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3472; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9616 = 12'h190 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6544; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12688 = 12'h190 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9616; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15760 = 12'h190 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12688; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18832 = 12'h190 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15760; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21904 = 12'h190 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18832; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24976 = 12'h190 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21904; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_400 = io_valid_in ? _GEN_24976 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_400 = 12'h190 == _T_2[11:0] ? image_400 : _GEN_399; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3473 = 12'h191 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6545 = 12'h191 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3473; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9617 = 12'h191 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6545; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12689 = 12'h191 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9617; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15761 = 12'h191 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12689; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18833 = 12'h191 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15761; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21905 = 12'h191 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18833; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24977 = 12'h191 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21905; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_401 = io_valid_in ? _GEN_24977 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_401 = 12'h191 == _T_2[11:0] ? image_401 : _GEN_400; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3474 = 12'h192 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6546 = 12'h192 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3474; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9618 = 12'h192 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6546; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12690 = 12'h192 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9618; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15762 = 12'h192 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12690; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18834 = 12'h192 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15762; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21906 = 12'h192 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18834; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24978 = 12'h192 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21906; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_402 = io_valid_in ? _GEN_24978 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_402 = 12'h192 == _T_2[11:0] ? image_402 : _GEN_401; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3475 = 12'h193 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6547 = 12'h193 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3475; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9619 = 12'h193 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6547; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12691 = 12'h193 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9619; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15763 = 12'h193 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12691; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18835 = 12'h193 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15763; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21907 = 12'h193 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18835; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24979 = 12'h193 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21907; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_403 = io_valid_in ? _GEN_24979 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_403 = 12'h193 == _T_2[11:0] ? image_403 : _GEN_402; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3476 = 12'h194 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6548 = 12'h194 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3476; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9620 = 12'h194 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6548; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12692 = 12'h194 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9620; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15764 = 12'h194 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12692; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18836 = 12'h194 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15764; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21908 = 12'h194 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18836; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24980 = 12'h194 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21908; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_404 = io_valid_in ? _GEN_24980 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_404 = 12'h194 == _T_2[11:0] ? image_404 : _GEN_403; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3477 = 12'h195 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6549 = 12'h195 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3477; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9621 = 12'h195 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6549; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12693 = 12'h195 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9621; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15765 = 12'h195 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12693; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18837 = 12'h195 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15765; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21909 = 12'h195 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18837; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24981 = 12'h195 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21909; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_405 = io_valid_in ? _GEN_24981 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_405 = 12'h195 == _T_2[11:0] ? image_405 : _GEN_404; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3478 = 12'h196 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6550 = 12'h196 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3478; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9622 = 12'h196 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6550; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12694 = 12'h196 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9622; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15766 = 12'h196 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12694; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18838 = 12'h196 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15766; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21910 = 12'h196 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18838; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24982 = 12'h196 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21910; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_406 = io_valid_in ? _GEN_24982 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_406 = 12'h196 == _T_2[11:0] ? image_406 : _GEN_405; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3479 = 12'h197 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6551 = 12'h197 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3479; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9623 = 12'h197 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6551; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12695 = 12'h197 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9623; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15767 = 12'h197 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12695; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18839 = 12'h197 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15767; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21911 = 12'h197 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18839; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24983 = 12'h197 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21911; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_407 = io_valid_in ? _GEN_24983 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_407 = 12'h197 == _T_2[11:0] ? image_407 : _GEN_406; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3480 = 12'h198 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6552 = 12'h198 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3480; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9624 = 12'h198 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6552; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12696 = 12'h198 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9624; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15768 = 12'h198 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12696; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18840 = 12'h198 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15768; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21912 = 12'h198 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18840; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24984 = 12'h198 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21912; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_408 = io_valid_in ? _GEN_24984 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_408 = 12'h198 == _T_2[11:0] ? image_408 : _GEN_407; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3481 = 12'h199 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6553 = 12'h199 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3481; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9625 = 12'h199 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6553; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12697 = 12'h199 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9625; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15769 = 12'h199 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12697; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18841 = 12'h199 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15769; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21913 = 12'h199 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18841; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24985 = 12'h199 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21913; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_409 = io_valid_in ? _GEN_24985 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_409 = 12'h199 == _T_2[11:0] ? image_409 : _GEN_408; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3482 = 12'h19a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6554 = 12'h19a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3482; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9626 = 12'h19a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6554; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12698 = 12'h19a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9626; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15770 = 12'h19a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12698; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18842 = 12'h19a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15770; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21914 = 12'h19a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18842; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24986 = 12'h19a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21914; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_410 = io_valid_in ? _GEN_24986 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_410 = 12'h19a == _T_2[11:0] ? image_410 : _GEN_409; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3483 = 12'h19b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6555 = 12'h19b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3483; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9627 = 12'h19b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6555; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12699 = 12'h19b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9627; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15771 = 12'h19b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12699; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18843 = 12'h19b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15771; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21915 = 12'h19b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18843; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24987 = 12'h19b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21915; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_411 = io_valid_in ? _GEN_24987 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_411 = 12'h19b == _T_2[11:0] ? image_411 : _GEN_410; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3484 = 12'h19c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6556 = 12'h19c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3484; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9628 = 12'h19c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6556; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12700 = 12'h19c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9628; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15772 = 12'h19c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12700; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18844 = 12'h19c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15772; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21916 = 12'h19c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18844; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24988 = 12'h19c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21916; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_412 = io_valid_in ? _GEN_24988 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_412 = 12'h19c == _T_2[11:0] ? image_412 : _GEN_411; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3485 = 12'h19d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6557 = 12'h19d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3485; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9629 = 12'h19d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6557; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12701 = 12'h19d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9629; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15773 = 12'h19d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12701; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18845 = 12'h19d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15773; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21917 = 12'h19d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18845; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24989 = 12'h19d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21917; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_413 = io_valid_in ? _GEN_24989 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_413 = 12'h19d == _T_2[11:0] ? image_413 : _GEN_412; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3486 = 12'h19e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6558 = 12'h19e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3486; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9630 = 12'h19e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6558; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12702 = 12'h19e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9630; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15774 = 12'h19e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12702; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18846 = 12'h19e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15774; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21918 = 12'h19e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18846; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24990 = 12'h19e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21918; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_414 = io_valid_in ? _GEN_24990 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_414 = 12'h19e == _T_2[11:0] ? image_414 : _GEN_413; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3487 = 12'h19f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6559 = 12'h19f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3487; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9631 = 12'h19f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6559; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12703 = 12'h19f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9631; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15775 = 12'h19f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12703; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18847 = 12'h19f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15775; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21919 = 12'h19f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18847; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24991 = 12'h19f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21919; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_415 = io_valid_in ? _GEN_24991 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_415 = 12'h19f == _T_2[11:0] ? image_415 : _GEN_414; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3488 = 12'h1a0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6560 = 12'h1a0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3488; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9632 = 12'h1a0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6560; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12704 = 12'h1a0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9632; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15776 = 12'h1a0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12704; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18848 = 12'h1a0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15776; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21920 = 12'h1a0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18848; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24992 = 12'h1a0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21920; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_416 = io_valid_in ? _GEN_24992 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_416 = 12'h1a0 == _T_2[11:0] ? image_416 : _GEN_415; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3489 = 12'h1a1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6561 = 12'h1a1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3489; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9633 = 12'h1a1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6561; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12705 = 12'h1a1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9633; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15777 = 12'h1a1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12705; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18849 = 12'h1a1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15777; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21921 = 12'h1a1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18849; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24993 = 12'h1a1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21921; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_417 = io_valid_in ? _GEN_24993 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_417 = 12'h1a1 == _T_2[11:0] ? image_417 : _GEN_416; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3490 = 12'h1a2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6562 = 12'h1a2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3490; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9634 = 12'h1a2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6562; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12706 = 12'h1a2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9634; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15778 = 12'h1a2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12706; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18850 = 12'h1a2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15778; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21922 = 12'h1a2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18850; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24994 = 12'h1a2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21922; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_418 = io_valid_in ? _GEN_24994 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_418 = 12'h1a2 == _T_2[11:0] ? image_418 : _GEN_417; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3491 = 12'h1a3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6563 = 12'h1a3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3491; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9635 = 12'h1a3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6563; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12707 = 12'h1a3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9635; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15779 = 12'h1a3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12707; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18851 = 12'h1a3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15779; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21923 = 12'h1a3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18851; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24995 = 12'h1a3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21923; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_419 = io_valid_in ? _GEN_24995 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_419 = 12'h1a3 == _T_2[11:0] ? image_419 : _GEN_418; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3492 = 12'h1a4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6564 = 12'h1a4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3492; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9636 = 12'h1a4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6564; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12708 = 12'h1a4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9636; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15780 = 12'h1a4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12708; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18852 = 12'h1a4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15780; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21924 = 12'h1a4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18852; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24996 = 12'h1a4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21924; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_420 = io_valid_in ? _GEN_24996 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_420 = 12'h1a4 == _T_2[11:0] ? image_420 : _GEN_419; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3493 = 12'h1a5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6565 = 12'h1a5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3493; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9637 = 12'h1a5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6565; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12709 = 12'h1a5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9637; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15781 = 12'h1a5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12709; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18853 = 12'h1a5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15781; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21925 = 12'h1a5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18853; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24997 = 12'h1a5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21925; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_421 = io_valid_in ? _GEN_24997 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_421 = 12'h1a5 == _T_2[11:0] ? image_421 : _GEN_420; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3494 = 12'h1a6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6566 = 12'h1a6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3494; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9638 = 12'h1a6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6566; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12710 = 12'h1a6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9638; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15782 = 12'h1a6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12710; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18854 = 12'h1a6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15782; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21926 = 12'h1a6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18854; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24998 = 12'h1a6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21926; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_422 = io_valid_in ? _GEN_24998 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_422 = 12'h1a6 == _T_2[11:0] ? image_422 : _GEN_421; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3495 = 12'h1a7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6567 = 12'h1a7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3495; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9639 = 12'h1a7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6567; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12711 = 12'h1a7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9639; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15783 = 12'h1a7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12711; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18855 = 12'h1a7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15783; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21927 = 12'h1a7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18855; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24999 = 12'h1a7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21927; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_423 = io_valid_in ? _GEN_24999 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_423 = 12'h1a7 == _T_2[11:0] ? image_423 : _GEN_422; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3496 = 12'h1a8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6568 = 12'h1a8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3496; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9640 = 12'h1a8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6568; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12712 = 12'h1a8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9640; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15784 = 12'h1a8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12712; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18856 = 12'h1a8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15784; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21928 = 12'h1a8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18856; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25000 = 12'h1a8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21928; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_424 = io_valid_in ? _GEN_25000 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_424 = 12'h1a8 == _T_2[11:0] ? image_424 : _GEN_423; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3497 = 12'h1a9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6569 = 12'h1a9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3497; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9641 = 12'h1a9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6569; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12713 = 12'h1a9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9641; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15785 = 12'h1a9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12713; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18857 = 12'h1a9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15785; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21929 = 12'h1a9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18857; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25001 = 12'h1a9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21929; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_425 = io_valid_in ? _GEN_25001 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_425 = 12'h1a9 == _T_2[11:0] ? image_425 : _GEN_424; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3498 = 12'h1aa == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6570 = 12'h1aa == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3498; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9642 = 12'h1aa == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6570; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12714 = 12'h1aa == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9642; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15786 = 12'h1aa == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12714; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18858 = 12'h1aa == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15786; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21930 = 12'h1aa == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18858; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25002 = 12'h1aa == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21930; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_426 = io_valid_in ? _GEN_25002 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_426 = 12'h1aa == _T_2[11:0] ? image_426 : _GEN_425; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3499 = 12'h1ab == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6571 = 12'h1ab == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3499; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9643 = 12'h1ab == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6571; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12715 = 12'h1ab == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9643; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15787 = 12'h1ab == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12715; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18859 = 12'h1ab == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15787; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21931 = 12'h1ab == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18859; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25003 = 12'h1ab == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21931; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_427 = io_valid_in ? _GEN_25003 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_427 = 12'h1ab == _T_2[11:0] ? image_427 : _GEN_426; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3500 = 12'h1ac == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6572 = 12'h1ac == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3500; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9644 = 12'h1ac == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6572; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12716 = 12'h1ac == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9644; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15788 = 12'h1ac == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12716; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18860 = 12'h1ac == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15788; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21932 = 12'h1ac == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18860; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25004 = 12'h1ac == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21932; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_428 = io_valid_in ? _GEN_25004 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_428 = 12'h1ac == _T_2[11:0] ? image_428 : _GEN_427; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3501 = 12'h1ad == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6573 = 12'h1ad == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3501; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9645 = 12'h1ad == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6573; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12717 = 12'h1ad == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9645; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15789 = 12'h1ad == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12717; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18861 = 12'h1ad == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15789; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21933 = 12'h1ad == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18861; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25005 = 12'h1ad == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21933; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_429 = io_valid_in ? _GEN_25005 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_429 = 12'h1ad == _T_2[11:0] ? image_429 : _GEN_428; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3502 = 12'h1ae == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6574 = 12'h1ae == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3502; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9646 = 12'h1ae == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6574; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12718 = 12'h1ae == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9646; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15790 = 12'h1ae == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12718; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18862 = 12'h1ae == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15790; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21934 = 12'h1ae == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18862; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25006 = 12'h1ae == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21934; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_430 = io_valid_in ? _GEN_25006 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_430 = 12'h1ae == _T_2[11:0] ? image_430 : _GEN_429; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3503 = 12'h1af == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6575 = 12'h1af == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3503; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9647 = 12'h1af == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6575; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12719 = 12'h1af == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9647; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15791 = 12'h1af == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12719; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18863 = 12'h1af == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15791; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21935 = 12'h1af == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18863; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25007 = 12'h1af == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21935; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_431 = io_valid_in ? _GEN_25007 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_431 = 12'h1af == _T_2[11:0] ? image_431 : _GEN_430; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3504 = 12'h1b0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6576 = 12'h1b0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3504; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9648 = 12'h1b0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6576; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12720 = 12'h1b0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9648; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15792 = 12'h1b0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12720; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18864 = 12'h1b0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15792; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21936 = 12'h1b0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18864; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25008 = 12'h1b0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21936; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_432 = io_valid_in ? _GEN_25008 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_432 = 12'h1b0 == _T_2[11:0] ? image_432 : _GEN_431; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3505 = 12'h1b1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6577 = 12'h1b1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3505; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9649 = 12'h1b1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6577; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12721 = 12'h1b1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9649; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15793 = 12'h1b1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12721; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18865 = 12'h1b1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15793; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21937 = 12'h1b1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18865; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25009 = 12'h1b1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21937; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_433 = io_valid_in ? _GEN_25009 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_433 = 12'h1b1 == _T_2[11:0] ? image_433 : _GEN_432; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3506 = 12'h1b2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6578 = 12'h1b2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3506; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9650 = 12'h1b2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6578; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12722 = 12'h1b2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9650; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15794 = 12'h1b2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12722; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18866 = 12'h1b2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15794; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21938 = 12'h1b2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18866; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25010 = 12'h1b2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21938; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_434 = io_valid_in ? _GEN_25010 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_434 = 12'h1b2 == _T_2[11:0] ? image_434 : _GEN_433; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3507 = 12'h1b3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6579 = 12'h1b3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3507; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9651 = 12'h1b3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6579; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12723 = 12'h1b3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9651; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15795 = 12'h1b3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12723; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18867 = 12'h1b3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15795; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21939 = 12'h1b3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18867; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25011 = 12'h1b3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21939; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_435 = io_valid_in ? _GEN_25011 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_435 = 12'h1b3 == _T_2[11:0] ? image_435 : _GEN_434; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3508 = 12'h1b4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6580 = 12'h1b4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3508; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9652 = 12'h1b4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6580; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12724 = 12'h1b4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9652; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15796 = 12'h1b4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12724; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18868 = 12'h1b4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15796; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21940 = 12'h1b4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18868; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25012 = 12'h1b4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21940; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_436 = io_valid_in ? _GEN_25012 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_436 = 12'h1b4 == _T_2[11:0] ? image_436 : _GEN_435; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3509 = 12'h1b5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6581 = 12'h1b5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3509; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9653 = 12'h1b5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6581; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12725 = 12'h1b5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9653; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15797 = 12'h1b5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12725; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18869 = 12'h1b5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15797; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21941 = 12'h1b5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18869; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25013 = 12'h1b5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21941; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_437 = io_valid_in ? _GEN_25013 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_437 = 12'h1b5 == _T_2[11:0] ? image_437 : _GEN_436; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3510 = 12'h1b6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6582 = 12'h1b6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3510; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9654 = 12'h1b6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6582; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12726 = 12'h1b6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9654; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15798 = 12'h1b6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12726; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18870 = 12'h1b6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15798; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21942 = 12'h1b6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18870; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25014 = 12'h1b6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21942; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_438 = io_valid_in ? _GEN_25014 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_438 = 12'h1b6 == _T_2[11:0] ? image_438 : _GEN_437; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3511 = 12'h1b7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6583 = 12'h1b7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3511; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9655 = 12'h1b7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6583; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12727 = 12'h1b7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9655; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15799 = 12'h1b7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12727; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18871 = 12'h1b7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15799; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21943 = 12'h1b7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18871; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25015 = 12'h1b7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21943; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_439 = io_valid_in ? _GEN_25015 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_439 = 12'h1b7 == _T_2[11:0] ? image_439 : _GEN_438; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3512 = 12'h1b8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6584 = 12'h1b8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3512; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9656 = 12'h1b8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6584; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12728 = 12'h1b8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9656; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15800 = 12'h1b8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12728; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18872 = 12'h1b8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15800; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21944 = 12'h1b8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18872; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25016 = 12'h1b8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21944; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_440 = io_valid_in ? _GEN_25016 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_440 = 12'h1b8 == _T_2[11:0] ? image_440 : _GEN_439; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3513 = 12'h1b9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6585 = 12'h1b9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3513; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9657 = 12'h1b9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6585; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12729 = 12'h1b9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9657; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15801 = 12'h1b9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12729; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18873 = 12'h1b9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15801; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21945 = 12'h1b9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18873; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25017 = 12'h1b9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21945; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_441 = io_valid_in ? _GEN_25017 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_441 = 12'h1b9 == _T_2[11:0] ? image_441 : _GEN_440; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3514 = 12'h1ba == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6586 = 12'h1ba == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3514; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9658 = 12'h1ba == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6586; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12730 = 12'h1ba == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9658; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15802 = 12'h1ba == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12730; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18874 = 12'h1ba == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15802; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21946 = 12'h1ba == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18874; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25018 = 12'h1ba == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21946; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_442 = io_valid_in ? _GEN_25018 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_442 = 12'h1ba == _T_2[11:0] ? image_442 : _GEN_441; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3515 = 12'h1bb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6587 = 12'h1bb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3515; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9659 = 12'h1bb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6587; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12731 = 12'h1bb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9659; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15803 = 12'h1bb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12731; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18875 = 12'h1bb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15803; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21947 = 12'h1bb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18875; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25019 = 12'h1bb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21947; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_443 = io_valid_in ? _GEN_25019 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_443 = 12'h1bb == _T_2[11:0] ? image_443 : _GEN_442; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3516 = 12'h1bc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6588 = 12'h1bc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3516; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9660 = 12'h1bc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6588; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12732 = 12'h1bc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9660; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15804 = 12'h1bc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12732; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18876 = 12'h1bc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15804; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21948 = 12'h1bc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18876; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25020 = 12'h1bc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21948; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_444 = io_valid_in ? _GEN_25020 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_444 = 12'h1bc == _T_2[11:0] ? image_444 : _GEN_443; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3517 = 12'h1bd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6589 = 12'h1bd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3517; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9661 = 12'h1bd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6589; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12733 = 12'h1bd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9661; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15805 = 12'h1bd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12733; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18877 = 12'h1bd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15805; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21949 = 12'h1bd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18877; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25021 = 12'h1bd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21949; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_445 = io_valid_in ? _GEN_25021 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_445 = 12'h1bd == _T_2[11:0] ? image_445 : _GEN_444; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3518 = 12'h1be == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6590 = 12'h1be == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3518; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9662 = 12'h1be == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6590; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12734 = 12'h1be == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9662; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15806 = 12'h1be == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12734; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18878 = 12'h1be == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15806; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21950 = 12'h1be == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18878; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25022 = 12'h1be == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21950; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_446 = io_valid_in ? _GEN_25022 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_446 = 12'h1be == _T_2[11:0] ? image_446 : _GEN_445; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3519 = 12'h1bf == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6591 = 12'h1bf == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3519; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9663 = 12'h1bf == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6591; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12735 = 12'h1bf == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9663; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15807 = 12'h1bf == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12735; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18879 = 12'h1bf == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15807; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21951 = 12'h1bf == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18879; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25023 = 12'h1bf == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21951; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_447 = io_valid_in ? _GEN_25023 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_447 = 12'h1bf == _T_2[11:0] ? image_447 : _GEN_446; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3520 = 12'h1c0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6592 = 12'h1c0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3520; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9664 = 12'h1c0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6592; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12736 = 12'h1c0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9664; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15808 = 12'h1c0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12736; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18880 = 12'h1c0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15808; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21952 = 12'h1c0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18880; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25024 = 12'h1c0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21952; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_448 = io_valid_in ? _GEN_25024 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_448 = 12'h1c0 == _T_2[11:0] ? image_448 : _GEN_447; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3521 = 12'h1c1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6593 = 12'h1c1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3521; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9665 = 12'h1c1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6593; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12737 = 12'h1c1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9665; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15809 = 12'h1c1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12737; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18881 = 12'h1c1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15809; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21953 = 12'h1c1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18881; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25025 = 12'h1c1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21953; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_449 = io_valid_in ? _GEN_25025 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_449 = 12'h1c1 == _T_2[11:0] ? image_449 : _GEN_448; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3522 = 12'h1c2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6594 = 12'h1c2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3522; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9666 = 12'h1c2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6594; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12738 = 12'h1c2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9666; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15810 = 12'h1c2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12738; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18882 = 12'h1c2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15810; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21954 = 12'h1c2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18882; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25026 = 12'h1c2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21954; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_450 = io_valid_in ? _GEN_25026 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_450 = 12'h1c2 == _T_2[11:0] ? image_450 : _GEN_449; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3523 = 12'h1c3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6595 = 12'h1c3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3523; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9667 = 12'h1c3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6595; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12739 = 12'h1c3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9667; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15811 = 12'h1c3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12739; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18883 = 12'h1c3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15811; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21955 = 12'h1c3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18883; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25027 = 12'h1c3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21955; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_451 = io_valid_in ? _GEN_25027 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_451 = 12'h1c3 == _T_2[11:0] ? image_451 : _GEN_450; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3524 = 12'h1c4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6596 = 12'h1c4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3524; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9668 = 12'h1c4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6596; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12740 = 12'h1c4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9668; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15812 = 12'h1c4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12740; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18884 = 12'h1c4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15812; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21956 = 12'h1c4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18884; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25028 = 12'h1c4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21956; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_452 = io_valid_in ? _GEN_25028 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_452 = 12'h1c4 == _T_2[11:0] ? image_452 : _GEN_451; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3525 = 12'h1c5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6597 = 12'h1c5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3525; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9669 = 12'h1c5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6597; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12741 = 12'h1c5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9669; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15813 = 12'h1c5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12741; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18885 = 12'h1c5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15813; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21957 = 12'h1c5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18885; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25029 = 12'h1c5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21957; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_453 = io_valid_in ? _GEN_25029 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_453 = 12'h1c5 == _T_2[11:0] ? image_453 : _GEN_452; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3526 = 12'h1c6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6598 = 12'h1c6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3526; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9670 = 12'h1c6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6598; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12742 = 12'h1c6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9670; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15814 = 12'h1c6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12742; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18886 = 12'h1c6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15814; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21958 = 12'h1c6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18886; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25030 = 12'h1c6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21958; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_454 = io_valid_in ? _GEN_25030 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_454 = 12'h1c6 == _T_2[11:0] ? image_454 : _GEN_453; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3527 = 12'h1c7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6599 = 12'h1c7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3527; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9671 = 12'h1c7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6599; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12743 = 12'h1c7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9671; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15815 = 12'h1c7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12743; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18887 = 12'h1c7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15815; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21959 = 12'h1c7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18887; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25031 = 12'h1c7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21959; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_455 = io_valid_in ? _GEN_25031 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_455 = 12'h1c7 == _T_2[11:0] ? image_455 : _GEN_454; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3528 = 12'h1c8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6600 = 12'h1c8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3528; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9672 = 12'h1c8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6600; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12744 = 12'h1c8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9672; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15816 = 12'h1c8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12744; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18888 = 12'h1c8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15816; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21960 = 12'h1c8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18888; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25032 = 12'h1c8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21960; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_456 = io_valid_in ? _GEN_25032 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_456 = 12'h1c8 == _T_2[11:0] ? image_456 : _GEN_455; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3529 = 12'h1c9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6601 = 12'h1c9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3529; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9673 = 12'h1c9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6601; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12745 = 12'h1c9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9673; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15817 = 12'h1c9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12745; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18889 = 12'h1c9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15817; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21961 = 12'h1c9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18889; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25033 = 12'h1c9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21961; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_457 = io_valid_in ? _GEN_25033 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_457 = 12'h1c9 == _T_2[11:0] ? image_457 : _GEN_456; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3530 = 12'h1ca == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6602 = 12'h1ca == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3530; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9674 = 12'h1ca == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6602; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12746 = 12'h1ca == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9674; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15818 = 12'h1ca == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12746; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18890 = 12'h1ca == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15818; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21962 = 12'h1ca == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18890; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25034 = 12'h1ca == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21962; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_458 = io_valid_in ? _GEN_25034 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_458 = 12'h1ca == _T_2[11:0] ? image_458 : _GEN_457; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3531 = 12'h1cb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6603 = 12'h1cb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3531; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9675 = 12'h1cb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6603; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12747 = 12'h1cb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9675; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15819 = 12'h1cb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12747; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18891 = 12'h1cb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15819; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21963 = 12'h1cb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18891; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25035 = 12'h1cb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21963; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_459 = io_valid_in ? _GEN_25035 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_459 = 12'h1cb == _T_2[11:0] ? image_459 : _GEN_458; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3532 = 12'h1cc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6604 = 12'h1cc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3532; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9676 = 12'h1cc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6604; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12748 = 12'h1cc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9676; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15820 = 12'h1cc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12748; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18892 = 12'h1cc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15820; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21964 = 12'h1cc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18892; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25036 = 12'h1cc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21964; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_460 = io_valid_in ? _GEN_25036 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_460 = 12'h1cc == _T_2[11:0] ? image_460 : _GEN_459; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3533 = 12'h1cd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6605 = 12'h1cd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3533; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9677 = 12'h1cd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6605; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12749 = 12'h1cd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9677; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15821 = 12'h1cd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12749; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18893 = 12'h1cd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15821; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21965 = 12'h1cd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18893; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25037 = 12'h1cd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21965; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_461 = io_valid_in ? _GEN_25037 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_461 = 12'h1cd == _T_2[11:0] ? image_461 : _GEN_460; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3534 = 12'h1ce == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6606 = 12'h1ce == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3534; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9678 = 12'h1ce == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6606; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12750 = 12'h1ce == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9678; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15822 = 12'h1ce == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12750; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18894 = 12'h1ce == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15822; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21966 = 12'h1ce == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18894; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25038 = 12'h1ce == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21966; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_462 = io_valid_in ? _GEN_25038 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_462 = 12'h1ce == _T_2[11:0] ? image_462 : _GEN_461; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3535 = 12'h1cf == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6607 = 12'h1cf == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3535; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9679 = 12'h1cf == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6607; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12751 = 12'h1cf == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9679; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15823 = 12'h1cf == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12751; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18895 = 12'h1cf == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15823; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21967 = 12'h1cf == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18895; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25039 = 12'h1cf == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21967; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_463 = io_valid_in ? _GEN_25039 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_463 = 12'h1cf == _T_2[11:0] ? image_463 : _GEN_462; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3536 = 12'h1d0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6608 = 12'h1d0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3536; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9680 = 12'h1d0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6608; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12752 = 12'h1d0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9680; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15824 = 12'h1d0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12752; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18896 = 12'h1d0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15824; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21968 = 12'h1d0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18896; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25040 = 12'h1d0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21968; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_464 = io_valid_in ? _GEN_25040 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_464 = 12'h1d0 == _T_2[11:0] ? image_464 : _GEN_463; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3537 = 12'h1d1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6609 = 12'h1d1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3537; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9681 = 12'h1d1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6609; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12753 = 12'h1d1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9681; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15825 = 12'h1d1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12753; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18897 = 12'h1d1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15825; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21969 = 12'h1d1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18897; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25041 = 12'h1d1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21969; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_465 = io_valid_in ? _GEN_25041 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_465 = 12'h1d1 == _T_2[11:0] ? image_465 : _GEN_464; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3538 = 12'h1d2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6610 = 12'h1d2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3538; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9682 = 12'h1d2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6610; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12754 = 12'h1d2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9682; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15826 = 12'h1d2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12754; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18898 = 12'h1d2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15826; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21970 = 12'h1d2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18898; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25042 = 12'h1d2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21970; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_466 = io_valid_in ? _GEN_25042 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_466 = 12'h1d2 == _T_2[11:0] ? image_466 : _GEN_465; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3539 = 12'h1d3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6611 = 12'h1d3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3539; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9683 = 12'h1d3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6611; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12755 = 12'h1d3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9683; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15827 = 12'h1d3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12755; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18899 = 12'h1d3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15827; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21971 = 12'h1d3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18899; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25043 = 12'h1d3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21971; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_467 = io_valid_in ? _GEN_25043 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_467 = 12'h1d3 == _T_2[11:0] ? image_467 : _GEN_466; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3540 = 12'h1d4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6612 = 12'h1d4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3540; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9684 = 12'h1d4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6612; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12756 = 12'h1d4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9684; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15828 = 12'h1d4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12756; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18900 = 12'h1d4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15828; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21972 = 12'h1d4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18900; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25044 = 12'h1d4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21972; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_468 = io_valid_in ? _GEN_25044 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_468 = 12'h1d4 == _T_2[11:0] ? image_468 : _GEN_467; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3541 = 12'h1d5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6613 = 12'h1d5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3541; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9685 = 12'h1d5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6613; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12757 = 12'h1d5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9685; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15829 = 12'h1d5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12757; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18901 = 12'h1d5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15829; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21973 = 12'h1d5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18901; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25045 = 12'h1d5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21973; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_469 = io_valid_in ? _GEN_25045 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_469 = 12'h1d5 == _T_2[11:0] ? image_469 : _GEN_468; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3542 = 12'h1d6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6614 = 12'h1d6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3542; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9686 = 12'h1d6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6614; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12758 = 12'h1d6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9686; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15830 = 12'h1d6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12758; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18902 = 12'h1d6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15830; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21974 = 12'h1d6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18902; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25046 = 12'h1d6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21974; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_470 = io_valid_in ? _GEN_25046 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_470 = 12'h1d6 == _T_2[11:0] ? image_470 : _GEN_469; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3543 = 12'h1d7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6615 = 12'h1d7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3543; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9687 = 12'h1d7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6615; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12759 = 12'h1d7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9687; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15831 = 12'h1d7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12759; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18903 = 12'h1d7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15831; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21975 = 12'h1d7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18903; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25047 = 12'h1d7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21975; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_471 = io_valid_in ? _GEN_25047 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_471 = 12'h1d7 == _T_2[11:0] ? image_471 : _GEN_470; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3544 = 12'h1d8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6616 = 12'h1d8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3544; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9688 = 12'h1d8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6616; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12760 = 12'h1d8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9688; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15832 = 12'h1d8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12760; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18904 = 12'h1d8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15832; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21976 = 12'h1d8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18904; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25048 = 12'h1d8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21976; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_472 = io_valid_in ? _GEN_25048 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_472 = 12'h1d8 == _T_2[11:0] ? image_472 : _GEN_471; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3545 = 12'h1d9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6617 = 12'h1d9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3545; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9689 = 12'h1d9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6617; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12761 = 12'h1d9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9689; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15833 = 12'h1d9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12761; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18905 = 12'h1d9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15833; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21977 = 12'h1d9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18905; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25049 = 12'h1d9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21977; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_473 = io_valid_in ? _GEN_25049 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_473 = 12'h1d9 == _T_2[11:0] ? image_473 : _GEN_472; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3546 = 12'h1da == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6618 = 12'h1da == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3546; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9690 = 12'h1da == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6618; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12762 = 12'h1da == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9690; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15834 = 12'h1da == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12762; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18906 = 12'h1da == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15834; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21978 = 12'h1da == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18906; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25050 = 12'h1da == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21978; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_474 = io_valid_in ? _GEN_25050 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_474 = 12'h1da == _T_2[11:0] ? image_474 : _GEN_473; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3547 = 12'h1db == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6619 = 12'h1db == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3547; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9691 = 12'h1db == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6619; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12763 = 12'h1db == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9691; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15835 = 12'h1db == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12763; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18907 = 12'h1db == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15835; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21979 = 12'h1db == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18907; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25051 = 12'h1db == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21979; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_475 = io_valid_in ? _GEN_25051 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_475 = 12'h1db == _T_2[11:0] ? image_475 : _GEN_474; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3548 = 12'h1dc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6620 = 12'h1dc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3548; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9692 = 12'h1dc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6620; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12764 = 12'h1dc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9692; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15836 = 12'h1dc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12764; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18908 = 12'h1dc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15836; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21980 = 12'h1dc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18908; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25052 = 12'h1dc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21980; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_476 = io_valid_in ? _GEN_25052 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_476 = 12'h1dc == _T_2[11:0] ? image_476 : _GEN_475; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3549 = 12'h1dd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6621 = 12'h1dd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3549; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9693 = 12'h1dd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6621; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12765 = 12'h1dd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9693; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15837 = 12'h1dd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12765; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18909 = 12'h1dd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15837; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21981 = 12'h1dd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18909; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25053 = 12'h1dd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21981; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_477 = io_valid_in ? _GEN_25053 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_477 = 12'h1dd == _T_2[11:0] ? image_477 : _GEN_476; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3550 = 12'h1de == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6622 = 12'h1de == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3550; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9694 = 12'h1de == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6622; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12766 = 12'h1de == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9694; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15838 = 12'h1de == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12766; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18910 = 12'h1de == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15838; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21982 = 12'h1de == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18910; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25054 = 12'h1de == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21982; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_478 = io_valid_in ? _GEN_25054 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_478 = 12'h1de == _T_2[11:0] ? image_478 : _GEN_477; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3551 = 12'h1df == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6623 = 12'h1df == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3551; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9695 = 12'h1df == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6623; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12767 = 12'h1df == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9695; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15839 = 12'h1df == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12767; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18911 = 12'h1df == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15839; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21983 = 12'h1df == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18911; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25055 = 12'h1df == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21983; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_479 = io_valid_in ? _GEN_25055 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_479 = 12'h1df == _T_2[11:0] ? image_479 : _GEN_478; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3552 = 12'h1e0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6624 = 12'h1e0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3552; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9696 = 12'h1e0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6624; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12768 = 12'h1e0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9696; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15840 = 12'h1e0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12768; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18912 = 12'h1e0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15840; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21984 = 12'h1e0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18912; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25056 = 12'h1e0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21984; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_480 = io_valid_in ? _GEN_25056 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_480 = 12'h1e0 == _T_2[11:0] ? image_480 : _GEN_479; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3553 = 12'h1e1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6625 = 12'h1e1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3553; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9697 = 12'h1e1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6625; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12769 = 12'h1e1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9697; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15841 = 12'h1e1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12769; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18913 = 12'h1e1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15841; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21985 = 12'h1e1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18913; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25057 = 12'h1e1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21985; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_481 = io_valid_in ? _GEN_25057 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_481 = 12'h1e1 == _T_2[11:0] ? image_481 : _GEN_480; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3554 = 12'h1e2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6626 = 12'h1e2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3554; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9698 = 12'h1e2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6626; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12770 = 12'h1e2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9698; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15842 = 12'h1e2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12770; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18914 = 12'h1e2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15842; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21986 = 12'h1e2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18914; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25058 = 12'h1e2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21986; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_482 = io_valid_in ? _GEN_25058 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_482 = 12'h1e2 == _T_2[11:0] ? image_482 : _GEN_481; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3555 = 12'h1e3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6627 = 12'h1e3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3555; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9699 = 12'h1e3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6627; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12771 = 12'h1e3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9699; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15843 = 12'h1e3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12771; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18915 = 12'h1e3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15843; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21987 = 12'h1e3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18915; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25059 = 12'h1e3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21987; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_483 = io_valid_in ? _GEN_25059 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_483 = 12'h1e3 == _T_2[11:0] ? image_483 : _GEN_482; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3556 = 12'h1e4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6628 = 12'h1e4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3556; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9700 = 12'h1e4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6628; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12772 = 12'h1e4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9700; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15844 = 12'h1e4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12772; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18916 = 12'h1e4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15844; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21988 = 12'h1e4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18916; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25060 = 12'h1e4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21988; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_484 = io_valid_in ? _GEN_25060 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_484 = 12'h1e4 == _T_2[11:0] ? image_484 : _GEN_483; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3557 = 12'h1e5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6629 = 12'h1e5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3557; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9701 = 12'h1e5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6629; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12773 = 12'h1e5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9701; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15845 = 12'h1e5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12773; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18917 = 12'h1e5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15845; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21989 = 12'h1e5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18917; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25061 = 12'h1e5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21989; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_485 = io_valid_in ? _GEN_25061 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_485 = 12'h1e5 == _T_2[11:0] ? image_485 : _GEN_484; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3558 = 12'h1e6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6630 = 12'h1e6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3558; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9702 = 12'h1e6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6630; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12774 = 12'h1e6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9702; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15846 = 12'h1e6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12774; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18918 = 12'h1e6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15846; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21990 = 12'h1e6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18918; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25062 = 12'h1e6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21990; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_486 = io_valid_in ? _GEN_25062 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_486 = 12'h1e6 == _T_2[11:0] ? image_486 : _GEN_485; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3559 = 12'h1e7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6631 = 12'h1e7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3559; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9703 = 12'h1e7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6631; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12775 = 12'h1e7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9703; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15847 = 12'h1e7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12775; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18919 = 12'h1e7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15847; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21991 = 12'h1e7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18919; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25063 = 12'h1e7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21991; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_487 = io_valid_in ? _GEN_25063 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_487 = 12'h1e7 == _T_2[11:0] ? image_487 : _GEN_486; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3560 = 12'h1e8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6632 = 12'h1e8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3560; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9704 = 12'h1e8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6632; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12776 = 12'h1e8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9704; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15848 = 12'h1e8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12776; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18920 = 12'h1e8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15848; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21992 = 12'h1e8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18920; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25064 = 12'h1e8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21992; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_488 = io_valid_in ? _GEN_25064 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_488 = 12'h1e8 == _T_2[11:0] ? image_488 : _GEN_487; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3561 = 12'h1e9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6633 = 12'h1e9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3561; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9705 = 12'h1e9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6633; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12777 = 12'h1e9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9705; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15849 = 12'h1e9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12777; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18921 = 12'h1e9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15849; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21993 = 12'h1e9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18921; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25065 = 12'h1e9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21993; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_489 = io_valid_in ? _GEN_25065 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_489 = 12'h1e9 == _T_2[11:0] ? image_489 : _GEN_488; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3562 = 12'h1ea == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6634 = 12'h1ea == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3562; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9706 = 12'h1ea == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6634; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12778 = 12'h1ea == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9706; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15850 = 12'h1ea == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12778; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18922 = 12'h1ea == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15850; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21994 = 12'h1ea == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18922; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25066 = 12'h1ea == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21994; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_490 = io_valid_in ? _GEN_25066 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_490 = 12'h1ea == _T_2[11:0] ? image_490 : _GEN_489; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3563 = 12'h1eb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6635 = 12'h1eb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3563; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9707 = 12'h1eb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6635; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12779 = 12'h1eb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9707; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15851 = 12'h1eb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12779; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18923 = 12'h1eb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15851; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21995 = 12'h1eb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18923; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25067 = 12'h1eb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21995; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_491 = io_valid_in ? _GEN_25067 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_491 = 12'h1eb == _T_2[11:0] ? image_491 : _GEN_490; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3564 = 12'h1ec == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6636 = 12'h1ec == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3564; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9708 = 12'h1ec == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6636; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12780 = 12'h1ec == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9708; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15852 = 12'h1ec == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12780; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18924 = 12'h1ec == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15852; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21996 = 12'h1ec == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18924; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25068 = 12'h1ec == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21996; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_492 = io_valid_in ? _GEN_25068 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_492 = 12'h1ec == _T_2[11:0] ? image_492 : _GEN_491; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3565 = 12'h1ed == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6637 = 12'h1ed == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3565; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9709 = 12'h1ed == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6637; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12781 = 12'h1ed == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9709; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15853 = 12'h1ed == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12781; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18925 = 12'h1ed == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15853; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21997 = 12'h1ed == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18925; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25069 = 12'h1ed == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21997; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_493 = io_valid_in ? _GEN_25069 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_493 = 12'h1ed == _T_2[11:0] ? image_493 : _GEN_492; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3566 = 12'h1ee == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6638 = 12'h1ee == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3566; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9710 = 12'h1ee == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6638; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12782 = 12'h1ee == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9710; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15854 = 12'h1ee == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12782; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18926 = 12'h1ee == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15854; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21998 = 12'h1ee == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18926; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25070 = 12'h1ee == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21998; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_494 = io_valid_in ? _GEN_25070 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_494 = 12'h1ee == _T_2[11:0] ? image_494 : _GEN_493; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3567 = 12'h1ef == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6639 = 12'h1ef == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3567; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9711 = 12'h1ef == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6639; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12783 = 12'h1ef == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9711; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15855 = 12'h1ef == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12783; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18927 = 12'h1ef == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15855; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21999 = 12'h1ef == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18927; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25071 = 12'h1ef == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_21999; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_495 = io_valid_in ? _GEN_25071 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_495 = 12'h1ef == _T_2[11:0] ? image_495 : _GEN_494; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3568 = 12'h1f0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6640 = 12'h1f0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3568; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9712 = 12'h1f0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6640; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12784 = 12'h1f0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9712; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15856 = 12'h1f0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12784; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18928 = 12'h1f0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15856; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22000 = 12'h1f0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18928; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25072 = 12'h1f0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22000; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_496 = io_valid_in ? _GEN_25072 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_496 = 12'h1f0 == _T_2[11:0] ? image_496 : _GEN_495; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3569 = 12'h1f1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6641 = 12'h1f1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3569; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9713 = 12'h1f1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6641; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12785 = 12'h1f1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9713; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15857 = 12'h1f1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12785; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18929 = 12'h1f1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15857; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22001 = 12'h1f1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18929; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25073 = 12'h1f1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22001; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_497 = io_valid_in ? _GEN_25073 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_497 = 12'h1f1 == _T_2[11:0] ? image_497 : _GEN_496; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3570 = 12'h1f2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6642 = 12'h1f2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3570; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9714 = 12'h1f2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6642; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12786 = 12'h1f2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9714; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15858 = 12'h1f2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12786; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18930 = 12'h1f2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15858; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22002 = 12'h1f2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18930; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25074 = 12'h1f2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22002; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_498 = io_valid_in ? _GEN_25074 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_498 = 12'h1f2 == _T_2[11:0] ? image_498 : _GEN_497; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3571 = 12'h1f3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6643 = 12'h1f3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3571; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9715 = 12'h1f3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6643; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12787 = 12'h1f3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9715; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15859 = 12'h1f3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12787; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18931 = 12'h1f3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15859; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22003 = 12'h1f3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18931; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25075 = 12'h1f3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22003; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_499 = io_valid_in ? _GEN_25075 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_499 = 12'h1f3 == _T_2[11:0] ? image_499 : _GEN_498; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3572 = 12'h1f4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6644 = 12'h1f4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3572; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9716 = 12'h1f4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6644; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12788 = 12'h1f4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9716; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15860 = 12'h1f4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12788; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18932 = 12'h1f4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15860; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22004 = 12'h1f4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18932; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25076 = 12'h1f4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22004; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_500 = io_valid_in ? _GEN_25076 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_500 = 12'h1f4 == _T_2[11:0] ? image_500 : _GEN_499; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3573 = 12'h1f5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6645 = 12'h1f5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3573; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9717 = 12'h1f5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6645; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12789 = 12'h1f5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9717; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15861 = 12'h1f5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12789; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18933 = 12'h1f5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15861; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22005 = 12'h1f5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18933; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25077 = 12'h1f5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22005; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_501 = io_valid_in ? _GEN_25077 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_501 = 12'h1f5 == _T_2[11:0] ? image_501 : _GEN_500; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3574 = 12'h1f6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6646 = 12'h1f6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3574; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9718 = 12'h1f6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6646; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12790 = 12'h1f6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9718; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15862 = 12'h1f6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12790; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18934 = 12'h1f6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15862; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22006 = 12'h1f6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18934; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25078 = 12'h1f6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22006; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_502 = io_valid_in ? _GEN_25078 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_502 = 12'h1f6 == _T_2[11:0] ? image_502 : _GEN_501; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3575 = 12'h1f7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6647 = 12'h1f7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3575; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9719 = 12'h1f7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6647; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12791 = 12'h1f7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9719; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15863 = 12'h1f7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12791; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18935 = 12'h1f7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15863; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22007 = 12'h1f7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18935; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25079 = 12'h1f7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22007; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_503 = io_valid_in ? _GEN_25079 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_503 = 12'h1f7 == _T_2[11:0] ? image_503 : _GEN_502; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3576 = 12'h1f8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6648 = 12'h1f8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3576; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9720 = 12'h1f8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6648; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12792 = 12'h1f8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9720; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15864 = 12'h1f8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12792; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18936 = 12'h1f8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15864; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22008 = 12'h1f8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18936; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25080 = 12'h1f8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22008; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_504 = io_valid_in ? _GEN_25080 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_504 = 12'h1f8 == _T_2[11:0] ? image_504 : _GEN_503; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3577 = 12'h1f9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6649 = 12'h1f9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3577; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9721 = 12'h1f9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6649; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12793 = 12'h1f9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9721; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15865 = 12'h1f9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12793; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18937 = 12'h1f9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15865; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22009 = 12'h1f9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18937; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25081 = 12'h1f9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22009; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_505 = io_valid_in ? _GEN_25081 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_505 = 12'h1f9 == _T_2[11:0] ? image_505 : _GEN_504; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3578 = 12'h1fa == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6650 = 12'h1fa == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3578; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9722 = 12'h1fa == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6650; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12794 = 12'h1fa == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9722; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15866 = 12'h1fa == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12794; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18938 = 12'h1fa == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15866; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22010 = 12'h1fa == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18938; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25082 = 12'h1fa == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22010; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_506 = io_valid_in ? _GEN_25082 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_506 = 12'h1fa == _T_2[11:0] ? image_506 : _GEN_505; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3579 = 12'h1fb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6651 = 12'h1fb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3579; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9723 = 12'h1fb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6651; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12795 = 12'h1fb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9723; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15867 = 12'h1fb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12795; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18939 = 12'h1fb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15867; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22011 = 12'h1fb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18939; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25083 = 12'h1fb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22011; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_507 = io_valid_in ? _GEN_25083 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_507 = 12'h1fb == _T_2[11:0] ? image_507 : _GEN_506; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3580 = 12'h1fc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6652 = 12'h1fc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3580; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9724 = 12'h1fc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6652; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12796 = 12'h1fc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9724; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15868 = 12'h1fc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12796; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18940 = 12'h1fc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15868; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22012 = 12'h1fc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18940; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25084 = 12'h1fc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22012; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_508 = io_valid_in ? _GEN_25084 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_508 = 12'h1fc == _T_2[11:0] ? image_508 : _GEN_507; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3581 = 12'h1fd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6653 = 12'h1fd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3581; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9725 = 12'h1fd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6653; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12797 = 12'h1fd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9725; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15869 = 12'h1fd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12797; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18941 = 12'h1fd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15869; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22013 = 12'h1fd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18941; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25085 = 12'h1fd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22013; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_509 = io_valid_in ? _GEN_25085 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_509 = 12'h1fd == _T_2[11:0] ? image_509 : _GEN_508; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3582 = 12'h1fe == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6654 = 12'h1fe == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3582; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9726 = 12'h1fe == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6654; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12798 = 12'h1fe == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9726; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15870 = 12'h1fe == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12798; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18942 = 12'h1fe == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15870; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22014 = 12'h1fe == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18942; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25086 = 12'h1fe == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22014; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_510 = io_valid_in ? _GEN_25086 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_510 = 12'h1fe == _T_2[11:0] ? image_510 : _GEN_509; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3583 = 12'h1ff == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6655 = 12'h1ff == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3583; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9727 = 12'h1ff == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6655; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12799 = 12'h1ff == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9727; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15871 = 12'h1ff == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12799; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18943 = 12'h1ff == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15871; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22015 = 12'h1ff == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18943; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25087 = 12'h1ff == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22015; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_511 = io_valid_in ? _GEN_25087 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_511 = 12'h1ff == _T_2[11:0] ? image_511 : _GEN_510; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3584 = 12'h200 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6656 = 12'h200 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3584; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9728 = 12'h200 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6656; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12800 = 12'h200 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9728; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15872 = 12'h200 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12800; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18944 = 12'h200 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15872; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22016 = 12'h200 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18944; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25088 = 12'h200 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22016; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_512 = io_valid_in ? _GEN_25088 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_512 = 12'h200 == _T_2[11:0] ? image_512 : _GEN_511; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3585 = 12'h201 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6657 = 12'h201 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3585; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9729 = 12'h201 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6657; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12801 = 12'h201 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9729; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15873 = 12'h201 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12801; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18945 = 12'h201 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15873; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22017 = 12'h201 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18945; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25089 = 12'h201 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22017; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_513 = io_valid_in ? _GEN_25089 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_513 = 12'h201 == _T_2[11:0] ? image_513 : _GEN_512; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3586 = 12'h202 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6658 = 12'h202 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3586; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9730 = 12'h202 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6658; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12802 = 12'h202 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9730; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15874 = 12'h202 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12802; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18946 = 12'h202 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15874; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22018 = 12'h202 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18946; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25090 = 12'h202 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22018; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_514 = io_valid_in ? _GEN_25090 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_514 = 12'h202 == _T_2[11:0] ? image_514 : _GEN_513; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3587 = 12'h203 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6659 = 12'h203 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3587; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9731 = 12'h203 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6659; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12803 = 12'h203 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9731; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15875 = 12'h203 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12803; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18947 = 12'h203 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15875; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22019 = 12'h203 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18947; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25091 = 12'h203 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22019; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_515 = io_valid_in ? _GEN_25091 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_515 = 12'h203 == _T_2[11:0] ? image_515 : _GEN_514; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3588 = 12'h204 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6660 = 12'h204 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3588; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9732 = 12'h204 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6660; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12804 = 12'h204 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9732; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15876 = 12'h204 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12804; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18948 = 12'h204 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15876; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22020 = 12'h204 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18948; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25092 = 12'h204 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22020; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_516 = io_valid_in ? _GEN_25092 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_516 = 12'h204 == _T_2[11:0] ? image_516 : _GEN_515; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3589 = 12'h205 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6661 = 12'h205 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3589; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9733 = 12'h205 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6661; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12805 = 12'h205 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9733; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15877 = 12'h205 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12805; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18949 = 12'h205 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15877; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22021 = 12'h205 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18949; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25093 = 12'h205 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22021; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_517 = io_valid_in ? _GEN_25093 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_517 = 12'h205 == _T_2[11:0] ? image_517 : _GEN_516; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3590 = 12'h206 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6662 = 12'h206 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3590; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9734 = 12'h206 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6662; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12806 = 12'h206 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9734; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15878 = 12'h206 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12806; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18950 = 12'h206 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15878; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22022 = 12'h206 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18950; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25094 = 12'h206 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22022; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_518 = io_valid_in ? _GEN_25094 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_518 = 12'h206 == _T_2[11:0] ? image_518 : _GEN_517; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3591 = 12'h207 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6663 = 12'h207 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3591; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9735 = 12'h207 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6663; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12807 = 12'h207 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9735; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15879 = 12'h207 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12807; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18951 = 12'h207 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15879; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22023 = 12'h207 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18951; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25095 = 12'h207 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22023; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_519 = io_valid_in ? _GEN_25095 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_519 = 12'h207 == _T_2[11:0] ? image_519 : _GEN_518; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3592 = 12'h208 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6664 = 12'h208 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3592; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9736 = 12'h208 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6664; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12808 = 12'h208 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9736; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15880 = 12'h208 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12808; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18952 = 12'h208 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15880; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22024 = 12'h208 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18952; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25096 = 12'h208 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22024; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_520 = io_valid_in ? _GEN_25096 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_520 = 12'h208 == _T_2[11:0] ? image_520 : _GEN_519; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3593 = 12'h209 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6665 = 12'h209 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3593; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9737 = 12'h209 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6665; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12809 = 12'h209 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9737; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15881 = 12'h209 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12809; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18953 = 12'h209 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15881; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22025 = 12'h209 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18953; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25097 = 12'h209 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22025; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_521 = io_valid_in ? _GEN_25097 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_521 = 12'h209 == _T_2[11:0] ? image_521 : _GEN_520; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3594 = 12'h20a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6666 = 12'h20a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3594; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9738 = 12'h20a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6666; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12810 = 12'h20a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9738; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15882 = 12'h20a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12810; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18954 = 12'h20a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15882; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22026 = 12'h20a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18954; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25098 = 12'h20a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22026; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_522 = io_valid_in ? _GEN_25098 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_522 = 12'h20a == _T_2[11:0] ? image_522 : _GEN_521; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3595 = 12'h20b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6667 = 12'h20b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3595; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9739 = 12'h20b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6667; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12811 = 12'h20b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9739; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15883 = 12'h20b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12811; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18955 = 12'h20b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15883; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22027 = 12'h20b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18955; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25099 = 12'h20b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22027; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_523 = io_valid_in ? _GEN_25099 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_523 = 12'h20b == _T_2[11:0] ? image_523 : _GEN_522; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3596 = 12'h20c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6668 = 12'h20c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3596; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9740 = 12'h20c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6668; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12812 = 12'h20c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9740; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15884 = 12'h20c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12812; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18956 = 12'h20c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15884; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22028 = 12'h20c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18956; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25100 = 12'h20c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22028; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_524 = io_valid_in ? _GEN_25100 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_524 = 12'h20c == _T_2[11:0] ? image_524 : _GEN_523; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3597 = 12'h20d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6669 = 12'h20d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3597; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9741 = 12'h20d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6669; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12813 = 12'h20d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9741; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15885 = 12'h20d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12813; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18957 = 12'h20d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15885; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22029 = 12'h20d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18957; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25101 = 12'h20d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22029; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_525 = io_valid_in ? _GEN_25101 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_525 = 12'h20d == _T_2[11:0] ? image_525 : _GEN_524; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3598 = 12'h20e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6670 = 12'h20e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3598; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9742 = 12'h20e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6670; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12814 = 12'h20e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9742; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15886 = 12'h20e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12814; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18958 = 12'h20e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15886; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22030 = 12'h20e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18958; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25102 = 12'h20e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22030; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_526 = io_valid_in ? _GEN_25102 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_526 = 12'h20e == _T_2[11:0] ? image_526 : _GEN_525; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3599 = 12'h20f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6671 = 12'h20f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3599; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9743 = 12'h20f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6671; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12815 = 12'h20f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9743; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15887 = 12'h20f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12815; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18959 = 12'h20f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15887; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22031 = 12'h20f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18959; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25103 = 12'h20f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22031; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_527 = io_valid_in ? _GEN_25103 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_527 = 12'h20f == _T_2[11:0] ? image_527 : _GEN_526; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3600 = 12'h210 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6672 = 12'h210 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3600; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9744 = 12'h210 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6672; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12816 = 12'h210 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9744; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15888 = 12'h210 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12816; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18960 = 12'h210 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15888; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22032 = 12'h210 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18960; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25104 = 12'h210 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22032; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_528 = io_valid_in ? _GEN_25104 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_528 = 12'h210 == _T_2[11:0] ? image_528 : _GEN_527; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3601 = 12'h211 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6673 = 12'h211 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3601; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9745 = 12'h211 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6673; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12817 = 12'h211 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9745; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15889 = 12'h211 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12817; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18961 = 12'h211 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15889; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22033 = 12'h211 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18961; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25105 = 12'h211 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22033; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_529 = io_valid_in ? _GEN_25105 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_529 = 12'h211 == _T_2[11:0] ? image_529 : _GEN_528; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3602 = 12'h212 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6674 = 12'h212 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3602; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9746 = 12'h212 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6674; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12818 = 12'h212 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9746; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15890 = 12'h212 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12818; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18962 = 12'h212 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15890; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22034 = 12'h212 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18962; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25106 = 12'h212 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22034; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_530 = io_valid_in ? _GEN_25106 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_530 = 12'h212 == _T_2[11:0] ? image_530 : _GEN_529; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3603 = 12'h213 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6675 = 12'h213 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3603; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9747 = 12'h213 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6675; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12819 = 12'h213 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9747; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15891 = 12'h213 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12819; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18963 = 12'h213 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15891; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22035 = 12'h213 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18963; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25107 = 12'h213 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22035; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_531 = io_valid_in ? _GEN_25107 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_531 = 12'h213 == _T_2[11:0] ? image_531 : _GEN_530; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3604 = 12'h214 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6676 = 12'h214 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3604; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9748 = 12'h214 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6676; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12820 = 12'h214 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9748; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15892 = 12'h214 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12820; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18964 = 12'h214 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15892; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22036 = 12'h214 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18964; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25108 = 12'h214 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22036; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_532 = io_valid_in ? _GEN_25108 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_532 = 12'h214 == _T_2[11:0] ? image_532 : _GEN_531; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3605 = 12'h215 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6677 = 12'h215 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3605; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9749 = 12'h215 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6677; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12821 = 12'h215 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9749; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15893 = 12'h215 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12821; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18965 = 12'h215 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15893; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22037 = 12'h215 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18965; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25109 = 12'h215 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22037; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_533 = io_valid_in ? _GEN_25109 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_533 = 12'h215 == _T_2[11:0] ? image_533 : _GEN_532; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3606 = 12'h216 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6678 = 12'h216 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3606; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9750 = 12'h216 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6678; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12822 = 12'h216 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9750; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15894 = 12'h216 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12822; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18966 = 12'h216 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15894; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22038 = 12'h216 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18966; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25110 = 12'h216 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22038; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_534 = io_valid_in ? _GEN_25110 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_534 = 12'h216 == _T_2[11:0] ? image_534 : _GEN_533; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3607 = 12'h217 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6679 = 12'h217 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3607; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9751 = 12'h217 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6679; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12823 = 12'h217 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9751; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15895 = 12'h217 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12823; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18967 = 12'h217 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15895; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22039 = 12'h217 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18967; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25111 = 12'h217 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22039; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_535 = io_valid_in ? _GEN_25111 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_535 = 12'h217 == _T_2[11:0] ? image_535 : _GEN_534; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3608 = 12'h218 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6680 = 12'h218 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3608; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9752 = 12'h218 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6680; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12824 = 12'h218 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9752; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15896 = 12'h218 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12824; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18968 = 12'h218 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15896; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22040 = 12'h218 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18968; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25112 = 12'h218 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22040; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_536 = io_valid_in ? _GEN_25112 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_536 = 12'h218 == _T_2[11:0] ? image_536 : _GEN_535; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3609 = 12'h219 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6681 = 12'h219 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3609; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9753 = 12'h219 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6681; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12825 = 12'h219 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9753; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15897 = 12'h219 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12825; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18969 = 12'h219 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15897; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22041 = 12'h219 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18969; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25113 = 12'h219 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22041; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_537 = io_valid_in ? _GEN_25113 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_537 = 12'h219 == _T_2[11:0] ? image_537 : _GEN_536; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3610 = 12'h21a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6682 = 12'h21a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3610; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9754 = 12'h21a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6682; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12826 = 12'h21a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9754; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15898 = 12'h21a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12826; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18970 = 12'h21a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15898; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22042 = 12'h21a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18970; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25114 = 12'h21a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22042; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_538 = io_valid_in ? _GEN_25114 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_538 = 12'h21a == _T_2[11:0] ? image_538 : _GEN_537; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3611 = 12'h21b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6683 = 12'h21b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3611; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9755 = 12'h21b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6683; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12827 = 12'h21b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9755; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15899 = 12'h21b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12827; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18971 = 12'h21b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15899; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22043 = 12'h21b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18971; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25115 = 12'h21b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22043; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_539 = io_valid_in ? _GEN_25115 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_539 = 12'h21b == _T_2[11:0] ? image_539 : _GEN_538; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3612 = 12'h21c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6684 = 12'h21c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3612; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9756 = 12'h21c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6684; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12828 = 12'h21c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9756; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15900 = 12'h21c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12828; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18972 = 12'h21c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15900; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22044 = 12'h21c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18972; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25116 = 12'h21c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22044; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_540 = io_valid_in ? _GEN_25116 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_540 = 12'h21c == _T_2[11:0] ? image_540 : _GEN_539; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3613 = 12'h21d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6685 = 12'h21d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3613; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9757 = 12'h21d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6685; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12829 = 12'h21d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9757; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15901 = 12'h21d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12829; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18973 = 12'h21d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15901; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22045 = 12'h21d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18973; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25117 = 12'h21d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22045; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_541 = io_valid_in ? _GEN_25117 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_541 = 12'h21d == _T_2[11:0] ? image_541 : _GEN_540; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3614 = 12'h21e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6686 = 12'h21e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3614; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9758 = 12'h21e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6686; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12830 = 12'h21e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9758; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15902 = 12'h21e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12830; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18974 = 12'h21e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15902; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22046 = 12'h21e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18974; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25118 = 12'h21e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22046; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_542 = io_valid_in ? _GEN_25118 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_542 = 12'h21e == _T_2[11:0] ? image_542 : _GEN_541; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3615 = 12'h21f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6687 = 12'h21f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3615; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9759 = 12'h21f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6687; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12831 = 12'h21f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9759; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15903 = 12'h21f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12831; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18975 = 12'h21f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15903; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22047 = 12'h21f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18975; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25119 = 12'h21f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22047; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_543 = io_valid_in ? _GEN_25119 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_543 = 12'h21f == _T_2[11:0] ? image_543 : _GEN_542; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3616 = 12'h220 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6688 = 12'h220 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3616; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9760 = 12'h220 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6688; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12832 = 12'h220 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9760; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15904 = 12'h220 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12832; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18976 = 12'h220 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15904; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22048 = 12'h220 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18976; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25120 = 12'h220 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22048; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_544 = io_valid_in ? _GEN_25120 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_544 = 12'h220 == _T_2[11:0] ? image_544 : _GEN_543; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3617 = 12'h221 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6689 = 12'h221 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3617; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9761 = 12'h221 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6689; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12833 = 12'h221 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9761; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15905 = 12'h221 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12833; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18977 = 12'h221 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15905; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22049 = 12'h221 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18977; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25121 = 12'h221 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22049; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_545 = io_valid_in ? _GEN_25121 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_545 = 12'h221 == _T_2[11:0] ? image_545 : _GEN_544; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3618 = 12'h222 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6690 = 12'h222 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3618; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9762 = 12'h222 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6690; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12834 = 12'h222 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9762; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15906 = 12'h222 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12834; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18978 = 12'h222 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15906; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22050 = 12'h222 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18978; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25122 = 12'h222 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22050; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_546 = io_valid_in ? _GEN_25122 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_546 = 12'h222 == _T_2[11:0] ? image_546 : _GEN_545; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3619 = 12'h223 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6691 = 12'h223 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3619; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9763 = 12'h223 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6691; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12835 = 12'h223 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9763; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15907 = 12'h223 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12835; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18979 = 12'h223 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15907; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22051 = 12'h223 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18979; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25123 = 12'h223 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22051; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_547 = io_valid_in ? _GEN_25123 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_547 = 12'h223 == _T_2[11:0] ? image_547 : _GEN_546; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3620 = 12'h224 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6692 = 12'h224 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3620; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9764 = 12'h224 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6692; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12836 = 12'h224 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9764; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15908 = 12'h224 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12836; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18980 = 12'h224 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15908; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22052 = 12'h224 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18980; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25124 = 12'h224 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22052; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_548 = io_valid_in ? _GEN_25124 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_548 = 12'h224 == _T_2[11:0] ? image_548 : _GEN_547; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3621 = 12'h225 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6693 = 12'h225 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3621; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9765 = 12'h225 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6693; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12837 = 12'h225 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9765; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15909 = 12'h225 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12837; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18981 = 12'h225 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15909; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22053 = 12'h225 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18981; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25125 = 12'h225 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22053; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_549 = io_valid_in ? _GEN_25125 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_549 = 12'h225 == _T_2[11:0] ? image_549 : _GEN_548; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3622 = 12'h226 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6694 = 12'h226 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3622; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9766 = 12'h226 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6694; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12838 = 12'h226 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9766; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15910 = 12'h226 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12838; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18982 = 12'h226 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15910; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22054 = 12'h226 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18982; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25126 = 12'h226 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22054; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_550 = io_valid_in ? _GEN_25126 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_550 = 12'h226 == _T_2[11:0] ? image_550 : _GEN_549; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3623 = 12'h227 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6695 = 12'h227 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3623; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9767 = 12'h227 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6695; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12839 = 12'h227 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9767; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15911 = 12'h227 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12839; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18983 = 12'h227 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15911; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22055 = 12'h227 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18983; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25127 = 12'h227 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22055; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_551 = io_valid_in ? _GEN_25127 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_551 = 12'h227 == _T_2[11:0] ? image_551 : _GEN_550; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3624 = 12'h228 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6696 = 12'h228 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3624; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9768 = 12'h228 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6696; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12840 = 12'h228 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9768; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15912 = 12'h228 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12840; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18984 = 12'h228 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15912; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22056 = 12'h228 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18984; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25128 = 12'h228 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22056; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_552 = io_valid_in ? _GEN_25128 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_552 = 12'h228 == _T_2[11:0] ? image_552 : _GEN_551; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3625 = 12'h229 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6697 = 12'h229 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3625; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9769 = 12'h229 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6697; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12841 = 12'h229 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9769; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15913 = 12'h229 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12841; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18985 = 12'h229 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15913; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22057 = 12'h229 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18985; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25129 = 12'h229 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22057; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_553 = io_valid_in ? _GEN_25129 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_553 = 12'h229 == _T_2[11:0] ? image_553 : _GEN_552; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3626 = 12'h22a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6698 = 12'h22a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3626; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9770 = 12'h22a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6698; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12842 = 12'h22a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9770; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15914 = 12'h22a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12842; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18986 = 12'h22a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15914; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22058 = 12'h22a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18986; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25130 = 12'h22a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22058; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_554 = io_valid_in ? _GEN_25130 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_554 = 12'h22a == _T_2[11:0] ? image_554 : _GEN_553; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3627 = 12'h22b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6699 = 12'h22b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3627; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9771 = 12'h22b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6699; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12843 = 12'h22b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9771; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15915 = 12'h22b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12843; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18987 = 12'h22b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15915; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22059 = 12'h22b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18987; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25131 = 12'h22b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22059; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_555 = io_valid_in ? _GEN_25131 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_555 = 12'h22b == _T_2[11:0] ? image_555 : _GEN_554; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3628 = 12'h22c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6700 = 12'h22c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3628; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9772 = 12'h22c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6700; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12844 = 12'h22c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9772; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15916 = 12'h22c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12844; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18988 = 12'h22c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15916; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22060 = 12'h22c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18988; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25132 = 12'h22c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22060; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_556 = io_valid_in ? _GEN_25132 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_556 = 12'h22c == _T_2[11:0] ? image_556 : _GEN_555; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3629 = 12'h22d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6701 = 12'h22d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3629; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9773 = 12'h22d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6701; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12845 = 12'h22d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9773; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15917 = 12'h22d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12845; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18989 = 12'h22d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15917; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22061 = 12'h22d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18989; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25133 = 12'h22d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22061; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_557 = io_valid_in ? _GEN_25133 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_557 = 12'h22d == _T_2[11:0] ? image_557 : _GEN_556; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3630 = 12'h22e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6702 = 12'h22e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3630; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9774 = 12'h22e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6702; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12846 = 12'h22e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9774; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15918 = 12'h22e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12846; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18990 = 12'h22e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15918; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22062 = 12'h22e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18990; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25134 = 12'h22e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22062; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_558 = io_valid_in ? _GEN_25134 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_558 = 12'h22e == _T_2[11:0] ? image_558 : _GEN_557; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3631 = 12'h22f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6703 = 12'h22f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3631; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9775 = 12'h22f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6703; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12847 = 12'h22f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9775; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15919 = 12'h22f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12847; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18991 = 12'h22f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15919; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22063 = 12'h22f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18991; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25135 = 12'h22f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22063; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_559 = io_valid_in ? _GEN_25135 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_559 = 12'h22f == _T_2[11:0] ? image_559 : _GEN_558; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3632 = 12'h230 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6704 = 12'h230 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3632; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9776 = 12'h230 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6704; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12848 = 12'h230 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9776; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15920 = 12'h230 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12848; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18992 = 12'h230 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15920; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22064 = 12'h230 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18992; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25136 = 12'h230 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22064; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_560 = io_valid_in ? _GEN_25136 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_560 = 12'h230 == _T_2[11:0] ? image_560 : _GEN_559; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3633 = 12'h231 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6705 = 12'h231 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3633; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9777 = 12'h231 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6705; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12849 = 12'h231 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9777; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15921 = 12'h231 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12849; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18993 = 12'h231 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15921; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22065 = 12'h231 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18993; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25137 = 12'h231 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22065; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_561 = io_valid_in ? _GEN_25137 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_561 = 12'h231 == _T_2[11:0] ? image_561 : _GEN_560; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3634 = 12'h232 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6706 = 12'h232 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3634; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9778 = 12'h232 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6706; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12850 = 12'h232 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9778; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15922 = 12'h232 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12850; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18994 = 12'h232 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15922; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22066 = 12'h232 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18994; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25138 = 12'h232 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22066; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_562 = io_valid_in ? _GEN_25138 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_562 = 12'h232 == _T_2[11:0] ? image_562 : _GEN_561; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3635 = 12'h233 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6707 = 12'h233 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3635; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9779 = 12'h233 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6707; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12851 = 12'h233 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9779; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15923 = 12'h233 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12851; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18995 = 12'h233 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15923; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22067 = 12'h233 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18995; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25139 = 12'h233 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22067; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_563 = io_valid_in ? _GEN_25139 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_563 = 12'h233 == _T_2[11:0] ? image_563 : _GEN_562; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3636 = 12'h234 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6708 = 12'h234 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3636; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9780 = 12'h234 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6708; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12852 = 12'h234 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9780; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15924 = 12'h234 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12852; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18996 = 12'h234 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15924; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22068 = 12'h234 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18996; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25140 = 12'h234 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22068; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_564 = io_valid_in ? _GEN_25140 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_564 = 12'h234 == _T_2[11:0] ? image_564 : _GEN_563; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3637 = 12'h235 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6709 = 12'h235 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3637; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9781 = 12'h235 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6709; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12853 = 12'h235 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9781; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15925 = 12'h235 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12853; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18997 = 12'h235 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15925; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22069 = 12'h235 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18997; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25141 = 12'h235 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22069; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_565 = io_valid_in ? _GEN_25141 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_565 = 12'h235 == _T_2[11:0] ? image_565 : _GEN_564; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3638 = 12'h236 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6710 = 12'h236 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3638; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9782 = 12'h236 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6710; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12854 = 12'h236 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9782; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15926 = 12'h236 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12854; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18998 = 12'h236 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15926; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22070 = 12'h236 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18998; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25142 = 12'h236 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22070; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_566 = io_valid_in ? _GEN_25142 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_566 = 12'h236 == _T_2[11:0] ? image_566 : _GEN_565; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3639 = 12'h237 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6711 = 12'h237 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3639; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9783 = 12'h237 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6711; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12855 = 12'h237 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9783; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15927 = 12'h237 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12855; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18999 = 12'h237 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15927; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22071 = 12'h237 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_18999; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25143 = 12'h237 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22071; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_567 = io_valid_in ? _GEN_25143 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_567 = 12'h237 == _T_2[11:0] ? image_567 : _GEN_566; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3640 = 12'h238 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6712 = 12'h238 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3640; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9784 = 12'h238 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6712; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12856 = 12'h238 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9784; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15928 = 12'h238 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12856; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19000 = 12'h238 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15928; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22072 = 12'h238 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19000; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25144 = 12'h238 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22072; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_568 = io_valid_in ? _GEN_25144 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_568 = 12'h238 == _T_2[11:0] ? image_568 : _GEN_567; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3641 = 12'h239 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6713 = 12'h239 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3641; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9785 = 12'h239 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6713; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12857 = 12'h239 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9785; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15929 = 12'h239 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12857; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19001 = 12'h239 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15929; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22073 = 12'h239 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19001; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25145 = 12'h239 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22073; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_569 = io_valid_in ? _GEN_25145 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_569 = 12'h239 == _T_2[11:0] ? image_569 : _GEN_568; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3642 = 12'h23a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6714 = 12'h23a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3642; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9786 = 12'h23a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6714; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12858 = 12'h23a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9786; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15930 = 12'h23a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12858; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19002 = 12'h23a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15930; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22074 = 12'h23a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19002; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25146 = 12'h23a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22074; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_570 = io_valid_in ? _GEN_25146 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_570 = 12'h23a == _T_2[11:0] ? image_570 : _GEN_569; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3643 = 12'h23b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6715 = 12'h23b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3643; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9787 = 12'h23b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6715; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12859 = 12'h23b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9787; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15931 = 12'h23b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12859; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19003 = 12'h23b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15931; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22075 = 12'h23b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19003; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25147 = 12'h23b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22075; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_571 = io_valid_in ? _GEN_25147 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_571 = 12'h23b == _T_2[11:0] ? image_571 : _GEN_570; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3644 = 12'h23c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6716 = 12'h23c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3644; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9788 = 12'h23c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6716; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12860 = 12'h23c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9788; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15932 = 12'h23c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12860; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19004 = 12'h23c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15932; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22076 = 12'h23c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19004; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25148 = 12'h23c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22076; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_572 = io_valid_in ? _GEN_25148 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_572 = 12'h23c == _T_2[11:0] ? image_572 : _GEN_571; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3645 = 12'h23d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6717 = 12'h23d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3645; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9789 = 12'h23d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6717; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12861 = 12'h23d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9789; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15933 = 12'h23d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12861; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19005 = 12'h23d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15933; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22077 = 12'h23d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19005; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25149 = 12'h23d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22077; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_573 = io_valid_in ? _GEN_25149 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_573 = 12'h23d == _T_2[11:0] ? image_573 : _GEN_572; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3646 = 12'h23e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6718 = 12'h23e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3646; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9790 = 12'h23e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6718; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12862 = 12'h23e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9790; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15934 = 12'h23e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12862; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19006 = 12'h23e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15934; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22078 = 12'h23e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19006; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25150 = 12'h23e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22078; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_574 = io_valid_in ? _GEN_25150 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_574 = 12'h23e == _T_2[11:0] ? image_574 : _GEN_573; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3647 = 12'h23f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6719 = 12'h23f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3647; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9791 = 12'h23f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6719; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12863 = 12'h23f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9791; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15935 = 12'h23f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12863; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19007 = 12'h23f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15935; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22079 = 12'h23f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19007; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25151 = 12'h23f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22079; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_575 = io_valid_in ? _GEN_25151 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_575 = 12'h23f == _T_2[11:0] ? image_575 : _GEN_574; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3648 = 12'h240 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6720 = 12'h240 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3648; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9792 = 12'h240 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6720; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12864 = 12'h240 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9792; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15936 = 12'h240 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12864; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19008 = 12'h240 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15936; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22080 = 12'h240 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19008; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25152 = 12'h240 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22080; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_576 = io_valid_in ? _GEN_25152 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_576 = 12'h240 == _T_2[11:0] ? image_576 : _GEN_575; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3649 = 12'h241 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6721 = 12'h241 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3649; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9793 = 12'h241 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6721; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12865 = 12'h241 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9793; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15937 = 12'h241 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12865; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19009 = 12'h241 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15937; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22081 = 12'h241 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19009; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25153 = 12'h241 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22081; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_577 = io_valid_in ? _GEN_25153 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_577 = 12'h241 == _T_2[11:0] ? image_577 : _GEN_576; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3650 = 12'h242 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6722 = 12'h242 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3650; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9794 = 12'h242 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6722; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12866 = 12'h242 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9794; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15938 = 12'h242 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12866; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19010 = 12'h242 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15938; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22082 = 12'h242 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19010; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25154 = 12'h242 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22082; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_578 = io_valid_in ? _GEN_25154 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_578 = 12'h242 == _T_2[11:0] ? image_578 : _GEN_577; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3651 = 12'h243 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6723 = 12'h243 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3651; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9795 = 12'h243 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6723; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12867 = 12'h243 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9795; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15939 = 12'h243 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12867; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19011 = 12'h243 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15939; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22083 = 12'h243 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19011; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25155 = 12'h243 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22083; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_579 = io_valid_in ? _GEN_25155 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_579 = 12'h243 == _T_2[11:0] ? image_579 : _GEN_578; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3652 = 12'h244 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6724 = 12'h244 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3652; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9796 = 12'h244 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6724; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12868 = 12'h244 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9796; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15940 = 12'h244 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12868; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19012 = 12'h244 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15940; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22084 = 12'h244 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19012; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25156 = 12'h244 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22084; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_580 = io_valid_in ? _GEN_25156 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_580 = 12'h244 == _T_2[11:0] ? image_580 : _GEN_579; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3653 = 12'h245 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6725 = 12'h245 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3653; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9797 = 12'h245 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6725; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12869 = 12'h245 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9797; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15941 = 12'h245 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12869; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19013 = 12'h245 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15941; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22085 = 12'h245 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19013; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25157 = 12'h245 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22085; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_581 = io_valid_in ? _GEN_25157 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_581 = 12'h245 == _T_2[11:0] ? image_581 : _GEN_580; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3654 = 12'h246 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6726 = 12'h246 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3654; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9798 = 12'h246 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6726; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12870 = 12'h246 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9798; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15942 = 12'h246 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12870; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19014 = 12'h246 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15942; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22086 = 12'h246 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19014; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25158 = 12'h246 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22086; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_582 = io_valid_in ? _GEN_25158 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_582 = 12'h246 == _T_2[11:0] ? image_582 : _GEN_581; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3655 = 12'h247 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6727 = 12'h247 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3655; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9799 = 12'h247 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6727; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12871 = 12'h247 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9799; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15943 = 12'h247 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12871; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19015 = 12'h247 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15943; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22087 = 12'h247 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19015; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25159 = 12'h247 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22087; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_583 = io_valid_in ? _GEN_25159 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_583 = 12'h247 == _T_2[11:0] ? image_583 : _GEN_582; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3656 = 12'h248 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6728 = 12'h248 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3656; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9800 = 12'h248 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6728; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12872 = 12'h248 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9800; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15944 = 12'h248 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12872; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19016 = 12'h248 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15944; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22088 = 12'h248 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19016; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25160 = 12'h248 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22088; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_584 = io_valid_in ? _GEN_25160 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_584 = 12'h248 == _T_2[11:0] ? image_584 : _GEN_583; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3657 = 12'h249 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6729 = 12'h249 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3657; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9801 = 12'h249 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6729; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12873 = 12'h249 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9801; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15945 = 12'h249 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12873; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19017 = 12'h249 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15945; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22089 = 12'h249 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19017; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25161 = 12'h249 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22089; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_585 = io_valid_in ? _GEN_25161 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_585 = 12'h249 == _T_2[11:0] ? image_585 : _GEN_584; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3658 = 12'h24a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6730 = 12'h24a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3658; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9802 = 12'h24a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6730; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12874 = 12'h24a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9802; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15946 = 12'h24a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12874; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19018 = 12'h24a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15946; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22090 = 12'h24a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19018; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25162 = 12'h24a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22090; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_586 = io_valid_in ? _GEN_25162 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_586 = 12'h24a == _T_2[11:0] ? image_586 : _GEN_585; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3659 = 12'h24b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6731 = 12'h24b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3659; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9803 = 12'h24b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6731; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12875 = 12'h24b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9803; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15947 = 12'h24b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12875; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19019 = 12'h24b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15947; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22091 = 12'h24b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19019; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25163 = 12'h24b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22091; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_587 = io_valid_in ? _GEN_25163 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_587 = 12'h24b == _T_2[11:0] ? image_587 : _GEN_586; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3660 = 12'h24c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6732 = 12'h24c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3660; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9804 = 12'h24c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6732; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12876 = 12'h24c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9804; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15948 = 12'h24c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12876; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19020 = 12'h24c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15948; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22092 = 12'h24c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19020; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25164 = 12'h24c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22092; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_588 = io_valid_in ? _GEN_25164 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_588 = 12'h24c == _T_2[11:0] ? image_588 : _GEN_587; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3661 = 12'h24d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6733 = 12'h24d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3661; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9805 = 12'h24d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6733; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12877 = 12'h24d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9805; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15949 = 12'h24d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12877; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19021 = 12'h24d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15949; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22093 = 12'h24d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19021; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25165 = 12'h24d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22093; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_589 = io_valid_in ? _GEN_25165 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_589 = 12'h24d == _T_2[11:0] ? image_589 : _GEN_588; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3662 = 12'h24e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6734 = 12'h24e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3662; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9806 = 12'h24e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6734; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12878 = 12'h24e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9806; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15950 = 12'h24e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12878; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19022 = 12'h24e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15950; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22094 = 12'h24e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19022; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25166 = 12'h24e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22094; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_590 = io_valid_in ? _GEN_25166 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_590 = 12'h24e == _T_2[11:0] ? image_590 : _GEN_589; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3663 = 12'h24f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6735 = 12'h24f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3663; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9807 = 12'h24f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6735; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12879 = 12'h24f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9807; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15951 = 12'h24f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12879; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19023 = 12'h24f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15951; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22095 = 12'h24f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19023; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25167 = 12'h24f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22095; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_591 = io_valid_in ? _GEN_25167 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_591 = 12'h24f == _T_2[11:0] ? image_591 : _GEN_590; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3664 = 12'h250 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6736 = 12'h250 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3664; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9808 = 12'h250 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6736; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12880 = 12'h250 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9808; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15952 = 12'h250 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12880; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19024 = 12'h250 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15952; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22096 = 12'h250 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19024; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25168 = 12'h250 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22096; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_592 = io_valid_in ? _GEN_25168 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_592 = 12'h250 == _T_2[11:0] ? image_592 : _GEN_591; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3665 = 12'h251 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6737 = 12'h251 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3665; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9809 = 12'h251 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6737; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12881 = 12'h251 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9809; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15953 = 12'h251 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12881; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19025 = 12'h251 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15953; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22097 = 12'h251 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19025; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25169 = 12'h251 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22097; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_593 = io_valid_in ? _GEN_25169 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_593 = 12'h251 == _T_2[11:0] ? image_593 : _GEN_592; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3666 = 12'h252 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6738 = 12'h252 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3666; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9810 = 12'h252 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6738; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12882 = 12'h252 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9810; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15954 = 12'h252 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12882; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19026 = 12'h252 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15954; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22098 = 12'h252 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19026; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25170 = 12'h252 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22098; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_594 = io_valid_in ? _GEN_25170 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_594 = 12'h252 == _T_2[11:0] ? image_594 : _GEN_593; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3667 = 12'h253 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6739 = 12'h253 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3667; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9811 = 12'h253 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6739; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12883 = 12'h253 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9811; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15955 = 12'h253 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12883; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19027 = 12'h253 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15955; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22099 = 12'h253 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19027; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25171 = 12'h253 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22099; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_595 = io_valid_in ? _GEN_25171 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_595 = 12'h253 == _T_2[11:0] ? image_595 : _GEN_594; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3668 = 12'h254 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6740 = 12'h254 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3668; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9812 = 12'h254 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6740; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12884 = 12'h254 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9812; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15956 = 12'h254 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12884; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19028 = 12'h254 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15956; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22100 = 12'h254 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19028; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25172 = 12'h254 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22100; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_596 = io_valid_in ? _GEN_25172 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_596 = 12'h254 == _T_2[11:0] ? image_596 : _GEN_595; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3669 = 12'h255 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6741 = 12'h255 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3669; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9813 = 12'h255 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6741; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12885 = 12'h255 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9813; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15957 = 12'h255 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12885; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19029 = 12'h255 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15957; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22101 = 12'h255 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19029; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25173 = 12'h255 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22101; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_597 = io_valid_in ? _GEN_25173 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_597 = 12'h255 == _T_2[11:0] ? image_597 : _GEN_596; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3670 = 12'h256 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6742 = 12'h256 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3670; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9814 = 12'h256 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6742; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12886 = 12'h256 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9814; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15958 = 12'h256 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12886; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19030 = 12'h256 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15958; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22102 = 12'h256 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19030; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25174 = 12'h256 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22102; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_598 = io_valid_in ? _GEN_25174 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_598 = 12'h256 == _T_2[11:0] ? image_598 : _GEN_597; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3671 = 12'h257 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6743 = 12'h257 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3671; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9815 = 12'h257 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6743; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12887 = 12'h257 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9815; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15959 = 12'h257 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12887; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19031 = 12'h257 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15959; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22103 = 12'h257 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19031; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25175 = 12'h257 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22103; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_599 = io_valid_in ? _GEN_25175 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_599 = 12'h257 == _T_2[11:0] ? image_599 : _GEN_598; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3672 = 12'h258 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6744 = 12'h258 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3672; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9816 = 12'h258 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6744; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12888 = 12'h258 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9816; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15960 = 12'h258 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12888; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19032 = 12'h258 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15960; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22104 = 12'h258 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19032; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25176 = 12'h258 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22104; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_600 = io_valid_in ? _GEN_25176 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_600 = 12'h258 == _T_2[11:0] ? image_600 : _GEN_599; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3673 = 12'h259 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6745 = 12'h259 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3673; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9817 = 12'h259 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6745; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12889 = 12'h259 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9817; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15961 = 12'h259 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12889; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19033 = 12'h259 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15961; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22105 = 12'h259 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19033; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25177 = 12'h259 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22105; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_601 = io_valid_in ? _GEN_25177 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_601 = 12'h259 == _T_2[11:0] ? image_601 : _GEN_600; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3674 = 12'h25a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6746 = 12'h25a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3674; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9818 = 12'h25a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6746; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12890 = 12'h25a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9818; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15962 = 12'h25a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12890; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19034 = 12'h25a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15962; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22106 = 12'h25a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19034; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25178 = 12'h25a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22106; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_602 = io_valid_in ? _GEN_25178 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_602 = 12'h25a == _T_2[11:0] ? image_602 : _GEN_601; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3675 = 12'h25b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6747 = 12'h25b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3675; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9819 = 12'h25b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6747; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12891 = 12'h25b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9819; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15963 = 12'h25b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12891; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19035 = 12'h25b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15963; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22107 = 12'h25b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19035; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25179 = 12'h25b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22107; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_603 = io_valid_in ? _GEN_25179 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_603 = 12'h25b == _T_2[11:0] ? image_603 : _GEN_602; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3676 = 12'h25c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6748 = 12'h25c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3676; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9820 = 12'h25c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6748; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12892 = 12'h25c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9820; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15964 = 12'h25c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12892; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19036 = 12'h25c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15964; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22108 = 12'h25c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19036; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25180 = 12'h25c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22108; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_604 = io_valid_in ? _GEN_25180 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_604 = 12'h25c == _T_2[11:0] ? image_604 : _GEN_603; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3677 = 12'h25d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6749 = 12'h25d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3677; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9821 = 12'h25d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6749; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12893 = 12'h25d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9821; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15965 = 12'h25d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12893; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19037 = 12'h25d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15965; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22109 = 12'h25d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19037; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25181 = 12'h25d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22109; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_605 = io_valid_in ? _GEN_25181 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_605 = 12'h25d == _T_2[11:0] ? image_605 : _GEN_604; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3678 = 12'h25e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6750 = 12'h25e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3678; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9822 = 12'h25e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6750; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12894 = 12'h25e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9822; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15966 = 12'h25e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12894; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19038 = 12'h25e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15966; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22110 = 12'h25e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19038; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25182 = 12'h25e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22110; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_606 = io_valid_in ? _GEN_25182 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_606 = 12'h25e == _T_2[11:0] ? image_606 : _GEN_605; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3679 = 12'h25f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6751 = 12'h25f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3679; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9823 = 12'h25f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6751; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12895 = 12'h25f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9823; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15967 = 12'h25f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12895; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19039 = 12'h25f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15967; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22111 = 12'h25f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19039; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25183 = 12'h25f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22111; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_607 = io_valid_in ? _GEN_25183 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_607 = 12'h25f == _T_2[11:0] ? image_607 : _GEN_606; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3680 = 12'h260 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6752 = 12'h260 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3680; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9824 = 12'h260 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6752; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12896 = 12'h260 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9824; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15968 = 12'h260 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12896; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19040 = 12'h260 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15968; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22112 = 12'h260 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19040; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25184 = 12'h260 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22112; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_608 = io_valid_in ? _GEN_25184 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_608 = 12'h260 == _T_2[11:0] ? image_608 : _GEN_607; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3681 = 12'h261 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6753 = 12'h261 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3681; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9825 = 12'h261 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6753; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12897 = 12'h261 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9825; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15969 = 12'h261 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12897; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19041 = 12'h261 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15969; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22113 = 12'h261 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19041; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25185 = 12'h261 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22113; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_609 = io_valid_in ? _GEN_25185 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_609 = 12'h261 == _T_2[11:0] ? image_609 : _GEN_608; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3682 = 12'h262 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6754 = 12'h262 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3682; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9826 = 12'h262 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6754; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12898 = 12'h262 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9826; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15970 = 12'h262 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12898; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19042 = 12'h262 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15970; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22114 = 12'h262 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19042; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25186 = 12'h262 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22114; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_610 = io_valid_in ? _GEN_25186 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_610 = 12'h262 == _T_2[11:0] ? image_610 : _GEN_609; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3683 = 12'h263 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6755 = 12'h263 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3683; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9827 = 12'h263 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6755; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12899 = 12'h263 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9827; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15971 = 12'h263 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12899; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19043 = 12'h263 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15971; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22115 = 12'h263 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19043; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25187 = 12'h263 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22115; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_611 = io_valid_in ? _GEN_25187 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_611 = 12'h263 == _T_2[11:0] ? image_611 : _GEN_610; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3684 = 12'h264 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6756 = 12'h264 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3684; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9828 = 12'h264 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6756; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12900 = 12'h264 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9828; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15972 = 12'h264 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12900; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19044 = 12'h264 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15972; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22116 = 12'h264 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19044; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25188 = 12'h264 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22116; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_612 = io_valid_in ? _GEN_25188 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_612 = 12'h264 == _T_2[11:0] ? image_612 : _GEN_611; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3685 = 12'h265 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6757 = 12'h265 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3685; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9829 = 12'h265 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6757; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12901 = 12'h265 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9829; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15973 = 12'h265 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12901; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19045 = 12'h265 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15973; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22117 = 12'h265 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19045; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25189 = 12'h265 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22117; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_613 = io_valid_in ? _GEN_25189 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_613 = 12'h265 == _T_2[11:0] ? image_613 : _GEN_612; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3686 = 12'h266 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6758 = 12'h266 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3686; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9830 = 12'h266 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6758; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12902 = 12'h266 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9830; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15974 = 12'h266 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12902; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19046 = 12'h266 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15974; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22118 = 12'h266 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19046; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25190 = 12'h266 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22118; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_614 = io_valid_in ? _GEN_25190 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_614 = 12'h266 == _T_2[11:0] ? image_614 : _GEN_613; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3687 = 12'h267 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6759 = 12'h267 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3687; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9831 = 12'h267 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6759; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12903 = 12'h267 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9831; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15975 = 12'h267 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12903; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19047 = 12'h267 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15975; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22119 = 12'h267 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19047; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25191 = 12'h267 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22119; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_615 = io_valid_in ? _GEN_25191 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_615 = 12'h267 == _T_2[11:0] ? image_615 : _GEN_614; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3688 = 12'h268 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6760 = 12'h268 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3688; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9832 = 12'h268 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6760; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12904 = 12'h268 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9832; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15976 = 12'h268 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12904; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19048 = 12'h268 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15976; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22120 = 12'h268 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19048; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25192 = 12'h268 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22120; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_616 = io_valid_in ? _GEN_25192 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_616 = 12'h268 == _T_2[11:0] ? image_616 : _GEN_615; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3689 = 12'h269 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6761 = 12'h269 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3689; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9833 = 12'h269 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6761; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12905 = 12'h269 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9833; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15977 = 12'h269 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12905; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19049 = 12'h269 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15977; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22121 = 12'h269 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19049; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25193 = 12'h269 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22121; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_617 = io_valid_in ? _GEN_25193 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_617 = 12'h269 == _T_2[11:0] ? image_617 : _GEN_616; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3690 = 12'h26a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6762 = 12'h26a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3690; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9834 = 12'h26a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6762; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12906 = 12'h26a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9834; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15978 = 12'h26a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12906; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19050 = 12'h26a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15978; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22122 = 12'h26a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19050; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25194 = 12'h26a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22122; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_618 = io_valid_in ? _GEN_25194 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_618 = 12'h26a == _T_2[11:0] ? image_618 : _GEN_617; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3691 = 12'h26b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6763 = 12'h26b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3691; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9835 = 12'h26b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6763; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12907 = 12'h26b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9835; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15979 = 12'h26b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12907; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19051 = 12'h26b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15979; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22123 = 12'h26b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19051; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25195 = 12'h26b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22123; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_619 = io_valid_in ? _GEN_25195 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_619 = 12'h26b == _T_2[11:0] ? image_619 : _GEN_618; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3692 = 12'h26c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6764 = 12'h26c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3692; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9836 = 12'h26c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6764; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12908 = 12'h26c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9836; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15980 = 12'h26c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12908; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19052 = 12'h26c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15980; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22124 = 12'h26c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19052; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25196 = 12'h26c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22124; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_620 = io_valid_in ? _GEN_25196 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_620 = 12'h26c == _T_2[11:0] ? image_620 : _GEN_619; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3693 = 12'h26d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6765 = 12'h26d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3693; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9837 = 12'h26d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6765; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12909 = 12'h26d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9837; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15981 = 12'h26d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12909; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19053 = 12'h26d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15981; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22125 = 12'h26d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19053; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25197 = 12'h26d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22125; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_621 = io_valid_in ? _GEN_25197 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_621 = 12'h26d == _T_2[11:0] ? image_621 : _GEN_620; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3694 = 12'h26e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6766 = 12'h26e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3694; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9838 = 12'h26e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6766; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12910 = 12'h26e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9838; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15982 = 12'h26e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12910; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19054 = 12'h26e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15982; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22126 = 12'h26e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19054; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25198 = 12'h26e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22126; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_622 = io_valid_in ? _GEN_25198 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_622 = 12'h26e == _T_2[11:0] ? image_622 : _GEN_621; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3695 = 12'h26f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6767 = 12'h26f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3695; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9839 = 12'h26f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6767; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12911 = 12'h26f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9839; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15983 = 12'h26f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12911; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19055 = 12'h26f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15983; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22127 = 12'h26f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19055; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25199 = 12'h26f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22127; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_623 = io_valid_in ? _GEN_25199 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_623 = 12'h26f == _T_2[11:0] ? image_623 : _GEN_622; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3696 = 12'h270 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6768 = 12'h270 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3696; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9840 = 12'h270 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6768; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12912 = 12'h270 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9840; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15984 = 12'h270 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12912; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19056 = 12'h270 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15984; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22128 = 12'h270 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19056; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25200 = 12'h270 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22128; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_624 = io_valid_in ? _GEN_25200 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_624 = 12'h270 == _T_2[11:0] ? image_624 : _GEN_623; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3697 = 12'h271 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6769 = 12'h271 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3697; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9841 = 12'h271 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6769; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12913 = 12'h271 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9841; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15985 = 12'h271 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12913; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19057 = 12'h271 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15985; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22129 = 12'h271 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19057; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25201 = 12'h271 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22129; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_625 = io_valid_in ? _GEN_25201 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_625 = 12'h271 == _T_2[11:0] ? image_625 : _GEN_624; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3698 = 12'h272 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6770 = 12'h272 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3698; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9842 = 12'h272 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6770; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12914 = 12'h272 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9842; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15986 = 12'h272 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12914; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19058 = 12'h272 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15986; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22130 = 12'h272 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19058; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25202 = 12'h272 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22130; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_626 = io_valid_in ? _GEN_25202 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_626 = 12'h272 == _T_2[11:0] ? image_626 : _GEN_625; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3699 = 12'h273 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6771 = 12'h273 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3699; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9843 = 12'h273 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6771; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12915 = 12'h273 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9843; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15987 = 12'h273 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12915; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19059 = 12'h273 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15987; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22131 = 12'h273 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19059; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25203 = 12'h273 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22131; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_627 = io_valid_in ? _GEN_25203 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_627 = 12'h273 == _T_2[11:0] ? image_627 : _GEN_626; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3700 = 12'h274 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6772 = 12'h274 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3700; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9844 = 12'h274 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6772; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12916 = 12'h274 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9844; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15988 = 12'h274 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12916; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19060 = 12'h274 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15988; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22132 = 12'h274 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19060; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25204 = 12'h274 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22132; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_628 = io_valid_in ? _GEN_25204 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_628 = 12'h274 == _T_2[11:0] ? image_628 : _GEN_627; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3701 = 12'h275 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6773 = 12'h275 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3701; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9845 = 12'h275 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6773; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12917 = 12'h275 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9845; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15989 = 12'h275 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12917; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19061 = 12'h275 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15989; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22133 = 12'h275 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19061; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25205 = 12'h275 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22133; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_629 = io_valid_in ? _GEN_25205 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_629 = 12'h275 == _T_2[11:0] ? image_629 : _GEN_628; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3702 = 12'h276 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6774 = 12'h276 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3702; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9846 = 12'h276 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6774; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12918 = 12'h276 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9846; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15990 = 12'h276 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12918; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19062 = 12'h276 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15990; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22134 = 12'h276 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19062; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25206 = 12'h276 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22134; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_630 = io_valid_in ? _GEN_25206 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_630 = 12'h276 == _T_2[11:0] ? image_630 : _GEN_629; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3703 = 12'h277 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6775 = 12'h277 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3703; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9847 = 12'h277 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6775; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12919 = 12'h277 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9847; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15991 = 12'h277 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12919; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19063 = 12'h277 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15991; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22135 = 12'h277 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19063; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25207 = 12'h277 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22135; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_631 = io_valid_in ? _GEN_25207 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_631 = 12'h277 == _T_2[11:0] ? image_631 : _GEN_630; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3704 = 12'h278 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6776 = 12'h278 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3704; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9848 = 12'h278 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6776; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12920 = 12'h278 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9848; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15992 = 12'h278 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12920; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19064 = 12'h278 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15992; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22136 = 12'h278 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19064; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25208 = 12'h278 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22136; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_632 = io_valid_in ? _GEN_25208 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_632 = 12'h278 == _T_2[11:0] ? image_632 : _GEN_631; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3705 = 12'h279 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6777 = 12'h279 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3705; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9849 = 12'h279 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6777; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12921 = 12'h279 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9849; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15993 = 12'h279 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12921; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19065 = 12'h279 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15993; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22137 = 12'h279 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19065; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25209 = 12'h279 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22137; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_633 = io_valid_in ? _GEN_25209 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_633 = 12'h279 == _T_2[11:0] ? image_633 : _GEN_632; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3706 = 12'h27a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6778 = 12'h27a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3706; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9850 = 12'h27a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6778; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12922 = 12'h27a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9850; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15994 = 12'h27a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12922; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19066 = 12'h27a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15994; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22138 = 12'h27a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19066; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25210 = 12'h27a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22138; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_634 = io_valid_in ? _GEN_25210 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_634 = 12'h27a == _T_2[11:0] ? image_634 : _GEN_633; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3707 = 12'h27b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6779 = 12'h27b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3707; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9851 = 12'h27b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6779; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12923 = 12'h27b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9851; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15995 = 12'h27b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12923; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19067 = 12'h27b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15995; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22139 = 12'h27b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19067; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25211 = 12'h27b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22139; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_635 = io_valid_in ? _GEN_25211 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_635 = 12'h27b == _T_2[11:0] ? image_635 : _GEN_634; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3708 = 12'h27c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6780 = 12'h27c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3708; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9852 = 12'h27c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6780; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12924 = 12'h27c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9852; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15996 = 12'h27c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12924; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19068 = 12'h27c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15996; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22140 = 12'h27c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19068; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25212 = 12'h27c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22140; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_636 = io_valid_in ? _GEN_25212 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_636 = 12'h27c == _T_2[11:0] ? image_636 : _GEN_635; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3709 = 12'h27d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6781 = 12'h27d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3709; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9853 = 12'h27d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6781; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12925 = 12'h27d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9853; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15997 = 12'h27d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12925; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19069 = 12'h27d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15997; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22141 = 12'h27d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19069; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25213 = 12'h27d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22141; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_637 = io_valid_in ? _GEN_25213 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_637 = 12'h27d == _T_2[11:0] ? image_637 : _GEN_636; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3710 = 12'h27e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6782 = 12'h27e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3710; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9854 = 12'h27e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6782; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12926 = 12'h27e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9854; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15998 = 12'h27e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12926; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19070 = 12'h27e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15998; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22142 = 12'h27e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19070; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25214 = 12'h27e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22142; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_638 = io_valid_in ? _GEN_25214 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_638 = 12'h27e == _T_2[11:0] ? image_638 : _GEN_637; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3711 = 12'h27f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6783 = 12'h27f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3711; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9855 = 12'h27f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6783; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12927 = 12'h27f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9855; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15999 = 12'h27f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12927; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19071 = 12'h27f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_15999; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22143 = 12'h27f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19071; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25215 = 12'h27f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22143; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_639 = io_valid_in ? _GEN_25215 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_639 = 12'h27f == _T_2[11:0] ? image_639 : _GEN_638; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3712 = 12'h280 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6784 = 12'h280 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3712; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9856 = 12'h280 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6784; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12928 = 12'h280 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9856; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16000 = 12'h280 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12928; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19072 = 12'h280 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16000; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22144 = 12'h280 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19072; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25216 = 12'h280 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22144; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_640 = io_valid_in ? _GEN_25216 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_640 = 12'h280 == _T_2[11:0] ? image_640 : _GEN_639; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3713 = 12'h281 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6785 = 12'h281 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3713; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9857 = 12'h281 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6785; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12929 = 12'h281 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9857; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16001 = 12'h281 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12929; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19073 = 12'h281 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16001; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22145 = 12'h281 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19073; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25217 = 12'h281 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22145; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_641 = io_valid_in ? _GEN_25217 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_641 = 12'h281 == _T_2[11:0] ? image_641 : _GEN_640; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3714 = 12'h282 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6786 = 12'h282 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3714; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9858 = 12'h282 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6786; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12930 = 12'h282 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9858; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16002 = 12'h282 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12930; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19074 = 12'h282 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16002; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22146 = 12'h282 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19074; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25218 = 12'h282 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22146; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_642 = io_valid_in ? _GEN_25218 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_642 = 12'h282 == _T_2[11:0] ? image_642 : _GEN_641; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3715 = 12'h283 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6787 = 12'h283 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3715; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9859 = 12'h283 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6787; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12931 = 12'h283 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9859; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16003 = 12'h283 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12931; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19075 = 12'h283 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16003; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22147 = 12'h283 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19075; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25219 = 12'h283 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22147; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_643 = io_valid_in ? _GEN_25219 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_643 = 12'h283 == _T_2[11:0] ? image_643 : _GEN_642; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3716 = 12'h284 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6788 = 12'h284 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3716; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9860 = 12'h284 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6788; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12932 = 12'h284 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9860; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16004 = 12'h284 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12932; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19076 = 12'h284 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16004; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22148 = 12'h284 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19076; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25220 = 12'h284 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22148; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_644 = io_valid_in ? _GEN_25220 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_644 = 12'h284 == _T_2[11:0] ? image_644 : _GEN_643; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3717 = 12'h285 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6789 = 12'h285 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3717; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9861 = 12'h285 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6789; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12933 = 12'h285 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9861; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16005 = 12'h285 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12933; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19077 = 12'h285 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16005; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22149 = 12'h285 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19077; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25221 = 12'h285 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22149; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_645 = io_valid_in ? _GEN_25221 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_645 = 12'h285 == _T_2[11:0] ? image_645 : _GEN_644; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3718 = 12'h286 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6790 = 12'h286 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3718; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9862 = 12'h286 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6790; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12934 = 12'h286 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9862; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16006 = 12'h286 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12934; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19078 = 12'h286 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16006; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22150 = 12'h286 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19078; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25222 = 12'h286 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22150; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_646 = io_valid_in ? _GEN_25222 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_646 = 12'h286 == _T_2[11:0] ? image_646 : _GEN_645; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3719 = 12'h287 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6791 = 12'h287 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3719; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9863 = 12'h287 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6791; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12935 = 12'h287 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9863; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16007 = 12'h287 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12935; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19079 = 12'h287 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16007; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22151 = 12'h287 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19079; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25223 = 12'h287 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22151; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_647 = io_valid_in ? _GEN_25223 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_647 = 12'h287 == _T_2[11:0] ? image_647 : _GEN_646; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3720 = 12'h288 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6792 = 12'h288 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3720; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9864 = 12'h288 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6792; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12936 = 12'h288 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9864; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16008 = 12'h288 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12936; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19080 = 12'h288 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16008; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22152 = 12'h288 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19080; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25224 = 12'h288 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22152; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_648 = io_valid_in ? _GEN_25224 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_648 = 12'h288 == _T_2[11:0] ? image_648 : _GEN_647; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3721 = 12'h289 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6793 = 12'h289 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3721; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9865 = 12'h289 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6793; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12937 = 12'h289 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9865; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16009 = 12'h289 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12937; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19081 = 12'h289 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16009; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22153 = 12'h289 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19081; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25225 = 12'h289 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22153; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_649 = io_valid_in ? _GEN_25225 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_649 = 12'h289 == _T_2[11:0] ? image_649 : _GEN_648; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3722 = 12'h28a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6794 = 12'h28a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3722; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9866 = 12'h28a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6794; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12938 = 12'h28a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9866; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16010 = 12'h28a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12938; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19082 = 12'h28a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16010; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22154 = 12'h28a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19082; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25226 = 12'h28a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22154; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_650 = io_valid_in ? _GEN_25226 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_650 = 12'h28a == _T_2[11:0] ? image_650 : _GEN_649; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3723 = 12'h28b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6795 = 12'h28b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3723; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9867 = 12'h28b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6795; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12939 = 12'h28b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9867; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16011 = 12'h28b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12939; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19083 = 12'h28b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16011; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22155 = 12'h28b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19083; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25227 = 12'h28b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22155; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_651 = io_valid_in ? _GEN_25227 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_651 = 12'h28b == _T_2[11:0] ? image_651 : _GEN_650; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3724 = 12'h28c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6796 = 12'h28c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3724; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9868 = 12'h28c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6796; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12940 = 12'h28c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9868; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16012 = 12'h28c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12940; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19084 = 12'h28c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16012; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22156 = 12'h28c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19084; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25228 = 12'h28c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22156; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_652 = io_valid_in ? _GEN_25228 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_652 = 12'h28c == _T_2[11:0] ? image_652 : _GEN_651; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3725 = 12'h28d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6797 = 12'h28d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3725; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9869 = 12'h28d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6797; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12941 = 12'h28d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9869; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16013 = 12'h28d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12941; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19085 = 12'h28d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16013; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22157 = 12'h28d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19085; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25229 = 12'h28d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22157; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_653 = io_valid_in ? _GEN_25229 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_653 = 12'h28d == _T_2[11:0] ? image_653 : _GEN_652; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3726 = 12'h28e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6798 = 12'h28e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3726; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9870 = 12'h28e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6798; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12942 = 12'h28e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9870; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16014 = 12'h28e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12942; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19086 = 12'h28e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16014; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22158 = 12'h28e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19086; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25230 = 12'h28e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22158; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_654 = io_valid_in ? _GEN_25230 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_654 = 12'h28e == _T_2[11:0] ? image_654 : _GEN_653; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3727 = 12'h28f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6799 = 12'h28f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3727; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9871 = 12'h28f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6799; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12943 = 12'h28f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9871; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16015 = 12'h28f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12943; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19087 = 12'h28f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16015; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22159 = 12'h28f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19087; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25231 = 12'h28f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22159; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_655 = io_valid_in ? _GEN_25231 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_655 = 12'h28f == _T_2[11:0] ? image_655 : _GEN_654; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3728 = 12'h290 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6800 = 12'h290 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3728; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9872 = 12'h290 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6800; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12944 = 12'h290 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9872; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16016 = 12'h290 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12944; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19088 = 12'h290 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16016; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22160 = 12'h290 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19088; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25232 = 12'h290 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22160; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_656 = io_valid_in ? _GEN_25232 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_656 = 12'h290 == _T_2[11:0] ? image_656 : _GEN_655; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3729 = 12'h291 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6801 = 12'h291 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3729; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9873 = 12'h291 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6801; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12945 = 12'h291 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9873; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16017 = 12'h291 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12945; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19089 = 12'h291 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16017; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22161 = 12'h291 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19089; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25233 = 12'h291 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22161; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_657 = io_valid_in ? _GEN_25233 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_657 = 12'h291 == _T_2[11:0] ? image_657 : _GEN_656; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3730 = 12'h292 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6802 = 12'h292 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3730; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9874 = 12'h292 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6802; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12946 = 12'h292 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9874; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16018 = 12'h292 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12946; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19090 = 12'h292 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16018; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22162 = 12'h292 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19090; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25234 = 12'h292 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22162; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_658 = io_valid_in ? _GEN_25234 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_658 = 12'h292 == _T_2[11:0] ? image_658 : _GEN_657; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3731 = 12'h293 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6803 = 12'h293 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3731; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9875 = 12'h293 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6803; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12947 = 12'h293 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9875; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16019 = 12'h293 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12947; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19091 = 12'h293 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16019; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22163 = 12'h293 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19091; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25235 = 12'h293 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22163; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_659 = io_valid_in ? _GEN_25235 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_659 = 12'h293 == _T_2[11:0] ? image_659 : _GEN_658; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3732 = 12'h294 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6804 = 12'h294 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3732; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9876 = 12'h294 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6804; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12948 = 12'h294 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9876; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16020 = 12'h294 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12948; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19092 = 12'h294 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16020; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22164 = 12'h294 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19092; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25236 = 12'h294 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22164; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_660 = io_valid_in ? _GEN_25236 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_660 = 12'h294 == _T_2[11:0] ? image_660 : _GEN_659; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3733 = 12'h295 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6805 = 12'h295 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3733; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9877 = 12'h295 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6805; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12949 = 12'h295 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9877; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16021 = 12'h295 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12949; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19093 = 12'h295 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16021; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22165 = 12'h295 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19093; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25237 = 12'h295 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22165; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_661 = io_valid_in ? _GEN_25237 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_661 = 12'h295 == _T_2[11:0] ? image_661 : _GEN_660; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3734 = 12'h296 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6806 = 12'h296 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3734; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9878 = 12'h296 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6806; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12950 = 12'h296 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9878; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16022 = 12'h296 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12950; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19094 = 12'h296 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16022; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22166 = 12'h296 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19094; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25238 = 12'h296 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22166; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_662 = io_valid_in ? _GEN_25238 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_662 = 12'h296 == _T_2[11:0] ? image_662 : _GEN_661; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3735 = 12'h297 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6807 = 12'h297 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3735; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9879 = 12'h297 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6807; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12951 = 12'h297 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9879; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16023 = 12'h297 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12951; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19095 = 12'h297 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16023; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22167 = 12'h297 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19095; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25239 = 12'h297 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22167; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_663 = io_valid_in ? _GEN_25239 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_663 = 12'h297 == _T_2[11:0] ? image_663 : _GEN_662; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3736 = 12'h298 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6808 = 12'h298 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3736; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9880 = 12'h298 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6808; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12952 = 12'h298 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9880; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16024 = 12'h298 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12952; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19096 = 12'h298 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16024; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22168 = 12'h298 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19096; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25240 = 12'h298 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22168; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_664 = io_valid_in ? _GEN_25240 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_664 = 12'h298 == _T_2[11:0] ? image_664 : _GEN_663; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3737 = 12'h299 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6809 = 12'h299 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3737; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9881 = 12'h299 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6809; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12953 = 12'h299 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9881; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16025 = 12'h299 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12953; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19097 = 12'h299 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16025; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22169 = 12'h299 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19097; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25241 = 12'h299 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22169; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_665 = io_valid_in ? _GEN_25241 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_665 = 12'h299 == _T_2[11:0] ? image_665 : _GEN_664; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3738 = 12'h29a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6810 = 12'h29a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3738; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9882 = 12'h29a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6810; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12954 = 12'h29a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9882; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16026 = 12'h29a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12954; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19098 = 12'h29a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16026; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22170 = 12'h29a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19098; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25242 = 12'h29a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22170; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_666 = io_valid_in ? _GEN_25242 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_666 = 12'h29a == _T_2[11:0] ? image_666 : _GEN_665; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3739 = 12'h29b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6811 = 12'h29b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3739; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9883 = 12'h29b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6811; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12955 = 12'h29b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9883; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16027 = 12'h29b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12955; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19099 = 12'h29b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16027; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22171 = 12'h29b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19099; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25243 = 12'h29b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22171; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_667 = io_valid_in ? _GEN_25243 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_667 = 12'h29b == _T_2[11:0] ? image_667 : _GEN_666; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3740 = 12'h29c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6812 = 12'h29c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3740; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9884 = 12'h29c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6812; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12956 = 12'h29c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9884; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16028 = 12'h29c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12956; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19100 = 12'h29c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16028; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22172 = 12'h29c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19100; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25244 = 12'h29c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22172; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_668 = io_valid_in ? _GEN_25244 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_668 = 12'h29c == _T_2[11:0] ? image_668 : _GEN_667; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3741 = 12'h29d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6813 = 12'h29d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3741; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9885 = 12'h29d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6813; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12957 = 12'h29d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9885; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16029 = 12'h29d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12957; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19101 = 12'h29d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16029; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22173 = 12'h29d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19101; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25245 = 12'h29d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22173; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_669 = io_valid_in ? _GEN_25245 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_669 = 12'h29d == _T_2[11:0] ? image_669 : _GEN_668; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3742 = 12'h29e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6814 = 12'h29e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3742; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9886 = 12'h29e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6814; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12958 = 12'h29e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9886; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16030 = 12'h29e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12958; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19102 = 12'h29e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16030; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22174 = 12'h29e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19102; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25246 = 12'h29e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22174; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_670 = io_valid_in ? _GEN_25246 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_670 = 12'h29e == _T_2[11:0] ? image_670 : _GEN_669; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3743 = 12'h29f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6815 = 12'h29f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3743; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9887 = 12'h29f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6815; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12959 = 12'h29f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9887; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16031 = 12'h29f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12959; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19103 = 12'h29f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16031; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22175 = 12'h29f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19103; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25247 = 12'h29f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22175; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_671 = io_valid_in ? _GEN_25247 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_671 = 12'h29f == _T_2[11:0] ? image_671 : _GEN_670; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3744 = 12'h2a0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6816 = 12'h2a0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3744; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9888 = 12'h2a0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6816; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12960 = 12'h2a0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9888; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16032 = 12'h2a0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12960; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19104 = 12'h2a0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16032; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22176 = 12'h2a0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19104; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25248 = 12'h2a0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22176; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_672 = io_valid_in ? _GEN_25248 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_672 = 12'h2a0 == _T_2[11:0] ? image_672 : _GEN_671; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3745 = 12'h2a1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6817 = 12'h2a1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3745; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9889 = 12'h2a1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6817; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12961 = 12'h2a1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9889; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16033 = 12'h2a1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12961; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19105 = 12'h2a1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16033; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22177 = 12'h2a1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19105; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25249 = 12'h2a1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22177; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_673 = io_valid_in ? _GEN_25249 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_673 = 12'h2a1 == _T_2[11:0] ? image_673 : _GEN_672; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3746 = 12'h2a2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6818 = 12'h2a2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3746; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9890 = 12'h2a2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6818; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12962 = 12'h2a2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9890; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16034 = 12'h2a2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12962; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19106 = 12'h2a2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16034; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22178 = 12'h2a2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19106; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25250 = 12'h2a2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22178; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_674 = io_valid_in ? _GEN_25250 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_674 = 12'h2a2 == _T_2[11:0] ? image_674 : _GEN_673; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3747 = 12'h2a3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6819 = 12'h2a3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3747; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9891 = 12'h2a3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6819; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12963 = 12'h2a3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9891; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16035 = 12'h2a3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12963; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19107 = 12'h2a3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16035; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22179 = 12'h2a3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19107; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25251 = 12'h2a3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22179; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_675 = io_valid_in ? _GEN_25251 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_675 = 12'h2a3 == _T_2[11:0] ? image_675 : _GEN_674; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3748 = 12'h2a4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6820 = 12'h2a4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3748; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9892 = 12'h2a4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6820; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12964 = 12'h2a4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9892; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16036 = 12'h2a4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12964; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19108 = 12'h2a4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16036; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22180 = 12'h2a4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19108; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25252 = 12'h2a4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22180; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_676 = io_valid_in ? _GEN_25252 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_676 = 12'h2a4 == _T_2[11:0] ? image_676 : _GEN_675; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3749 = 12'h2a5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6821 = 12'h2a5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3749; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9893 = 12'h2a5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6821; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12965 = 12'h2a5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9893; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16037 = 12'h2a5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12965; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19109 = 12'h2a5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16037; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22181 = 12'h2a5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19109; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25253 = 12'h2a5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22181; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_677 = io_valid_in ? _GEN_25253 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_677 = 12'h2a5 == _T_2[11:0] ? image_677 : _GEN_676; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3750 = 12'h2a6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6822 = 12'h2a6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3750; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9894 = 12'h2a6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6822; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12966 = 12'h2a6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9894; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16038 = 12'h2a6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12966; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19110 = 12'h2a6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16038; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22182 = 12'h2a6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19110; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25254 = 12'h2a6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22182; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_678 = io_valid_in ? _GEN_25254 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_678 = 12'h2a6 == _T_2[11:0] ? image_678 : _GEN_677; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3751 = 12'h2a7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6823 = 12'h2a7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3751; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9895 = 12'h2a7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6823; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12967 = 12'h2a7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9895; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16039 = 12'h2a7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12967; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19111 = 12'h2a7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16039; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22183 = 12'h2a7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19111; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25255 = 12'h2a7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22183; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_679 = io_valid_in ? _GEN_25255 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_679 = 12'h2a7 == _T_2[11:0] ? image_679 : _GEN_678; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3752 = 12'h2a8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6824 = 12'h2a8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3752; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9896 = 12'h2a8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6824; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12968 = 12'h2a8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9896; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16040 = 12'h2a8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12968; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19112 = 12'h2a8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16040; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22184 = 12'h2a8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19112; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25256 = 12'h2a8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22184; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_680 = io_valid_in ? _GEN_25256 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_680 = 12'h2a8 == _T_2[11:0] ? image_680 : _GEN_679; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3753 = 12'h2a9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6825 = 12'h2a9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3753; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9897 = 12'h2a9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6825; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12969 = 12'h2a9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9897; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16041 = 12'h2a9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12969; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19113 = 12'h2a9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16041; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22185 = 12'h2a9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19113; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25257 = 12'h2a9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22185; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_681 = io_valid_in ? _GEN_25257 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_681 = 12'h2a9 == _T_2[11:0] ? image_681 : _GEN_680; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3754 = 12'h2aa == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6826 = 12'h2aa == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3754; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9898 = 12'h2aa == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6826; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12970 = 12'h2aa == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9898; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16042 = 12'h2aa == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12970; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19114 = 12'h2aa == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16042; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22186 = 12'h2aa == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19114; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25258 = 12'h2aa == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22186; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_682 = io_valid_in ? _GEN_25258 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_682 = 12'h2aa == _T_2[11:0] ? image_682 : _GEN_681; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3755 = 12'h2ab == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6827 = 12'h2ab == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3755; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9899 = 12'h2ab == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6827; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12971 = 12'h2ab == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9899; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16043 = 12'h2ab == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12971; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19115 = 12'h2ab == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16043; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22187 = 12'h2ab == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19115; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25259 = 12'h2ab == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22187; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_683 = io_valid_in ? _GEN_25259 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_683 = 12'h2ab == _T_2[11:0] ? image_683 : _GEN_682; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3756 = 12'h2ac == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6828 = 12'h2ac == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3756; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9900 = 12'h2ac == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6828; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12972 = 12'h2ac == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9900; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16044 = 12'h2ac == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12972; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19116 = 12'h2ac == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16044; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22188 = 12'h2ac == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19116; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25260 = 12'h2ac == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22188; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_684 = io_valid_in ? _GEN_25260 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_684 = 12'h2ac == _T_2[11:0] ? image_684 : _GEN_683; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3757 = 12'h2ad == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6829 = 12'h2ad == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3757; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9901 = 12'h2ad == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6829; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12973 = 12'h2ad == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9901; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16045 = 12'h2ad == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12973; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19117 = 12'h2ad == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16045; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22189 = 12'h2ad == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19117; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25261 = 12'h2ad == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22189; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_685 = io_valid_in ? _GEN_25261 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_685 = 12'h2ad == _T_2[11:0] ? image_685 : _GEN_684; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3758 = 12'h2ae == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6830 = 12'h2ae == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3758; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9902 = 12'h2ae == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6830; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12974 = 12'h2ae == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9902; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16046 = 12'h2ae == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12974; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19118 = 12'h2ae == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16046; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22190 = 12'h2ae == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19118; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25262 = 12'h2ae == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22190; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_686 = io_valid_in ? _GEN_25262 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_686 = 12'h2ae == _T_2[11:0] ? image_686 : _GEN_685; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3759 = 12'h2af == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6831 = 12'h2af == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3759; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9903 = 12'h2af == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6831; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12975 = 12'h2af == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9903; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16047 = 12'h2af == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12975; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19119 = 12'h2af == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16047; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22191 = 12'h2af == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19119; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25263 = 12'h2af == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22191; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_687 = io_valid_in ? _GEN_25263 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_687 = 12'h2af == _T_2[11:0] ? image_687 : _GEN_686; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3760 = 12'h2b0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6832 = 12'h2b0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3760; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9904 = 12'h2b0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6832; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12976 = 12'h2b0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9904; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16048 = 12'h2b0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12976; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19120 = 12'h2b0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16048; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22192 = 12'h2b0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19120; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25264 = 12'h2b0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22192; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_688 = io_valid_in ? _GEN_25264 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_688 = 12'h2b0 == _T_2[11:0] ? image_688 : _GEN_687; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3761 = 12'h2b1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6833 = 12'h2b1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3761; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9905 = 12'h2b1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6833; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12977 = 12'h2b1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9905; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16049 = 12'h2b1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12977; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19121 = 12'h2b1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16049; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22193 = 12'h2b1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19121; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25265 = 12'h2b1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22193; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_689 = io_valid_in ? _GEN_25265 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_689 = 12'h2b1 == _T_2[11:0] ? image_689 : _GEN_688; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3762 = 12'h2b2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6834 = 12'h2b2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3762; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9906 = 12'h2b2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6834; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12978 = 12'h2b2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9906; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16050 = 12'h2b2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12978; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19122 = 12'h2b2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16050; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22194 = 12'h2b2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19122; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25266 = 12'h2b2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22194; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_690 = io_valid_in ? _GEN_25266 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_690 = 12'h2b2 == _T_2[11:0] ? image_690 : _GEN_689; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3763 = 12'h2b3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6835 = 12'h2b3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3763; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9907 = 12'h2b3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6835; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12979 = 12'h2b3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9907; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16051 = 12'h2b3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12979; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19123 = 12'h2b3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16051; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22195 = 12'h2b3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19123; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25267 = 12'h2b3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22195; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_691 = io_valid_in ? _GEN_25267 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_691 = 12'h2b3 == _T_2[11:0] ? image_691 : _GEN_690; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3764 = 12'h2b4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6836 = 12'h2b4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3764; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9908 = 12'h2b4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6836; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12980 = 12'h2b4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9908; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16052 = 12'h2b4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12980; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19124 = 12'h2b4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16052; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22196 = 12'h2b4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19124; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25268 = 12'h2b4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22196; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_692 = io_valid_in ? _GEN_25268 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_692 = 12'h2b4 == _T_2[11:0] ? image_692 : _GEN_691; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3765 = 12'h2b5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6837 = 12'h2b5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3765; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9909 = 12'h2b5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6837; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12981 = 12'h2b5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9909; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16053 = 12'h2b5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12981; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19125 = 12'h2b5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16053; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22197 = 12'h2b5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19125; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25269 = 12'h2b5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22197; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_693 = io_valid_in ? _GEN_25269 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_693 = 12'h2b5 == _T_2[11:0] ? image_693 : _GEN_692; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3766 = 12'h2b6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6838 = 12'h2b6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3766; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9910 = 12'h2b6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6838; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12982 = 12'h2b6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9910; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16054 = 12'h2b6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12982; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19126 = 12'h2b6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16054; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22198 = 12'h2b6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19126; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25270 = 12'h2b6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22198; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_694 = io_valid_in ? _GEN_25270 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_694 = 12'h2b6 == _T_2[11:0] ? image_694 : _GEN_693; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3767 = 12'h2b7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6839 = 12'h2b7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3767; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9911 = 12'h2b7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6839; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12983 = 12'h2b7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9911; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16055 = 12'h2b7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12983; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19127 = 12'h2b7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16055; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22199 = 12'h2b7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19127; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25271 = 12'h2b7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22199; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_695 = io_valid_in ? _GEN_25271 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_695 = 12'h2b7 == _T_2[11:0] ? image_695 : _GEN_694; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3768 = 12'h2b8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6840 = 12'h2b8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3768; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9912 = 12'h2b8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6840; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12984 = 12'h2b8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9912; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16056 = 12'h2b8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12984; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19128 = 12'h2b8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16056; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22200 = 12'h2b8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19128; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25272 = 12'h2b8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22200; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_696 = io_valid_in ? _GEN_25272 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_696 = 12'h2b8 == _T_2[11:0] ? image_696 : _GEN_695; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3769 = 12'h2b9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6841 = 12'h2b9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3769; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9913 = 12'h2b9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6841; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12985 = 12'h2b9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9913; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16057 = 12'h2b9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12985; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19129 = 12'h2b9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16057; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22201 = 12'h2b9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19129; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25273 = 12'h2b9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22201; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_697 = io_valid_in ? _GEN_25273 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_697 = 12'h2b9 == _T_2[11:0] ? image_697 : _GEN_696; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3770 = 12'h2ba == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6842 = 12'h2ba == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3770; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9914 = 12'h2ba == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6842; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12986 = 12'h2ba == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9914; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16058 = 12'h2ba == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12986; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19130 = 12'h2ba == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16058; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22202 = 12'h2ba == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19130; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25274 = 12'h2ba == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22202; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_698 = io_valid_in ? _GEN_25274 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_698 = 12'h2ba == _T_2[11:0] ? image_698 : _GEN_697; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3771 = 12'h2bb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6843 = 12'h2bb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3771; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9915 = 12'h2bb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6843; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12987 = 12'h2bb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9915; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16059 = 12'h2bb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12987; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19131 = 12'h2bb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16059; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22203 = 12'h2bb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19131; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25275 = 12'h2bb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22203; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_699 = io_valid_in ? _GEN_25275 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_699 = 12'h2bb == _T_2[11:0] ? image_699 : _GEN_698; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3772 = 12'h2bc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6844 = 12'h2bc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3772; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9916 = 12'h2bc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6844; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12988 = 12'h2bc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9916; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16060 = 12'h2bc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12988; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19132 = 12'h2bc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16060; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22204 = 12'h2bc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19132; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25276 = 12'h2bc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22204; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_700 = io_valid_in ? _GEN_25276 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_700 = 12'h2bc == _T_2[11:0] ? image_700 : _GEN_699; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3773 = 12'h2bd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6845 = 12'h2bd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3773; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9917 = 12'h2bd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6845; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12989 = 12'h2bd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9917; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16061 = 12'h2bd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12989; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19133 = 12'h2bd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16061; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22205 = 12'h2bd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19133; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25277 = 12'h2bd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22205; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_701 = io_valid_in ? _GEN_25277 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_701 = 12'h2bd == _T_2[11:0] ? image_701 : _GEN_700; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3774 = 12'h2be == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6846 = 12'h2be == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3774; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9918 = 12'h2be == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6846; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12990 = 12'h2be == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9918; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16062 = 12'h2be == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12990; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19134 = 12'h2be == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16062; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22206 = 12'h2be == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19134; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25278 = 12'h2be == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22206; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_702 = io_valid_in ? _GEN_25278 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_702 = 12'h2be == _T_2[11:0] ? image_702 : _GEN_701; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3775 = 12'h2bf == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6847 = 12'h2bf == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3775; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9919 = 12'h2bf == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6847; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12991 = 12'h2bf == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9919; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16063 = 12'h2bf == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12991; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19135 = 12'h2bf == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16063; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22207 = 12'h2bf == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19135; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25279 = 12'h2bf == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22207; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_703 = io_valid_in ? _GEN_25279 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_703 = 12'h2bf == _T_2[11:0] ? image_703 : _GEN_702; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3776 = 12'h2c0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6848 = 12'h2c0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3776; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9920 = 12'h2c0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6848; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12992 = 12'h2c0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9920; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16064 = 12'h2c0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12992; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19136 = 12'h2c0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16064; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22208 = 12'h2c0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19136; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25280 = 12'h2c0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22208; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_704 = io_valid_in ? _GEN_25280 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_704 = 12'h2c0 == _T_2[11:0] ? image_704 : _GEN_703; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3777 = 12'h2c1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6849 = 12'h2c1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3777; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9921 = 12'h2c1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6849; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12993 = 12'h2c1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9921; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16065 = 12'h2c1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12993; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19137 = 12'h2c1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16065; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22209 = 12'h2c1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19137; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25281 = 12'h2c1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22209; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_705 = io_valid_in ? _GEN_25281 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_705 = 12'h2c1 == _T_2[11:0] ? image_705 : _GEN_704; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3778 = 12'h2c2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6850 = 12'h2c2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3778; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9922 = 12'h2c2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6850; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12994 = 12'h2c2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9922; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16066 = 12'h2c2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12994; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19138 = 12'h2c2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16066; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22210 = 12'h2c2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19138; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25282 = 12'h2c2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22210; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_706 = io_valid_in ? _GEN_25282 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_706 = 12'h2c2 == _T_2[11:0] ? image_706 : _GEN_705; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3779 = 12'h2c3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6851 = 12'h2c3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3779; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9923 = 12'h2c3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6851; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12995 = 12'h2c3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9923; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16067 = 12'h2c3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12995; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19139 = 12'h2c3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16067; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22211 = 12'h2c3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19139; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25283 = 12'h2c3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22211; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_707 = io_valid_in ? _GEN_25283 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_707 = 12'h2c3 == _T_2[11:0] ? image_707 : _GEN_706; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3780 = 12'h2c4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6852 = 12'h2c4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3780; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9924 = 12'h2c4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6852; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12996 = 12'h2c4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9924; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16068 = 12'h2c4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12996; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19140 = 12'h2c4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16068; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22212 = 12'h2c4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19140; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25284 = 12'h2c4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22212; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_708 = io_valid_in ? _GEN_25284 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_708 = 12'h2c4 == _T_2[11:0] ? image_708 : _GEN_707; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3781 = 12'h2c5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6853 = 12'h2c5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3781; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9925 = 12'h2c5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6853; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12997 = 12'h2c5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9925; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16069 = 12'h2c5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12997; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19141 = 12'h2c5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16069; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22213 = 12'h2c5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19141; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25285 = 12'h2c5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22213; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_709 = io_valid_in ? _GEN_25285 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_709 = 12'h2c5 == _T_2[11:0] ? image_709 : _GEN_708; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3782 = 12'h2c6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6854 = 12'h2c6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3782; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9926 = 12'h2c6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6854; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12998 = 12'h2c6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9926; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16070 = 12'h2c6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12998; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19142 = 12'h2c6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16070; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22214 = 12'h2c6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19142; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25286 = 12'h2c6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22214; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_710 = io_valid_in ? _GEN_25286 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_710 = 12'h2c6 == _T_2[11:0] ? image_710 : _GEN_709; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3783 = 12'h2c7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6855 = 12'h2c7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3783; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9927 = 12'h2c7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6855; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12999 = 12'h2c7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9927; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16071 = 12'h2c7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_12999; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19143 = 12'h2c7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16071; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22215 = 12'h2c7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19143; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25287 = 12'h2c7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22215; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_711 = io_valid_in ? _GEN_25287 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_711 = 12'h2c7 == _T_2[11:0] ? image_711 : _GEN_710; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3784 = 12'h2c8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6856 = 12'h2c8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3784; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9928 = 12'h2c8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6856; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13000 = 12'h2c8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9928; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16072 = 12'h2c8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13000; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19144 = 12'h2c8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16072; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22216 = 12'h2c8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19144; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25288 = 12'h2c8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22216; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_712 = io_valid_in ? _GEN_25288 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_712 = 12'h2c8 == _T_2[11:0] ? image_712 : _GEN_711; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3785 = 12'h2c9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6857 = 12'h2c9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3785; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9929 = 12'h2c9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6857; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13001 = 12'h2c9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9929; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16073 = 12'h2c9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13001; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19145 = 12'h2c9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16073; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22217 = 12'h2c9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19145; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25289 = 12'h2c9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22217; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_713 = io_valid_in ? _GEN_25289 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_713 = 12'h2c9 == _T_2[11:0] ? image_713 : _GEN_712; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3786 = 12'h2ca == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6858 = 12'h2ca == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3786; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9930 = 12'h2ca == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6858; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13002 = 12'h2ca == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9930; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16074 = 12'h2ca == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13002; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19146 = 12'h2ca == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16074; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22218 = 12'h2ca == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19146; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25290 = 12'h2ca == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22218; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_714 = io_valid_in ? _GEN_25290 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_714 = 12'h2ca == _T_2[11:0] ? image_714 : _GEN_713; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3787 = 12'h2cb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6859 = 12'h2cb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3787; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9931 = 12'h2cb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6859; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13003 = 12'h2cb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9931; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16075 = 12'h2cb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13003; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19147 = 12'h2cb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16075; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22219 = 12'h2cb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19147; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25291 = 12'h2cb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22219; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_715 = io_valid_in ? _GEN_25291 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_715 = 12'h2cb == _T_2[11:0] ? image_715 : _GEN_714; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3788 = 12'h2cc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6860 = 12'h2cc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3788; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9932 = 12'h2cc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6860; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13004 = 12'h2cc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9932; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16076 = 12'h2cc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13004; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19148 = 12'h2cc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16076; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22220 = 12'h2cc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19148; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25292 = 12'h2cc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22220; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_716 = io_valid_in ? _GEN_25292 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_716 = 12'h2cc == _T_2[11:0] ? image_716 : _GEN_715; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3789 = 12'h2cd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6861 = 12'h2cd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3789; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9933 = 12'h2cd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6861; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13005 = 12'h2cd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9933; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16077 = 12'h2cd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13005; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19149 = 12'h2cd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16077; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22221 = 12'h2cd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19149; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25293 = 12'h2cd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22221; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_717 = io_valid_in ? _GEN_25293 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_717 = 12'h2cd == _T_2[11:0] ? image_717 : _GEN_716; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3790 = 12'h2ce == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6862 = 12'h2ce == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3790; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9934 = 12'h2ce == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6862; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13006 = 12'h2ce == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9934; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16078 = 12'h2ce == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13006; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19150 = 12'h2ce == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16078; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22222 = 12'h2ce == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19150; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25294 = 12'h2ce == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22222; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_718 = io_valid_in ? _GEN_25294 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_718 = 12'h2ce == _T_2[11:0] ? image_718 : _GEN_717; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3791 = 12'h2cf == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6863 = 12'h2cf == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3791; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9935 = 12'h2cf == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6863; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13007 = 12'h2cf == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9935; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16079 = 12'h2cf == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13007; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19151 = 12'h2cf == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16079; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22223 = 12'h2cf == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19151; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25295 = 12'h2cf == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22223; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_719 = io_valid_in ? _GEN_25295 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_719 = 12'h2cf == _T_2[11:0] ? image_719 : _GEN_718; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3792 = 12'h2d0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6864 = 12'h2d0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3792; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9936 = 12'h2d0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6864; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13008 = 12'h2d0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9936; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16080 = 12'h2d0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13008; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19152 = 12'h2d0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16080; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22224 = 12'h2d0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19152; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25296 = 12'h2d0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22224; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_720 = io_valid_in ? _GEN_25296 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_720 = 12'h2d0 == _T_2[11:0] ? image_720 : _GEN_719; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3793 = 12'h2d1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6865 = 12'h2d1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3793; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9937 = 12'h2d1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6865; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13009 = 12'h2d1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9937; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16081 = 12'h2d1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13009; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19153 = 12'h2d1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16081; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22225 = 12'h2d1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19153; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25297 = 12'h2d1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22225; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_721 = io_valid_in ? _GEN_25297 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_721 = 12'h2d1 == _T_2[11:0] ? image_721 : _GEN_720; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3794 = 12'h2d2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6866 = 12'h2d2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3794; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9938 = 12'h2d2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6866; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13010 = 12'h2d2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9938; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16082 = 12'h2d2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13010; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19154 = 12'h2d2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16082; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22226 = 12'h2d2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19154; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25298 = 12'h2d2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22226; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_722 = io_valid_in ? _GEN_25298 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_722 = 12'h2d2 == _T_2[11:0] ? image_722 : _GEN_721; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3795 = 12'h2d3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6867 = 12'h2d3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3795; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9939 = 12'h2d3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6867; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13011 = 12'h2d3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9939; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16083 = 12'h2d3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13011; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19155 = 12'h2d3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16083; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22227 = 12'h2d3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19155; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25299 = 12'h2d3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22227; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_723 = io_valid_in ? _GEN_25299 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_723 = 12'h2d3 == _T_2[11:0] ? image_723 : _GEN_722; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3796 = 12'h2d4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6868 = 12'h2d4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3796; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9940 = 12'h2d4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6868; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13012 = 12'h2d4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9940; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16084 = 12'h2d4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13012; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19156 = 12'h2d4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16084; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22228 = 12'h2d4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19156; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25300 = 12'h2d4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22228; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_724 = io_valid_in ? _GEN_25300 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_724 = 12'h2d4 == _T_2[11:0] ? image_724 : _GEN_723; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3797 = 12'h2d5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6869 = 12'h2d5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3797; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9941 = 12'h2d5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6869; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13013 = 12'h2d5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9941; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16085 = 12'h2d5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13013; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19157 = 12'h2d5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16085; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22229 = 12'h2d5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19157; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25301 = 12'h2d5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22229; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_725 = io_valid_in ? _GEN_25301 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_725 = 12'h2d5 == _T_2[11:0] ? image_725 : _GEN_724; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3798 = 12'h2d6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6870 = 12'h2d6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3798; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9942 = 12'h2d6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6870; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13014 = 12'h2d6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9942; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16086 = 12'h2d6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13014; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19158 = 12'h2d6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16086; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22230 = 12'h2d6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19158; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25302 = 12'h2d6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22230; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_726 = io_valid_in ? _GEN_25302 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_726 = 12'h2d6 == _T_2[11:0] ? image_726 : _GEN_725; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3799 = 12'h2d7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6871 = 12'h2d7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3799; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9943 = 12'h2d7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6871; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13015 = 12'h2d7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9943; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16087 = 12'h2d7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13015; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19159 = 12'h2d7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16087; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22231 = 12'h2d7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19159; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25303 = 12'h2d7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22231; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_727 = io_valid_in ? _GEN_25303 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_727 = 12'h2d7 == _T_2[11:0] ? image_727 : _GEN_726; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3800 = 12'h2d8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6872 = 12'h2d8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3800; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9944 = 12'h2d8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6872; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13016 = 12'h2d8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9944; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16088 = 12'h2d8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13016; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19160 = 12'h2d8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16088; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22232 = 12'h2d8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19160; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25304 = 12'h2d8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22232; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_728 = io_valid_in ? _GEN_25304 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_728 = 12'h2d8 == _T_2[11:0] ? image_728 : _GEN_727; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3801 = 12'h2d9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6873 = 12'h2d9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3801; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9945 = 12'h2d9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6873; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13017 = 12'h2d9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9945; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16089 = 12'h2d9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13017; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19161 = 12'h2d9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16089; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22233 = 12'h2d9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19161; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25305 = 12'h2d9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22233; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_729 = io_valid_in ? _GEN_25305 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_729 = 12'h2d9 == _T_2[11:0] ? image_729 : _GEN_728; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3802 = 12'h2da == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6874 = 12'h2da == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3802; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9946 = 12'h2da == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6874; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13018 = 12'h2da == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9946; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16090 = 12'h2da == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13018; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19162 = 12'h2da == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16090; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22234 = 12'h2da == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19162; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25306 = 12'h2da == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22234; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_730 = io_valid_in ? _GEN_25306 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_730 = 12'h2da == _T_2[11:0] ? image_730 : _GEN_729; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3803 = 12'h2db == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6875 = 12'h2db == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3803; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9947 = 12'h2db == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6875; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13019 = 12'h2db == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9947; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16091 = 12'h2db == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13019; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19163 = 12'h2db == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16091; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22235 = 12'h2db == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19163; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25307 = 12'h2db == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22235; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_731 = io_valid_in ? _GEN_25307 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_731 = 12'h2db == _T_2[11:0] ? image_731 : _GEN_730; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3804 = 12'h2dc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6876 = 12'h2dc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3804; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9948 = 12'h2dc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6876; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13020 = 12'h2dc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9948; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16092 = 12'h2dc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13020; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19164 = 12'h2dc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16092; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22236 = 12'h2dc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19164; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25308 = 12'h2dc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22236; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_732 = io_valid_in ? _GEN_25308 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_732 = 12'h2dc == _T_2[11:0] ? image_732 : _GEN_731; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3805 = 12'h2dd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6877 = 12'h2dd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3805; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9949 = 12'h2dd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6877; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13021 = 12'h2dd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9949; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16093 = 12'h2dd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13021; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19165 = 12'h2dd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16093; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22237 = 12'h2dd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19165; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25309 = 12'h2dd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22237; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_733 = io_valid_in ? _GEN_25309 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_733 = 12'h2dd == _T_2[11:0] ? image_733 : _GEN_732; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3806 = 12'h2de == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6878 = 12'h2de == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3806; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9950 = 12'h2de == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6878; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13022 = 12'h2de == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9950; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16094 = 12'h2de == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13022; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19166 = 12'h2de == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16094; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22238 = 12'h2de == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19166; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25310 = 12'h2de == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22238; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_734 = io_valid_in ? _GEN_25310 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_734 = 12'h2de == _T_2[11:0] ? image_734 : _GEN_733; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3807 = 12'h2df == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6879 = 12'h2df == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3807; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9951 = 12'h2df == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6879; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13023 = 12'h2df == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9951; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16095 = 12'h2df == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13023; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19167 = 12'h2df == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16095; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22239 = 12'h2df == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19167; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25311 = 12'h2df == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22239; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_735 = io_valid_in ? _GEN_25311 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_735 = 12'h2df == _T_2[11:0] ? image_735 : _GEN_734; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3808 = 12'h2e0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6880 = 12'h2e0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3808; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9952 = 12'h2e0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6880; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13024 = 12'h2e0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9952; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16096 = 12'h2e0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13024; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19168 = 12'h2e0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16096; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22240 = 12'h2e0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19168; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25312 = 12'h2e0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22240; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_736 = io_valid_in ? _GEN_25312 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_736 = 12'h2e0 == _T_2[11:0] ? image_736 : _GEN_735; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3809 = 12'h2e1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6881 = 12'h2e1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3809; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9953 = 12'h2e1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6881; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13025 = 12'h2e1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9953; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16097 = 12'h2e1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13025; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19169 = 12'h2e1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16097; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22241 = 12'h2e1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19169; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25313 = 12'h2e1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22241; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_737 = io_valid_in ? _GEN_25313 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_737 = 12'h2e1 == _T_2[11:0] ? image_737 : _GEN_736; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3810 = 12'h2e2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6882 = 12'h2e2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3810; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9954 = 12'h2e2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6882; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13026 = 12'h2e2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9954; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16098 = 12'h2e2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13026; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19170 = 12'h2e2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16098; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22242 = 12'h2e2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19170; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25314 = 12'h2e2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22242; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_738 = io_valid_in ? _GEN_25314 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_738 = 12'h2e2 == _T_2[11:0] ? image_738 : _GEN_737; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3811 = 12'h2e3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6883 = 12'h2e3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3811; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9955 = 12'h2e3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6883; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13027 = 12'h2e3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9955; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16099 = 12'h2e3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13027; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19171 = 12'h2e3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16099; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22243 = 12'h2e3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19171; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25315 = 12'h2e3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22243; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_739 = io_valid_in ? _GEN_25315 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_739 = 12'h2e3 == _T_2[11:0] ? image_739 : _GEN_738; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3812 = 12'h2e4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6884 = 12'h2e4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3812; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9956 = 12'h2e4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6884; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13028 = 12'h2e4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9956; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16100 = 12'h2e4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13028; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19172 = 12'h2e4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16100; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22244 = 12'h2e4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19172; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25316 = 12'h2e4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22244; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_740 = io_valid_in ? _GEN_25316 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_740 = 12'h2e4 == _T_2[11:0] ? image_740 : _GEN_739; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3813 = 12'h2e5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6885 = 12'h2e5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3813; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9957 = 12'h2e5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6885; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13029 = 12'h2e5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9957; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16101 = 12'h2e5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13029; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19173 = 12'h2e5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16101; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22245 = 12'h2e5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19173; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25317 = 12'h2e5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22245; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_741 = io_valid_in ? _GEN_25317 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_741 = 12'h2e5 == _T_2[11:0] ? image_741 : _GEN_740; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3814 = 12'h2e6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6886 = 12'h2e6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3814; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9958 = 12'h2e6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6886; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13030 = 12'h2e6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9958; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16102 = 12'h2e6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13030; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19174 = 12'h2e6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16102; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22246 = 12'h2e6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19174; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25318 = 12'h2e6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22246; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_742 = io_valid_in ? _GEN_25318 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_742 = 12'h2e6 == _T_2[11:0] ? image_742 : _GEN_741; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3815 = 12'h2e7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6887 = 12'h2e7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3815; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9959 = 12'h2e7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6887; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13031 = 12'h2e7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9959; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16103 = 12'h2e7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13031; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19175 = 12'h2e7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16103; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22247 = 12'h2e7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19175; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25319 = 12'h2e7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22247; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_743 = io_valid_in ? _GEN_25319 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_743 = 12'h2e7 == _T_2[11:0] ? image_743 : _GEN_742; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3816 = 12'h2e8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6888 = 12'h2e8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3816; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9960 = 12'h2e8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6888; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13032 = 12'h2e8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9960; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16104 = 12'h2e8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13032; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19176 = 12'h2e8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16104; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22248 = 12'h2e8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19176; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25320 = 12'h2e8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22248; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_744 = io_valid_in ? _GEN_25320 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_744 = 12'h2e8 == _T_2[11:0] ? image_744 : _GEN_743; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3817 = 12'h2e9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6889 = 12'h2e9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3817; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9961 = 12'h2e9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6889; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13033 = 12'h2e9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9961; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16105 = 12'h2e9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13033; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19177 = 12'h2e9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16105; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22249 = 12'h2e9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19177; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25321 = 12'h2e9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22249; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_745 = io_valid_in ? _GEN_25321 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_745 = 12'h2e9 == _T_2[11:0] ? image_745 : _GEN_744; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3818 = 12'h2ea == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6890 = 12'h2ea == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3818; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9962 = 12'h2ea == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6890; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13034 = 12'h2ea == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9962; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16106 = 12'h2ea == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13034; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19178 = 12'h2ea == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16106; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22250 = 12'h2ea == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19178; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25322 = 12'h2ea == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22250; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_746 = io_valid_in ? _GEN_25322 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_746 = 12'h2ea == _T_2[11:0] ? image_746 : _GEN_745; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3819 = 12'h2eb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6891 = 12'h2eb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3819; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9963 = 12'h2eb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6891; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13035 = 12'h2eb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9963; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16107 = 12'h2eb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13035; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19179 = 12'h2eb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16107; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22251 = 12'h2eb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19179; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25323 = 12'h2eb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22251; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_747 = io_valid_in ? _GEN_25323 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_747 = 12'h2eb == _T_2[11:0] ? image_747 : _GEN_746; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3820 = 12'h2ec == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6892 = 12'h2ec == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3820; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9964 = 12'h2ec == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6892; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13036 = 12'h2ec == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9964; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16108 = 12'h2ec == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13036; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19180 = 12'h2ec == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16108; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22252 = 12'h2ec == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19180; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25324 = 12'h2ec == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22252; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_748 = io_valid_in ? _GEN_25324 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_748 = 12'h2ec == _T_2[11:0] ? image_748 : _GEN_747; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3821 = 12'h2ed == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6893 = 12'h2ed == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3821; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9965 = 12'h2ed == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6893; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13037 = 12'h2ed == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9965; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16109 = 12'h2ed == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13037; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19181 = 12'h2ed == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16109; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22253 = 12'h2ed == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19181; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25325 = 12'h2ed == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22253; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_749 = io_valid_in ? _GEN_25325 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_749 = 12'h2ed == _T_2[11:0] ? image_749 : _GEN_748; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3822 = 12'h2ee == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6894 = 12'h2ee == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3822; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9966 = 12'h2ee == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6894; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13038 = 12'h2ee == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9966; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16110 = 12'h2ee == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13038; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19182 = 12'h2ee == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16110; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22254 = 12'h2ee == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19182; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25326 = 12'h2ee == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22254; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_750 = io_valid_in ? _GEN_25326 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_750 = 12'h2ee == _T_2[11:0] ? image_750 : _GEN_749; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3823 = 12'h2ef == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6895 = 12'h2ef == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3823; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9967 = 12'h2ef == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6895; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13039 = 12'h2ef == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9967; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16111 = 12'h2ef == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13039; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19183 = 12'h2ef == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16111; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22255 = 12'h2ef == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19183; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25327 = 12'h2ef == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22255; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_751 = io_valid_in ? _GEN_25327 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_751 = 12'h2ef == _T_2[11:0] ? image_751 : _GEN_750; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3824 = 12'h2f0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6896 = 12'h2f0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3824; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9968 = 12'h2f0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6896; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13040 = 12'h2f0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9968; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16112 = 12'h2f0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13040; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19184 = 12'h2f0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16112; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22256 = 12'h2f0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19184; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25328 = 12'h2f0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22256; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_752 = io_valid_in ? _GEN_25328 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_752 = 12'h2f0 == _T_2[11:0] ? image_752 : _GEN_751; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3825 = 12'h2f1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6897 = 12'h2f1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3825; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9969 = 12'h2f1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6897; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13041 = 12'h2f1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9969; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16113 = 12'h2f1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13041; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19185 = 12'h2f1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16113; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22257 = 12'h2f1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19185; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25329 = 12'h2f1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22257; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_753 = io_valid_in ? _GEN_25329 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_753 = 12'h2f1 == _T_2[11:0] ? image_753 : _GEN_752; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3826 = 12'h2f2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6898 = 12'h2f2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3826; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9970 = 12'h2f2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6898; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13042 = 12'h2f2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9970; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16114 = 12'h2f2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13042; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19186 = 12'h2f2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16114; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22258 = 12'h2f2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19186; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25330 = 12'h2f2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22258; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_754 = io_valid_in ? _GEN_25330 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_754 = 12'h2f2 == _T_2[11:0] ? image_754 : _GEN_753; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3827 = 12'h2f3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6899 = 12'h2f3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3827; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9971 = 12'h2f3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6899; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13043 = 12'h2f3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9971; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16115 = 12'h2f3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13043; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19187 = 12'h2f3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16115; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22259 = 12'h2f3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19187; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25331 = 12'h2f3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22259; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_755 = io_valid_in ? _GEN_25331 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_755 = 12'h2f3 == _T_2[11:0] ? image_755 : _GEN_754; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3828 = 12'h2f4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6900 = 12'h2f4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3828; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9972 = 12'h2f4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6900; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13044 = 12'h2f4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9972; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16116 = 12'h2f4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13044; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19188 = 12'h2f4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16116; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22260 = 12'h2f4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19188; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25332 = 12'h2f4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22260; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_756 = io_valid_in ? _GEN_25332 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_756 = 12'h2f4 == _T_2[11:0] ? image_756 : _GEN_755; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3829 = 12'h2f5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6901 = 12'h2f5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3829; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9973 = 12'h2f5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6901; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13045 = 12'h2f5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9973; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16117 = 12'h2f5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13045; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19189 = 12'h2f5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16117; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22261 = 12'h2f5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19189; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25333 = 12'h2f5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22261; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_757 = io_valid_in ? _GEN_25333 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_757 = 12'h2f5 == _T_2[11:0] ? image_757 : _GEN_756; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3830 = 12'h2f6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6902 = 12'h2f6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3830; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9974 = 12'h2f6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6902; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13046 = 12'h2f6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9974; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16118 = 12'h2f6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13046; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19190 = 12'h2f6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16118; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22262 = 12'h2f6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19190; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25334 = 12'h2f6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22262; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_758 = io_valid_in ? _GEN_25334 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_758 = 12'h2f6 == _T_2[11:0] ? image_758 : _GEN_757; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3831 = 12'h2f7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6903 = 12'h2f7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3831; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9975 = 12'h2f7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6903; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13047 = 12'h2f7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9975; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16119 = 12'h2f7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13047; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19191 = 12'h2f7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16119; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22263 = 12'h2f7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19191; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25335 = 12'h2f7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22263; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_759 = io_valid_in ? _GEN_25335 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_759 = 12'h2f7 == _T_2[11:0] ? image_759 : _GEN_758; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3832 = 12'h2f8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6904 = 12'h2f8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3832; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9976 = 12'h2f8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6904; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13048 = 12'h2f8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9976; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16120 = 12'h2f8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13048; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19192 = 12'h2f8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16120; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22264 = 12'h2f8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19192; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25336 = 12'h2f8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22264; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_760 = io_valid_in ? _GEN_25336 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_760 = 12'h2f8 == _T_2[11:0] ? image_760 : _GEN_759; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3833 = 12'h2f9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6905 = 12'h2f9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3833; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9977 = 12'h2f9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6905; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13049 = 12'h2f9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9977; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16121 = 12'h2f9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13049; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19193 = 12'h2f9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16121; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22265 = 12'h2f9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19193; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25337 = 12'h2f9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22265; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_761 = io_valid_in ? _GEN_25337 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_761 = 12'h2f9 == _T_2[11:0] ? image_761 : _GEN_760; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3834 = 12'h2fa == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6906 = 12'h2fa == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3834; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9978 = 12'h2fa == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6906; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13050 = 12'h2fa == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9978; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16122 = 12'h2fa == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13050; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19194 = 12'h2fa == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16122; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22266 = 12'h2fa == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19194; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25338 = 12'h2fa == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22266; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_762 = io_valid_in ? _GEN_25338 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_762 = 12'h2fa == _T_2[11:0] ? image_762 : _GEN_761; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3835 = 12'h2fb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6907 = 12'h2fb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3835; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9979 = 12'h2fb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6907; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13051 = 12'h2fb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9979; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16123 = 12'h2fb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13051; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19195 = 12'h2fb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16123; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22267 = 12'h2fb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19195; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25339 = 12'h2fb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22267; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_763 = io_valid_in ? _GEN_25339 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_763 = 12'h2fb == _T_2[11:0] ? image_763 : _GEN_762; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3836 = 12'h2fc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6908 = 12'h2fc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3836; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9980 = 12'h2fc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6908; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13052 = 12'h2fc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9980; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16124 = 12'h2fc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13052; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19196 = 12'h2fc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16124; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22268 = 12'h2fc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19196; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25340 = 12'h2fc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22268; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_764 = io_valid_in ? _GEN_25340 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_764 = 12'h2fc == _T_2[11:0] ? image_764 : _GEN_763; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3837 = 12'h2fd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6909 = 12'h2fd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3837; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9981 = 12'h2fd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6909; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13053 = 12'h2fd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9981; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16125 = 12'h2fd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13053; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19197 = 12'h2fd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16125; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22269 = 12'h2fd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19197; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25341 = 12'h2fd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22269; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_765 = io_valid_in ? _GEN_25341 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_765 = 12'h2fd == _T_2[11:0] ? image_765 : _GEN_764; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3838 = 12'h2fe == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6910 = 12'h2fe == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3838; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9982 = 12'h2fe == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6910; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13054 = 12'h2fe == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9982; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16126 = 12'h2fe == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13054; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19198 = 12'h2fe == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16126; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22270 = 12'h2fe == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19198; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25342 = 12'h2fe == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22270; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_766 = io_valid_in ? _GEN_25342 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_766 = 12'h2fe == _T_2[11:0] ? image_766 : _GEN_765; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3839 = 12'h2ff == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6911 = 12'h2ff == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3839; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9983 = 12'h2ff == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6911; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13055 = 12'h2ff == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9983; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16127 = 12'h2ff == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13055; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19199 = 12'h2ff == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16127; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22271 = 12'h2ff == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19199; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25343 = 12'h2ff == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22271; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_767 = io_valid_in ? _GEN_25343 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_767 = 12'h2ff == _T_2[11:0] ? image_767 : _GEN_766; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3840 = 12'h300 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6912 = 12'h300 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3840; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9984 = 12'h300 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6912; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13056 = 12'h300 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9984; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16128 = 12'h300 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13056; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19200 = 12'h300 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16128; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22272 = 12'h300 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19200; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25344 = 12'h300 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22272; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_768 = io_valid_in ? _GEN_25344 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_768 = 12'h300 == _T_2[11:0] ? image_768 : _GEN_767; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3841 = 12'h301 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6913 = 12'h301 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3841; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9985 = 12'h301 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6913; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13057 = 12'h301 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9985; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16129 = 12'h301 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13057; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19201 = 12'h301 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16129; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22273 = 12'h301 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19201; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25345 = 12'h301 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22273; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_769 = io_valid_in ? _GEN_25345 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_769 = 12'h301 == _T_2[11:0] ? image_769 : _GEN_768; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3842 = 12'h302 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6914 = 12'h302 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3842; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9986 = 12'h302 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6914; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13058 = 12'h302 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9986; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16130 = 12'h302 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13058; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19202 = 12'h302 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16130; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22274 = 12'h302 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19202; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25346 = 12'h302 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22274; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_770 = io_valid_in ? _GEN_25346 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_770 = 12'h302 == _T_2[11:0] ? image_770 : _GEN_769; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3843 = 12'h303 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6915 = 12'h303 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3843; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9987 = 12'h303 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6915; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13059 = 12'h303 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9987; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16131 = 12'h303 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13059; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19203 = 12'h303 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16131; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22275 = 12'h303 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19203; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25347 = 12'h303 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22275; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_771 = io_valid_in ? _GEN_25347 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_771 = 12'h303 == _T_2[11:0] ? image_771 : _GEN_770; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3844 = 12'h304 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6916 = 12'h304 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3844; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9988 = 12'h304 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6916; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13060 = 12'h304 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9988; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16132 = 12'h304 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13060; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19204 = 12'h304 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16132; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22276 = 12'h304 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19204; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25348 = 12'h304 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22276; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_772 = io_valid_in ? _GEN_25348 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_772 = 12'h304 == _T_2[11:0] ? image_772 : _GEN_771; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3845 = 12'h305 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6917 = 12'h305 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3845; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9989 = 12'h305 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6917; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13061 = 12'h305 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9989; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16133 = 12'h305 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13061; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19205 = 12'h305 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16133; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22277 = 12'h305 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19205; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25349 = 12'h305 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22277; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_773 = io_valid_in ? _GEN_25349 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_773 = 12'h305 == _T_2[11:0] ? image_773 : _GEN_772; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3846 = 12'h306 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6918 = 12'h306 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3846; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9990 = 12'h306 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6918; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13062 = 12'h306 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9990; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16134 = 12'h306 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13062; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19206 = 12'h306 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16134; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22278 = 12'h306 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19206; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25350 = 12'h306 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22278; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_774 = io_valid_in ? _GEN_25350 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_774 = 12'h306 == _T_2[11:0] ? image_774 : _GEN_773; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3847 = 12'h307 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6919 = 12'h307 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3847; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9991 = 12'h307 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6919; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13063 = 12'h307 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9991; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16135 = 12'h307 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13063; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19207 = 12'h307 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16135; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22279 = 12'h307 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19207; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25351 = 12'h307 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22279; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_775 = io_valid_in ? _GEN_25351 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_775 = 12'h307 == _T_2[11:0] ? image_775 : _GEN_774; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3848 = 12'h308 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6920 = 12'h308 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3848; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9992 = 12'h308 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6920; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13064 = 12'h308 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9992; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16136 = 12'h308 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13064; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19208 = 12'h308 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16136; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22280 = 12'h308 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19208; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25352 = 12'h308 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22280; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_776 = io_valid_in ? _GEN_25352 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_776 = 12'h308 == _T_2[11:0] ? image_776 : _GEN_775; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3849 = 12'h309 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6921 = 12'h309 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3849; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9993 = 12'h309 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6921; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13065 = 12'h309 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9993; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16137 = 12'h309 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13065; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19209 = 12'h309 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16137; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22281 = 12'h309 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19209; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25353 = 12'h309 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22281; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_777 = io_valid_in ? _GEN_25353 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_777 = 12'h309 == _T_2[11:0] ? image_777 : _GEN_776; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3850 = 12'h30a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6922 = 12'h30a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3850; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9994 = 12'h30a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6922; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13066 = 12'h30a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9994; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16138 = 12'h30a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13066; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19210 = 12'h30a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16138; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22282 = 12'h30a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19210; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25354 = 12'h30a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22282; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_778 = io_valid_in ? _GEN_25354 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_778 = 12'h30a == _T_2[11:0] ? image_778 : _GEN_777; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3851 = 12'h30b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6923 = 12'h30b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3851; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9995 = 12'h30b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6923; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13067 = 12'h30b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9995; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16139 = 12'h30b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13067; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19211 = 12'h30b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16139; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22283 = 12'h30b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19211; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25355 = 12'h30b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22283; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_779 = io_valid_in ? _GEN_25355 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_779 = 12'h30b == _T_2[11:0] ? image_779 : _GEN_778; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3852 = 12'h30c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6924 = 12'h30c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3852; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9996 = 12'h30c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6924; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13068 = 12'h30c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9996; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16140 = 12'h30c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13068; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19212 = 12'h30c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16140; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22284 = 12'h30c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19212; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25356 = 12'h30c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22284; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_780 = io_valid_in ? _GEN_25356 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_780 = 12'h30c == _T_2[11:0] ? image_780 : _GEN_779; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3853 = 12'h30d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6925 = 12'h30d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3853; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9997 = 12'h30d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6925; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13069 = 12'h30d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9997; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16141 = 12'h30d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13069; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19213 = 12'h30d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16141; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22285 = 12'h30d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19213; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25357 = 12'h30d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22285; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_781 = io_valid_in ? _GEN_25357 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_781 = 12'h30d == _T_2[11:0] ? image_781 : _GEN_780; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3854 = 12'h30e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6926 = 12'h30e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3854; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9998 = 12'h30e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6926; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13070 = 12'h30e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9998; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16142 = 12'h30e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13070; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19214 = 12'h30e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16142; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22286 = 12'h30e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19214; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25358 = 12'h30e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22286; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_782 = io_valid_in ? _GEN_25358 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_782 = 12'h30e == _T_2[11:0] ? image_782 : _GEN_781; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3855 = 12'h30f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6927 = 12'h30f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3855; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9999 = 12'h30f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6927; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13071 = 12'h30f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_9999; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16143 = 12'h30f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13071; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19215 = 12'h30f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16143; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22287 = 12'h30f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19215; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25359 = 12'h30f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22287; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_783 = io_valid_in ? _GEN_25359 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_783 = 12'h30f == _T_2[11:0] ? image_783 : _GEN_782; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3856 = 12'h310 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6928 = 12'h310 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3856; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10000 = 12'h310 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6928; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13072 = 12'h310 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10000; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16144 = 12'h310 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13072; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19216 = 12'h310 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16144; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22288 = 12'h310 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19216; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25360 = 12'h310 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22288; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_784 = io_valid_in ? _GEN_25360 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_784 = 12'h310 == _T_2[11:0] ? image_784 : _GEN_783; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3857 = 12'h311 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6929 = 12'h311 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3857; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10001 = 12'h311 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6929; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13073 = 12'h311 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10001; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16145 = 12'h311 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13073; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19217 = 12'h311 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16145; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22289 = 12'h311 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19217; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25361 = 12'h311 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22289; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_785 = io_valid_in ? _GEN_25361 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_785 = 12'h311 == _T_2[11:0] ? image_785 : _GEN_784; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3858 = 12'h312 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6930 = 12'h312 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3858; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10002 = 12'h312 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6930; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13074 = 12'h312 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10002; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16146 = 12'h312 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13074; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19218 = 12'h312 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16146; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22290 = 12'h312 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19218; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25362 = 12'h312 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22290; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_786 = io_valid_in ? _GEN_25362 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_786 = 12'h312 == _T_2[11:0] ? image_786 : _GEN_785; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3859 = 12'h313 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6931 = 12'h313 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3859; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10003 = 12'h313 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6931; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13075 = 12'h313 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10003; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16147 = 12'h313 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13075; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19219 = 12'h313 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16147; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22291 = 12'h313 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19219; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25363 = 12'h313 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22291; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_787 = io_valid_in ? _GEN_25363 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_787 = 12'h313 == _T_2[11:0] ? image_787 : _GEN_786; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3860 = 12'h314 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6932 = 12'h314 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3860; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10004 = 12'h314 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6932; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13076 = 12'h314 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10004; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16148 = 12'h314 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13076; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19220 = 12'h314 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16148; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22292 = 12'h314 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19220; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25364 = 12'h314 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22292; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_788 = io_valid_in ? _GEN_25364 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_788 = 12'h314 == _T_2[11:0] ? image_788 : _GEN_787; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3861 = 12'h315 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6933 = 12'h315 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3861; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10005 = 12'h315 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6933; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13077 = 12'h315 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10005; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16149 = 12'h315 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13077; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19221 = 12'h315 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16149; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22293 = 12'h315 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19221; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25365 = 12'h315 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22293; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_789 = io_valid_in ? _GEN_25365 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_789 = 12'h315 == _T_2[11:0] ? image_789 : _GEN_788; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3862 = 12'h316 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6934 = 12'h316 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3862; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10006 = 12'h316 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6934; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13078 = 12'h316 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10006; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16150 = 12'h316 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13078; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19222 = 12'h316 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16150; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22294 = 12'h316 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19222; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25366 = 12'h316 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22294; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_790 = io_valid_in ? _GEN_25366 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_790 = 12'h316 == _T_2[11:0] ? image_790 : _GEN_789; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3863 = 12'h317 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6935 = 12'h317 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3863; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10007 = 12'h317 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6935; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13079 = 12'h317 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10007; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16151 = 12'h317 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13079; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19223 = 12'h317 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16151; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22295 = 12'h317 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19223; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25367 = 12'h317 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22295; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_791 = io_valid_in ? _GEN_25367 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_791 = 12'h317 == _T_2[11:0] ? image_791 : _GEN_790; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3864 = 12'h318 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6936 = 12'h318 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3864; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10008 = 12'h318 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6936; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13080 = 12'h318 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10008; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16152 = 12'h318 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13080; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19224 = 12'h318 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16152; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22296 = 12'h318 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19224; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25368 = 12'h318 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22296; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_792 = io_valid_in ? _GEN_25368 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_792 = 12'h318 == _T_2[11:0] ? image_792 : _GEN_791; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3865 = 12'h319 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6937 = 12'h319 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3865; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10009 = 12'h319 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6937; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13081 = 12'h319 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10009; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16153 = 12'h319 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13081; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19225 = 12'h319 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16153; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22297 = 12'h319 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19225; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25369 = 12'h319 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22297; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_793 = io_valid_in ? _GEN_25369 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_793 = 12'h319 == _T_2[11:0] ? image_793 : _GEN_792; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3866 = 12'h31a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6938 = 12'h31a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3866; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10010 = 12'h31a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6938; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13082 = 12'h31a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10010; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16154 = 12'h31a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13082; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19226 = 12'h31a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16154; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22298 = 12'h31a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19226; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25370 = 12'h31a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22298; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_794 = io_valid_in ? _GEN_25370 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_794 = 12'h31a == _T_2[11:0] ? image_794 : _GEN_793; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3867 = 12'h31b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6939 = 12'h31b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3867; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10011 = 12'h31b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6939; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13083 = 12'h31b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10011; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16155 = 12'h31b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13083; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19227 = 12'h31b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16155; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22299 = 12'h31b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19227; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25371 = 12'h31b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22299; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_795 = io_valid_in ? _GEN_25371 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_795 = 12'h31b == _T_2[11:0] ? image_795 : _GEN_794; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3868 = 12'h31c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6940 = 12'h31c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3868; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10012 = 12'h31c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6940; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13084 = 12'h31c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10012; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16156 = 12'h31c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13084; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19228 = 12'h31c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16156; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22300 = 12'h31c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19228; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25372 = 12'h31c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22300; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_796 = io_valid_in ? _GEN_25372 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_796 = 12'h31c == _T_2[11:0] ? image_796 : _GEN_795; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3869 = 12'h31d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6941 = 12'h31d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3869; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10013 = 12'h31d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6941; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13085 = 12'h31d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10013; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16157 = 12'h31d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13085; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19229 = 12'h31d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16157; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22301 = 12'h31d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19229; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25373 = 12'h31d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22301; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_797 = io_valid_in ? _GEN_25373 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_797 = 12'h31d == _T_2[11:0] ? image_797 : _GEN_796; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3870 = 12'h31e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6942 = 12'h31e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3870; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10014 = 12'h31e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6942; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13086 = 12'h31e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10014; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16158 = 12'h31e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13086; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19230 = 12'h31e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16158; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22302 = 12'h31e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19230; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25374 = 12'h31e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22302; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_798 = io_valid_in ? _GEN_25374 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_798 = 12'h31e == _T_2[11:0] ? image_798 : _GEN_797; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3871 = 12'h31f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6943 = 12'h31f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3871; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10015 = 12'h31f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6943; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13087 = 12'h31f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10015; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16159 = 12'h31f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13087; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19231 = 12'h31f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16159; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22303 = 12'h31f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19231; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25375 = 12'h31f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22303; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_799 = io_valid_in ? _GEN_25375 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_799 = 12'h31f == _T_2[11:0] ? image_799 : _GEN_798; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3872 = 12'h320 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6944 = 12'h320 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3872; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10016 = 12'h320 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6944; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13088 = 12'h320 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10016; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16160 = 12'h320 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13088; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19232 = 12'h320 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16160; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22304 = 12'h320 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19232; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25376 = 12'h320 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22304; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_800 = io_valid_in ? _GEN_25376 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_800 = 12'h320 == _T_2[11:0] ? image_800 : _GEN_799; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3873 = 12'h321 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6945 = 12'h321 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3873; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10017 = 12'h321 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6945; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13089 = 12'h321 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10017; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16161 = 12'h321 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13089; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19233 = 12'h321 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16161; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22305 = 12'h321 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19233; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25377 = 12'h321 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22305; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_801 = io_valid_in ? _GEN_25377 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_801 = 12'h321 == _T_2[11:0] ? image_801 : _GEN_800; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3874 = 12'h322 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6946 = 12'h322 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3874; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10018 = 12'h322 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6946; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13090 = 12'h322 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10018; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16162 = 12'h322 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13090; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19234 = 12'h322 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16162; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22306 = 12'h322 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19234; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25378 = 12'h322 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22306; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_802 = io_valid_in ? _GEN_25378 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_802 = 12'h322 == _T_2[11:0] ? image_802 : _GEN_801; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3875 = 12'h323 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6947 = 12'h323 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3875; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10019 = 12'h323 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6947; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13091 = 12'h323 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10019; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16163 = 12'h323 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13091; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19235 = 12'h323 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16163; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22307 = 12'h323 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19235; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25379 = 12'h323 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22307; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_803 = io_valid_in ? _GEN_25379 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_803 = 12'h323 == _T_2[11:0] ? image_803 : _GEN_802; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3876 = 12'h324 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6948 = 12'h324 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3876; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10020 = 12'h324 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6948; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13092 = 12'h324 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10020; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16164 = 12'h324 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13092; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19236 = 12'h324 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16164; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22308 = 12'h324 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19236; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25380 = 12'h324 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22308; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_804 = io_valid_in ? _GEN_25380 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_804 = 12'h324 == _T_2[11:0] ? image_804 : _GEN_803; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3877 = 12'h325 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6949 = 12'h325 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3877; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10021 = 12'h325 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6949; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13093 = 12'h325 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10021; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16165 = 12'h325 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13093; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19237 = 12'h325 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16165; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22309 = 12'h325 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19237; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25381 = 12'h325 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22309; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_805 = io_valid_in ? _GEN_25381 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_805 = 12'h325 == _T_2[11:0] ? image_805 : _GEN_804; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3878 = 12'h326 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6950 = 12'h326 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3878; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10022 = 12'h326 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6950; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13094 = 12'h326 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10022; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16166 = 12'h326 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13094; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19238 = 12'h326 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16166; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22310 = 12'h326 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19238; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25382 = 12'h326 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22310; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_806 = io_valid_in ? _GEN_25382 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_806 = 12'h326 == _T_2[11:0] ? image_806 : _GEN_805; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3879 = 12'h327 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6951 = 12'h327 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3879; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10023 = 12'h327 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6951; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13095 = 12'h327 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10023; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16167 = 12'h327 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13095; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19239 = 12'h327 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16167; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22311 = 12'h327 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19239; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25383 = 12'h327 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22311; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_807 = io_valid_in ? _GEN_25383 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_807 = 12'h327 == _T_2[11:0] ? image_807 : _GEN_806; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3880 = 12'h328 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6952 = 12'h328 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3880; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10024 = 12'h328 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6952; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13096 = 12'h328 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10024; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16168 = 12'h328 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13096; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19240 = 12'h328 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16168; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22312 = 12'h328 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19240; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25384 = 12'h328 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22312; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_808 = io_valid_in ? _GEN_25384 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_808 = 12'h328 == _T_2[11:0] ? image_808 : _GEN_807; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3881 = 12'h329 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6953 = 12'h329 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3881; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10025 = 12'h329 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6953; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13097 = 12'h329 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10025; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16169 = 12'h329 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13097; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19241 = 12'h329 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16169; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22313 = 12'h329 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19241; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25385 = 12'h329 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22313; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_809 = io_valid_in ? _GEN_25385 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_809 = 12'h329 == _T_2[11:0] ? image_809 : _GEN_808; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3882 = 12'h32a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6954 = 12'h32a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3882; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10026 = 12'h32a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6954; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13098 = 12'h32a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10026; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16170 = 12'h32a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13098; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19242 = 12'h32a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16170; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22314 = 12'h32a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19242; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25386 = 12'h32a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22314; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_810 = io_valid_in ? _GEN_25386 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_810 = 12'h32a == _T_2[11:0] ? image_810 : _GEN_809; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3883 = 12'h32b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6955 = 12'h32b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3883; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10027 = 12'h32b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6955; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13099 = 12'h32b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10027; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16171 = 12'h32b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13099; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19243 = 12'h32b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16171; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22315 = 12'h32b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19243; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25387 = 12'h32b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22315; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_811 = io_valid_in ? _GEN_25387 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_811 = 12'h32b == _T_2[11:0] ? image_811 : _GEN_810; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3884 = 12'h32c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6956 = 12'h32c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3884; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10028 = 12'h32c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6956; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13100 = 12'h32c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10028; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16172 = 12'h32c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13100; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19244 = 12'h32c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16172; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22316 = 12'h32c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19244; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25388 = 12'h32c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22316; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_812 = io_valid_in ? _GEN_25388 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_812 = 12'h32c == _T_2[11:0] ? image_812 : _GEN_811; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3885 = 12'h32d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6957 = 12'h32d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3885; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10029 = 12'h32d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6957; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13101 = 12'h32d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10029; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16173 = 12'h32d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13101; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19245 = 12'h32d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16173; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22317 = 12'h32d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19245; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25389 = 12'h32d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22317; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_813 = io_valid_in ? _GEN_25389 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_813 = 12'h32d == _T_2[11:0] ? image_813 : _GEN_812; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3886 = 12'h32e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6958 = 12'h32e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3886; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10030 = 12'h32e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6958; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13102 = 12'h32e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10030; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16174 = 12'h32e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13102; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19246 = 12'h32e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16174; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22318 = 12'h32e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19246; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25390 = 12'h32e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22318; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_814 = io_valid_in ? _GEN_25390 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_814 = 12'h32e == _T_2[11:0] ? image_814 : _GEN_813; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3887 = 12'h32f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6959 = 12'h32f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3887; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10031 = 12'h32f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6959; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13103 = 12'h32f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10031; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16175 = 12'h32f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13103; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19247 = 12'h32f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16175; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22319 = 12'h32f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19247; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25391 = 12'h32f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22319; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_815 = io_valid_in ? _GEN_25391 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_815 = 12'h32f == _T_2[11:0] ? image_815 : _GEN_814; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3888 = 12'h330 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6960 = 12'h330 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3888; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10032 = 12'h330 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6960; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13104 = 12'h330 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10032; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16176 = 12'h330 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13104; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19248 = 12'h330 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16176; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22320 = 12'h330 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19248; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25392 = 12'h330 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22320; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_816 = io_valid_in ? _GEN_25392 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_816 = 12'h330 == _T_2[11:0] ? image_816 : _GEN_815; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3889 = 12'h331 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6961 = 12'h331 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3889; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10033 = 12'h331 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6961; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13105 = 12'h331 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10033; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16177 = 12'h331 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13105; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19249 = 12'h331 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16177; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22321 = 12'h331 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19249; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25393 = 12'h331 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22321; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_817 = io_valid_in ? _GEN_25393 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_817 = 12'h331 == _T_2[11:0] ? image_817 : _GEN_816; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3890 = 12'h332 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6962 = 12'h332 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3890; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10034 = 12'h332 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6962; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13106 = 12'h332 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10034; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16178 = 12'h332 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13106; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19250 = 12'h332 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16178; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22322 = 12'h332 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19250; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25394 = 12'h332 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22322; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_818 = io_valid_in ? _GEN_25394 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_818 = 12'h332 == _T_2[11:0] ? image_818 : _GEN_817; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3891 = 12'h333 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6963 = 12'h333 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3891; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10035 = 12'h333 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6963; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13107 = 12'h333 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10035; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16179 = 12'h333 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13107; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19251 = 12'h333 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16179; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22323 = 12'h333 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19251; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25395 = 12'h333 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22323; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_819 = io_valid_in ? _GEN_25395 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_819 = 12'h333 == _T_2[11:0] ? image_819 : _GEN_818; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3892 = 12'h334 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6964 = 12'h334 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3892; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10036 = 12'h334 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6964; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13108 = 12'h334 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10036; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16180 = 12'h334 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13108; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19252 = 12'h334 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16180; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22324 = 12'h334 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19252; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25396 = 12'h334 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22324; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_820 = io_valid_in ? _GEN_25396 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_820 = 12'h334 == _T_2[11:0] ? image_820 : _GEN_819; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3893 = 12'h335 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6965 = 12'h335 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3893; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10037 = 12'h335 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6965; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13109 = 12'h335 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10037; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16181 = 12'h335 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13109; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19253 = 12'h335 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16181; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22325 = 12'h335 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19253; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25397 = 12'h335 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22325; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_821 = io_valid_in ? _GEN_25397 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_821 = 12'h335 == _T_2[11:0] ? image_821 : _GEN_820; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3894 = 12'h336 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6966 = 12'h336 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3894; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10038 = 12'h336 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6966; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13110 = 12'h336 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10038; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16182 = 12'h336 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13110; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19254 = 12'h336 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16182; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22326 = 12'h336 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19254; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25398 = 12'h336 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22326; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_822 = io_valid_in ? _GEN_25398 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_822 = 12'h336 == _T_2[11:0] ? image_822 : _GEN_821; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3895 = 12'h337 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6967 = 12'h337 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3895; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10039 = 12'h337 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6967; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13111 = 12'h337 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10039; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16183 = 12'h337 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13111; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19255 = 12'h337 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16183; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22327 = 12'h337 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19255; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25399 = 12'h337 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22327; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_823 = io_valid_in ? _GEN_25399 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_823 = 12'h337 == _T_2[11:0] ? image_823 : _GEN_822; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3896 = 12'h338 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6968 = 12'h338 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3896; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10040 = 12'h338 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6968; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13112 = 12'h338 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10040; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16184 = 12'h338 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13112; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19256 = 12'h338 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16184; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22328 = 12'h338 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19256; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25400 = 12'h338 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22328; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_824 = io_valid_in ? _GEN_25400 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_824 = 12'h338 == _T_2[11:0] ? image_824 : _GEN_823; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3897 = 12'h339 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6969 = 12'h339 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3897; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10041 = 12'h339 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6969; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13113 = 12'h339 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10041; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16185 = 12'h339 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13113; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19257 = 12'h339 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16185; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22329 = 12'h339 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19257; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25401 = 12'h339 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22329; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_825 = io_valid_in ? _GEN_25401 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_825 = 12'h339 == _T_2[11:0] ? image_825 : _GEN_824; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3898 = 12'h33a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6970 = 12'h33a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3898; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10042 = 12'h33a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6970; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13114 = 12'h33a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10042; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16186 = 12'h33a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13114; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19258 = 12'h33a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16186; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22330 = 12'h33a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19258; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25402 = 12'h33a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22330; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_826 = io_valid_in ? _GEN_25402 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_826 = 12'h33a == _T_2[11:0] ? image_826 : _GEN_825; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3899 = 12'h33b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6971 = 12'h33b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3899; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10043 = 12'h33b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6971; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13115 = 12'h33b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10043; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16187 = 12'h33b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13115; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19259 = 12'h33b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16187; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22331 = 12'h33b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19259; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25403 = 12'h33b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22331; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_827 = io_valid_in ? _GEN_25403 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_827 = 12'h33b == _T_2[11:0] ? image_827 : _GEN_826; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3900 = 12'h33c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6972 = 12'h33c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3900; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10044 = 12'h33c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6972; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13116 = 12'h33c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10044; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16188 = 12'h33c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13116; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19260 = 12'h33c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16188; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22332 = 12'h33c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19260; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25404 = 12'h33c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22332; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_828 = io_valid_in ? _GEN_25404 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_828 = 12'h33c == _T_2[11:0] ? image_828 : _GEN_827; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3901 = 12'h33d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6973 = 12'h33d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3901; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10045 = 12'h33d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6973; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13117 = 12'h33d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10045; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16189 = 12'h33d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13117; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19261 = 12'h33d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16189; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22333 = 12'h33d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19261; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25405 = 12'h33d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22333; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_829 = io_valid_in ? _GEN_25405 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_829 = 12'h33d == _T_2[11:0] ? image_829 : _GEN_828; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3902 = 12'h33e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6974 = 12'h33e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3902; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10046 = 12'h33e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6974; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13118 = 12'h33e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10046; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16190 = 12'h33e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13118; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19262 = 12'h33e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16190; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22334 = 12'h33e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19262; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25406 = 12'h33e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22334; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_830 = io_valid_in ? _GEN_25406 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_830 = 12'h33e == _T_2[11:0] ? image_830 : _GEN_829; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3903 = 12'h33f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6975 = 12'h33f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3903; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10047 = 12'h33f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6975; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13119 = 12'h33f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10047; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16191 = 12'h33f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13119; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19263 = 12'h33f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16191; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22335 = 12'h33f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19263; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25407 = 12'h33f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22335; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_831 = io_valid_in ? _GEN_25407 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_831 = 12'h33f == _T_2[11:0] ? image_831 : _GEN_830; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3904 = 12'h340 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6976 = 12'h340 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3904; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10048 = 12'h340 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6976; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13120 = 12'h340 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10048; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16192 = 12'h340 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13120; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19264 = 12'h340 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16192; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22336 = 12'h340 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19264; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25408 = 12'h340 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22336; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_832 = io_valid_in ? _GEN_25408 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_832 = 12'h340 == _T_2[11:0] ? image_832 : _GEN_831; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3905 = 12'h341 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6977 = 12'h341 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3905; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10049 = 12'h341 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6977; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13121 = 12'h341 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10049; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16193 = 12'h341 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13121; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19265 = 12'h341 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16193; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22337 = 12'h341 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19265; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25409 = 12'h341 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22337; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_833 = io_valid_in ? _GEN_25409 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_833 = 12'h341 == _T_2[11:0] ? image_833 : _GEN_832; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3906 = 12'h342 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6978 = 12'h342 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3906; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10050 = 12'h342 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6978; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13122 = 12'h342 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10050; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16194 = 12'h342 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13122; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19266 = 12'h342 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16194; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22338 = 12'h342 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19266; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25410 = 12'h342 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22338; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_834 = io_valid_in ? _GEN_25410 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_834 = 12'h342 == _T_2[11:0] ? image_834 : _GEN_833; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3907 = 12'h343 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6979 = 12'h343 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3907; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10051 = 12'h343 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6979; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13123 = 12'h343 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10051; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16195 = 12'h343 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13123; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19267 = 12'h343 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16195; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22339 = 12'h343 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19267; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25411 = 12'h343 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22339; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_835 = io_valid_in ? _GEN_25411 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_835 = 12'h343 == _T_2[11:0] ? image_835 : _GEN_834; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3908 = 12'h344 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6980 = 12'h344 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3908; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10052 = 12'h344 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6980; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13124 = 12'h344 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10052; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16196 = 12'h344 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13124; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19268 = 12'h344 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16196; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22340 = 12'h344 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19268; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25412 = 12'h344 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22340; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_836 = io_valid_in ? _GEN_25412 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_836 = 12'h344 == _T_2[11:0] ? image_836 : _GEN_835; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3909 = 12'h345 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6981 = 12'h345 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3909; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10053 = 12'h345 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6981; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13125 = 12'h345 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10053; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16197 = 12'h345 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13125; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19269 = 12'h345 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16197; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22341 = 12'h345 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19269; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25413 = 12'h345 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22341; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_837 = io_valid_in ? _GEN_25413 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_837 = 12'h345 == _T_2[11:0] ? image_837 : _GEN_836; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3910 = 12'h346 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6982 = 12'h346 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3910; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10054 = 12'h346 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6982; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13126 = 12'h346 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10054; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16198 = 12'h346 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13126; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19270 = 12'h346 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16198; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22342 = 12'h346 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19270; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25414 = 12'h346 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22342; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_838 = io_valid_in ? _GEN_25414 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_838 = 12'h346 == _T_2[11:0] ? image_838 : _GEN_837; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3911 = 12'h347 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6983 = 12'h347 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3911; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10055 = 12'h347 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6983; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13127 = 12'h347 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10055; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16199 = 12'h347 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13127; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19271 = 12'h347 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16199; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22343 = 12'h347 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19271; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25415 = 12'h347 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22343; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_839 = io_valid_in ? _GEN_25415 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_839 = 12'h347 == _T_2[11:0] ? image_839 : _GEN_838; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3912 = 12'h348 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6984 = 12'h348 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3912; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10056 = 12'h348 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6984; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13128 = 12'h348 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10056; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16200 = 12'h348 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13128; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19272 = 12'h348 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16200; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22344 = 12'h348 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19272; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25416 = 12'h348 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22344; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_840 = io_valid_in ? _GEN_25416 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_840 = 12'h348 == _T_2[11:0] ? image_840 : _GEN_839; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3913 = 12'h349 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6985 = 12'h349 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3913; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10057 = 12'h349 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6985; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13129 = 12'h349 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10057; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16201 = 12'h349 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13129; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19273 = 12'h349 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16201; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22345 = 12'h349 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19273; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25417 = 12'h349 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22345; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_841 = io_valid_in ? _GEN_25417 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_841 = 12'h349 == _T_2[11:0] ? image_841 : _GEN_840; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3914 = 12'h34a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6986 = 12'h34a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3914; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10058 = 12'h34a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6986; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13130 = 12'h34a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10058; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16202 = 12'h34a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13130; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19274 = 12'h34a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16202; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22346 = 12'h34a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19274; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25418 = 12'h34a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22346; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_842 = io_valid_in ? _GEN_25418 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_842 = 12'h34a == _T_2[11:0] ? image_842 : _GEN_841; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3915 = 12'h34b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6987 = 12'h34b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3915; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10059 = 12'h34b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6987; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13131 = 12'h34b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10059; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16203 = 12'h34b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13131; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19275 = 12'h34b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16203; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22347 = 12'h34b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19275; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25419 = 12'h34b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22347; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_843 = io_valid_in ? _GEN_25419 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_843 = 12'h34b == _T_2[11:0] ? image_843 : _GEN_842; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3916 = 12'h34c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6988 = 12'h34c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3916; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10060 = 12'h34c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6988; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13132 = 12'h34c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10060; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16204 = 12'h34c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13132; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19276 = 12'h34c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16204; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22348 = 12'h34c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19276; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25420 = 12'h34c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22348; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_844 = io_valid_in ? _GEN_25420 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_844 = 12'h34c == _T_2[11:0] ? image_844 : _GEN_843; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3917 = 12'h34d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6989 = 12'h34d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3917; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10061 = 12'h34d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6989; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13133 = 12'h34d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10061; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16205 = 12'h34d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13133; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19277 = 12'h34d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16205; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22349 = 12'h34d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19277; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25421 = 12'h34d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22349; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_845 = io_valid_in ? _GEN_25421 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_845 = 12'h34d == _T_2[11:0] ? image_845 : _GEN_844; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3918 = 12'h34e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6990 = 12'h34e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3918; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10062 = 12'h34e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6990; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13134 = 12'h34e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10062; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16206 = 12'h34e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13134; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19278 = 12'h34e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16206; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22350 = 12'h34e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19278; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25422 = 12'h34e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22350; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_846 = io_valid_in ? _GEN_25422 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_846 = 12'h34e == _T_2[11:0] ? image_846 : _GEN_845; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3919 = 12'h34f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6991 = 12'h34f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3919; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10063 = 12'h34f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6991; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13135 = 12'h34f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10063; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16207 = 12'h34f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13135; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19279 = 12'h34f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16207; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22351 = 12'h34f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19279; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25423 = 12'h34f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22351; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_847 = io_valid_in ? _GEN_25423 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_847 = 12'h34f == _T_2[11:0] ? image_847 : _GEN_846; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3920 = 12'h350 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6992 = 12'h350 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3920; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10064 = 12'h350 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6992; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13136 = 12'h350 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10064; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16208 = 12'h350 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13136; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19280 = 12'h350 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16208; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22352 = 12'h350 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19280; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25424 = 12'h350 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22352; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_848 = io_valid_in ? _GEN_25424 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_848 = 12'h350 == _T_2[11:0] ? image_848 : _GEN_847; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3921 = 12'h351 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6993 = 12'h351 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3921; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10065 = 12'h351 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6993; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13137 = 12'h351 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10065; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16209 = 12'h351 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13137; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19281 = 12'h351 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16209; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22353 = 12'h351 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19281; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25425 = 12'h351 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22353; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_849 = io_valid_in ? _GEN_25425 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_849 = 12'h351 == _T_2[11:0] ? image_849 : _GEN_848; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3922 = 12'h352 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6994 = 12'h352 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3922; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10066 = 12'h352 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6994; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13138 = 12'h352 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10066; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16210 = 12'h352 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13138; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19282 = 12'h352 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16210; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22354 = 12'h352 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19282; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25426 = 12'h352 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22354; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_850 = io_valid_in ? _GEN_25426 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_850 = 12'h352 == _T_2[11:0] ? image_850 : _GEN_849; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3923 = 12'h353 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6995 = 12'h353 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3923; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10067 = 12'h353 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6995; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13139 = 12'h353 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10067; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16211 = 12'h353 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13139; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19283 = 12'h353 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16211; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22355 = 12'h353 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19283; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25427 = 12'h353 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22355; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_851 = io_valid_in ? _GEN_25427 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_851 = 12'h353 == _T_2[11:0] ? image_851 : _GEN_850; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3924 = 12'h354 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6996 = 12'h354 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3924; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10068 = 12'h354 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6996; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13140 = 12'h354 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10068; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16212 = 12'h354 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13140; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19284 = 12'h354 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16212; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22356 = 12'h354 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19284; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25428 = 12'h354 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22356; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_852 = io_valid_in ? _GEN_25428 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_852 = 12'h354 == _T_2[11:0] ? image_852 : _GEN_851; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3925 = 12'h355 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6997 = 12'h355 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3925; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10069 = 12'h355 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6997; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13141 = 12'h355 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10069; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16213 = 12'h355 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13141; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19285 = 12'h355 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16213; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22357 = 12'h355 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19285; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25429 = 12'h355 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22357; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_853 = io_valid_in ? _GEN_25429 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_853 = 12'h355 == _T_2[11:0] ? image_853 : _GEN_852; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3926 = 12'h356 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6998 = 12'h356 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3926; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10070 = 12'h356 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6998; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13142 = 12'h356 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10070; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16214 = 12'h356 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13142; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19286 = 12'h356 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16214; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22358 = 12'h356 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19286; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25430 = 12'h356 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22358; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_854 = io_valid_in ? _GEN_25430 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_854 = 12'h356 == _T_2[11:0] ? image_854 : _GEN_853; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3927 = 12'h357 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_6999 = 12'h357 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3927; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10071 = 12'h357 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_6999; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13143 = 12'h357 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10071; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16215 = 12'h357 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13143; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19287 = 12'h357 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16215; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22359 = 12'h357 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19287; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25431 = 12'h357 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22359; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_855 = io_valid_in ? _GEN_25431 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_855 = 12'h357 == _T_2[11:0] ? image_855 : _GEN_854; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3928 = 12'h358 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7000 = 12'h358 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3928; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10072 = 12'h358 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7000; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13144 = 12'h358 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10072; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16216 = 12'h358 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13144; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19288 = 12'h358 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16216; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22360 = 12'h358 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19288; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25432 = 12'h358 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22360; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_856 = io_valid_in ? _GEN_25432 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_856 = 12'h358 == _T_2[11:0] ? image_856 : _GEN_855; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3929 = 12'h359 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7001 = 12'h359 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3929; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10073 = 12'h359 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7001; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13145 = 12'h359 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10073; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16217 = 12'h359 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13145; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19289 = 12'h359 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16217; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22361 = 12'h359 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19289; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25433 = 12'h359 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22361; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_857 = io_valid_in ? _GEN_25433 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_857 = 12'h359 == _T_2[11:0] ? image_857 : _GEN_856; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3930 = 12'h35a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7002 = 12'h35a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3930; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10074 = 12'h35a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7002; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13146 = 12'h35a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10074; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16218 = 12'h35a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13146; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19290 = 12'h35a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16218; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22362 = 12'h35a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19290; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25434 = 12'h35a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22362; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_858 = io_valid_in ? _GEN_25434 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_858 = 12'h35a == _T_2[11:0] ? image_858 : _GEN_857; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3931 = 12'h35b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7003 = 12'h35b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3931; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10075 = 12'h35b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7003; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13147 = 12'h35b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10075; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16219 = 12'h35b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13147; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19291 = 12'h35b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16219; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22363 = 12'h35b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19291; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25435 = 12'h35b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22363; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_859 = io_valid_in ? _GEN_25435 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_859 = 12'h35b == _T_2[11:0] ? image_859 : _GEN_858; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3932 = 12'h35c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7004 = 12'h35c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3932; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10076 = 12'h35c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7004; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13148 = 12'h35c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10076; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16220 = 12'h35c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13148; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19292 = 12'h35c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16220; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22364 = 12'h35c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19292; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25436 = 12'h35c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22364; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_860 = io_valid_in ? _GEN_25436 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_860 = 12'h35c == _T_2[11:0] ? image_860 : _GEN_859; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3933 = 12'h35d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7005 = 12'h35d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3933; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10077 = 12'h35d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7005; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13149 = 12'h35d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10077; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16221 = 12'h35d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13149; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19293 = 12'h35d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16221; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22365 = 12'h35d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19293; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25437 = 12'h35d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22365; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_861 = io_valid_in ? _GEN_25437 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_861 = 12'h35d == _T_2[11:0] ? image_861 : _GEN_860; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3934 = 12'h35e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7006 = 12'h35e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3934; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10078 = 12'h35e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7006; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13150 = 12'h35e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10078; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16222 = 12'h35e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13150; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19294 = 12'h35e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16222; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22366 = 12'h35e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19294; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25438 = 12'h35e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22366; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_862 = io_valid_in ? _GEN_25438 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_862 = 12'h35e == _T_2[11:0] ? image_862 : _GEN_861; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3935 = 12'h35f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7007 = 12'h35f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3935; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10079 = 12'h35f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7007; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13151 = 12'h35f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10079; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16223 = 12'h35f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13151; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19295 = 12'h35f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16223; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22367 = 12'h35f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19295; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25439 = 12'h35f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22367; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_863 = io_valid_in ? _GEN_25439 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_863 = 12'h35f == _T_2[11:0] ? image_863 : _GEN_862; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3936 = 12'h360 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7008 = 12'h360 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3936; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10080 = 12'h360 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7008; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13152 = 12'h360 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10080; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16224 = 12'h360 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13152; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19296 = 12'h360 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16224; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22368 = 12'h360 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19296; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25440 = 12'h360 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22368; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_864 = io_valid_in ? _GEN_25440 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_864 = 12'h360 == _T_2[11:0] ? image_864 : _GEN_863; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3937 = 12'h361 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7009 = 12'h361 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3937; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10081 = 12'h361 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7009; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13153 = 12'h361 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10081; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16225 = 12'h361 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13153; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19297 = 12'h361 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16225; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22369 = 12'h361 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19297; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25441 = 12'h361 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22369; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_865 = io_valid_in ? _GEN_25441 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_865 = 12'h361 == _T_2[11:0] ? image_865 : _GEN_864; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3938 = 12'h362 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7010 = 12'h362 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3938; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10082 = 12'h362 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7010; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13154 = 12'h362 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10082; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16226 = 12'h362 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13154; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19298 = 12'h362 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16226; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22370 = 12'h362 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19298; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25442 = 12'h362 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22370; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_866 = io_valid_in ? _GEN_25442 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_866 = 12'h362 == _T_2[11:0] ? image_866 : _GEN_865; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3939 = 12'h363 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7011 = 12'h363 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3939; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10083 = 12'h363 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7011; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13155 = 12'h363 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10083; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16227 = 12'h363 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13155; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19299 = 12'h363 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16227; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22371 = 12'h363 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19299; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25443 = 12'h363 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22371; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_867 = io_valid_in ? _GEN_25443 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_867 = 12'h363 == _T_2[11:0] ? image_867 : _GEN_866; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3940 = 12'h364 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7012 = 12'h364 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3940; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10084 = 12'h364 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7012; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13156 = 12'h364 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10084; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16228 = 12'h364 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13156; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19300 = 12'h364 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16228; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22372 = 12'h364 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19300; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25444 = 12'h364 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22372; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_868 = io_valid_in ? _GEN_25444 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_868 = 12'h364 == _T_2[11:0] ? image_868 : _GEN_867; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3941 = 12'h365 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7013 = 12'h365 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3941; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10085 = 12'h365 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7013; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13157 = 12'h365 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10085; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16229 = 12'h365 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13157; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19301 = 12'h365 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16229; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22373 = 12'h365 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19301; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25445 = 12'h365 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22373; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_869 = io_valid_in ? _GEN_25445 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_869 = 12'h365 == _T_2[11:0] ? image_869 : _GEN_868; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3942 = 12'h366 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7014 = 12'h366 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3942; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10086 = 12'h366 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7014; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13158 = 12'h366 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10086; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16230 = 12'h366 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13158; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19302 = 12'h366 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16230; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22374 = 12'h366 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19302; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25446 = 12'h366 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22374; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_870 = io_valid_in ? _GEN_25446 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_870 = 12'h366 == _T_2[11:0] ? image_870 : _GEN_869; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3943 = 12'h367 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7015 = 12'h367 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3943; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10087 = 12'h367 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7015; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13159 = 12'h367 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10087; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16231 = 12'h367 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13159; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19303 = 12'h367 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16231; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22375 = 12'h367 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19303; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25447 = 12'h367 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22375; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_871 = io_valid_in ? _GEN_25447 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_871 = 12'h367 == _T_2[11:0] ? image_871 : _GEN_870; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3944 = 12'h368 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7016 = 12'h368 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3944; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10088 = 12'h368 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7016; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13160 = 12'h368 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10088; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16232 = 12'h368 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13160; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19304 = 12'h368 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16232; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22376 = 12'h368 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19304; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25448 = 12'h368 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22376; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_872 = io_valid_in ? _GEN_25448 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_872 = 12'h368 == _T_2[11:0] ? image_872 : _GEN_871; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3945 = 12'h369 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7017 = 12'h369 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3945; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10089 = 12'h369 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7017; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13161 = 12'h369 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10089; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16233 = 12'h369 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13161; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19305 = 12'h369 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16233; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22377 = 12'h369 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19305; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25449 = 12'h369 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22377; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_873 = io_valid_in ? _GEN_25449 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_873 = 12'h369 == _T_2[11:0] ? image_873 : _GEN_872; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3946 = 12'h36a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7018 = 12'h36a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3946; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10090 = 12'h36a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7018; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13162 = 12'h36a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10090; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16234 = 12'h36a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13162; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19306 = 12'h36a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16234; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22378 = 12'h36a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19306; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25450 = 12'h36a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22378; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_874 = io_valid_in ? _GEN_25450 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_874 = 12'h36a == _T_2[11:0] ? image_874 : _GEN_873; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3947 = 12'h36b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7019 = 12'h36b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3947; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10091 = 12'h36b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7019; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13163 = 12'h36b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10091; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16235 = 12'h36b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13163; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19307 = 12'h36b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16235; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22379 = 12'h36b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19307; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25451 = 12'h36b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22379; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_875 = io_valid_in ? _GEN_25451 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_875 = 12'h36b == _T_2[11:0] ? image_875 : _GEN_874; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3948 = 12'h36c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7020 = 12'h36c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3948; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10092 = 12'h36c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7020; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13164 = 12'h36c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10092; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16236 = 12'h36c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13164; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19308 = 12'h36c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16236; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22380 = 12'h36c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19308; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25452 = 12'h36c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22380; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_876 = io_valid_in ? _GEN_25452 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_876 = 12'h36c == _T_2[11:0] ? image_876 : _GEN_875; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3949 = 12'h36d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7021 = 12'h36d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3949; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10093 = 12'h36d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7021; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13165 = 12'h36d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10093; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16237 = 12'h36d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13165; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19309 = 12'h36d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16237; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22381 = 12'h36d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19309; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25453 = 12'h36d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22381; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_877 = io_valid_in ? _GEN_25453 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_877 = 12'h36d == _T_2[11:0] ? image_877 : _GEN_876; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3950 = 12'h36e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7022 = 12'h36e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3950; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10094 = 12'h36e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7022; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13166 = 12'h36e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10094; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16238 = 12'h36e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13166; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19310 = 12'h36e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16238; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22382 = 12'h36e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19310; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25454 = 12'h36e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22382; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_878 = io_valid_in ? _GEN_25454 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_878 = 12'h36e == _T_2[11:0] ? image_878 : _GEN_877; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3951 = 12'h36f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7023 = 12'h36f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3951; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10095 = 12'h36f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7023; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13167 = 12'h36f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10095; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16239 = 12'h36f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13167; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19311 = 12'h36f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16239; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22383 = 12'h36f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19311; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25455 = 12'h36f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22383; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_879 = io_valid_in ? _GEN_25455 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_879 = 12'h36f == _T_2[11:0] ? image_879 : _GEN_878; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3952 = 12'h370 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7024 = 12'h370 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3952; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10096 = 12'h370 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7024; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13168 = 12'h370 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10096; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16240 = 12'h370 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13168; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19312 = 12'h370 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16240; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22384 = 12'h370 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19312; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25456 = 12'h370 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22384; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_880 = io_valid_in ? _GEN_25456 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_880 = 12'h370 == _T_2[11:0] ? image_880 : _GEN_879; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3953 = 12'h371 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7025 = 12'h371 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3953; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10097 = 12'h371 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7025; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13169 = 12'h371 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10097; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16241 = 12'h371 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13169; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19313 = 12'h371 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16241; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22385 = 12'h371 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19313; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25457 = 12'h371 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22385; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_881 = io_valid_in ? _GEN_25457 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_881 = 12'h371 == _T_2[11:0] ? image_881 : _GEN_880; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3954 = 12'h372 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7026 = 12'h372 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3954; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10098 = 12'h372 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7026; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13170 = 12'h372 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10098; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16242 = 12'h372 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13170; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19314 = 12'h372 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16242; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22386 = 12'h372 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19314; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25458 = 12'h372 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22386; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_882 = io_valid_in ? _GEN_25458 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_882 = 12'h372 == _T_2[11:0] ? image_882 : _GEN_881; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3955 = 12'h373 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7027 = 12'h373 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3955; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10099 = 12'h373 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7027; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13171 = 12'h373 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10099; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16243 = 12'h373 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13171; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19315 = 12'h373 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16243; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22387 = 12'h373 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19315; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25459 = 12'h373 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22387; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_883 = io_valid_in ? _GEN_25459 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_883 = 12'h373 == _T_2[11:0] ? image_883 : _GEN_882; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3956 = 12'h374 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7028 = 12'h374 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3956; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10100 = 12'h374 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7028; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13172 = 12'h374 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10100; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16244 = 12'h374 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13172; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19316 = 12'h374 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16244; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22388 = 12'h374 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19316; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25460 = 12'h374 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22388; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_884 = io_valid_in ? _GEN_25460 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_884 = 12'h374 == _T_2[11:0] ? image_884 : _GEN_883; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3957 = 12'h375 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7029 = 12'h375 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3957; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10101 = 12'h375 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7029; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13173 = 12'h375 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10101; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16245 = 12'h375 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13173; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19317 = 12'h375 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16245; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22389 = 12'h375 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19317; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25461 = 12'h375 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22389; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_885 = io_valid_in ? _GEN_25461 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_885 = 12'h375 == _T_2[11:0] ? image_885 : _GEN_884; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3958 = 12'h376 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7030 = 12'h376 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3958; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10102 = 12'h376 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7030; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13174 = 12'h376 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10102; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16246 = 12'h376 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13174; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19318 = 12'h376 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16246; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22390 = 12'h376 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19318; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25462 = 12'h376 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22390; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_886 = io_valid_in ? _GEN_25462 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_886 = 12'h376 == _T_2[11:0] ? image_886 : _GEN_885; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3959 = 12'h377 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7031 = 12'h377 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3959; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10103 = 12'h377 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7031; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13175 = 12'h377 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10103; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16247 = 12'h377 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13175; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19319 = 12'h377 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16247; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22391 = 12'h377 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19319; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25463 = 12'h377 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22391; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_887 = io_valid_in ? _GEN_25463 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_887 = 12'h377 == _T_2[11:0] ? image_887 : _GEN_886; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3960 = 12'h378 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7032 = 12'h378 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3960; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10104 = 12'h378 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7032; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13176 = 12'h378 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10104; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16248 = 12'h378 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13176; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19320 = 12'h378 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16248; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22392 = 12'h378 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19320; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25464 = 12'h378 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22392; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_888 = io_valid_in ? _GEN_25464 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_888 = 12'h378 == _T_2[11:0] ? image_888 : _GEN_887; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3961 = 12'h379 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7033 = 12'h379 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3961; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10105 = 12'h379 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7033; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13177 = 12'h379 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10105; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16249 = 12'h379 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13177; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19321 = 12'h379 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16249; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22393 = 12'h379 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19321; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25465 = 12'h379 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22393; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_889 = io_valid_in ? _GEN_25465 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_889 = 12'h379 == _T_2[11:0] ? image_889 : _GEN_888; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3962 = 12'h37a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7034 = 12'h37a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3962; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10106 = 12'h37a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7034; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13178 = 12'h37a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10106; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16250 = 12'h37a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13178; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19322 = 12'h37a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16250; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22394 = 12'h37a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19322; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25466 = 12'h37a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22394; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_890 = io_valid_in ? _GEN_25466 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_890 = 12'h37a == _T_2[11:0] ? image_890 : _GEN_889; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3963 = 12'h37b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7035 = 12'h37b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3963; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10107 = 12'h37b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7035; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13179 = 12'h37b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10107; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16251 = 12'h37b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13179; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19323 = 12'h37b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16251; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22395 = 12'h37b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19323; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25467 = 12'h37b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22395; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_891 = io_valid_in ? _GEN_25467 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_891 = 12'h37b == _T_2[11:0] ? image_891 : _GEN_890; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3964 = 12'h37c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7036 = 12'h37c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3964; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10108 = 12'h37c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7036; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13180 = 12'h37c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10108; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16252 = 12'h37c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13180; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19324 = 12'h37c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16252; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22396 = 12'h37c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19324; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25468 = 12'h37c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22396; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_892 = io_valid_in ? _GEN_25468 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_892 = 12'h37c == _T_2[11:0] ? image_892 : _GEN_891; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3965 = 12'h37d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7037 = 12'h37d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3965; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10109 = 12'h37d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7037; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13181 = 12'h37d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10109; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16253 = 12'h37d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13181; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19325 = 12'h37d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16253; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22397 = 12'h37d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19325; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25469 = 12'h37d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22397; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_893 = io_valid_in ? _GEN_25469 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_893 = 12'h37d == _T_2[11:0] ? image_893 : _GEN_892; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3966 = 12'h37e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7038 = 12'h37e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3966; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10110 = 12'h37e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7038; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13182 = 12'h37e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10110; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16254 = 12'h37e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13182; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19326 = 12'h37e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16254; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22398 = 12'h37e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19326; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25470 = 12'h37e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22398; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_894 = io_valid_in ? _GEN_25470 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_894 = 12'h37e == _T_2[11:0] ? image_894 : _GEN_893; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3967 = 12'h37f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7039 = 12'h37f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3967; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10111 = 12'h37f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7039; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13183 = 12'h37f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10111; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16255 = 12'h37f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13183; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19327 = 12'h37f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16255; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22399 = 12'h37f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19327; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25471 = 12'h37f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22399; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_895 = io_valid_in ? _GEN_25471 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_895 = 12'h37f == _T_2[11:0] ? image_895 : _GEN_894; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3968 = 12'h380 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7040 = 12'h380 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3968; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10112 = 12'h380 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7040; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13184 = 12'h380 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10112; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16256 = 12'h380 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13184; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19328 = 12'h380 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16256; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22400 = 12'h380 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19328; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25472 = 12'h380 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22400; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_896 = io_valid_in ? _GEN_25472 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_896 = 12'h380 == _T_2[11:0] ? image_896 : _GEN_895; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3969 = 12'h381 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7041 = 12'h381 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3969; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10113 = 12'h381 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7041; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13185 = 12'h381 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10113; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16257 = 12'h381 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13185; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19329 = 12'h381 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16257; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22401 = 12'h381 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19329; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25473 = 12'h381 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22401; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_897 = io_valid_in ? _GEN_25473 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_897 = 12'h381 == _T_2[11:0] ? image_897 : _GEN_896; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3970 = 12'h382 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7042 = 12'h382 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3970; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10114 = 12'h382 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7042; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13186 = 12'h382 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10114; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16258 = 12'h382 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13186; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19330 = 12'h382 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16258; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22402 = 12'h382 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19330; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25474 = 12'h382 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22402; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_898 = io_valid_in ? _GEN_25474 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_898 = 12'h382 == _T_2[11:0] ? image_898 : _GEN_897; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3971 = 12'h383 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7043 = 12'h383 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3971; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10115 = 12'h383 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7043; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13187 = 12'h383 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10115; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16259 = 12'h383 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13187; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19331 = 12'h383 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16259; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22403 = 12'h383 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19331; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25475 = 12'h383 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22403; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_899 = io_valid_in ? _GEN_25475 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_899 = 12'h383 == _T_2[11:0] ? image_899 : _GEN_898; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3972 = 12'h384 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7044 = 12'h384 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3972; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10116 = 12'h384 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7044; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13188 = 12'h384 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10116; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16260 = 12'h384 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13188; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19332 = 12'h384 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16260; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22404 = 12'h384 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19332; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25476 = 12'h384 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22404; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_900 = io_valid_in ? _GEN_25476 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_900 = 12'h384 == _T_2[11:0] ? image_900 : _GEN_899; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3973 = 12'h385 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7045 = 12'h385 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3973; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10117 = 12'h385 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7045; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13189 = 12'h385 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10117; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16261 = 12'h385 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13189; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19333 = 12'h385 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16261; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22405 = 12'h385 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19333; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25477 = 12'h385 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22405; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_901 = io_valid_in ? _GEN_25477 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_901 = 12'h385 == _T_2[11:0] ? image_901 : _GEN_900; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3974 = 12'h386 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7046 = 12'h386 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3974; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10118 = 12'h386 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7046; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13190 = 12'h386 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10118; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16262 = 12'h386 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13190; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19334 = 12'h386 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16262; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22406 = 12'h386 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19334; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25478 = 12'h386 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22406; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_902 = io_valid_in ? _GEN_25478 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_902 = 12'h386 == _T_2[11:0] ? image_902 : _GEN_901; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3975 = 12'h387 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7047 = 12'h387 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3975; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10119 = 12'h387 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7047; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13191 = 12'h387 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10119; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16263 = 12'h387 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13191; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19335 = 12'h387 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16263; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22407 = 12'h387 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19335; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25479 = 12'h387 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22407; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_903 = io_valid_in ? _GEN_25479 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_903 = 12'h387 == _T_2[11:0] ? image_903 : _GEN_902; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3976 = 12'h388 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7048 = 12'h388 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3976; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10120 = 12'h388 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7048; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13192 = 12'h388 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10120; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16264 = 12'h388 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13192; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19336 = 12'h388 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16264; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22408 = 12'h388 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19336; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25480 = 12'h388 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22408; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_904 = io_valid_in ? _GEN_25480 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_904 = 12'h388 == _T_2[11:0] ? image_904 : _GEN_903; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3977 = 12'h389 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7049 = 12'h389 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3977; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10121 = 12'h389 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7049; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13193 = 12'h389 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10121; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16265 = 12'h389 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13193; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19337 = 12'h389 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16265; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22409 = 12'h389 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19337; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25481 = 12'h389 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22409; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_905 = io_valid_in ? _GEN_25481 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_905 = 12'h389 == _T_2[11:0] ? image_905 : _GEN_904; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3978 = 12'h38a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7050 = 12'h38a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3978; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10122 = 12'h38a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7050; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13194 = 12'h38a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10122; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16266 = 12'h38a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13194; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19338 = 12'h38a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16266; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22410 = 12'h38a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19338; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25482 = 12'h38a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22410; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_906 = io_valid_in ? _GEN_25482 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_906 = 12'h38a == _T_2[11:0] ? image_906 : _GEN_905; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3979 = 12'h38b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7051 = 12'h38b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3979; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10123 = 12'h38b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7051; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13195 = 12'h38b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10123; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16267 = 12'h38b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13195; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19339 = 12'h38b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16267; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22411 = 12'h38b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19339; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25483 = 12'h38b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22411; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_907 = io_valid_in ? _GEN_25483 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_907 = 12'h38b == _T_2[11:0] ? image_907 : _GEN_906; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3980 = 12'h38c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7052 = 12'h38c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3980; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10124 = 12'h38c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7052; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13196 = 12'h38c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10124; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16268 = 12'h38c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13196; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19340 = 12'h38c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16268; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22412 = 12'h38c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19340; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25484 = 12'h38c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22412; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_908 = io_valid_in ? _GEN_25484 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_908 = 12'h38c == _T_2[11:0] ? image_908 : _GEN_907; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3981 = 12'h38d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7053 = 12'h38d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3981; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10125 = 12'h38d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7053; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13197 = 12'h38d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10125; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16269 = 12'h38d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13197; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19341 = 12'h38d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16269; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22413 = 12'h38d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19341; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25485 = 12'h38d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22413; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_909 = io_valid_in ? _GEN_25485 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_909 = 12'h38d == _T_2[11:0] ? image_909 : _GEN_908; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3982 = 12'h38e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7054 = 12'h38e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3982; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10126 = 12'h38e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7054; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13198 = 12'h38e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10126; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16270 = 12'h38e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13198; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19342 = 12'h38e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16270; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22414 = 12'h38e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19342; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25486 = 12'h38e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22414; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_910 = io_valid_in ? _GEN_25486 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_910 = 12'h38e == _T_2[11:0] ? image_910 : _GEN_909; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3983 = 12'h38f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7055 = 12'h38f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3983; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10127 = 12'h38f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7055; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13199 = 12'h38f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10127; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16271 = 12'h38f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13199; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19343 = 12'h38f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16271; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22415 = 12'h38f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19343; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25487 = 12'h38f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22415; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_911 = io_valid_in ? _GEN_25487 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_911 = 12'h38f == _T_2[11:0] ? image_911 : _GEN_910; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3984 = 12'h390 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7056 = 12'h390 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3984; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10128 = 12'h390 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7056; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13200 = 12'h390 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10128; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16272 = 12'h390 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13200; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19344 = 12'h390 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16272; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22416 = 12'h390 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19344; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25488 = 12'h390 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22416; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_912 = io_valid_in ? _GEN_25488 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_912 = 12'h390 == _T_2[11:0] ? image_912 : _GEN_911; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3985 = 12'h391 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7057 = 12'h391 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3985; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10129 = 12'h391 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7057; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13201 = 12'h391 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10129; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16273 = 12'h391 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13201; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19345 = 12'h391 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16273; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22417 = 12'h391 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19345; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25489 = 12'h391 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22417; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_913 = io_valid_in ? _GEN_25489 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_913 = 12'h391 == _T_2[11:0] ? image_913 : _GEN_912; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3986 = 12'h392 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7058 = 12'h392 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3986; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10130 = 12'h392 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7058; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13202 = 12'h392 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10130; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16274 = 12'h392 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13202; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19346 = 12'h392 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16274; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22418 = 12'h392 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19346; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25490 = 12'h392 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22418; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_914 = io_valid_in ? _GEN_25490 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_914 = 12'h392 == _T_2[11:0] ? image_914 : _GEN_913; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3987 = 12'h393 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7059 = 12'h393 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3987; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10131 = 12'h393 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7059; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13203 = 12'h393 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10131; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16275 = 12'h393 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13203; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19347 = 12'h393 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16275; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22419 = 12'h393 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19347; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25491 = 12'h393 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22419; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_915 = io_valid_in ? _GEN_25491 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_915 = 12'h393 == _T_2[11:0] ? image_915 : _GEN_914; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3988 = 12'h394 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7060 = 12'h394 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3988; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10132 = 12'h394 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7060; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13204 = 12'h394 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10132; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16276 = 12'h394 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13204; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19348 = 12'h394 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16276; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22420 = 12'h394 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19348; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25492 = 12'h394 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22420; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_916 = io_valid_in ? _GEN_25492 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_916 = 12'h394 == _T_2[11:0] ? image_916 : _GEN_915; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3989 = 12'h395 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7061 = 12'h395 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3989; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10133 = 12'h395 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7061; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13205 = 12'h395 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10133; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16277 = 12'h395 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13205; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19349 = 12'h395 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16277; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22421 = 12'h395 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19349; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25493 = 12'h395 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22421; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_917 = io_valid_in ? _GEN_25493 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_917 = 12'h395 == _T_2[11:0] ? image_917 : _GEN_916; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3990 = 12'h396 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7062 = 12'h396 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3990; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10134 = 12'h396 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7062; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13206 = 12'h396 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10134; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16278 = 12'h396 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13206; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19350 = 12'h396 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16278; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22422 = 12'h396 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19350; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25494 = 12'h396 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22422; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_918 = io_valid_in ? _GEN_25494 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_918 = 12'h396 == _T_2[11:0] ? image_918 : _GEN_917; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3991 = 12'h397 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7063 = 12'h397 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3991; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10135 = 12'h397 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7063; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13207 = 12'h397 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10135; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16279 = 12'h397 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13207; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19351 = 12'h397 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16279; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22423 = 12'h397 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19351; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25495 = 12'h397 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22423; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_919 = io_valid_in ? _GEN_25495 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_919 = 12'h397 == _T_2[11:0] ? image_919 : _GEN_918; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3992 = 12'h398 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7064 = 12'h398 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3992; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10136 = 12'h398 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7064; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13208 = 12'h398 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10136; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16280 = 12'h398 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13208; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19352 = 12'h398 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16280; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22424 = 12'h398 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19352; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25496 = 12'h398 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22424; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_920 = io_valid_in ? _GEN_25496 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_920 = 12'h398 == _T_2[11:0] ? image_920 : _GEN_919; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3993 = 12'h399 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7065 = 12'h399 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3993; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10137 = 12'h399 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7065; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13209 = 12'h399 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10137; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16281 = 12'h399 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13209; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19353 = 12'h399 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16281; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22425 = 12'h399 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19353; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25497 = 12'h399 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22425; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_921 = io_valid_in ? _GEN_25497 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_921 = 12'h399 == _T_2[11:0] ? image_921 : _GEN_920; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3994 = 12'h39a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7066 = 12'h39a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3994; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10138 = 12'h39a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7066; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13210 = 12'h39a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10138; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16282 = 12'h39a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13210; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19354 = 12'h39a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16282; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22426 = 12'h39a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19354; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25498 = 12'h39a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22426; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_922 = io_valid_in ? _GEN_25498 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_922 = 12'h39a == _T_2[11:0] ? image_922 : _GEN_921; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3995 = 12'h39b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7067 = 12'h39b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3995; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10139 = 12'h39b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7067; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13211 = 12'h39b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10139; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16283 = 12'h39b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13211; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19355 = 12'h39b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16283; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22427 = 12'h39b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19355; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25499 = 12'h39b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22427; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_923 = io_valid_in ? _GEN_25499 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_923 = 12'h39b == _T_2[11:0] ? image_923 : _GEN_922; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3996 = 12'h39c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7068 = 12'h39c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3996; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10140 = 12'h39c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7068; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13212 = 12'h39c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10140; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16284 = 12'h39c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13212; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19356 = 12'h39c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16284; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22428 = 12'h39c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19356; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25500 = 12'h39c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22428; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_924 = io_valid_in ? _GEN_25500 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_924 = 12'h39c == _T_2[11:0] ? image_924 : _GEN_923; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3997 = 12'h39d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7069 = 12'h39d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3997; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10141 = 12'h39d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7069; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13213 = 12'h39d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10141; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16285 = 12'h39d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13213; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19357 = 12'h39d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16285; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22429 = 12'h39d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19357; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25501 = 12'h39d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22429; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_925 = io_valid_in ? _GEN_25501 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_925 = 12'h39d == _T_2[11:0] ? image_925 : _GEN_924; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3998 = 12'h39e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7070 = 12'h39e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3998; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10142 = 12'h39e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7070; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13214 = 12'h39e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10142; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16286 = 12'h39e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13214; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19358 = 12'h39e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16286; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22430 = 12'h39e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19358; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25502 = 12'h39e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22430; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_926 = io_valid_in ? _GEN_25502 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_926 = 12'h39e == _T_2[11:0] ? image_926 : _GEN_925; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_3999 = 12'h39f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7071 = 12'h39f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_3999; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10143 = 12'h39f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7071; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13215 = 12'h39f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10143; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16287 = 12'h39f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13215; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19359 = 12'h39f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16287; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22431 = 12'h39f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19359; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25503 = 12'h39f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22431; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_927 = io_valid_in ? _GEN_25503 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_927 = 12'h39f == _T_2[11:0] ? image_927 : _GEN_926; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4000 = 12'h3a0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7072 = 12'h3a0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4000; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10144 = 12'h3a0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7072; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13216 = 12'h3a0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10144; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16288 = 12'h3a0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13216; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19360 = 12'h3a0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16288; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22432 = 12'h3a0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19360; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25504 = 12'h3a0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22432; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_928 = io_valid_in ? _GEN_25504 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_928 = 12'h3a0 == _T_2[11:0] ? image_928 : _GEN_927; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4001 = 12'h3a1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7073 = 12'h3a1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4001; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10145 = 12'h3a1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7073; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13217 = 12'h3a1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10145; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16289 = 12'h3a1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13217; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19361 = 12'h3a1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16289; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22433 = 12'h3a1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19361; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25505 = 12'h3a1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22433; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_929 = io_valid_in ? _GEN_25505 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_929 = 12'h3a1 == _T_2[11:0] ? image_929 : _GEN_928; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4002 = 12'h3a2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7074 = 12'h3a2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4002; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10146 = 12'h3a2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7074; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13218 = 12'h3a2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10146; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16290 = 12'h3a2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13218; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19362 = 12'h3a2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16290; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22434 = 12'h3a2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19362; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25506 = 12'h3a2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22434; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_930 = io_valid_in ? _GEN_25506 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_930 = 12'h3a2 == _T_2[11:0] ? image_930 : _GEN_929; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4003 = 12'h3a3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7075 = 12'h3a3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4003; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10147 = 12'h3a3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7075; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13219 = 12'h3a3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10147; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16291 = 12'h3a3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13219; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19363 = 12'h3a3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16291; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22435 = 12'h3a3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19363; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25507 = 12'h3a3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22435; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_931 = io_valid_in ? _GEN_25507 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_931 = 12'h3a3 == _T_2[11:0] ? image_931 : _GEN_930; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4004 = 12'h3a4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7076 = 12'h3a4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4004; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10148 = 12'h3a4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7076; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13220 = 12'h3a4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10148; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16292 = 12'h3a4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13220; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19364 = 12'h3a4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16292; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22436 = 12'h3a4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19364; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25508 = 12'h3a4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22436; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_932 = io_valid_in ? _GEN_25508 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_932 = 12'h3a4 == _T_2[11:0] ? image_932 : _GEN_931; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4005 = 12'h3a5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7077 = 12'h3a5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4005; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10149 = 12'h3a5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7077; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13221 = 12'h3a5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10149; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16293 = 12'h3a5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13221; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19365 = 12'h3a5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16293; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22437 = 12'h3a5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19365; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25509 = 12'h3a5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22437; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_933 = io_valid_in ? _GEN_25509 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_933 = 12'h3a5 == _T_2[11:0] ? image_933 : _GEN_932; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4006 = 12'h3a6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7078 = 12'h3a6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4006; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10150 = 12'h3a6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7078; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13222 = 12'h3a6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10150; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16294 = 12'h3a6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13222; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19366 = 12'h3a6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16294; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22438 = 12'h3a6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19366; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25510 = 12'h3a6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22438; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_934 = io_valid_in ? _GEN_25510 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_934 = 12'h3a6 == _T_2[11:0] ? image_934 : _GEN_933; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4007 = 12'h3a7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7079 = 12'h3a7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4007; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10151 = 12'h3a7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7079; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13223 = 12'h3a7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10151; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16295 = 12'h3a7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13223; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19367 = 12'h3a7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16295; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22439 = 12'h3a7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19367; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25511 = 12'h3a7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22439; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_935 = io_valid_in ? _GEN_25511 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_935 = 12'h3a7 == _T_2[11:0] ? image_935 : _GEN_934; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4008 = 12'h3a8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7080 = 12'h3a8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4008; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10152 = 12'h3a8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7080; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13224 = 12'h3a8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10152; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16296 = 12'h3a8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13224; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19368 = 12'h3a8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16296; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22440 = 12'h3a8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19368; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25512 = 12'h3a8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22440; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_936 = io_valid_in ? _GEN_25512 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_936 = 12'h3a8 == _T_2[11:0] ? image_936 : _GEN_935; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4009 = 12'h3a9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7081 = 12'h3a9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4009; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10153 = 12'h3a9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7081; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13225 = 12'h3a9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10153; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16297 = 12'h3a9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13225; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19369 = 12'h3a9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16297; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22441 = 12'h3a9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19369; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25513 = 12'h3a9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22441; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_937 = io_valid_in ? _GEN_25513 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_937 = 12'h3a9 == _T_2[11:0] ? image_937 : _GEN_936; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4010 = 12'h3aa == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7082 = 12'h3aa == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4010; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10154 = 12'h3aa == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7082; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13226 = 12'h3aa == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10154; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16298 = 12'h3aa == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13226; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19370 = 12'h3aa == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16298; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22442 = 12'h3aa == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19370; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25514 = 12'h3aa == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22442; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_938 = io_valid_in ? _GEN_25514 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_938 = 12'h3aa == _T_2[11:0] ? image_938 : _GEN_937; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4011 = 12'h3ab == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7083 = 12'h3ab == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4011; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10155 = 12'h3ab == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7083; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13227 = 12'h3ab == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10155; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16299 = 12'h3ab == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13227; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19371 = 12'h3ab == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16299; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22443 = 12'h3ab == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19371; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25515 = 12'h3ab == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22443; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_939 = io_valid_in ? _GEN_25515 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_939 = 12'h3ab == _T_2[11:0] ? image_939 : _GEN_938; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4012 = 12'h3ac == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7084 = 12'h3ac == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4012; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10156 = 12'h3ac == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7084; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13228 = 12'h3ac == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10156; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16300 = 12'h3ac == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13228; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19372 = 12'h3ac == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16300; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22444 = 12'h3ac == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19372; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25516 = 12'h3ac == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22444; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_940 = io_valid_in ? _GEN_25516 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_940 = 12'h3ac == _T_2[11:0] ? image_940 : _GEN_939; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4013 = 12'h3ad == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7085 = 12'h3ad == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4013; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10157 = 12'h3ad == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7085; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13229 = 12'h3ad == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10157; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16301 = 12'h3ad == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13229; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19373 = 12'h3ad == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16301; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22445 = 12'h3ad == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19373; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25517 = 12'h3ad == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22445; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_941 = io_valid_in ? _GEN_25517 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_941 = 12'h3ad == _T_2[11:0] ? image_941 : _GEN_940; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4014 = 12'h3ae == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7086 = 12'h3ae == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4014; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10158 = 12'h3ae == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7086; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13230 = 12'h3ae == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10158; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16302 = 12'h3ae == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13230; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19374 = 12'h3ae == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16302; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22446 = 12'h3ae == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19374; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25518 = 12'h3ae == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22446; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_942 = io_valid_in ? _GEN_25518 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_942 = 12'h3ae == _T_2[11:0] ? image_942 : _GEN_941; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4015 = 12'h3af == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7087 = 12'h3af == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4015; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10159 = 12'h3af == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7087; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13231 = 12'h3af == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10159; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16303 = 12'h3af == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13231; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19375 = 12'h3af == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16303; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22447 = 12'h3af == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19375; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25519 = 12'h3af == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22447; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_943 = io_valid_in ? _GEN_25519 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_943 = 12'h3af == _T_2[11:0] ? image_943 : _GEN_942; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4016 = 12'h3b0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7088 = 12'h3b0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4016; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10160 = 12'h3b0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7088; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13232 = 12'h3b0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10160; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16304 = 12'h3b0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13232; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19376 = 12'h3b0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16304; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22448 = 12'h3b0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19376; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25520 = 12'h3b0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22448; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_944 = io_valid_in ? _GEN_25520 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_944 = 12'h3b0 == _T_2[11:0] ? image_944 : _GEN_943; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4017 = 12'h3b1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7089 = 12'h3b1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4017; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10161 = 12'h3b1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7089; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13233 = 12'h3b1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10161; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16305 = 12'h3b1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13233; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19377 = 12'h3b1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16305; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22449 = 12'h3b1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19377; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25521 = 12'h3b1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22449; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_945 = io_valid_in ? _GEN_25521 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_945 = 12'h3b1 == _T_2[11:0] ? image_945 : _GEN_944; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4018 = 12'h3b2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7090 = 12'h3b2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4018; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10162 = 12'h3b2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7090; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13234 = 12'h3b2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10162; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16306 = 12'h3b2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13234; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19378 = 12'h3b2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16306; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22450 = 12'h3b2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19378; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25522 = 12'h3b2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22450; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_946 = io_valid_in ? _GEN_25522 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_946 = 12'h3b2 == _T_2[11:0] ? image_946 : _GEN_945; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4019 = 12'h3b3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7091 = 12'h3b3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4019; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10163 = 12'h3b3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7091; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13235 = 12'h3b3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10163; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16307 = 12'h3b3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13235; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19379 = 12'h3b3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16307; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22451 = 12'h3b3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19379; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25523 = 12'h3b3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22451; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_947 = io_valid_in ? _GEN_25523 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_947 = 12'h3b3 == _T_2[11:0] ? image_947 : _GEN_946; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4020 = 12'h3b4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7092 = 12'h3b4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4020; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10164 = 12'h3b4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7092; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13236 = 12'h3b4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10164; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16308 = 12'h3b4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13236; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19380 = 12'h3b4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16308; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22452 = 12'h3b4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19380; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25524 = 12'h3b4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22452; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_948 = io_valid_in ? _GEN_25524 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_948 = 12'h3b4 == _T_2[11:0] ? image_948 : _GEN_947; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4021 = 12'h3b5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7093 = 12'h3b5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4021; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10165 = 12'h3b5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7093; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13237 = 12'h3b5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10165; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16309 = 12'h3b5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13237; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19381 = 12'h3b5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16309; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22453 = 12'h3b5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19381; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25525 = 12'h3b5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22453; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_949 = io_valid_in ? _GEN_25525 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_949 = 12'h3b5 == _T_2[11:0] ? image_949 : _GEN_948; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4022 = 12'h3b6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7094 = 12'h3b6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4022; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10166 = 12'h3b6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7094; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13238 = 12'h3b6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10166; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16310 = 12'h3b6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13238; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19382 = 12'h3b6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16310; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22454 = 12'h3b6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19382; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25526 = 12'h3b6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22454; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_950 = io_valid_in ? _GEN_25526 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_950 = 12'h3b6 == _T_2[11:0] ? image_950 : _GEN_949; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4023 = 12'h3b7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7095 = 12'h3b7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4023; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10167 = 12'h3b7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7095; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13239 = 12'h3b7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10167; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16311 = 12'h3b7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13239; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19383 = 12'h3b7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16311; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22455 = 12'h3b7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19383; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25527 = 12'h3b7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22455; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_951 = io_valid_in ? _GEN_25527 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_951 = 12'h3b7 == _T_2[11:0] ? image_951 : _GEN_950; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4024 = 12'h3b8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7096 = 12'h3b8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4024; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10168 = 12'h3b8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7096; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13240 = 12'h3b8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10168; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16312 = 12'h3b8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13240; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19384 = 12'h3b8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16312; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22456 = 12'h3b8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19384; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25528 = 12'h3b8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22456; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_952 = io_valid_in ? _GEN_25528 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_952 = 12'h3b8 == _T_2[11:0] ? image_952 : _GEN_951; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4025 = 12'h3b9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7097 = 12'h3b9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4025; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10169 = 12'h3b9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7097; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13241 = 12'h3b9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10169; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16313 = 12'h3b9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13241; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19385 = 12'h3b9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16313; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22457 = 12'h3b9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19385; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25529 = 12'h3b9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22457; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_953 = io_valid_in ? _GEN_25529 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_953 = 12'h3b9 == _T_2[11:0] ? image_953 : _GEN_952; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4026 = 12'h3ba == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7098 = 12'h3ba == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4026; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10170 = 12'h3ba == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7098; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13242 = 12'h3ba == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10170; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16314 = 12'h3ba == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13242; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19386 = 12'h3ba == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16314; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22458 = 12'h3ba == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19386; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25530 = 12'h3ba == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22458; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_954 = io_valid_in ? _GEN_25530 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_954 = 12'h3ba == _T_2[11:0] ? image_954 : _GEN_953; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4027 = 12'h3bb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7099 = 12'h3bb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4027; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10171 = 12'h3bb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7099; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13243 = 12'h3bb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10171; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16315 = 12'h3bb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13243; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19387 = 12'h3bb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16315; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22459 = 12'h3bb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19387; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25531 = 12'h3bb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22459; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_955 = io_valid_in ? _GEN_25531 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_955 = 12'h3bb == _T_2[11:0] ? image_955 : _GEN_954; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4028 = 12'h3bc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7100 = 12'h3bc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4028; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10172 = 12'h3bc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7100; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13244 = 12'h3bc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10172; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16316 = 12'h3bc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13244; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19388 = 12'h3bc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16316; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22460 = 12'h3bc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19388; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25532 = 12'h3bc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22460; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_956 = io_valid_in ? _GEN_25532 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_956 = 12'h3bc == _T_2[11:0] ? image_956 : _GEN_955; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4029 = 12'h3bd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7101 = 12'h3bd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4029; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10173 = 12'h3bd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7101; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13245 = 12'h3bd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10173; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16317 = 12'h3bd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13245; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19389 = 12'h3bd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16317; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22461 = 12'h3bd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19389; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25533 = 12'h3bd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22461; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_957 = io_valid_in ? _GEN_25533 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_957 = 12'h3bd == _T_2[11:0] ? image_957 : _GEN_956; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4030 = 12'h3be == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7102 = 12'h3be == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4030; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10174 = 12'h3be == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7102; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13246 = 12'h3be == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10174; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16318 = 12'h3be == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13246; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19390 = 12'h3be == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16318; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22462 = 12'h3be == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19390; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25534 = 12'h3be == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22462; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_958 = io_valid_in ? _GEN_25534 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_958 = 12'h3be == _T_2[11:0] ? image_958 : _GEN_957; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4031 = 12'h3bf == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7103 = 12'h3bf == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4031; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10175 = 12'h3bf == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7103; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13247 = 12'h3bf == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10175; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16319 = 12'h3bf == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13247; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19391 = 12'h3bf == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16319; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22463 = 12'h3bf == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19391; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25535 = 12'h3bf == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22463; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_959 = io_valid_in ? _GEN_25535 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_959 = 12'h3bf == _T_2[11:0] ? image_959 : _GEN_958; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4032 = 12'h3c0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7104 = 12'h3c0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4032; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10176 = 12'h3c0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7104; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13248 = 12'h3c0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10176; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16320 = 12'h3c0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13248; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19392 = 12'h3c0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16320; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22464 = 12'h3c0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19392; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25536 = 12'h3c0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22464; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_960 = io_valid_in ? _GEN_25536 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_960 = 12'h3c0 == _T_2[11:0] ? image_960 : _GEN_959; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4033 = 12'h3c1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7105 = 12'h3c1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4033; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10177 = 12'h3c1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7105; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13249 = 12'h3c1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10177; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16321 = 12'h3c1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13249; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19393 = 12'h3c1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16321; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22465 = 12'h3c1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19393; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25537 = 12'h3c1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22465; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_961 = io_valid_in ? _GEN_25537 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_961 = 12'h3c1 == _T_2[11:0] ? image_961 : _GEN_960; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4034 = 12'h3c2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7106 = 12'h3c2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4034; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10178 = 12'h3c2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7106; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13250 = 12'h3c2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10178; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16322 = 12'h3c2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13250; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19394 = 12'h3c2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16322; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22466 = 12'h3c2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19394; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25538 = 12'h3c2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22466; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_962 = io_valid_in ? _GEN_25538 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_962 = 12'h3c2 == _T_2[11:0] ? image_962 : _GEN_961; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4035 = 12'h3c3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7107 = 12'h3c3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4035; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10179 = 12'h3c3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7107; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13251 = 12'h3c3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10179; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16323 = 12'h3c3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13251; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19395 = 12'h3c3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16323; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22467 = 12'h3c3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19395; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25539 = 12'h3c3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22467; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_963 = io_valid_in ? _GEN_25539 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_963 = 12'h3c3 == _T_2[11:0] ? image_963 : _GEN_962; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4036 = 12'h3c4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7108 = 12'h3c4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4036; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10180 = 12'h3c4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7108; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13252 = 12'h3c4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10180; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16324 = 12'h3c4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13252; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19396 = 12'h3c4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16324; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22468 = 12'h3c4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19396; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25540 = 12'h3c4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22468; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_964 = io_valid_in ? _GEN_25540 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_964 = 12'h3c4 == _T_2[11:0] ? image_964 : _GEN_963; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4037 = 12'h3c5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7109 = 12'h3c5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4037; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10181 = 12'h3c5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7109; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13253 = 12'h3c5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10181; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16325 = 12'h3c5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13253; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19397 = 12'h3c5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16325; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22469 = 12'h3c5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19397; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25541 = 12'h3c5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22469; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_965 = io_valid_in ? _GEN_25541 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_965 = 12'h3c5 == _T_2[11:0] ? image_965 : _GEN_964; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4038 = 12'h3c6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7110 = 12'h3c6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4038; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10182 = 12'h3c6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7110; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13254 = 12'h3c6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10182; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16326 = 12'h3c6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13254; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19398 = 12'h3c6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16326; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22470 = 12'h3c6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19398; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25542 = 12'h3c6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22470; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_966 = io_valid_in ? _GEN_25542 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_966 = 12'h3c6 == _T_2[11:0] ? image_966 : _GEN_965; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4039 = 12'h3c7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7111 = 12'h3c7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4039; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10183 = 12'h3c7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7111; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13255 = 12'h3c7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10183; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16327 = 12'h3c7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13255; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19399 = 12'h3c7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16327; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22471 = 12'h3c7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19399; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25543 = 12'h3c7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22471; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_967 = io_valid_in ? _GEN_25543 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_967 = 12'h3c7 == _T_2[11:0] ? image_967 : _GEN_966; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4040 = 12'h3c8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7112 = 12'h3c8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4040; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10184 = 12'h3c8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7112; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13256 = 12'h3c8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10184; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16328 = 12'h3c8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13256; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19400 = 12'h3c8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16328; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22472 = 12'h3c8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19400; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25544 = 12'h3c8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22472; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_968 = io_valid_in ? _GEN_25544 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_968 = 12'h3c8 == _T_2[11:0] ? image_968 : _GEN_967; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4041 = 12'h3c9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7113 = 12'h3c9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4041; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10185 = 12'h3c9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7113; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13257 = 12'h3c9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10185; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16329 = 12'h3c9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13257; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19401 = 12'h3c9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16329; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22473 = 12'h3c9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19401; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25545 = 12'h3c9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22473; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_969 = io_valid_in ? _GEN_25545 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_969 = 12'h3c9 == _T_2[11:0] ? image_969 : _GEN_968; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4042 = 12'h3ca == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7114 = 12'h3ca == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4042; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10186 = 12'h3ca == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7114; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13258 = 12'h3ca == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10186; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16330 = 12'h3ca == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13258; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19402 = 12'h3ca == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16330; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22474 = 12'h3ca == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19402; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25546 = 12'h3ca == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22474; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_970 = io_valid_in ? _GEN_25546 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_970 = 12'h3ca == _T_2[11:0] ? image_970 : _GEN_969; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4043 = 12'h3cb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7115 = 12'h3cb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4043; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10187 = 12'h3cb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7115; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13259 = 12'h3cb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10187; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16331 = 12'h3cb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13259; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19403 = 12'h3cb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16331; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22475 = 12'h3cb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19403; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25547 = 12'h3cb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22475; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_971 = io_valid_in ? _GEN_25547 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_971 = 12'h3cb == _T_2[11:0] ? image_971 : _GEN_970; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4044 = 12'h3cc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7116 = 12'h3cc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4044; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10188 = 12'h3cc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7116; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13260 = 12'h3cc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10188; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16332 = 12'h3cc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13260; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19404 = 12'h3cc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16332; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22476 = 12'h3cc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19404; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25548 = 12'h3cc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22476; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_972 = io_valid_in ? _GEN_25548 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_972 = 12'h3cc == _T_2[11:0] ? image_972 : _GEN_971; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4045 = 12'h3cd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7117 = 12'h3cd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4045; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10189 = 12'h3cd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7117; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13261 = 12'h3cd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10189; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16333 = 12'h3cd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13261; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19405 = 12'h3cd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16333; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22477 = 12'h3cd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19405; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25549 = 12'h3cd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22477; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_973 = io_valid_in ? _GEN_25549 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_973 = 12'h3cd == _T_2[11:0] ? image_973 : _GEN_972; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4046 = 12'h3ce == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7118 = 12'h3ce == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4046; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10190 = 12'h3ce == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7118; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13262 = 12'h3ce == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10190; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16334 = 12'h3ce == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13262; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19406 = 12'h3ce == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16334; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22478 = 12'h3ce == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19406; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25550 = 12'h3ce == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22478; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_974 = io_valid_in ? _GEN_25550 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_974 = 12'h3ce == _T_2[11:0] ? image_974 : _GEN_973; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4047 = 12'h3cf == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7119 = 12'h3cf == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4047; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10191 = 12'h3cf == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7119; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13263 = 12'h3cf == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10191; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16335 = 12'h3cf == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13263; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19407 = 12'h3cf == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16335; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22479 = 12'h3cf == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19407; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25551 = 12'h3cf == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22479; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_975 = io_valid_in ? _GEN_25551 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_975 = 12'h3cf == _T_2[11:0] ? image_975 : _GEN_974; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4048 = 12'h3d0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7120 = 12'h3d0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4048; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10192 = 12'h3d0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7120; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13264 = 12'h3d0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10192; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16336 = 12'h3d0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13264; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19408 = 12'h3d0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16336; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22480 = 12'h3d0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19408; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25552 = 12'h3d0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22480; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_976 = io_valid_in ? _GEN_25552 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_976 = 12'h3d0 == _T_2[11:0] ? image_976 : _GEN_975; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4049 = 12'h3d1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7121 = 12'h3d1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4049; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10193 = 12'h3d1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7121; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13265 = 12'h3d1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10193; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16337 = 12'h3d1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13265; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19409 = 12'h3d1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16337; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22481 = 12'h3d1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19409; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25553 = 12'h3d1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22481; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_977 = io_valid_in ? _GEN_25553 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_977 = 12'h3d1 == _T_2[11:0] ? image_977 : _GEN_976; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4050 = 12'h3d2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7122 = 12'h3d2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4050; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10194 = 12'h3d2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7122; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13266 = 12'h3d2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10194; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16338 = 12'h3d2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13266; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19410 = 12'h3d2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16338; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22482 = 12'h3d2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19410; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25554 = 12'h3d2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22482; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_978 = io_valid_in ? _GEN_25554 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_978 = 12'h3d2 == _T_2[11:0] ? image_978 : _GEN_977; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4051 = 12'h3d3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7123 = 12'h3d3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4051; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10195 = 12'h3d3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7123; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13267 = 12'h3d3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10195; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16339 = 12'h3d3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13267; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19411 = 12'h3d3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16339; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22483 = 12'h3d3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19411; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25555 = 12'h3d3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22483; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_979 = io_valid_in ? _GEN_25555 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_979 = 12'h3d3 == _T_2[11:0] ? image_979 : _GEN_978; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4052 = 12'h3d4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7124 = 12'h3d4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4052; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10196 = 12'h3d4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7124; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13268 = 12'h3d4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10196; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16340 = 12'h3d4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13268; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19412 = 12'h3d4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16340; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22484 = 12'h3d4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19412; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25556 = 12'h3d4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22484; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_980 = io_valid_in ? _GEN_25556 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_980 = 12'h3d4 == _T_2[11:0] ? image_980 : _GEN_979; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4053 = 12'h3d5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7125 = 12'h3d5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4053; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10197 = 12'h3d5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7125; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13269 = 12'h3d5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10197; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16341 = 12'h3d5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13269; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19413 = 12'h3d5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16341; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22485 = 12'h3d5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19413; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25557 = 12'h3d5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22485; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_981 = io_valid_in ? _GEN_25557 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_981 = 12'h3d5 == _T_2[11:0] ? image_981 : _GEN_980; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4054 = 12'h3d6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7126 = 12'h3d6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4054; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10198 = 12'h3d6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7126; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13270 = 12'h3d6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10198; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16342 = 12'h3d6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13270; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19414 = 12'h3d6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16342; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22486 = 12'h3d6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19414; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25558 = 12'h3d6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22486; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_982 = io_valid_in ? _GEN_25558 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_982 = 12'h3d6 == _T_2[11:0] ? image_982 : _GEN_981; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4055 = 12'h3d7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7127 = 12'h3d7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4055; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10199 = 12'h3d7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7127; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13271 = 12'h3d7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10199; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16343 = 12'h3d7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13271; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19415 = 12'h3d7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16343; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22487 = 12'h3d7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19415; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25559 = 12'h3d7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22487; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_983 = io_valid_in ? _GEN_25559 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_983 = 12'h3d7 == _T_2[11:0] ? image_983 : _GEN_982; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4056 = 12'h3d8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7128 = 12'h3d8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4056; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10200 = 12'h3d8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7128; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13272 = 12'h3d8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10200; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16344 = 12'h3d8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13272; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19416 = 12'h3d8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16344; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22488 = 12'h3d8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19416; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25560 = 12'h3d8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22488; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_984 = io_valid_in ? _GEN_25560 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_984 = 12'h3d8 == _T_2[11:0] ? image_984 : _GEN_983; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4057 = 12'h3d9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7129 = 12'h3d9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4057; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10201 = 12'h3d9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7129; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13273 = 12'h3d9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10201; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16345 = 12'h3d9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13273; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19417 = 12'h3d9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16345; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22489 = 12'h3d9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19417; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25561 = 12'h3d9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22489; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_985 = io_valid_in ? _GEN_25561 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_985 = 12'h3d9 == _T_2[11:0] ? image_985 : _GEN_984; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4058 = 12'h3da == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7130 = 12'h3da == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4058; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10202 = 12'h3da == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7130; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13274 = 12'h3da == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10202; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16346 = 12'h3da == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13274; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19418 = 12'h3da == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16346; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22490 = 12'h3da == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19418; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25562 = 12'h3da == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22490; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_986 = io_valid_in ? _GEN_25562 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_986 = 12'h3da == _T_2[11:0] ? image_986 : _GEN_985; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4059 = 12'h3db == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7131 = 12'h3db == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4059; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10203 = 12'h3db == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7131; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13275 = 12'h3db == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10203; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16347 = 12'h3db == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13275; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19419 = 12'h3db == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16347; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22491 = 12'h3db == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19419; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25563 = 12'h3db == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22491; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_987 = io_valid_in ? _GEN_25563 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_987 = 12'h3db == _T_2[11:0] ? image_987 : _GEN_986; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4060 = 12'h3dc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7132 = 12'h3dc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4060; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10204 = 12'h3dc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7132; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13276 = 12'h3dc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10204; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16348 = 12'h3dc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13276; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19420 = 12'h3dc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16348; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22492 = 12'h3dc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19420; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25564 = 12'h3dc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22492; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_988 = io_valid_in ? _GEN_25564 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_988 = 12'h3dc == _T_2[11:0] ? image_988 : _GEN_987; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4061 = 12'h3dd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7133 = 12'h3dd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4061; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10205 = 12'h3dd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7133; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13277 = 12'h3dd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10205; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16349 = 12'h3dd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13277; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19421 = 12'h3dd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16349; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22493 = 12'h3dd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19421; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25565 = 12'h3dd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22493; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_989 = io_valid_in ? _GEN_25565 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_989 = 12'h3dd == _T_2[11:0] ? image_989 : _GEN_988; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4062 = 12'h3de == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7134 = 12'h3de == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4062; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10206 = 12'h3de == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7134; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13278 = 12'h3de == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10206; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16350 = 12'h3de == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13278; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19422 = 12'h3de == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16350; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22494 = 12'h3de == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19422; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25566 = 12'h3de == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22494; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_990 = io_valid_in ? _GEN_25566 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_990 = 12'h3de == _T_2[11:0] ? image_990 : _GEN_989; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4063 = 12'h3df == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7135 = 12'h3df == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4063; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10207 = 12'h3df == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7135; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13279 = 12'h3df == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10207; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16351 = 12'h3df == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13279; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19423 = 12'h3df == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16351; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22495 = 12'h3df == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19423; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25567 = 12'h3df == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22495; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_991 = io_valid_in ? _GEN_25567 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_991 = 12'h3df == _T_2[11:0] ? image_991 : _GEN_990; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4064 = 12'h3e0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7136 = 12'h3e0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4064; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10208 = 12'h3e0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7136; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13280 = 12'h3e0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10208; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16352 = 12'h3e0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13280; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19424 = 12'h3e0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16352; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22496 = 12'h3e0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19424; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25568 = 12'h3e0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22496; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_992 = io_valid_in ? _GEN_25568 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_992 = 12'h3e0 == _T_2[11:0] ? image_992 : _GEN_991; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4065 = 12'h3e1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7137 = 12'h3e1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4065; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10209 = 12'h3e1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7137; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13281 = 12'h3e1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10209; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16353 = 12'h3e1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13281; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19425 = 12'h3e1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16353; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22497 = 12'h3e1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19425; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25569 = 12'h3e1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22497; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_993 = io_valid_in ? _GEN_25569 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_993 = 12'h3e1 == _T_2[11:0] ? image_993 : _GEN_992; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4066 = 12'h3e2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7138 = 12'h3e2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4066; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10210 = 12'h3e2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7138; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13282 = 12'h3e2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10210; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16354 = 12'h3e2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13282; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19426 = 12'h3e2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16354; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22498 = 12'h3e2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19426; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25570 = 12'h3e2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22498; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_994 = io_valid_in ? _GEN_25570 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_994 = 12'h3e2 == _T_2[11:0] ? image_994 : _GEN_993; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4067 = 12'h3e3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7139 = 12'h3e3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4067; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10211 = 12'h3e3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7139; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13283 = 12'h3e3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10211; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16355 = 12'h3e3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13283; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19427 = 12'h3e3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16355; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22499 = 12'h3e3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19427; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25571 = 12'h3e3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22499; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_995 = io_valid_in ? _GEN_25571 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_995 = 12'h3e3 == _T_2[11:0] ? image_995 : _GEN_994; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4068 = 12'h3e4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7140 = 12'h3e4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4068; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10212 = 12'h3e4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7140; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13284 = 12'h3e4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10212; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16356 = 12'h3e4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13284; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19428 = 12'h3e4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16356; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22500 = 12'h3e4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19428; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25572 = 12'h3e4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22500; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_996 = io_valid_in ? _GEN_25572 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_996 = 12'h3e4 == _T_2[11:0] ? image_996 : _GEN_995; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4069 = 12'h3e5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7141 = 12'h3e5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4069; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10213 = 12'h3e5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7141; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13285 = 12'h3e5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10213; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16357 = 12'h3e5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13285; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19429 = 12'h3e5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16357; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22501 = 12'h3e5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19429; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25573 = 12'h3e5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22501; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_997 = io_valid_in ? _GEN_25573 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_997 = 12'h3e5 == _T_2[11:0] ? image_997 : _GEN_996; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4070 = 12'h3e6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7142 = 12'h3e6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4070; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10214 = 12'h3e6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7142; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13286 = 12'h3e6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10214; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16358 = 12'h3e6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13286; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19430 = 12'h3e6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16358; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22502 = 12'h3e6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19430; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25574 = 12'h3e6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22502; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_998 = io_valid_in ? _GEN_25574 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_998 = 12'h3e6 == _T_2[11:0] ? image_998 : _GEN_997; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4071 = 12'h3e7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7143 = 12'h3e7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4071; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10215 = 12'h3e7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7143; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13287 = 12'h3e7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10215; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16359 = 12'h3e7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13287; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19431 = 12'h3e7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16359; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22503 = 12'h3e7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19431; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25575 = 12'h3e7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22503; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_999 = io_valid_in ? _GEN_25575 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_999 = 12'h3e7 == _T_2[11:0] ? image_999 : _GEN_998; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4072 = 12'h3e8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7144 = 12'h3e8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4072; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10216 = 12'h3e8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7144; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13288 = 12'h3e8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10216; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16360 = 12'h3e8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13288; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19432 = 12'h3e8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16360; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22504 = 12'h3e8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19432; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25576 = 12'h3e8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22504; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1000 = io_valid_in ? _GEN_25576 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1000 = 12'h3e8 == _T_2[11:0] ? image_1000 : _GEN_999; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4073 = 12'h3e9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7145 = 12'h3e9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4073; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10217 = 12'h3e9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7145; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13289 = 12'h3e9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10217; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16361 = 12'h3e9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13289; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19433 = 12'h3e9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16361; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22505 = 12'h3e9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19433; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25577 = 12'h3e9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22505; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1001 = io_valid_in ? _GEN_25577 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1001 = 12'h3e9 == _T_2[11:0] ? image_1001 : _GEN_1000; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4074 = 12'h3ea == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7146 = 12'h3ea == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4074; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10218 = 12'h3ea == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7146; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13290 = 12'h3ea == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10218; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16362 = 12'h3ea == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13290; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19434 = 12'h3ea == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16362; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22506 = 12'h3ea == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19434; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25578 = 12'h3ea == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22506; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1002 = io_valid_in ? _GEN_25578 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1002 = 12'h3ea == _T_2[11:0] ? image_1002 : _GEN_1001; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4075 = 12'h3eb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7147 = 12'h3eb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4075; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10219 = 12'h3eb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7147; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13291 = 12'h3eb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10219; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16363 = 12'h3eb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13291; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19435 = 12'h3eb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16363; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22507 = 12'h3eb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19435; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25579 = 12'h3eb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22507; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1003 = io_valid_in ? _GEN_25579 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1003 = 12'h3eb == _T_2[11:0] ? image_1003 : _GEN_1002; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4076 = 12'h3ec == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7148 = 12'h3ec == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4076; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10220 = 12'h3ec == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7148; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13292 = 12'h3ec == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10220; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16364 = 12'h3ec == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13292; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19436 = 12'h3ec == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16364; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22508 = 12'h3ec == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19436; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25580 = 12'h3ec == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22508; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1004 = io_valid_in ? _GEN_25580 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1004 = 12'h3ec == _T_2[11:0] ? image_1004 : _GEN_1003; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4077 = 12'h3ed == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7149 = 12'h3ed == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4077; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10221 = 12'h3ed == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7149; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13293 = 12'h3ed == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10221; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16365 = 12'h3ed == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13293; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19437 = 12'h3ed == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16365; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22509 = 12'h3ed == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19437; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25581 = 12'h3ed == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22509; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1005 = io_valid_in ? _GEN_25581 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1005 = 12'h3ed == _T_2[11:0] ? image_1005 : _GEN_1004; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4078 = 12'h3ee == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7150 = 12'h3ee == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4078; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10222 = 12'h3ee == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7150; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13294 = 12'h3ee == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10222; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16366 = 12'h3ee == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13294; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19438 = 12'h3ee == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16366; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22510 = 12'h3ee == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19438; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25582 = 12'h3ee == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22510; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1006 = io_valid_in ? _GEN_25582 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1006 = 12'h3ee == _T_2[11:0] ? image_1006 : _GEN_1005; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4079 = 12'h3ef == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7151 = 12'h3ef == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4079; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10223 = 12'h3ef == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7151; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13295 = 12'h3ef == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10223; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16367 = 12'h3ef == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13295; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19439 = 12'h3ef == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16367; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22511 = 12'h3ef == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19439; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25583 = 12'h3ef == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22511; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1007 = io_valid_in ? _GEN_25583 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1007 = 12'h3ef == _T_2[11:0] ? image_1007 : _GEN_1006; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4080 = 12'h3f0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7152 = 12'h3f0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4080; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10224 = 12'h3f0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7152; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13296 = 12'h3f0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10224; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16368 = 12'h3f0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13296; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19440 = 12'h3f0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16368; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22512 = 12'h3f0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19440; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25584 = 12'h3f0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22512; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1008 = io_valid_in ? _GEN_25584 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1008 = 12'h3f0 == _T_2[11:0] ? image_1008 : _GEN_1007; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4081 = 12'h3f1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7153 = 12'h3f1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4081; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10225 = 12'h3f1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7153; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13297 = 12'h3f1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10225; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16369 = 12'h3f1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13297; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19441 = 12'h3f1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16369; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22513 = 12'h3f1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19441; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25585 = 12'h3f1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22513; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1009 = io_valid_in ? _GEN_25585 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1009 = 12'h3f1 == _T_2[11:0] ? image_1009 : _GEN_1008; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4082 = 12'h3f2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7154 = 12'h3f2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4082; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10226 = 12'h3f2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7154; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13298 = 12'h3f2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10226; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16370 = 12'h3f2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13298; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19442 = 12'h3f2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16370; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22514 = 12'h3f2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19442; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25586 = 12'h3f2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22514; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1010 = io_valid_in ? _GEN_25586 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1010 = 12'h3f2 == _T_2[11:0] ? image_1010 : _GEN_1009; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4083 = 12'h3f3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7155 = 12'h3f3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4083; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10227 = 12'h3f3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7155; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13299 = 12'h3f3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10227; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16371 = 12'h3f3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13299; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19443 = 12'h3f3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16371; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22515 = 12'h3f3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19443; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25587 = 12'h3f3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22515; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1011 = io_valid_in ? _GEN_25587 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1011 = 12'h3f3 == _T_2[11:0] ? image_1011 : _GEN_1010; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4084 = 12'h3f4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7156 = 12'h3f4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4084; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10228 = 12'h3f4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7156; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13300 = 12'h3f4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10228; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16372 = 12'h3f4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13300; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19444 = 12'h3f4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16372; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22516 = 12'h3f4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19444; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25588 = 12'h3f4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22516; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1012 = io_valid_in ? _GEN_25588 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1012 = 12'h3f4 == _T_2[11:0] ? image_1012 : _GEN_1011; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4085 = 12'h3f5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7157 = 12'h3f5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4085; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10229 = 12'h3f5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7157; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13301 = 12'h3f5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10229; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16373 = 12'h3f5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13301; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19445 = 12'h3f5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16373; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22517 = 12'h3f5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19445; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25589 = 12'h3f5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22517; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1013 = io_valid_in ? _GEN_25589 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1013 = 12'h3f5 == _T_2[11:0] ? image_1013 : _GEN_1012; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4086 = 12'h3f6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7158 = 12'h3f6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4086; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10230 = 12'h3f6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7158; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13302 = 12'h3f6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10230; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16374 = 12'h3f6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13302; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19446 = 12'h3f6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16374; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22518 = 12'h3f6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19446; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25590 = 12'h3f6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22518; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1014 = io_valid_in ? _GEN_25590 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1014 = 12'h3f6 == _T_2[11:0] ? image_1014 : _GEN_1013; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4087 = 12'h3f7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7159 = 12'h3f7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4087; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10231 = 12'h3f7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7159; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13303 = 12'h3f7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10231; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16375 = 12'h3f7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13303; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19447 = 12'h3f7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16375; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22519 = 12'h3f7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19447; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25591 = 12'h3f7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22519; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1015 = io_valid_in ? _GEN_25591 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1015 = 12'h3f7 == _T_2[11:0] ? image_1015 : _GEN_1014; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4088 = 12'h3f8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7160 = 12'h3f8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4088; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10232 = 12'h3f8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7160; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13304 = 12'h3f8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10232; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16376 = 12'h3f8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13304; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19448 = 12'h3f8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16376; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22520 = 12'h3f8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19448; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25592 = 12'h3f8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22520; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1016 = io_valid_in ? _GEN_25592 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1016 = 12'h3f8 == _T_2[11:0] ? image_1016 : _GEN_1015; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4089 = 12'h3f9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7161 = 12'h3f9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4089; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10233 = 12'h3f9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7161; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13305 = 12'h3f9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10233; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16377 = 12'h3f9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13305; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19449 = 12'h3f9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16377; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22521 = 12'h3f9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19449; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25593 = 12'h3f9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22521; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1017 = io_valid_in ? _GEN_25593 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1017 = 12'h3f9 == _T_2[11:0] ? image_1017 : _GEN_1016; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4090 = 12'h3fa == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7162 = 12'h3fa == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4090; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10234 = 12'h3fa == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7162; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13306 = 12'h3fa == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10234; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16378 = 12'h3fa == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13306; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19450 = 12'h3fa == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16378; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22522 = 12'h3fa == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19450; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25594 = 12'h3fa == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22522; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1018 = io_valid_in ? _GEN_25594 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1018 = 12'h3fa == _T_2[11:0] ? image_1018 : _GEN_1017; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4091 = 12'h3fb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7163 = 12'h3fb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4091; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10235 = 12'h3fb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7163; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13307 = 12'h3fb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10235; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16379 = 12'h3fb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13307; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19451 = 12'h3fb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16379; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22523 = 12'h3fb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19451; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25595 = 12'h3fb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22523; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1019 = io_valid_in ? _GEN_25595 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1019 = 12'h3fb == _T_2[11:0] ? image_1019 : _GEN_1018; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4092 = 12'h3fc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7164 = 12'h3fc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4092; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10236 = 12'h3fc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7164; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13308 = 12'h3fc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10236; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16380 = 12'h3fc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13308; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19452 = 12'h3fc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16380; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22524 = 12'h3fc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19452; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25596 = 12'h3fc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22524; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1020 = io_valid_in ? _GEN_25596 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1020 = 12'h3fc == _T_2[11:0] ? image_1020 : _GEN_1019; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4093 = 12'h3fd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7165 = 12'h3fd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4093; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10237 = 12'h3fd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7165; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13309 = 12'h3fd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10237; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16381 = 12'h3fd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13309; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19453 = 12'h3fd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16381; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22525 = 12'h3fd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19453; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25597 = 12'h3fd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22525; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1021 = io_valid_in ? _GEN_25597 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1021 = 12'h3fd == _T_2[11:0] ? image_1021 : _GEN_1020; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4094 = 12'h3fe == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7166 = 12'h3fe == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4094; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10238 = 12'h3fe == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7166; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13310 = 12'h3fe == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10238; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16382 = 12'h3fe == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13310; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19454 = 12'h3fe == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16382; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22526 = 12'h3fe == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19454; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25598 = 12'h3fe == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22526; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1022 = io_valid_in ? _GEN_25598 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1022 = 12'h3fe == _T_2[11:0] ? image_1022 : _GEN_1021; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4095 = 12'h3ff == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7167 = 12'h3ff == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4095; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10239 = 12'h3ff == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7167; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13311 = 12'h3ff == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10239; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16383 = 12'h3ff == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13311; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19455 = 12'h3ff == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16383; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22527 = 12'h3ff == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19455; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25599 = 12'h3ff == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22527; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1023 = io_valid_in ? _GEN_25599 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1023 = 12'h3ff == _T_2[11:0] ? image_1023 : _GEN_1022; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4096 = 12'h400 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7168 = 12'h400 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4096; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10240 = 12'h400 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7168; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13312 = 12'h400 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10240; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16384 = 12'h400 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13312; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19456 = 12'h400 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16384; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22528 = 12'h400 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19456; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25600 = 12'h400 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22528; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1024 = io_valid_in ? _GEN_25600 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1024 = 12'h400 == _T_2[11:0] ? image_1024 : _GEN_1023; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4097 = 12'h401 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7169 = 12'h401 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4097; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10241 = 12'h401 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7169; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13313 = 12'h401 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10241; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16385 = 12'h401 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13313; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19457 = 12'h401 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16385; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22529 = 12'h401 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19457; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25601 = 12'h401 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22529; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1025 = io_valid_in ? _GEN_25601 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1025 = 12'h401 == _T_2[11:0] ? image_1025 : _GEN_1024; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4098 = 12'h402 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7170 = 12'h402 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4098; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10242 = 12'h402 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7170; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13314 = 12'h402 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10242; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16386 = 12'h402 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13314; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19458 = 12'h402 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16386; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22530 = 12'h402 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19458; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25602 = 12'h402 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22530; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1026 = io_valid_in ? _GEN_25602 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1026 = 12'h402 == _T_2[11:0] ? image_1026 : _GEN_1025; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4099 = 12'h403 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7171 = 12'h403 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4099; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10243 = 12'h403 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7171; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13315 = 12'h403 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10243; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16387 = 12'h403 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13315; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19459 = 12'h403 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16387; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22531 = 12'h403 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19459; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25603 = 12'h403 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22531; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1027 = io_valid_in ? _GEN_25603 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1027 = 12'h403 == _T_2[11:0] ? image_1027 : _GEN_1026; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4100 = 12'h404 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7172 = 12'h404 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4100; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10244 = 12'h404 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7172; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13316 = 12'h404 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10244; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16388 = 12'h404 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13316; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19460 = 12'h404 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16388; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22532 = 12'h404 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19460; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25604 = 12'h404 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22532; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1028 = io_valid_in ? _GEN_25604 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1028 = 12'h404 == _T_2[11:0] ? image_1028 : _GEN_1027; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4101 = 12'h405 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7173 = 12'h405 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4101; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10245 = 12'h405 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7173; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13317 = 12'h405 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10245; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16389 = 12'h405 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13317; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19461 = 12'h405 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16389; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22533 = 12'h405 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19461; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25605 = 12'h405 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22533; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1029 = io_valid_in ? _GEN_25605 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1029 = 12'h405 == _T_2[11:0] ? image_1029 : _GEN_1028; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4102 = 12'h406 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7174 = 12'h406 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4102; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10246 = 12'h406 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7174; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13318 = 12'h406 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10246; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16390 = 12'h406 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13318; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19462 = 12'h406 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16390; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22534 = 12'h406 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19462; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25606 = 12'h406 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22534; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1030 = io_valid_in ? _GEN_25606 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1030 = 12'h406 == _T_2[11:0] ? image_1030 : _GEN_1029; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4103 = 12'h407 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7175 = 12'h407 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4103; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10247 = 12'h407 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7175; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13319 = 12'h407 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10247; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16391 = 12'h407 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13319; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19463 = 12'h407 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16391; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22535 = 12'h407 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19463; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25607 = 12'h407 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22535; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1031 = io_valid_in ? _GEN_25607 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1031 = 12'h407 == _T_2[11:0] ? image_1031 : _GEN_1030; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4104 = 12'h408 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7176 = 12'h408 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4104; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10248 = 12'h408 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7176; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13320 = 12'h408 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10248; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16392 = 12'h408 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13320; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19464 = 12'h408 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16392; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22536 = 12'h408 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19464; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25608 = 12'h408 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22536; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1032 = io_valid_in ? _GEN_25608 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1032 = 12'h408 == _T_2[11:0] ? image_1032 : _GEN_1031; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4105 = 12'h409 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7177 = 12'h409 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4105; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10249 = 12'h409 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7177; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13321 = 12'h409 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10249; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16393 = 12'h409 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13321; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19465 = 12'h409 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16393; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22537 = 12'h409 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19465; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25609 = 12'h409 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22537; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1033 = io_valid_in ? _GEN_25609 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1033 = 12'h409 == _T_2[11:0] ? image_1033 : _GEN_1032; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4106 = 12'h40a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7178 = 12'h40a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4106; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10250 = 12'h40a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7178; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13322 = 12'h40a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10250; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16394 = 12'h40a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13322; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19466 = 12'h40a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16394; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22538 = 12'h40a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19466; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25610 = 12'h40a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22538; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1034 = io_valid_in ? _GEN_25610 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1034 = 12'h40a == _T_2[11:0] ? image_1034 : _GEN_1033; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4107 = 12'h40b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7179 = 12'h40b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4107; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10251 = 12'h40b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7179; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13323 = 12'h40b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10251; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16395 = 12'h40b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13323; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19467 = 12'h40b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16395; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22539 = 12'h40b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19467; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25611 = 12'h40b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22539; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1035 = io_valid_in ? _GEN_25611 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1035 = 12'h40b == _T_2[11:0] ? image_1035 : _GEN_1034; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4108 = 12'h40c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7180 = 12'h40c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4108; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10252 = 12'h40c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7180; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13324 = 12'h40c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10252; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16396 = 12'h40c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13324; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19468 = 12'h40c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16396; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22540 = 12'h40c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19468; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25612 = 12'h40c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22540; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1036 = io_valid_in ? _GEN_25612 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1036 = 12'h40c == _T_2[11:0] ? image_1036 : _GEN_1035; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4109 = 12'h40d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7181 = 12'h40d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4109; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10253 = 12'h40d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7181; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13325 = 12'h40d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10253; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16397 = 12'h40d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13325; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19469 = 12'h40d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16397; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22541 = 12'h40d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19469; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25613 = 12'h40d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22541; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1037 = io_valid_in ? _GEN_25613 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1037 = 12'h40d == _T_2[11:0] ? image_1037 : _GEN_1036; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4110 = 12'h40e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7182 = 12'h40e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4110; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10254 = 12'h40e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7182; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13326 = 12'h40e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10254; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16398 = 12'h40e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13326; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19470 = 12'h40e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16398; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22542 = 12'h40e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19470; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25614 = 12'h40e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22542; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1038 = io_valid_in ? _GEN_25614 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1038 = 12'h40e == _T_2[11:0] ? image_1038 : _GEN_1037; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4111 = 12'h40f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7183 = 12'h40f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4111; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10255 = 12'h40f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7183; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13327 = 12'h40f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10255; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16399 = 12'h40f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13327; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19471 = 12'h40f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16399; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22543 = 12'h40f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19471; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25615 = 12'h40f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22543; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1039 = io_valid_in ? _GEN_25615 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1039 = 12'h40f == _T_2[11:0] ? image_1039 : _GEN_1038; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4112 = 12'h410 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7184 = 12'h410 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4112; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10256 = 12'h410 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7184; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13328 = 12'h410 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10256; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16400 = 12'h410 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13328; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19472 = 12'h410 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16400; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22544 = 12'h410 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19472; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25616 = 12'h410 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22544; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1040 = io_valid_in ? _GEN_25616 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1040 = 12'h410 == _T_2[11:0] ? image_1040 : _GEN_1039; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4113 = 12'h411 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7185 = 12'h411 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4113; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10257 = 12'h411 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7185; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13329 = 12'h411 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10257; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16401 = 12'h411 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13329; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19473 = 12'h411 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16401; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22545 = 12'h411 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19473; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25617 = 12'h411 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22545; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1041 = io_valid_in ? _GEN_25617 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1041 = 12'h411 == _T_2[11:0] ? image_1041 : _GEN_1040; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4114 = 12'h412 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7186 = 12'h412 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4114; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10258 = 12'h412 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7186; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13330 = 12'h412 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10258; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16402 = 12'h412 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13330; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19474 = 12'h412 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16402; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22546 = 12'h412 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19474; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25618 = 12'h412 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22546; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1042 = io_valid_in ? _GEN_25618 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1042 = 12'h412 == _T_2[11:0] ? image_1042 : _GEN_1041; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4115 = 12'h413 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7187 = 12'h413 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4115; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10259 = 12'h413 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7187; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13331 = 12'h413 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10259; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16403 = 12'h413 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13331; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19475 = 12'h413 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16403; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22547 = 12'h413 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19475; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25619 = 12'h413 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22547; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1043 = io_valid_in ? _GEN_25619 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1043 = 12'h413 == _T_2[11:0] ? image_1043 : _GEN_1042; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4116 = 12'h414 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7188 = 12'h414 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4116; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10260 = 12'h414 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7188; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13332 = 12'h414 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10260; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16404 = 12'h414 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13332; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19476 = 12'h414 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16404; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22548 = 12'h414 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19476; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25620 = 12'h414 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22548; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1044 = io_valid_in ? _GEN_25620 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1044 = 12'h414 == _T_2[11:0] ? image_1044 : _GEN_1043; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4117 = 12'h415 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7189 = 12'h415 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4117; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10261 = 12'h415 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7189; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13333 = 12'h415 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10261; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16405 = 12'h415 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13333; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19477 = 12'h415 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16405; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22549 = 12'h415 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19477; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25621 = 12'h415 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22549; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1045 = io_valid_in ? _GEN_25621 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1045 = 12'h415 == _T_2[11:0] ? image_1045 : _GEN_1044; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4118 = 12'h416 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7190 = 12'h416 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4118; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10262 = 12'h416 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7190; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13334 = 12'h416 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10262; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16406 = 12'h416 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13334; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19478 = 12'h416 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16406; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22550 = 12'h416 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19478; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25622 = 12'h416 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22550; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1046 = io_valid_in ? _GEN_25622 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1046 = 12'h416 == _T_2[11:0] ? image_1046 : _GEN_1045; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4119 = 12'h417 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7191 = 12'h417 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4119; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10263 = 12'h417 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7191; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13335 = 12'h417 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10263; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16407 = 12'h417 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13335; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19479 = 12'h417 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16407; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22551 = 12'h417 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19479; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25623 = 12'h417 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22551; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1047 = io_valid_in ? _GEN_25623 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1047 = 12'h417 == _T_2[11:0] ? image_1047 : _GEN_1046; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4120 = 12'h418 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7192 = 12'h418 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4120; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10264 = 12'h418 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7192; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13336 = 12'h418 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10264; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16408 = 12'h418 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13336; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19480 = 12'h418 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16408; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22552 = 12'h418 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19480; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25624 = 12'h418 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22552; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1048 = io_valid_in ? _GEN_25624 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1048 = 12'h418 == _T_2[11:0] ? image_1048 : _GEN_1047; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4121 = 12'h419 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7193 = 12'h419 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4121; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10265 = 12'h419 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7193; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13337 = 12'h419 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10265; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16409 = 12'h419 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13337; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19481 = 12'h419 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16409; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22553 = 12'h419 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19481; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25625 = 12'h419 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22553; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1049 = io_valid_in ? _GEN_25625 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1049 = 12'h419 == _T_2[11:0] ? image_1049 : _GEN_1048; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4122 = 12'h41a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7194 = 12'h41a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4122; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10266 = 12'h41a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7194; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13338 = 12'h41a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10266; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16410 = 12'h41a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13338; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19482 = 12'h41a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16410; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22554 = 12'h41a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19482; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25626 = 12'h41a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22554; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1050 = io_valid_in ? _GEN_25626 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1050 = 12'h41a == _T_2[11:0] ? image_1050 : _GEN_1049; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4123 = 12'h41b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7195 = 12'h41b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4123; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10267 = 12'h41b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7195; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13339 = 12'h41b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10267; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16411 = 12'h41b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13339; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19483 = 12'h41b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16411; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22555 = 12'h41b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19483; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25627 = 12'h41b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22555; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1051 = io_valid_in ? _GEN_25627 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1051 = 12'h41b == _T_2[11:0] ? image_1051 : _GEN_1050; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4124 = 12'h41c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7196 = 12'h41c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4124; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10268 = 12'h41c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7196; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13340 = 12'h41c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10268; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16412 = 12'h41c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13340; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19484 = 12'h41c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16412; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22556 = 12'h41c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19484; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25628 = 12'h41c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22556; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1052 = io_valid_in ? _GEN_25628 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1052 = 12'h41c == _T_2[11:0] ? image_1052 : _GEN_1051; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4125 = 12'h41d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7197 = 12'h41d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4125; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10269 = 12'h41d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7197; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13341 = 12'h41d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10269; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16413 = 12'h41d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13341; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19485 = 12'h41d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16413; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22557 = 12'h41d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19485; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25629 = 12'h41d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22557; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1053 = io_valid_in ? _GEN_25629 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1053 = 12'h41d == _T_2[11:0] ? image_1053 : _GEN_1052; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4126 = 12'h41e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7198 = 12'h41e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4126; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10270 = 12'h41e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7198; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13342 = 12'h41e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10270; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16414 = 12'h41e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13342; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19486 = 12'h41e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16414; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22558 = 12'h41e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19486; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25630 = 12'h41e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22558; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1054 = io_valid_in ? _GEN_25630 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1054 = 12'h41e == _T_2[11:0] ? image_1054 : _GEN_1053; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4127 = 12'h41f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7199 = 12'h41f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4127; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10271 = 12'h41f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7199; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13343 = 12'h41f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10271; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16415 = 12'h41f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13343; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19487 = 12'h41f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16415; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22559 = 12'h41f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19487; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25631 = 12'h41f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22559; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1055 = io_valid_in ? _GEN_25631 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1055 = 12'h41f == _T_2[11:0] ? image_1055 : _GEN_1054; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4128 = 12'h420 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7200 = 12'h420 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4128; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10272 = 12'h420 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7200; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13344 = 12'h420 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10272; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16416 = 12'h420 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13344; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19488 = 12'h420 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16416; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22560 = 12'h420 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19488; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25632 = 12'h420 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22560; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1056 = io_valid_in ? _GEN_25632 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1056 = 12'h420 == _T_2[11:0] ? image_1056 : _GEN_1055; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4129 = 12'h421 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7201 = 12'h421 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4129; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10273 = 12'h421 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7201; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13345 = 12'h421 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10273; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16417 = 12'h421 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13345; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19489 = 12'h421 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16417; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22561 = 12'h421 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19489; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25633 = 12'h421 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22561; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1057 = io_valid_in ? _GEN_25633 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1057 = 12'h421 == _T_2[11:0] ? image_1057 : _GEN_1056; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4130 = 12'h422 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7202 = 12'h422 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4130; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10274 = 12'h422 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7202; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13346 = 12'h422 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10274; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16418 = 12'h422 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13346; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19490 = 12'h422 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16418; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22562 = 12'h422 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19490; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25634 = 12'h422 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22562; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1058 = io_valid_in ? _GEN_25634 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1058 = 12'h422 == _T_2[11:0] ? image_1058 : _GEN_1057; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4131 = 12'h423 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7203 = 12'h423 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4131; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10275 = 12'h423 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7203; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13347 = 12'h423 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10275; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16419 = 12'h423 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13347; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19491 = 12'h423 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16419; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22563 = 12'h423 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19491; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25635 = 12'h423 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22563; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1059 = io_valid_in ? _GEN_25635 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1059 = 12'h423 == _T_2[11:0] ? image_1059 : _GEN_1058; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4132 = 12'h424 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7204 = 12'h424 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4132; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10276 = 12'h424 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7204; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13348 = 12'h424 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10276; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16420 = 12'h424 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13348; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19492 = 12'h424 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16420; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22564 = 12'h424 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19492; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25636 = 12'h424 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22564; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1060 = io_valid_in ? _GEN_25636 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1060 = 12'h424 == _T_2[11:0] ? image_1060 : _GEN_1059; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4133 = 12'h425 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7205 = 12'h425 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4133; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10277 = 12'h425 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7205; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13349 = 12'h425 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10277; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16421 = 12'h425 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13349; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19493 = 12'h425 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16421; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22565 = 12'h425 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19493; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25637 = 12'h425 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22565; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1061 = io_valid_in ? _GEN_25637 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1061 = 12'h425 == _T_2[11:0] ? image_1061 : _GEN_1060; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4134 = 12'h426 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7206 = 12'h426 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4134; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10278 = 12'h426 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7206; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13350 = 12'h426 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10278; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16422 = 12'h426 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13350; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19494 = 12'h426 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16422; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22566 = 12'h426 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19494; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25638 = 12'h426 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22566; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1062 = io_valid_in ? _GEN_25638 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1062 = 12'h426 == _T_2[11:0] ? image_1062 : _GEN_1061; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4135 = 12'h427 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7207 = 12'h427 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4135; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10279 = 12'h427 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7207; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13351 = 12'h427 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10279; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16423 = 12'h427 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13351; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19495 = 12'h427 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16423; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22567 = 12'h427 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19495; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25639 = 12'h427 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22567; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1063 = io_valid_in ? _GEN_25639 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1063 = 12'h427 == _T_2[11:0] ? image_1063 : _GEN_1062; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4136 = 12'h428 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7208 = 12'h428 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4136; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10280 = 12'h428 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7208; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13352 = 12'h428 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10280; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16424 = 12'h428 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13352; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19496 = 12'h428 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16424; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22568 = 12'h428 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19496; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25640 = 12'h428 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22568; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1064 = io_valid_in ? _GEN_25640 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1064 = 12'h428 == _T_2[11:0] ? image_1064 : _GEN_1063; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4137 = 12'h429 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7209 = 12'h429 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4137; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10281 = 12'h429 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7209; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13353 = 12'h429 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10281; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16425 = 12'h429 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13353; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19497 = 12'h429 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16425; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22569 = 12'h429 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19497; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25641 = 12'h429 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22569; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1065 = io_valid_in ? _GEN_25641 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1065 = 12'h429 == _T_2[11:0] ? image_1065 : _GEN_1064; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4138 = 12'h42a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7210 = 12'h42a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4138; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10282 = 12'h42a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7210; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13354 = 12'h42a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10282; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16426 = 12'h42a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13354; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19498 = 12'h42a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16426; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22570 = 12'h42a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19498; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25642 = 12'h42a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22570; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1066 = io_valid_in ? _GEN_25642 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1066 = 12'h42a == _T_2[11:0] ? image_1066 : _GEN_1065; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4139 = 12'h42b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7211 = 12'h42b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4139; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10283 = 12'h42b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7211; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13355 = 12'h42b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10283; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16427 = 12'h42b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13355; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19499 = 12'h42b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16427; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22571 = 12'h42b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19499; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25643 = 12'h42b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22571; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1067 = io_valid_in ? _GEN_25643 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1067 = 12'h42b == _T_2[11:0] ? image_1067 : _GEN_1066; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4140 = 12'h42c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7212 = 12'h42c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4140; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10284 = 12'h42c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7212; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13356 = 12'h42c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10284; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16428 = 12'h42c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13356; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19500 = 12'h42c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16428; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22572 = 12'h42c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19500; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25644 = 12'h42c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22572; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1068 = io_valid_in ? _GEN_25644 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1068 = 12'h42c == _T_2[11:0] ? image_1068 : _GEN_1067; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4141 = 12'h42d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7213 = 12'h42d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4141; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10285 = 12'h42d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7213; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13357 = 12'h42d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10285; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16429 = 12'h42d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13357; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19501 = 12'h42d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16429; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22573 = 12'h42d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19501; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25645 = 12'h42d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22573; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1069 = io_valid_in ? _GEN_25645 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1069 = 12'h42d == _T_2[11:0] ? image_1069 : _GEN_1068; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4142 = 12'h42e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7214 = 12'h42e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4142; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10286 = 12'h42e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7214; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13358 = 12'h42e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10286; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16430 = 12'h42e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13358; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19502 = 12'h42e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16430; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22574 = 12'h42e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19502; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25646 = 12'h42e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22574; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1070 = io_valid_in ? _GEN_25646 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1070 = 12'h42e == _T_2[11:0] ? image_1070 : _GEN_1069; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4143 = 12'h42f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7215 = 12'h42f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4143; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10287 = 12'h42f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7215; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13359 = 12'h42f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10287; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16431 = 12'h42f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13359; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19503 = 12'h42f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16431; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22575 = 12'h42f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19503; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25647 = 12'h42f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22575; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1071 = io_valid_in ? _GEN_25647 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1071 = 12'h42f == _T_2[11:0] ? image_1071 : _GEN_1070; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4144 = 12'h430 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7216 = 12'h430 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4144; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10288 = 12'h430 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7216; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13360 = 12'h430 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10288; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16432 = 12'h430 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13360; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19504 = 12'h430 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16432; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22576 = 12'h430 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19504; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25648 = 12'h430 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22576; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1072 = io_valid_in ? _GEN_25648 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1072 = 12'h430 == _T_2[11:0] ? image_1072 : _GEN_1071; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4145 = 12'h431 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7217 = 12'h431 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4145; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10289 = 12'h431 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7217; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13361 = 12'h431 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10289; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16433 = 12'h431 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13361; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19505 = 12'h431 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16433; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22577 = 12'h431 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19505; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25649 = 12'h431 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22577; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1073 = io_valid_in ? _GEN_25649 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1073 = 12'h431 == _T_2[11:0] ? image_1073 : _GEN_1072; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4146 = 12'h432 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7218 = 12'h432 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4146; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10290 = 12'h432 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7218; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13362 = 12'h432 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10290; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16434 = 12'h432 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13362; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19506 = 12'h432 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16434; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22578 = 12'h432 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19506; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25650 = 12'h432 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22578; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1074 = io_valid_in ? _GEN_25650 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1074 = 12'h432 == _T_2[11:0] ? image_1074 : _GEN_1073; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4147 = 12'h433 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7219 = 12'h433 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4147; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10291 = 12'h433 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7219; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13363 = 12'h433 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10291; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16435 = 12'h433 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13363; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19507 = 12'h433 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16435; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22579 = 12'h433 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19507; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25651 = 12'h433 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22579; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1075 = io_valid_in ? _GEN_25651 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1075 = 12'h433 == _T_2[11:0] ? image_1075 : _GEN_1074; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4148 = 12'h434 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7220 = 12'h434 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4148; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10292 = 12'h434 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7220; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13364 = 12'h434 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10292; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16436 = 12'h434 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13364; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19508 = 12'h434 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16436; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22580 = 12'h434 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19508; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25652 = 12'h434 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22580; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1076 = io_valid_in ? _GEN_25652 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1076 = 12'h434 == _T_2[11:0] ? image_1076 : _GEN_1075; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4149 = 12'h435 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7221 = 12'h435 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4149; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10293 = 12'h435 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7221; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13365 = 12'h435 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10293; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16437 = 12'h435 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13365; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19509 = 12'h435 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16437; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22581 = 12'h435 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19509; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25653 = 12'h435 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22581; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1077 = io_valid_in ? _GEN_25653 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1077 = 12'h435 == _T_2[11:0] ? image_1077 : _GEN_1076; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4150 = 12'h436 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7222 = 12'h436 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4150; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10294 = 12'h436 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7222; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13366 = 12'h436 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10294; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16438 = 12'h436 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13366; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19510 = 12'h436 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16438; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22582 = 12'h436 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19510; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25654 = 12'h436 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22582; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1078 = io_valid_in ? _GEN_25654 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1078 = 12'h436 == _T_2[11:0] ? image_1078 : _GEN_1077; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4151 = 12'h437 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7223 = 12'h437 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4151; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10295 = 12'h437 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7223; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13367 = 12'h437 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10295; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16439 = 12'h437 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13367; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19511 = 12'h437 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16439; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22583 = 12'h437 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19511; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25655 = 12'h437 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22583; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1079 = io_valid_in ? _GEN_25655 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1079 = 12'h437 == _T_2[11:0] ? image_1079 : _GEN_1078; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4152 = 12'h438 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7224 = 12'h438 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4152; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10296 = 12'h438 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7224; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13368 = 12'h438 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10296; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16440 = 12'h438 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13368; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19512 = 12'h438 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16440; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22584 = 12'h438 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19512; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25656 = 12'h438 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22584; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1080 = io_valid_in ? _GEN_25656 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1080 = 12'h438 == _T_2[11:0] ? image_1080 : _GEN_1079; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4153 = 12'h439 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7225 = 12'h439 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4153; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10297 = 12'h439 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7225; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13369 = 12'h439 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10297; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16441 = 12'h439 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13369; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19513 = 12'h439 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16441; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22585 = 12'h439 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19513; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25657 = 12'h439 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22585; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1081 = io_valid_in ? _GEN_25657 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1081 = 12'h439 == _T_2[11:0] ? image_1081 : _GEN_1080; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4154 = 12'h43a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7226 = 12'h43a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4154; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10298 = 12'h43a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7226; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13370 = 12'h43a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10298; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16442 = 12'h43a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13370; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19514 = 12'h43a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16442; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22586 = 12'h43a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19514; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25658 = 12'h43a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22586; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1082 = io_valid_in ? _GEN_25658 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1082 = 12'h43a == _T_2[11:0] ? image_1082 : _GEN_1081; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4155 = 12'h43b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7227 = 12'h43b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4155; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10299 = 12'h43b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7227; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13371 = 12'h43b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10299; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16443 = 12'h43b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13371; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19515 = 12'h43b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16443; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22587 = 12'h43b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19515; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25659 = 12'h43b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22587; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1083 = io_valid_in ? _GEN_25659 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1083 = 12'h43b == _T_2[11:0] ? image_1083 : _GEN_1082; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4156 = 12'h43c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7228 = 12'h43c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4156; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10300 = 12'h43c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7228; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13372 = 12'h43c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10300; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16444 = 12'h43c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13372; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19516 = 12'h43c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16444; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22588 = 12'h43c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19516; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25660 = 12'h43c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22588; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1084 = io_valid_in ? _GEN_25660 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1084 = 12'h43c == _T_2[11:0] ? image_1084 : _GEN_1083; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4157 = 12'h43d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7229 = 12'h43d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4157; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10301 = 12'h43d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7229; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13373 = 12'h43d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10301; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16445 = 12'h43d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13373; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19517 = 12'h43d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16445; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22589 = 12'h43d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19517; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25661 = 12'h43d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22589; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1085 = io_valid_in ? _GEN_25661 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1085 = 12'h43d == _T_2[11:0] ? image_1085 : _GEN_1084; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4158 = 12'h43e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7230 = 12'h43e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4158; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10302 = 12'h43e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7230; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13374 = 12'h43e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10302; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16446 = 12'h43e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13374; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19518 = 12'h43e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16446; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22590 = 12'h43e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19518; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25662 = 12'h43e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22590; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1086 = io_valid_in ? _GEN_25662 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1086 = 12'h43e == _T_2[11:0] ? image_1086 : _GEN_1085; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4159 = 12'h43f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7231 = 12'h43f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4159; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10303 = 12'h43f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7231; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13375 = 12'h43f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10303; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16447 = 12'h43f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13375; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19519 = 12'h43f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16447; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22591 = 12'h43f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19519; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25663 = 12'h43f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22591; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1087 = io_valid_in ? _GEN_25663 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1087 = 12'h43f == _T_2[11:0] ? image_1087 : _GEN_1086; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4160 = 12'h440 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7232 = 12'h440 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4160; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10304 = 12'h440 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7232; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13376 = 12'h440 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10304; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16448 = 12'h440 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13376; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19520 = 12'h440 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16448; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22592 = 12'h440 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19520; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25664 = 12'h440 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22592; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1088 = io_valid_in ? _GEN_25664 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1088 = 12'h440 == _T_2[11:0] ? image_1088 : _GEN_1087; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4161 = 12'h441 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7233 = 12'h441 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4161; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10305 = 12'h441 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7233; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13377 = 12'h441 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10305; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16449 = 12'h441 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13377; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19521 = 12'h441 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16449; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22593 = 12'h441 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19521; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25665 = 12'h441 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22593; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1089 = io_valid_in ? _GEN_25665 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1089 = 12'h441 == _T_2[11:0] ? image_1089 : _GEN_1088; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4162 = 12'h442 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7234 = 12'h442 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4162; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10306 = 12'h442 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7234; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13378 = 12'h442 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10306; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16450 = 12'h442 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13378; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19522 = 12'h442 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16450; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22594 = 12'h442 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19522; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25666 = 12'h442 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22594; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1090 = io_valid_in ? _GEN_25666 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1090 = 12'h442 == _T_2[11:0] ? image_1090 : _GEN_1089; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4163 = 12'h443 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7235 = 12'h443 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4163; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10307 = 12'h443 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7235; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13379 = 12'h443 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10307; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16451 = 12'h443 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13379; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19523 = 12'h443 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16451; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22595 = 12'h443 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19523; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25667 = 12'h443 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22595; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1091 = io_valid_in ? _GEN_25667 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1091 = 12'h443 == _T_2[11:0] ? image_1091 : _GEN_1090; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4164 = 12'h444 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7236 = 12'h444 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4164; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10308 = 12'h444 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7236; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13380 = 12'h444 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10308; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16452 = 12'h444 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13380; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19524 = 12'h444 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16452; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22596 = 12'h444 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19524; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25668 = 12'h444 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22596; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1092 = io_valid_in ? _GEN_25668 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1092 = 12'h444 == _T_2[11:0] ? image_1092 : _GEN_1091; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4165 = 12'h445 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7237 = 12'h445 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4165; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10309 = 12'h445 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7237; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13381 = 12'h445 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10309; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16453 = 12'h445 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13381; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19525 = 12'h445 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16453; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22597 = 12'h445 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19525; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25669 = 12'h445 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22597; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1093 = io_valid_in ? _GEN_25669 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1093 = 12'h445 == _T_2[11:0] ? image_1093 : _GEN_1092; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4166 = 12'h446 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7238 = 12'h446 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4166; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10310 = 12'h446 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7238; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13382 = 12'h446 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10310; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16454 = 12'h446 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13382; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19526 = 12'h446 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16454; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22598 = 12'h446 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19526; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25670 = 12'h446 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22598; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1094 = io_valid_in ? _GEN_25670 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1094 = 12'h446 == _T_2[11:0] ? image_1094 : _GEN_1093; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4167 = 12'h447 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7239 = 12'h447 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4167; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10311 = 12'h447 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7239; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13383 = 12'h447 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10311; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16455 = 12'h447 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13383; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19527 = 12'h447 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16455; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22599 = 12'h447 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19527; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25671 = 12'h447 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22599; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1095 = io_valid_in ? _GEN_25671 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1095 = 12'h447 == _T_2[11:0] ? image_1095 : _GEN_1094; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4168 = 12'h448 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7240 = 12'h448 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4168; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10312 = 12'h448 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7240; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13384 = 12'h448 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10312; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16456 = 12'h448 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13384; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19528 = 12'h448 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16456; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22600 = 12'h448 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19528; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25672 = 12'h448 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22600; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1096 = io_valid_in ? _GEN_25672 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1096 = 12'h448 == _T_2[11:0] ? image_1096 : _GEN_1095; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4169 = 12'h449 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7241 = 12'h449 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4169; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10313 = 12'h449 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7241; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13385 = 12'h449 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10313; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16457 = 12'h449 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13385; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19529 = 12'h449 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16457; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22601 = 12'h449 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19529; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25673 = 12'h449 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22601; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1097 = io_valid_in ? _GEN_25673 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1097 = 12'h449 == _T_2[11:0] ? image_1097 : _GEN_1096; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4170 = 12'h44a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7242 = 12'h44a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4170; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10314 = 12'h44a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7242; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13386 = 12'h44a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10314; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16458 = 12'h44a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13386; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19530 = 12'h44a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16458; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22602 = 12'h44a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19530; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25674 = 12'h44a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22602; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1098 = io_valid_in ? _GEN_25674 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1098 = 12'h44a == _T_2[11:0] ? image_1098 : _GEN_1097; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4171 = 12'h44b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7243 = 12'h44b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4171; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10315 = 12'h44b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7243; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13387 = 12'h44b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10315; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16459 = 12'h44b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13387; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19531 = 12'h44b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16459; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22603 = 12'h44b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19531; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25675 = 12'h44b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22603; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1099 = io_valid_in ? _GEN_25675 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1099 = 12'h44b == _T_2[11:0] ? image_1099 : _GEN_1098; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4172 = 12'h44c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7244 = 12'h44c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4172; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10316 = 12'h44c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7244; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13388 = 12'h44c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10316; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16460 = 12'h44c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13388; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19532 = 12'h44c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16460; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22604 = 12'h44c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19532; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25676 = 12'h44c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22604; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1100 = io_valid_in ? _GEN_25676 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1100 = 12'h44c == _T_2[11:0] ? image_1100 : _GEN_1099; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4173 = 12'h44d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7245 = 12'h44d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4173; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10317 = 12'h44d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7245; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13389 = 12'h44d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10317; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16461 = 12'h44d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13389; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19533 = 12'h44d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16461; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22605 = 12'h44d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19533; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25677 = 12'h44d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22605; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1101 = io_valid_in ? _GEN_25677 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1101 = 12'h44d == _T_2[11:0] ? image_1101 : _GEN_1100; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4174 = 12'h44e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7246 = 12'h44e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4174; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10318 = 12'h44e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7246; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13390 = 12'h44e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10318; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16462 = 12'h44e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13390; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19534 = 12'h44e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16462; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22606 = 12'h44e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19534; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25678 = 12'h44e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22606; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1102 = io_valid_in ? _GEN_25678 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1102 = 12'h44e == _T_2[11:0] ? image_1102 : _GEN_1101; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4175 = 12'h44f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7247 = 12'h44f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4175; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10319 = 12'h44f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7247; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13391 = 12'h44f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10319; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16463 = 12'h44f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13391; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19535 = 12'h44f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16463; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22607 = 12'h44f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19535; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25679 = 12'h44f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22607; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1103 = io_valid_in ? _GEN_25679 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1103 = 12'h44f == _T_2[11:0] ? image_1103 : _GEN_1102; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4176 = 12'h450 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7248 = 12'h450 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4176; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10320 = 12'h450 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7248; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13392 = 12'h450 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10320; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16464 = 12'h450 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13392; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19536 = 12'h450 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16464; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22608 = 12'h450 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19536; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25680 = 12'h450 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22608; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1104 = io_valid_in ? _GEN_25680 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1104 = 12'h450 == _T_2[11:0] ? image_1104 : _GEN_1103; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4177 = 12'h451 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7249 = 12'h451 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4177; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10321 = 12'h451 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7249; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13393 = 12'h451 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10321; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16465 = 12'h451 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13393; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19537 = 12'h451 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16465; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22609 = 12'h451 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19537; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25681 = 12'h451 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22609; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1105 = io_valid_in ? _GEN_25681 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1105 = 12'h451 == _T_2[11:0] ? image_1105 : _GEN_1104; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4178 = 12'h452 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7250 = 12'h452 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4178; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10322 = 12'h452 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7250; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13394 = 12'h452 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10322; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16466 = 12'h452 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13394; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19538 = 12'h452 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16466; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22610 = 12'h452 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19538; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25682 = 12'h452 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22610; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1106 = io_valid_in ? _GEN_25682 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1106 = 12'h452 == _T_2[11:0] ? image_1106 : _GEN_1105; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4179 = 12'h453 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7251 = 12'h453 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4179; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10323 = 12'h453 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7251; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13395 = 12'h453 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10323; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16467 = 12'h453 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13395; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19539 = 12'h453 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16467; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22611 = 12'h453 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19539; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25683 = 12'h453 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22611; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1107 = io_valid_in ? _GEN_25683 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1107 = 12'h453 == _T_2[11:0] ? image_1107 : _GEN_1106; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4180 = 12'h454 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7252 = 12'h454 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4180; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10324 = 12'h454 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7252; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13396 = 12'h454 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10324; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16468 = 12'h454 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13396; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19540 = 12'h454 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16468; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22612 = 12'h454 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19540; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25684 = 12'h454 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22612; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1108 = io_valid_in ? _GEN_25684 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1108 = 12'h454 == _T_2[11:0] ? image_1108 : _GEN_1107; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4181 = 12'h455 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7253 = 12'h455 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4181; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10325 = 12'h455 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7253; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13397 = 12'h455 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10325; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16469 = 12'h455 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13397; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19541 = 12'h455 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16469; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22613 = 12'h455 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19541; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25685 = 12'h455 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22613; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1109 = io_valid_in ? _GEN_25685 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1109 = 12'h455 == _T_2[11:0] ? image_1109 : _GEN_1108; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4182 = 12'h456 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7254 = 12'h456 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4182; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10326 = 12'h456 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7254; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13398 = 12'h456 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10326; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16470 = 12'h456 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13398; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19542 = 12'h456 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16470; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22614 = 12'h456 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19542; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25686 = 12'h456 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22614; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1110 = io_valid_in ? _GEN_25686 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1110 = 12'h456 == _T_2[11:0] ? image_1110 : _GEN_1109; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4183 = 12'h457 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7255 = 12'h457 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4183; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10327 = 12'h457 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7255; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13399 = 12'h457 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10327; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16471 = 12'h457 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13399; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19543 = 12'h457 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16471; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22615 = 12'h457 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19543; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25687 = 12'h457 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22615; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1111 = io_valid_in ? _GEN_25687 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1111 = 12'h457 == _T_2[11:0] ? image_1111 : _GEN_1110; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4184 = 12'h458 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7256 = 12'h458 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4184; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10328 = 12'h458 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7256; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13400 = 12'h458 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10328; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16472 = 12'h458 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13400; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19544 = 12'h458 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16472; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22616 = 12'h458 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19544; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25688 = 12'h458 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22616; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1112 = io_valid_in ? _GEN_25688 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1112 = 12'h458 == _T_2[11:0] ? image_1112 : _GEN_1111; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4185 = 12'h459 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7257 = 12'h459 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4185; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10329 = 12'h459 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7257; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13401 = 12'h459 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10329; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16473 = 12'h459 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13401; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19545 = 12'h459 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16473; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22617 = 12'h459 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19545; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25689 = 12'h459 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22617; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1113 = io_valid_in ? _GEN_25689 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1113 = 12'h459 == _T_2[11:0] ? image_1113 : _GEN_1112; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4186 = 12'h45a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7258 = 12'h45a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4186; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10330 = 12'h45a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7258; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13402 = 12'h45a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10330; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16474 = 12'h45a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13402; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19546 = 12'h45a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16474; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22618 = 12'h45a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19546; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25690 = 12'h45a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22618; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1114 = io_valid_in ? _GEN_25690 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1114 = 12'h45a == _T_2[11:0] ? image_1114 : _GEN_1113; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4187 = 12'h45b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7259 = 12'h45b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4187; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10331 = 12'h45b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7259; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13403 = 12'h45b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10331; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16475 = 12'h45b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13403; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19547 = 12'h45b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16475; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22619 = 12'h45b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19547; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25691 = 12'h45b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22619; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1115 = io_valid_in ? _GEN_25691 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1115 = 12'h45b == _T_2[11:0] ? image_1115 : _GEN_1114; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4188 = 12'h45c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7260 = 12'h45c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4188; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10332 = 12'h45c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7260; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13404 = 12'h45c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10332; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16476 = 12'h45c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13404; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19548 = 12'h45c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16476; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22620 = 12'h45c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19548; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25692 = 12'h45c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22620; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1116 = io_valid_in ? _GEN_25692 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1116 = 12'h45c == _T_2[11:0] ? image_1116 : _GEN_1115; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4189 = 12'h45d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7261 = 12'h45d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4189; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10333 = 12'h45d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7261; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13405 = 12'h45d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10333; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16477 = 12'h45d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13405; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19549 = 12'h45d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16477; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22621 = 12'h45d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19549; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25693 = 12'h45d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22621; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1117 = io_valid_in ? _GEN_25693 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1117 = 12'h45d == _T_2[11:0] ? image_1117 : _GEN_1116; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4190 = 12'h45e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7262 = 12'h45e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4190; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10334 = 12'h45e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7262; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13406 = 12'h45e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10334; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16478 = 12'h45e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13406; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19550 = 12'h45e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16478; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22622 = 12'h45e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19550; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25694 = 12'h45e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22622; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1118 = io_valid_in ? _GEN_25694 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1118 = 12'h45e == _T_2[11:0] ? image_1118 : _GEN_1117; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4191 = 12'h45f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7263 = 12'h45f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4191; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10335 = 12'h45f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7263; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13407 = 12'h45f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10335; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16479 = 12'h45f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13407; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19551 = 12'h45f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16479; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22623 = 12'h45f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19551; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25695 = 12'h45f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22623; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1119 = io_valid_in ? _GEN_25695 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1119 = 12'h45f == _T_2[11:0] ? image_1119 : _GEN_1118; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4192 = 12'h460 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7264 = 12'h460 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4192; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10336 = 12'h460 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7264; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13408 = 12'h460 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10336; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16480 = 12'h460 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13408; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19552 = 12'h460 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16480; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22624 = 12'h460 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19552; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25696 = 12'h460 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22624; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1120 = io_valid_in ? _GEN_25696 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1120 = 12'h460 == _T_2[11:0] ? image_1120 : _GEN_1119; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4193 = 12'h461 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7265 = 12'h461 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4193; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10337 = 12'h461 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7265; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13409 = 12'h461 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10337; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16481 = 12'h461 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13409; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19553 = 12'h461 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16481; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22625 = 12'h461 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19553; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25697 = 12'h461 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22625; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1121 = io_valid_in ? _GEN_25697 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1121 = 12'h461 == _T_2[11:0] ? image_1121 : _GEN_1120; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4194 = 12'h462 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7266 = 12'h462 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4194; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10338 = 12'h462 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7266; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13410 = 12'h462 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10338; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16482 = 12'h462 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13410; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19554 = 12'h462 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16482; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22626 = 12'h462 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19554; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25698 = 12'h462 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22626; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1122 = io_valid_in ? _GEN_25698 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1122 = 12'h462 == _T_2[11:0] ? image_1122 : _GEN_1121; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4195 = 12'h463 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7267 = 12'h463 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4195; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10339 = 12'h463 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7267; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13411 = 12'h463 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10339; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16483 = 12'h463 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13411; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19555 = 12'h463 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16483; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22627 = 12'h463 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19555; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25699 = 12'h463 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22627; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1123 = io_valid_in ? _GEN_25699 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1123 = 12'h463 == _T_2[11:0] ? image_1123 : _GEN_1122; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4196 = 12'h464 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7268 = 12'h464 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4196; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10340 = 12'h464 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7268; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13412 = 12'h464 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10340; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16484 = 12'h464 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13412; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19556 = 12'h464 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16484; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22628 = 12'h464 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19556; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25700 = 12'h464 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22628; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1124 = io_valid_in ? _GEN_25700 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1124 = 12'h464 == _T_2[11:0] ? image_1124 : _GEN_1123; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4197 = 12'h465 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7269 = 12'h465 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4197; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10341 = 12'h465 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7269; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13413 = 12'h465 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10341; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16485 = 12'h465 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13413; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19557 = 12'h465 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16485; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22629 = 12'h465 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19557; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25701 = 12'h465 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22629; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1125 = io_valid_in ? _GEN_25701 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1125 = 12'h465 == _T_2[11:0] ? image_1125 : _GEN_1124; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4198 = 12'h466 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7270 = 12'h466 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4198; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10342 = 12'h466 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7270; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13414 = 12'h466 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10342; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16486 = 12'h466 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13414; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19558 = 12'h466 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16486; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22630 = 12'h466 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19558; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25702 = 12'h466 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22630; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1126 = io_valid_in ? _GEN_25702 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1126 = 12'h466 == _T_2[11:0] ? image_1126 : _GEN_1125; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4199 = 12'h467 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7271 = 12'h467 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4199; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10343 = 12'h467 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7271; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13415 = 12'h467 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10343; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16487 = 12'h467 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13415; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19559 = 12'h467 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16487; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22631 = 12'h467 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19559; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25703 = 12'h467 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22631; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1127 = io_valid_in ? _GEN_25703 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1127 = 12'h467 == _T_2[11:0] ? image_1127 : _GEN_1126; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4200 = 12'h468 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7272 = 12'h468 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4200; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10344 = 12'h468 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7272; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13416 = 12'h468 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10344; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16488 = 12'h468 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13416; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19560 = 12'h468 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16488; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22632 = 12'h468 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19560; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25704 = 12'h468 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22632; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1128 = io_valid_in ? _GEN_25704 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1128 = 12'h468 == _T_2[11:0] ? image_1128 : _GEN_1127; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4201 = 12'h469 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7273 = 12'h469 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4201; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10345 = 12'h469 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7273; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13417 = 12'h469 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10345; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16489 = 12'h469 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13417; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19561 = 12'h469 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16489; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22633 = 12'h469 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19561; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25705 = 12'h469 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22633; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1129 = io_valid_in ? _GEN_25705 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1129 = 12'h469 == _T_2[11:0] ? image_1129 : _GEN_1128; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4202 = 12'h46a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7274 = 12'h46a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4202; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10346 = 12'h46a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7274; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13418 = 12'h46a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10346; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16490 = 12'h46a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13418; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19562 = 12'h46a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16490; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22634 = 12'h46a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19562; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25706 = 12'h46a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22634; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1130 = io_valid_in ? _GEN_25706 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1130 = 12'h46a == _T_2[11:0] ? image_1130 : _GEN_1129; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4203 = 12'h46b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7275 = 12'h46b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4203; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10347 = 12'h46b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7275; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13419 = 12'h46b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10347; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16491 = 12'h46b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13419; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19563 = 12'h46b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16491; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22635 = 12'h46b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19563; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25707 = 12'h46b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22635; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1131 = io_valid_in ? _GEN_25707 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1131 = 12'h46b == _T_2[11:0] ? image_1131 : _GEN_1130; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4204 = 12'h46c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7276 = 12'h46c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4204; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10348 = 12'h46c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7276; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13420 = 12'h46c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10348; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16492 = 12'h46c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13420; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19564 = 12'h46c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16492; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22636 = 12'h46c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19564; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25708 = 12'h46c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22636; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1132 = io_valid_in ? _GEN_25708 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1132 = 12'h46c == _T_2[11:0] ? image_1132 : _GEN_1131; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4205 = 12'h46d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7277 = 12'h46d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4205; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10349 = 12'h46d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7277; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13421 = 12'h46d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10349; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16493 = 12'h46d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13421; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19565 = 12'h46d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16493; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22637 = 12'h46d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19565; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25709 = 12'h46d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22637; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1133 = io_valid_in ? _GEN_25709 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1133 = 12'h46d == _T_2[11:0] ? image_1133 : _GEN_1132; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4206 = 12'h46e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7278 = 12'h46e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4206; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10350 = 12'h46e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7278; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13422 = 12'h46e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10350; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16494 = 12'h46e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13422; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19566 = 12'h46e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16494; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22638 = 12'h46e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19566; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25710 = 12'h46e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22638; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1134 = io_valid_in ? _GEN_25710 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1134 = 12'h46e == _T_2[11:0] ? image_1134 : _GEN_1133; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4207 = 12'h46f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7279 = 12'h46f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4207; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10351 = 12'h46f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7279; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13423 = 12'h46f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10351; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16495 = 12'h46f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13423; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19567 = 12'h46f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16495; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22639 = 12'h46f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19567; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25711 = 12'h46f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22639; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1135 = io_valid_in ? _GEN_25711 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1135 = 12'h46f == _T_2[11:0] ? image_1135 : _GEN_1134; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4208 = 12'h470 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7280 = 12'h470 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4208; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10352 = 12'h470 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7280; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13424 = 12'h470 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10352; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16496 = 12'h470 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13424; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19568 = 12'h470 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16496; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22640 = 12'h470 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19568; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25712 = 12'h470 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22640; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1136 = io_valid_in ? _GEN_25712 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1136 = 12'h470 == _T_2[11:0] ? image_1136 : _GEN_1135; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4209 = 12'h471 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7281 = 12'h471 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4209; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10353 = 12'h471 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7281; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13425 = 12'h471 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10353; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16497 = 12'h471 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13425; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19569 = 12'h471 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16497; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22641 = 12'h471 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19569; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25713 = 12'h471 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22641; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1137 = io_valid_in ? _GEN_25713 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1137 = 12'h471 == _T_2[11:0] ? image_1137 : _GEN_1136; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4210 = 12'h472 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7282 = 12'h472 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4210; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10354 = 12'h472 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7282; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13426 = 12'h472 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10354; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16498 = 12'h472 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13426; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19570 = 12'h472 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16498; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22642 = 12'h472 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19570; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25714 = 12'h472 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22642; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1138 = io_valid_in ? _GEN_25714 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1138 = 12'h472 == _T_2[11:0] ? image_1138 : _GEN_1137; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4211 = 12'h473 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7283 = 12'h473 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4211; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10355 = 12'h473 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7283; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13427 = 12'h473 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10355; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16499 = 12'h473 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13427; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19571 = 12'h473 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16499; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22643 = 12'h473 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19571; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25715 = 12'h473 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22643; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1139 = io_valid_in ? _GEN_25715 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1139 = 12'h473 == _T_2[11:0] ? image_1139 : _GEN_1138; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4212 = 12'h474 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7284 = 12'h474 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4212; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10356 = 12'h474 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7284; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13428 = 12'h474 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10356; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16500 = 12'h474 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13428; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19572 = 12'h474 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16500; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22644 = 12'h474 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19572; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25716 = 12'h474 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22644; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1140 = io_valid_in ? _GEN_25716 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1140 = 12'h474 == _T_2[11:0] ? image_1140 : _GEN_1139; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4213 = 12'h475 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7285 = 12'h475 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4213; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10357 = 12'h475 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7285; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13429 = 12'h475 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10357; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16501 = 12'h475 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13429; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19573 = 12'h475 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16501; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22645 = 12'h475 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19573; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25717 = 12'h475 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22645; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1141 = io_valid_in ? _GEN_25717 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1141 = 12'h475 == _T_2[11:0] ? image_1141 : _GEN_1140; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4214 = 12'h476 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7286 = 12'h476 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4214; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10358 = 12'h476 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7286; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13430 = 12'h476 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10358; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16502 = 12'h476 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13430; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19574 = 12'h476 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16502; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22646 = 12'h476 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19574; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25718 = 12'h476 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22646; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1142 = io_valid_in ? _GEN_25718 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1142 = 12'h476 == _T_2[11:0] ? image_1142 : _GEN_1141; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4215 = 12'h477 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7287 = 12'h477 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4215; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10359 = 12'h477 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7287; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13431 = 12'h477 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10359; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16503 = 12'h477 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13431; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19575 = 12'h477 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16503; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22647 = 12'h477 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19575; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25719 = 12'h477 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22647; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1143 = io_valid_in ? _GEN_25719 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1143 = 12'h477 == _T_2[11:0] ? image_1143 : _GEN_1142; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4216 = 12'h478 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7288 = 12'h478 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4216; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10360 = 12'h478 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7288; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13432 = 12'h478 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10360; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16504 = 12'h478 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13432; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19576 = 12'h478 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16504; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22648 = 12'h478 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19576; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25720 = 12'h478 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22648; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1144 = io_valid_in ? _GEN_25720 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1144 = 12'h478 == _T_2[11:0] ? image_1144 : _GEN_1143; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4217 = 12'h479 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7289 = 12'h479 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4217; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10361 = 12'h479 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7289; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13433 = 12'h479 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10361; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16505 = 12'h479 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13433; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19577 = 12'h479 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16505; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22649 = 12'h479 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19577; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25721 = 12'h479 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22649; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1145 = io_valid_in ? _GEN_25721 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1145 = 12'h479 == _T_2[11:0] ? image_1145 : _GEN_1144; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4218 = 12'h47a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7290 = 12'h47a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4218; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10362 = 12'h47a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7290; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13434 = 12'h47a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10362; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16506 = 12'h47a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13434; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19578 = 12'h47a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16506; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22650 = 12'h47a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19578; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25722 = 12'h47a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22650; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1146 = io_valid_in ? _GEN_25722 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1146 = 12'h47a == _T_2[11:0] ? image_1146 : _GEN_1145; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4219 = 12'h47b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7291 = 12'h47b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4219; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10363 = 12'h47b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7291; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13435 = 12'h47b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10363; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16507 = 12'h47b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13435; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19579 = 12'h47b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16507; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22651 = 12'h47b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19579; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25723 = 12'h47b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22651; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1147 = io_valid_in ? _GEN_25723 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1147 = 12'h47b == _T_2[11:0] ? image_1147 : _GEN_1146; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4220 = 12'h47c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7292 = 12'h47c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4220; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10364 = 12'h47c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7292; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13436 = 12'h47c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10364; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16508 = 12'h47c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13436; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19580 = 12'h47c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16508; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22652 = 12'h47c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19580; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25724 = 12'h47c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22652; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1148 = io_valid_in ? _GEN_25724 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1148 = 12'h47c == _T_2[11:0] ? image_1148 : _GEN_1147; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4221 = 12'h47d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7293 = 12'h47d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4221; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10365 = 12'h47d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7293; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13437 = 12'h47d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10365; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16509 = 12'h47d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13437; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19581 = 12'h47d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16509; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22653 = 12'h47d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19581; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25725 = 12'h47d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22653; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1149 = io_valid_in ? _GEN_25725 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1149 = 12'h47d == _T_2[11:0] ? image_1149 : _GEN_1148; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4222 = 12'h47e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7294 = 12'h47e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4222; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10366 = 12'h47e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7294; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13438 = 12'h47e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10366; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16510 = 12'h47e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13438; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19582 = 12'h47e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16510; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22654 = 12'h47e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19582; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25726 = 12'h47e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22654; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1150 = io_valid_in ? _GEN_25726 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1150 = 12'h47e == _T_2[11:0] ? image_1150 : _GEN_1149; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4223 = 12'h47f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7295 = 12'h47f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4223; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10367 = 12'h47f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7295; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13439 = 12'h47f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10367; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16511 = 12'h47f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13439; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19583 = 12'h47f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16511; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22655 = 12'h47f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19583; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25727 = 12'h47f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22655; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1151 = io_valid_in ? _GEN_25727 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1151 = 12'h47f == _T_2[11:0] ? image_1151 : _GEN_1150; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4224 = 12'h480 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7296 = 12'h480 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4224; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10368 = 12'h480 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7296; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13440 = 12'h480 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10368; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16512 = 12'h480 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13440; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19584 = 12'h480 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16512; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22656 = 12'h480 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19584; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25728 = 12'h480 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22656; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1152 = io_valid_in ? _GEN_25728 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1152 = 12'h480 == _T_2[11:0] ? image_1152 : _GEN_1151; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4225 = 12'h481 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7297 = 12'h481 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4225; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10369 = 12'h481 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7297; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13441 = 12'h481 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10369; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16513 = 12'h481 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13441; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19585 = 12'h481 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16513; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22657 = 12'h481 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19585; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25729 = 12'h481 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22657; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1153 = io_valid_in ? _GEN_25729 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1153 = 12'h481 == _T_2[11:0] ? image_1153 : _GEN_1152; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4226 = 12'h482 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7298 = 12'h482 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4226; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10370 = 12'h482 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7298; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13442 = 12'h482 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10370; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16514 = 12'h482 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13442; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19586 = 12'h482 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16514; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22658 = 12'h482 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19586; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25730 = 12'h482 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22658; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1154 = io_valid_in ? _GEN_25730 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1154 = 12'h482 == _T_2[11:0] ? image_1154 : _GEN_1153; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4227 = 12'h483 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7299 = 12'h483 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4227; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10371 = 12'h483 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7299; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13443 = 12'h483 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10371; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16515 = 12'h483 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13443; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19587 = 12'h483 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16515; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22659 = 12'h483 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19587; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25731 = 12'h483 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22659; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1155 = io_valid_in ? _GEN_25731 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1155 = 12'h483 == _T_2[11:0] ? image_1155 : _GEN_1154; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4228 = 12'h484 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7300 = 12'h484 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4228; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10372 = 12'h484 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7300; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13444 = 12'h484 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10372; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16516 = 12'h484 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13444; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19588 = 12'h484 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16516; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22660 = 12'h484 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19588; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25732 = 12'h484 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22660; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1156 = io_valid_in ? _GEN_25732 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1156 = 12'h484 == _T_2[11:0] ? image_1156 : _GEN_1155; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4229 = 12'h485 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7301 = 12'h485 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4229; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10373 = 12'h485 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7301; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13445 = 12'h485 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10373; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16517 = 12'h485 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13445; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19589 = 12'h485 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16517; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22661 = 12'h485 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19589; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25733 = 12'h485 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22661; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1157 = io_valid_in ? _GEN_25733 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1157 = 12'h485 == _T_2[11:0] ? image_1157 : _GEN_1156; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4230 = 12'h486 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7302 = 12'h486 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4230; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10374 = 12'h486 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7302; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13446 = 12'h486 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10374; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16518 = 12'h486 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13446; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19590 = 12'h486 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16518; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22662 = 12'h486 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19590; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25734 = 12'h486 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22662; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1158 = io_valid_in ? _GEN_25734 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1158 = 12'h486 == _T_2[11:0] ? image_1158 : _GEN_1157; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4231 = 12'h487 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7303 = 12'h487 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4231; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10375 = 12'h487 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7303; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13447 = 12'h487 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10375; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16519 = 12'h487 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13447; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19591 = 12'h487 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16519; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22663 = 12'h487 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19591; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25735 = 12'h487 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22663; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1159 = io_valid_in ? _GEN_25735 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1159 = 12'h487 == _T_2[11:0] ? image_1159 : _GEN_1158; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4232 = 12'h488 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7304 = 12'h488 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4232; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10376 = 12'h488 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7304; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13448 = 12'h488 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10376; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16520 = 12'h488 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13448; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19592 = 12'h488 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16520; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22664 = 12'h488 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19592; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25736 = 12'h488 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22664; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1160 = io_valid_in ? _GEN_25736 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1160 = 12'h488 == _T_2[11:0] ? image_1160 : _GEN_1159; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4233 = 12'h489 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7305 = 12'h489 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4233; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10377 = 12'h489 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7305; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13449 = 12'h489 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10377; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16521 = 12'h489 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13449; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19593 = 12'h489 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16521; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22665 = 12'h489 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19593; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25737 = 12'h489 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22665; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1161 = io_valid_in ? _GEN_25737 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1161 = 12'h489 == _T_2[11:0] ? image_1161 : _GEN_1160; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4234 = 12'h48a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7306 = 12'h48a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4234; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10378 = 12'h48a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7306; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13450 = 12'h48a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10378; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16522 = 12'h48a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13450; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19594 = 12'h48a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16522; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22666 = 12'h48a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19594; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25738 = 12'h48a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22666; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1162 = io_valid_in ? _GEN_25738 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1162 = 12'h48a == _T_2[11:0] ? image_1162 : _GEN_1161; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4235 = 12'h48b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7307 = 12'h48b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4235; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10379 = 12'h48b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7307; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13451 = 12'h48b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10379; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16523 = 12'h48b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13451; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19595 = 12'h48b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16523; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22667 = 12'h48b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19595; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25739 = 12'h48b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22667; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1163 = io_valid_in ? _GEN_25739 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1163 = 12'h48b == _T_2[11:0] ? image_1163 : _GEN_1162; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4236 = 12'h48c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7308 = 12'h48c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4236; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10380 = 12'h48c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7308; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13452 = 12'h48c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10380; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16524 = 12'h48c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13452; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19596 = 12'h48c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16524; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22668 = 12'h48c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19596; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25740 = 12'h48c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22668; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1164 = io_valid_in ? _GEN_25740 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1164 = 12'h48c == _T_2[11:0] ? image_1164 : _GEN_1163; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4237 = 12'h48d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7309 = 12'h48d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4237; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10381 = 12'h48d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7309; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13453 = 12'h48d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10381; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16525 = 12'h48d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13453; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19597 = 12'h48d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16525; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22669 = 12'h48d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19597; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25741 = 12'h48d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22669; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1165 = io_valid_in ? _GEN_25741 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1165 = 12'h48d == _T_2[11:0] ? image_1165 : _GEN_1164; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4238 = 12'h48e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7310 = 12'h48e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4238; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10382 = 12'h48e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7310; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13454 = 12'h48e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10382; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16526 = 12'h48e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13454; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19598 = 12'h48e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16526; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22670 = 12'h48e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19598; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25742 = 12'h48e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22670; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1166 = io_valid_in ? _GEN_25742 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1166 = 12'h48e == _T_2[11:0] ? image_1166 : _GEN_1165; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4239 = 12'h48f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7311 = 12'h48f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4239; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10383 = 12'h48f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7311; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13455 = 12'h48f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10383; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16527 = 12'h48f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13455; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19599 = 12'h48f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16527; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22671 = 12'h48f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19599; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25743 = 12'h48f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22671; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1167 = io_valid_in ? _GEN_25743 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1167 = 12'h48f == _T_2[11:0] ? image_1167 : _GEN_1166; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4240 = 12'h490 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7312 = 12'h490 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4240; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10384 = 12'h490 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7312; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13456 = 12'h490 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10384; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16528 = 12'h490 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13456; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19600 = 12'h490 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16528; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22672 = 12'h490 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19600; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25744 = 12'h490 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22672; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1168 = io_valid_in ? _GEN_25744 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1168 = 12'h490 == _T_2[11:0] ? image_1168 : _GEN_1167; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4241 = 12'h491 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7313 = 12'h491 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4241; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10385 = 12'h491 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7313; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13457 = 12'h491 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10385; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16529 = 12'h491 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13457; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19601 = 12'h491 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16529; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22673 = 12'h491 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19601; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25745 = 12'h491 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22673; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1169 = io_valid_in ? _GEN_25745 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1169 = 12'h491 == _T_2[11:0] ? image_1169 : _GEN_1168; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4242 = 12'h492 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7314 = 12'h492 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4242; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10386 = 12'h492 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7314; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13458 = 12'h492 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10386; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16530 = 12'h492 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13458; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19602 = 12'h492 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16530; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22674 = 12'h492 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19602; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25746 = 12'h492 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22674; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1170 = io_valid_in ? _GEN_25746 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1170 = 12'h492 == _T_2[11:0] ? image_1170 : _GEN_1169; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4243 = 12'h493 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7315 = 12'h493 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4243; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10387 = 12'h493 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7315; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13459 = 12'h493 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10387; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16531 = 12'h493 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13459; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19603 = 12'h493 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16531; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22675 = 12'h493 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19603; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25747 = 12'h493 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22675; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1171 = io_valid_in ? _GEN_25747 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1171 = 12'h493 == _T_2[11:0] ? image_1171 : _GEN_1170; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4244 = 12'h494 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7316 = 12'h494 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4244; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10388 = 12'h494 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7316; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13460 = 12'h494 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10388; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16532 = 12'h494 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13460; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19604 = 12'h494 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16532; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22676 = 12'h494 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19604; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25748 = 12'h494 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22676; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1172 = io_valid_in ? _GEN_25748 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1172 = 12'h494 == _T_2[11:0] ? image_1172 : _GEN_1171; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4245 = 12'h495 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7317 = 12'h495 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4245; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10389 = 12'h495 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7317; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13461 = 12'h495 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10389; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16533 = 12'h495 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13461; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19605 = 12'h495 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16533; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22677 = 12'h495 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19605; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25749 = 12'h495 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22677; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1173 = io_valid_in ? _GEN_25749 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1173 = 12'h495 == _T_2[11:0] ? image_1173 : _GEN_1172; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4246 = 12'h496 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7318 = 12'h496 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4246; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10390 = 12'h496 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7318; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13462 = 12'h496 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10390; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16534 = 12'h496 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13462; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19606 = 12'h496 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16534; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22678 = 12'h496 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19606; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25750 = 12'h496 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22678; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1174 = io_valid_in ? _GEN_25750 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1174 = 12'h496 == _T_2[11:0] ? image_1174 : _GEN_1173; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4247 = 12'h497 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7319 = 12'h497 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4247; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10391 = 12'h497 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7319; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13463 = 12'h497 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10391; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16535 = 12'h497 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13463; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19607 = 12'h497 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16535; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22679 = 12'h497 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19607; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25751 = 12'h497 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22679; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1175 = io_valid_in ? _GEN_25751 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1175 = 12'h497 == _T_2[11:0] ? image_1175 : _GEN_1174; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4248 = 12'h498 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7320 = 12'h498 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4248; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10392 = 12'h498 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7320; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13464 = 12'h498 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10392; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16536 = 12'h498 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13464; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19608 = 12'h498 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16536; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22680 = 12'h498 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19608; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25752 = 12'h498 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22680; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1176 = io_valid_in ? _GEN_25752 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1176 = 12'h498 == _T_2[11:0] ? image_1176 : _GEN_1175; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4249 = 12'h499 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7321 = 12'h499 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4249; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10393 = 12'h499 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7321; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13465 = 12'h499 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10393; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16537 = 12'h499 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13465; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19609 = 12'h499 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16537; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22681 = 12'h499 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19609; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25753 = 12'h499 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22681; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1177 = io_valid_in ? _GEN_25753 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1177 = 12'h499 == _T_2[11:0] ? image_1177 : _GEN_1176; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4250 = 12'h49a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7322 = 12'h49a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4250; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10394 = 12'h49a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7322; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13466 = 12'h49a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10394; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16538 = 12'h49a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13466; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19610 = 12'h49a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16538; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22682 = 12'h49a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19610; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25754 = 12'h49a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22682; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1178 = io_valid_in ? _GEN_25754 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1178 = 12'h49a == _T_2[11:0] ? image_1178 : _GEN_1177; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4251 = 12'h49b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7323 = 12'h49b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4251; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10395 = 12'h49b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7323; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13467 = 12'h49b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10395; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16539 = 12'h49b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13467; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19611 = 12'h49b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16539; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22683 = 12'h49b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19611; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25755 = 12'h49b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22683; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1179 = io_valid_in ? _GEN_25755 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1179 = 12'h49b == _T_2[11:0] ? image_1179 : _GEN_1178; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4252 = 12'h49c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7324 = 12'h49c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4252; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10396 = 12'h49c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7324; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13468 = 12'h49c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10396; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16540 = 12'h49c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13468; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19612 = 12'h49c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16540; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22684 = 12'h49c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19612; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25756 = 12'h49c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22684; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1180 = io_valid_in ? _GEN_25756 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1180 = 12'h49c == _T_2[11:0] ? image_1180 : _GEN_1179; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4253 = 12'h49d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7325 = 12'h49d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4253; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10397 = 12'h49d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7325; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13469 = 12'h49d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10397; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16541 = 12'h49d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13469; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19613 = 12'h49d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16541; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22685 = 12'h49d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19613; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25757 = 12'h49d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22685; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1181 = io_valid_in ? _GEN_25757 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1181 = 12'h49d == _T_2[11:0] ? image_1181 : _GEN_1180; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4254 = 12'h49e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7326 = 12'h49e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4254; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10398 = 12'h49e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7326; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13470 = 12'h49e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10398; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16542 = 12'h49e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13470; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19614 = 12'h49e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16542; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22686 = 12'h49e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19614; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25758 = 12'h49e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22686; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1182 = io_valid_in ? _GEN_25758 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1182 = 12'h49e == _T_2[11:0] ? image_1182 : _GEN_1181; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4255 = 12'h49f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7327 = 12'h49f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4255; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10399 = 12'h49f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7327; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13471 = 12'h49f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10399; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16543 = 12'h49f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13471; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19615 = 12'h49f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16543; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22687 = 12'h49f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19615; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25759 = 12'h49f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22687; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1183 = io_valid_in ? _GEN_25759 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1183 = 12'h49f == _T_2[11:0] ? image_1183 : _GEN_1182; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4256 = 12'h4a0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7328 = 12'h4a0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4256; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10400 = 12'h4a0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7328; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13472 = 12'h4a0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10400; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16544 = 12'h4a0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13472; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19616 = 12'h4a0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16544; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22688 = 12'h4a0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19616; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25760 = 12'h4a0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22688; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1184 = io_valid_in ? _GEN_25760 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1184 = 12'h4a0 == _T_2[11:0] ? image_1184 : _GEN_1183; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4257 = 12'h4a1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7329 = 12'h4a1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4257; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10401 = 12'h4a1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7329; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13473 = 12'h4a1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10401; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16545 = 12'h4a1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13473; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19617 = 12'h4a1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16545; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22689 = 12'h4a1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19617; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25761 = 12'h4a1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22689; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1185 = io_valid_in ? _GEN_25761 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1185 = 12'h4a1 == _T_2[11:0] ? image_1185 : _GEN_1184; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4258 = 12'h4a2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7330 = 12'h4a2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4258; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10402 = 12'h4a2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7330; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13474 = 12'h4a2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10402; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16546 = 12'h4a2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13474; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19618 = 12'h4a2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16546; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22690 = 12'h4a2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19618; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25762 = 12'h4a2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22690; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1186 = io_valid_in ? _GEN_25762 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1186 = 12'h4a2 == _T_2[11:0] ? image_1186 : _GEN_1185; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4259 = 12'h4a3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7331 = 12'h4a3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4259; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10403 = 12'h4a3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7331; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13475 = 12'h4a3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10403; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16547 = 12'h4a3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13475; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19619 = 12'h4a3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16547; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22691 = 12'h4a3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19619; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25763 = 12'h4a3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22691; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1187 = io_valid_in ? _GEN_25763 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1187 = 12'h4a3 == _T_2[11:0] ? image_1187 : _GEN_1186; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4260 = 12'h4a4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7332 = 12'h4a4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4260; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10404 = 12'h4a4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7332; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13476 = 12'h4a4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10404; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16548 = 12'h4a4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13476; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19620 = 12'h4a4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16548; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22692 = 12'h4a4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19620; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25764 = 12'h4a4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22692; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1188 = io_valid_in ? _GEN_25764 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1188 = 12'h4a4 == _T_2[11:0] ? image_1188 : _GEN_1187; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4261 = 12'h4a5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7333 = 12'h4a5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4261; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10405 = 12'h4a5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7333; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13477 = 12'h4a5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10405; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16549 = 12'h4a5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13477; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19621 = 12'h4a5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16549; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22693 = 12'h4a5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19621; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25765 = 12'h4a5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22693; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1189 = io_valid_in ? _GEN_25765 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1189 = 12'h4a5 == _T_2[11:0] ? image_1189 : _GEN_1188; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4262 = 12'h4a6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7334 = 12'h4a6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4262; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10406 = 12'h4a6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7334; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13478 = 12'h4a6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10406; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16550 = 12'h4a6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13478; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19622 = 12'h4a6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16550; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22694 = 12'h4a6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19622; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25766 = 12'h4a6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22694; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1190 = io_valid_in ? _GEN_25766 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1190 = 12'h4a6 == _T_2[11:0] ? image_1190 : _GEN_1189; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4263 = 12'h4a7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7335 = 12'h4a7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4263; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10407 = 12'h4a7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7335; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13479 = 12'h4a7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10407; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16551 = 12'h4a7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13479; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19623 = 12'h4a7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16551; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22695 = 12'h4a7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19623; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25767 = 12'h4a7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22695; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1191 = io_valid_in ? _GEN_25767 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1191 = 12'h4a7 == _T_2[11:0] ? image_1191 : _GEN_1190; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4264 = 12'h4a8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7336 = 12'h4a8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4264; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10408 = 12'h4a8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7336; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13480 = 12'h4a8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10408; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16552 = 12'h4a8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13480; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19624 = 12'h4a8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16552; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22696 = 12'h4a8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19624; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25768 = 12'h4a8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22696; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1192 = io_valid_in ? _GEN_25768 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1192 = 12'h4a8 == _T_2[11:0] ? image_1192 : _GEN_1191; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4265 = 12'h4a9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7337 = 12'h4a9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4265; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10409 = 12'h4a9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7337; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13481 = 12'h4a9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10409; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16553 = 12'h4a9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13481; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19625 = 12'h4a9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16553; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22697 = 12'h4a9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19625; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25769 = 12'h4a9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22697; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1193 = io_valid_in ? _GEN_25769 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1193 = 12'h4a9 == _T_2[11:0] ? image_1193 : _GEN_1192; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4266 = 12'h4aa == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7338 = 12'h4aa == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4266; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10410 = 12'h4aa == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7338; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13482 = 12'h4aa == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10410; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16554 = 12'h4aa == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13482; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19626 = 12'h4aa == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16554; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22698 = 12'h4aa == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19626; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25770 = 12'h4aa == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22698; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1194 = io_valid_in ? _GEN_25770 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1194 = 12'h4aa == _T_2[11:0] ? image_1194 : _GEN_1193; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4267 = 12'h4ab == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7339 = 12'h4ab == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4267; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10411 = 12'h4ab == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7339; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13483 = 12'h4ab == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10411; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16555 = 12'h4ab == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13483; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19627 = 12'h4ab == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16555; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22699 = 12'h4ab == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19627; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25771 = 12'h4ab == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22699; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1195 = io_valid_in ? _GEN_25771 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1195 = 12'h4ab == _T_2[11:0] ? image_1195 : _GEN_1194; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4268 = 12'h4ac == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7340 = 12'h4ac == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4268; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10412 = 12'h4ac == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7340; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13484 = 12'h4ac == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10412; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16556 = 12'h4ac == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13484; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19628 = 12'h4ac == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16556; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22700 = 12'h4ac == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19628; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25772 = 12'h4ac == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22700; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1196 = io_valid_in ? _GEN_25772 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1196 = 12'h4ac == _T_2[11:0] ? image_1196 : _GEN_1195; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4269 = 12'h4ad == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7341 = 12'h4ad == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4269; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10413 = 12'h4ad == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7341; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13485 = 12'h4ad == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10413; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16557 = 12'h4ad == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13485; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19629 = 12'h4ad == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16557; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22701 = 12'h4ad == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19629; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25773 = 12'h4ad == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22701; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1197 = io_valid_in ? _GEN_25773 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1197 = 12'h4ad == _T_2[11:0] ? image_1197 : _GEN_1196; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4270 = 12'h4ae == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7342 = 12'h4ae == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4270; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10414 = 12'h4ae == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7342; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13486 = 12'h4ae == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10414; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16558 = 12'h4ae == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13486; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19630 = 12'h4ae == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16558; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22702 = 12'h4ae == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19630; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25774 = 12'h4ae == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22702; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1198 = io_valid_in ? _GEN_25774 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1198 = 12'h4ae == _T_2[11:0] ? image_1198 : _GEN_1197; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4271 = 12'h4af == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7343 = 12'h4af == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4271; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10415 = 12'h4af == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7343; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13487 = 12'h4af == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10415; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16559 = 12'h4af == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13487; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19631 = 12'h4af == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16559; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22703 = 12'h4af == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19631; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25775 = 12'h4af == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22703; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1199 = io_valid_in ? _GEN_25775 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1199 = 12'h4af == _T_2[11:0] ? image_1199 : _GEN_1198; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4272 = 12'h4b0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7344 = 12'h4b0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4272; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10416 = 12'h4b0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7344; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13488 = 12'h4b0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10416; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16560 = 12'h4b0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13488; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19632 = 12'h4b0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16560; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22704 = 12'h4b0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19632; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25776 = 12'h4b0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22704; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1200 = io_valid_in ? _GEN_25776 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1200 = 12'h4b0 == _T_2[11:0] ? image_1200 : _GEN_1199; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4273 = 12'h4b1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7345 = 12'h4b1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4273; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10417 = 12'h4b1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7345; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13489 = 12'h4b1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10417; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16561 = 12'h4b1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13489; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19633 = 12'h4b1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16561; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22705 = 12'h4b1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19633; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25777 = 12'h4b1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22705; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1201 = io_valid_in ? _GEN_25777 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1201 = 12'h4b1 == _T_2[11:0] ? image_1201 : _GEN_1200; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4274 = 12'h4b2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7346 = 12'h4b2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4274; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10418 = 12'h4b2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7346; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13490 = 12'h4b2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10418; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16562 = 12'h4b2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13490; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19634 = 12'h4b2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16562; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22706 = 12'h4b2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19634; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25778 = 12'h4b2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22706; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1202 = io_valid_in ? _GEN_25778 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1202 = 12'h4b2 == _T_2[11:0] ? image_1202 : _GEN_1201; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4275 = 12'h4b3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7347 = 12'h4b3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4275; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10419 = 12'h4b3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7347; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13491 = 12'h4b3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10419; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16563 = 12'h4b3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13491; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19635 = 12'h4b3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16563; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22707 = 12'h4b3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19635; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25779 = 12'h4b3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22707; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1203 = io_valid_in ? _GEN_25779 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1203 = 12'h4b3 == _T_2[11:0] ? image_1203 : _GEN_1202; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4276 = 12'h4b4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7348 = 12'h4b4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4276; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10420 = 12'h4b4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7348; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13492 = 12'h4b4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10420; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16564 = 12'h4b4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13492; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19636 = 12'h4b4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16564; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22708 = 12'h4b4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19636; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25780 = 12'h4b4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22708; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1204 = io_valid_in ? _GEN_25780 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1204 = 12'h4b4 == _T_2[11:0] ? image_1204 : _GEN_1203; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4277 = 12'h4b5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7349 = 12'h4b5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4277; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10421 = 12'h4b5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7349; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13493 = 12'h4b5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10421; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16565 = 12'h4b5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13493; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19637 = 12'h4b5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16565; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22709 = 12'h4b5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19637; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25781 = 12'h4b5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22709; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1205 = io_valid_in ? _GEN_25781 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1205 = 12'h4b5 == _T_2[11:0] ? image_1205 : _GEN_1204; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4278 = 12'h4b6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7350 = 12'h4b6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4278; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10422 = 12'h4b6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7350; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13494 = 12'h4b6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10422; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16566 = 12'h4b6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13494; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19638 = 12'h4b6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16566; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22710 = 12'h4b6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19638; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25782 = 12'h4b6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22710; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1206 = io_valid_in ? _GEN_25782 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1206 = 12'h4b6 == _T_2[11:0] ? image_1206 : _GEN_1205; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4279 = 12'h4b7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7351 = 12'h4b7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4279; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10423 = 12'h4b7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7351; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13495 = 12'h4b7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10423; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16567 = 12'h4b7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13495; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19639 = 12'h4b7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16567; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22711 = 12'h4b7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19639; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25783 = 12'h4b7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22711; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1207 = io_valid_in ? _GEN_25783 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1207 = 12'h4b7 == _T_2[11:0] ? image_1207 : _GEN_1206; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4280 = 12'h4b8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7352 = 12'h4b8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4280; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10424 = 12'h4b8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7352; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13496 = 12'h4b8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10424; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16568 = 12'h4b8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13496; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19640 = 12'h4b8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16568; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22712 = 12'h4b8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19640; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25784 = 12'h4b8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22712; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1208 = io_valid_in ? _GEN_25784 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1208 = 12'h4b8 == _T_2[11:0] ? image_1208 : _GEN_1207; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4281 = 12'h4b9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7353 = 12'h4b9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4281; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10425 = 12'h4b9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7353; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13497 = 12'h4b9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10425; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16569 = 12'h4b9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13497; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19641 = 12'h4b9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16569; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22713 = 12'h4b9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19641; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25785 = 12'h4b9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22713; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1209 = io_valid_in ? _GEN_25785 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1209 = 12'h4b9 == _T_2[11:0] ? image_1209 : _GEN_1208; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4282 = 12'h4ba == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7354 = 12'h4ba == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4282; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10426 = 12'h4ba == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7354; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13498 = 12'h4ba == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10426; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16570 = 12'h4ba == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13498; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19642 = 12'h4ba == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16570; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22714 = 12'h4ba == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19642; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25786 = 12'h4ba == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22714; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1210 = io_valid_in ? _GEN_25786 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1210 = 12'h4ba == _T_2[11:0] ? image_1210 : _GEN_1209; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4283 = 12'h4bb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7355 = 12'h4bb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4283; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10427 = 12'h4bb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7355; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13499 = 12'h4bb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10427; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16571 = 12'h4bb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13499; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19643 = 12'h4bb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16571; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22715 = 12'h4bb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19643; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25787 = 12'h4bb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22715; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1211 = io_valid_in ? _GEN_25787 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1211 = 12'h4bb == _T_2[11:0] ? image_1211 : _GEN_1210; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4284 = 12'h4bc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7356 = 12'h4bc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4284; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10428 = 12'h4bc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7356; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13500 = 12'h4bc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10428; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16572 = 12'h4bc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13500; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19644 = 12'h4bc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16572; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22716 = 12'h4bc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19644; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25788 = 12'h4bc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22716; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1212 = io_valid_in ? _GEN_25788 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1212 = 12'h4bc == _T_2[11:0] ? image_1212 : _GEN_1211; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4285 = 12'h4bd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7357 = 12'h4bd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4285; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10429 = 12'h4bd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7357; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13501 = 12'h4bd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10429; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16573 = 12'h4bd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13501; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19645 = 12'h4bd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16573; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22717 = 12'h4bd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19645; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25789 = 12'h4bd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22717; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1213 = io_valid_in ? _GEN_25789 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1213 = 12'h4bd == _T_2[11:0] ? image_1213 : _GEN_1212; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4286 = 12'h4be == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7358 = 12'h4be == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4286; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10430 = 12'h4be == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7358; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13502 = 12'h4be == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10430; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16574 = 12'h4be == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13502; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19646 = 12'h4be == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16574; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22718 = 12'h4be == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19646; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25790 = 12'h4be == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22718; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1214 = io_valid_in ? _GEN_25790 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1214 = 12'h4be == _T_2[11:0] ? image_1214 : _GEN_1213; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4287 = 12'h4bf == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7359 = 12'h4bf == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4287; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10431 = 12'h4bf == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7359; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13503 = 12'h4bf == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10431; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16575 = 12'h4bf == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13503; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19647 = 12'h4bf == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16575; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22719 = 12'h4bf == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19647; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25791 = 12'h4bf == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22719; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1215 = io_valid_in ? _GEN_25791 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1215 = 12'h4bf == _T_2[11:0] ? image_1215 : _GEN_1214; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4288 = 12'h4c0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7360 = 12'h4c0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4288; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10432 = 12'h4c0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7360; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13504 = 12'h4c0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10432; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16576 = 12'h4c0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13504; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19648 = 12'h4c0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16576; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22720 = 12'h4c0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19648; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25792 = 12'h4c0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22720; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1216 = io_valid_in ? _GEN_25792 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1216 = 12'h4c0 == _T_2[11:0] ? image_1216 : _GEN_1215; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4289 = 12'h4c1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7361 = 12'h4c1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4289; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10433 = 12'h4c1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7361; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13505 = 12'h4c1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10433; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16577 = 12'h4c1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13505; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19649 = 12'h4c1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16577; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22721 = 12'h4c1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19649; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25793 = 12'h4c1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22721; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1217 = io_valid_in ? _GEN_25793 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1217 = 12'h4c1 == _T_2[11:0] ? image_1217 : _GEN_1216; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4290 = 12'h4c2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7362 = 12'h4c2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4290; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10434 = 12'h4c2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7362; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13506 = 12'h4c2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10434; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16578 = 12'h4c2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13506; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19650 = 12'h4c2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16578; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22722 = 12'h4c2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19650; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25794 = 12'h4c2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22722; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1218 = io_valid_in ? _GEN_25794 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1218 = 12'h4c2 == _T_2[11:0] ? image_1218 : _GEN_1217; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4291 = 12'h4c3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7363 = 12'h4c3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4291; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10435 = 12'h4c3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7363; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13507 = 12'h4c3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10435; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16579 = 12'h4c3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13507; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19651 = 12'h4c3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16579; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22723 = 12'h4c3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19651; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25795 = 12'h4c3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22723; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1219 = io_valid_in ? _GEN_25795 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1219 = 12'h4c3 == _T_2[11:0] ? image_1219 : _GEN_1218; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4292 = 12'h4c4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7364 = 12'h4c4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4292; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10436 = 12'h4c4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7364; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13508 = 12'h4c4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10436; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16580 = 12'h4c4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13508; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19652 = 12'h4c4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16580; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22724 = 12'h4c4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19652; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25796 = 12'h4c4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22724; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1220 = io_valid_in ? _GEN_25796 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1220 = 12'h4c4 == _T_2[11:0] ? image_1220 : _GEN_1219; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4293 = 12'h4c5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7365 = 12'h4c5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4293; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10437 = 12'h4c5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7365; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13509 = 12'h4c5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10437; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16581 = 12'h4c5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13509; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19653 = 12'h4c5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16581; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22725 = 12'h4c5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19653; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25797 = 12'h4c5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22725; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1221 = io_valid_in ? _GEN_25797 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1221 = 12'h4c5 == _T_2[11:0] ? image_1221 : _GEN_1220; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4294 = 12'h4c6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7366 = 12'h4c6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4294; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10438 = 12'h4c6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7366; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13510 = 12'h4c6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10438; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16582 = 12'h4c6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13510; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19654 = 12'h4c6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16582; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22726 = 12'h4c6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19654; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25798 = 12'h4c6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22726; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1222 = io_valid_in ? _GEN_25798 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1222 = 12'h4c6 == _T_2[11:0] ? image_1222 : _GEN_1221; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4295 = 12'h4c7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7367 = 12'h4c7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4295; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10439 = 12'h4c7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7367; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13511 = 12'h4c7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10439; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16583 = 12'h4c7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13511; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19655 = 12'h4c7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16583; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22727 = 12'h4c7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19655; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25799 = 12'h4c7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22727; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1223 = io_valid_in ? _GEN_25799 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1223 = 12'h4c7 == _T_2[11:0] ? image_1223 : _GEN_1222; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4296 = 12'h4c8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7368 = 12'h4c8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4296; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10440 = 12'h4c8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7368; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13512 = 12'h4c8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10440; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16584 = 12'h4c8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13512; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19656 = 12'h4c8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16584; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22728 = 12'h4c8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19656; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25800 = 12'h4c8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22728; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1224 = io_valid_in ? _GEN_25800 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1224 = 12'h4c8 == _T_2[11:0] ? image_1224 : _GEN_1223; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4297 = 12'h4c9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7369 = 12'h4c9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4297; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10441 = 12'h4c9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7369; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13513 = 12'h4c9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10441; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16585 = 12'h4c9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13513; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19657 = 12'h4c9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16585; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22729 = 12'h4c9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19657; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25801 = 12'h4c9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22729; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1225 = io_valid_in ? _GEN_25801 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1225 = 12'h4c9 == _T_2[11:0] ? image_1225 : _GEN_1224; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4298 = 12'h4ca == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7370 = 12'h4ca == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4298; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10442 = 12'h4ca == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7370; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13514 = 12'h4ca == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10442; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16586 = 12'h4ca == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13514; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19658 = 12'h4ca == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16586; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22730 = 12'h4ca == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19658; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25802 = 12'h4ca == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22730; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1226 = io_valid_in ? _GEN_25802 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1226 = 12'h4ca == _T_2[11:0] ? image_1226 : _GEN_1225; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4299 = 12'h4cb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7371 = 12'h4cb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4299; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10443 = 12'h4cb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7371; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13515 = 12'h4cb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10443; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16587 = 12'h4cb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13515; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19659 = 12'h4cb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16587; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22731 = 12'h4cb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19659; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25803 = 12'h4cb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22731; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1227 = io_valid_in ? _GEN_25803 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1227 = 12'h4cb == _T_2[11:0] ? image_1227 : _GEN_1226; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4300 = 12'h4cc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7372 = 12'h4cc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4300; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10444 = 12'h4cc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7372; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13516 = 12'h4cc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10444; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16588 = 12'h4cc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13516; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19660 = 12'h4cc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16588; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22732 = 12'h4cc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19660; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25804 = 12'h4cc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22732; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1228 = io_valid_in ? _GEN_25804 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1228 = 12'h4cc == _T_2[11:0] ? image_1228 : _GEN_1227; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4301 = 12'h4cd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7373 = 12'h4cd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4301; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10445 = 12'h4cd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7373; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13517 = 12'h4cd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10445; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16589 = 12'h4cd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13517; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19661 = 12'h4cd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16589; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22733 = 12'h4cd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19661; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25805 = 12'h4cd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22733; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1229 = io_valid_in ? _GEN_25805 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1229 = 12'h4cd == _T_2[11:0] ? image_1229 : _GEN_1228; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4302 = 12'h4ce == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7374 = 12'h4ce == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4302; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10446 = 12'h4ce == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7374; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13518 = 12'h4ce == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10446; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16590 = 12'h4ce == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13518; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19662 = 12'h4ce == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16590; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22734 = 12'h4ce == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19662; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25806 = 12'h4ce == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22734; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1230 = io_valid_in ? _GEN_25806 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1230 = 12'h4ce == _T_2[11:0] ? image_1230 : _GEN_1229; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4303 = 12'h4cf == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7375 = 12'h4cf == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4303; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10447 = 12'h4cf == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7375; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13519 = 12'h4cf == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10447; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16591 = 12'h4cf == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13519; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19663 = 12'h4cf == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16591; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22735 = 12'h4cf == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19663; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25807 = 12'h4cf == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22735; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1231 = io_valid_in ? _GEN_25807 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1231 = 12'h4cf == _T_2[11:0] ? image_1231 : _GEN_1230; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4304 = 12'h4d0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7376 = 12'h4d0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4304; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10448 = 12'h4d0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7376; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13520 = 12'h4d0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10448; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16592 = 12'h4d0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13520; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19664 = 12'h4d0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16592; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22736 = 12'h4d0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19664; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25808 = 12'h4d0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22736; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1232 = io_valid_in ? _GEN_25808 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1232 = 12'h4d0 == _T_2[11:0] ? image_1232 : _GEN_1231; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4305 = 12'h4d1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7377 = 12'h4d1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4305; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10449 = 12'h4d1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7377; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13521 = 12'h4d1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10449; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16593 = 12'h4d1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13521; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19665 = 12'h4d1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16593; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22737 = 12'h4d1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19665; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25809 = 12'h4d1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22737; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1233 = io_valid_in ? _GEN_25809 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1233 = 12'h4d1 == _T_2[11:0] ? image_1233 : _GEN_1232; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4306 = 12'h4d2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7378 = 12'h4d2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4306; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10450 = 12'h4d2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7378; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13522 = 12'h4d2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10450; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16594 = 12'h4d2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13522; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19666 = 12'h4d2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16594; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22738 = 12'h4d2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19666; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25810 = 12'h4d2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22738; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1234 = io_valid_in ? _GEN_25810 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1234 = 12'h4d2 == _T_2[11:0] ? image_1234 : _GEN_1233; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4307 = 12'h4d3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7379 = 12'h4d3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4307; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10451 = 12'h4d3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7379; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13523 = 12'h4d3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10451; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16595 = 12'h4d3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13523; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19667 = 12'h4d3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16595; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22739 = 12'h4d3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19667; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25811 = 12'h4d3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22739; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1235 = io_valid_in ? _GEN_25811 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1235 = 12'h4d3 == _T_2[11:0] ? image_1235 : _GEN_1234; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4308 = 12'h4d4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7380 = 12'h4d4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4308; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10452 = 12'h4d4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7380; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13524 = 12'h4d4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10452; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16596 = 12'h4d4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13524; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19668 = 12'h4d4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16596; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22740 = 12'h4d4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19668; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25812 = 12'h4d4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22740; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1236 = io_valid_in ? _GEN_25812 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1236 = 12'h4d4 == _T_2[11:0] ? image_1236 : _GEN_1235; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4309 = 12'h4d5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7381 = 12'h4d5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4309; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10453 = 12'h4d5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7381; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13525 = 12'h4d5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10453; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16597 = 12'h4d5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13525; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19669 = 12'h4d5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16597; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22741 = 12'h4d5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19669; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25813 = 12'h4d5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22741; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1237 = io_valid_in ? _GEN_25813 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1237 = 12'h4d5 == _T_2[11:0] ? image_1237 : _GEN_1236; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4310 = 12'h4d6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7382 = 12'h4d6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4310; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10454 = 12'h4d6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7382; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13526 = 12'h4d6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10454; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16598 = 12'h4d6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13526; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19670 = 12'h4d6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16598; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22742 = 12'h4d6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19670; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25814 = 12'h4d6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22742; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1238 = io_valid_in ? _GEN_25814 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1238 = 12'h4d6 == _T_2[11:0] ? image_1238 : _GEN_1237; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4311 = 12'h4d7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7383 = 12'h4d7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4311; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10455 = 12'h4d7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7383; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13527 = 12'h4d7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10455; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16599 = 12'h4d7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13527; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19671 = 12'h4d7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16599; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22743 = 12'h4d7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19671; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25815 = 12'h4d7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22743; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1239 = io_valid_in ? _GEN_25815 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1239 = 12'h4d7 == _T_2[11:0] ? image_1239 : _GEN_1238; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4312 = 12'h4d8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7384 = 12'h4d8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4312; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10456 = 12'h4d8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7384; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13528 = 12'h4d8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10456; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16600 = 12'h4d8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13528; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19672 = 12'h4d8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16600; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22744 = 12'h4d8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19672; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25816 = 12'h4d8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22744; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1240 = io_valid_in ? _GEN_25816 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1240 = 12'h4d8 == _T_2[11:0] ? image_1240 : _GEN_1239; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4313 = 12'h4d9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7385 = 12'h4d9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4313; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10457 = 12'h4d9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7385; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13529 = 12'h4d9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10457; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16601 = 12'h4d9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13529; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19673 = 12'h4d9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16601; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22745 = 12'h4d9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19673; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25817 = 12'h4d9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22745; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1241 = io_valid_in ? _GEN_25817 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1241 = 12'h4d9 == _T_2[11:0] ? image_1241 : _GEN_1240; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4314 = 12'h4da == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7386 = 12'h4da == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4314; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10458 = 12'h4da == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7386; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13530 = 12'h4da == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10458; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16602 = 12'h4da == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13530; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19674 = 12'h4da == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16602; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22746 = 12'h4da == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19674; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25818 = 12'h4da == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22746; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1242 = io_valid_in ? _GEN_25818 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1242 = 12'h4da == _T_2[11:0] ? image_1242 : _GEN_1241; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4315 = 12'h4db == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7387 = 12'h4db == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4315; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10459 = 12'h4db == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7387; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13531 = 12'h4db == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10459; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16603 = 12'h4db == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13531; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19675 = 12'h4db == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16603; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22747 = 12'h4db == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19675; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25819 = 12'h4db == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22747; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1243 = io_valid_in ? _GEN_25819 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1243 = 12'h4db == _T_2[11:0] ? image_1243 : _GEN_1242; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4316 = 12'h4dc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7388 = 12'h4dc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4316; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10460 = 12'h4dc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7388; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13532 = 12'h4dc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10460; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16604 = 12'h4dc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13532; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19676 = 12'h4dc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16604; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22748 = 12'h4dc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19676; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25820 = 12'h4dc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22748; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1244 = io_valid_in ? _GEN_25820 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1244 = 12'h4dc == _T_2[11:0] ? image_1244 : _GEN_1243; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4317 = 12'h4dd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7389 = 12'h4dd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4317; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10461 = 12'h4dd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7389; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13533 = 12'h4dd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10461; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16605 = 12'h4dd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13533; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19677 = 12'h4dd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16605; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22749 = 12'h4dd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19677; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25821 = 12'h4dd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22749; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1245 = io_valid_in ? _GEN_25821 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1245 = 12'h4dd == _T_2[11:0] ? image_1245 : _GEN_1244; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4318 = 12'h4de == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7390 = 12'h4de == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4318; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10462 = 12'h4de == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7390; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13534 = 12'h4de == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10462; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16606 = 12'h4de == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13534; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19678 = 12'h4de == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16606; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22750 = 12'h4de == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19678; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25822 = 12'h4de == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22750; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1246 = io_valid_in ? _GEN_25822 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1246 = 12'h4de == _T_2[11:0] ? image_1246 : _GEN_1245; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4319 = 12'h4df == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7391 = 12'h4df == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4319; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10463 = 12'h4df == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7391; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13535 = 12'h4df == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10463; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16607 = 12'h4df == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13535; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19679 = 12'h4df == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16607; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22751 = 12'h4df == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19679; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25823 = 12'h4df == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22751; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1247 = io_valid_in ? _GEN_25823 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1247 = 12'h4df == _T_2[11:0] ? image_1247 : _GEN_1246; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4320 = 12'h4e0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7392 = 12'h4e0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4320; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10464 = 12'h4e0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7392; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13536 = 12'h4e0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10464; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16608 = 12'h4e0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13536; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19680 = 12'h4e0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16608; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22752 = 12'h4e0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19680; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25824 = 12'h4e0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22752; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1248 = io_valid_in ? _GEN_25824 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1248 = 12'h4e0 == _T_2[11:0] ? image_1248 : _GEN_1247; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4321 = 12'h4e1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7393 = 12'h4e1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4321; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10465 = 12'h4e1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7393; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13537 = 12'h4e1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10465; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16609 = 12'h4e1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13537; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19681 = 12'h4e1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16609; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22753 = 12'h4e1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19681; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25825 = 12'h4e1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22753; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1249 = io_valid_in ? _GEN_25825 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1249 = 12'h4e1 == _T_2[11:0] ? image_1249 : _GEN_1248; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4322 = 12'h4e2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7394 = 12'h4e2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4322; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10466 = 12'h4e2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7394; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13538 = 12'h4e2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10466; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16610 = 12'h4e2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13538; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19682 = 12'h4e2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16610; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22754 = 12'h4e2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19682; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25826 = 12'h4e2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22754; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1250 = io_valid_in ? _GEN_25826 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1250 = 12'h4e2 == _T_2[11:0] ? image_1250 : _GEN_1249; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4323 = 12'h4e3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7395 = 12'h4e3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4323; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10467 = 12'h4e3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7395; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13539 = 12'h4e3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10467; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16611 = 12'h4e3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13539; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19683 = 12'h4e3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16611; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22755 = 12'h4e3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19683; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25827 = 12'h4e3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22755; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1251 = io_valid_in ? _GEN_25827 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1251 = 12'h4e3 == _T_2[11:0] ? image_1251 : _GEN_1250; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4324 = 12'h4e4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7396 = 12'h4e4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4324; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10468 = 12'h4e4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7396; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13540 = 12'h4e4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10468; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16612 = 12'h4e4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13540; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19684 = 12'h4e4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16612; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22756 = 12'h4e4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19684; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25828 = 12'h4e4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22756; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1252 = io_valid_in ? _GEN_25828 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1252 = 12'h4e4 == _T_2[11:0] ? image_1252 : _GEN_1251; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4325 = 12'h4e5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7397 = 12'h4e5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4325; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10469 = 12'h4e5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7397; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13541 = 12'h4e5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10469; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16613 = 12'h4e5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13541; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19685 = 12'h4e5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16613; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22757 = 12'h4e5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19685; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25829 = 12'h4e5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22757; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1253 = io_valid_in ? _GEN_25829 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1253 = 12'h4e5 == _T_2[11:0] ? image_1253 : _GEN_1252; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4326 = 12'h4e6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7398 = 12'h4e6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4326; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10470 = 12'h4e6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7398; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13542 = 12'h4e6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10470; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16614 = 12'h4e6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13542; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19686 = 12'h4e6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16614; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22758 = 12'h4e6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19686; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25830 = 12'h4e6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22758; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1254 = io_valid_in ? _GEN_25830 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1254 = 12'h4e6 == _T_2[11:0] ? image_1254 : _GEN_1253; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4327 = 12'h4e7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7399 = 12'h4e7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4327; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10471 = 12'h4e7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7399; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13543 = 12'h4e7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10471; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16615 = 12'h4e7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13543; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19687 = 12'h4e7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16615; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22759 = 12'h4e7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19687; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25831 = 12'h4e7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22759; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1255 = io_valid_in ? _GEN_25831 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1255 = 12'h4e7 == _T_2[11:0] ? image_1255 : _GEN_1254; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4328 = 12'h4e8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7400 = 12'h4e8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4328; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10472 = 12'h4e8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7400; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13544 = 12'h4e8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10472; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16616 = 12'h4e8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13544; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19688 = 12'h4e8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16616; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22760 = 12'h4e8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19688; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25832 = 12'h4e8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22760; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1256 = io_valid_in ? _GEN_25832 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1256 = 12'h4e8 == _T_2[11:0] ? image_1256 : _GEN_1255; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4329 = 12'h4e9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7401 = 12'h4e9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4329; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10473 = 12'h4e9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7401; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13545 = 12'h4e9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10473; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16617 = 12'h4e9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13545; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19689 = 12'h4e9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16617; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22761 = 12'h4e9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19689; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25833 = 12'h4e9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22761; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1257 = io_valid_in ? _GEN_25833 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1257 = 12'h4e9 == _T_2[11:0] ? image_1257 : _GEN_1256; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4330 = 12'h4ea == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7402 = 12'h4ea == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4330; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10474 = 12'h4ea == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7402; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13546 = 12'h4ea == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10474; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16618 = 12'h4ea == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13546; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19690 = 12'h4ea == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16618; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22762 = 12'h4ea == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19690; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25834 = 12'h4ea == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22762; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1258 = io_valid_in ? _GEN_25834 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1258 = 12'h4ea == _T_2[11:0] ? image_1258 : _GEN_1257; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4331 = 12'h4eb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7403 = 12'h4eb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4331; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10475 = 12'h4eb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7403; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13547 = 12'h4eb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10475; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16619 = 12'h4eb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13547; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19691 = 12'h4eb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16619; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22763 = 12'h4eb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19691; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25835 = 12'h4eb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22763; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1259 = io_valid_in ? _GEN_25835 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1259 = 12'h4eb == _T_2[11:0] ? image_1259 : _GEN_1258; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4332 = 12'h4ec == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7404 = 12'h4ec == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4332; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10476 = 12'h4ec == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7404; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13548 = 12'h4ec == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10476; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16620 = 12'h4ec == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13548; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19692 = 12'h4ec == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16620; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22764 = 12'h4ec == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19692; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25836 = 12'h4ec == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22764; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1260 = io_valid_in ? _GEN_25836 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1260 = 12'h4ec == _T_2[11:0] ? image_1260 : _GEN_1259; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4333 = 12'h4ed == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7405 = 12'h4ed == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4333; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10477 = 12'h4ed == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7405; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13549 = 12'h4ed == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10477; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16621 = 12'h4ed == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13549; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19693 = 12'h4ed == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16621; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22765 = 12'h4ed == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19693; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25837 = 12'h4ed == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22765; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1261 = io_valid_in ? _GEN_25837 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1261 = 12'h4ed == _T_2[11:0] ? image_1261 : _GEN_1260; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4334 = 12'h4ee == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7406 = 12'h4ee == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4334; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10478 = 12'h4ee == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7406; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13550 = 12'h4ee == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10478; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16622 = 12'h4ee == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13550; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19694 = 12'h4ee == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16622; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22766 = 12'h4ee == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19694; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25838 = 12'h4ee == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22766; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1262 = io_valid_in ? _GEN_25838 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1262 = 12'h4ee == _T_2[11:0] ? image_1262 : _GEN_1261; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4335 = 12'h4ef == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7407 = 12'h4ef == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4335; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10479 = 12'h4ef == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7407; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13551 = 12'h4ef == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10479; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16623 = 12'h4ef == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13551; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19695 = 12'h4ef == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16623; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22767 = 12'h4ef == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19695; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25839 = 12'h4ef == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22767; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1263 = io_valid_in ? _GEN_25839 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1263 = 12'h4ef == _T_2[11:0] ? image_1263 : _GEN_1262; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4336 = 12'h4f0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7408 = 12'h4f0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4336; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10480 = 12'h4f0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7408; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13552 = 12'h4f0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10480; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16624 = 12'h4f0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13552; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19696 = 12'h4f0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16624; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22768 = 12'h4f0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19696; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25840 = 12'h4f0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22768; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1264 = io_valid_in ? _GEN_25840 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1264 = 12'h4f0 == _T_2[11:0] ? image_1264 : _GEN_1263; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4337 = 12'h4f1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7409 = 12'h4f1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4337; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10481 = 12'h4f1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7409; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13553 = 12'h4f1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10481; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16625 = 12'h4f1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13553; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19697 = 12'h4f1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16625; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22769 = 12'h4f1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19697; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25841 = 12'h4f1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22769; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1265 = io_valid_in ? _GEN_25841 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1265 = 12'h4f1 == _T_2[11:0] ? image_1265 : _GEN_1264; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4338 = 12'h4f2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7410 = 12'h4f2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4338; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10482 = 12'h4f2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7410; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13554 = 12'h4f2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10482; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16626 = 12'h4f2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13554; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19698 = 12'h4f2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16626; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22770 = 12'h4f2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19698; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25842 = 12'h4f2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22770; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1266 = io_valid_in ? _GEN_25842 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1266 = 12'h4f2 == _T_2[11:0] ? image_1266 : _GEN_1265; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4339 = 12'h4f3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7411 = 12'h4f3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4339; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10483 = 12'h4f3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7411; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13555 = 12'h4f3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10483; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16627 = 12'h4f3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13555; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19699 = 12'h4f3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16627; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22771 = 12'h4f3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19699; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25843 = 12'h4f3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22771; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1267 = io_valid_in ? _GEN_25843 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1267 = 12'h4f3 == _T_2[11:0] ? image_1267 : _GEN_1266; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4340 = 12'h4f4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7412 = 12'h4f4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4340; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10484 = 12'h4f4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7412; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13556 = 12'h4f4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10484; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16628 = 12'h4f4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13556; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19700 = 12'h4f4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16628; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22772 = 12'h4f4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19700; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25844 = 12'h4f4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22772; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1268 = io_valid_in ? _GEN_25844 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1268 = 12'h4f4 == _T_2[11:0] ? image_1268 : _GEN_1267; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4341 = 12'h4f5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7413 = 12'h4f5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4341; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10485 = 12'h4f5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7413; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13557 = 12'h4f5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10485; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16629 = 12'h4f5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13557; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19701 = 12'h4f5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16629; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22773 = 12'h4f5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19701; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25845 = 12'h4f5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22773; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1269 = io_valid_in ? _GEN_25845 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1269 = 12'h4f5 == _T_2[11:0] ? image_1269 : _GEN_1268; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4342 = 12'h4f6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7414 = 12'h4f6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4342; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10486 = 12'h4f6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7414; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13558 = 12'h4f6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10486; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16630 = 12'h4f6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13558; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19702 = 12'h4f6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16630; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22774 = 12'h4f6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19702; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25846 = 12'h4f6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22774; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1270 = io_valid_in ? _GEN_25846 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1270 = 12'h4f6 == _T_2[11:0] ? image_1270 : _GEN_1269; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4343 = 12'h4f7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7415 = 12'h4f7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4343; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10487 = 12'h4f7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7415; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13559 = 12'h4f7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10487; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16631 = 12'h4f7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13559; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19703 = 12'h4f7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16631; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22775 = 12'h4f7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19703; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25847 = 12'h4f7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22775; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1271 = io_valid_in ? _GEN_25847 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1271 = 12'h4f7 == _T_2[11:0] ? image_1271 : _GEN_1270; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4344 = 12'h4f8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7416 = 12'h4f8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4344; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10488 = 12'h4f8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7416; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13560 = 12'h4f8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10488; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16632 = 12'h4f8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13560; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19704 = 12'h4f8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16632; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22776 = 12'h4f8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19704; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25848 = 12'h4f8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22776; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1272 = io_valid_in ? _GEN_25848 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1272 = 12'h4f8 == _T_2[11:0] ? image_1272 : _GEN_1271; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4345 = 12'h4f9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7417 = 12'h4f9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4345; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10489 = 12'h4f9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7417; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13561 = 12'h4f9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10489; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16633 = 12'h4f9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13561; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19705 = 12'h4f9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16633; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22777 = 12'h4f9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19705; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25849 = 12'h4f9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22777; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1273 = io_valid_in ? _GEN_25849 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1273 = 12'h4f9 == _T_2[11:0] ? image_1273 : _GEN_1272; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4346 = 12'h4fa == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7418 = 12'h4fa == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4346; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10490 = 12'h4fa == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7418; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13562 = 12'h4fa == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10490; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16634 = 12'h4fa == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13562; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19706 = 12'h4fa == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16634; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22778 = 12'h4fa == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19706; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25850 = 12'h4fa == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22778; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1274 = io_valid_in ? _GEN_25850 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1274 = 12'h4fa == _T_2[11:0] ? image_1274 : _GEN_1273; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4347 = 12'h4fb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7419 = 12'h4fb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4347; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10491 = 12'h4fb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7419; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13563 = 12'h4fb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10491; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16635 = 12'h4fb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13563; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19707 = 12'h4fb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16635; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22779 = 12'h4fb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19707; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25851 = 12'h4fb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22779; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1275 = io_valid_in ? _GEN_25851 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1275 = 12'h4fb == _T_2[11:0] ? image_1275 : _GEN_1274; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4348 = 12'h4fc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7420 = 12'h4fc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4348; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10492 = 12'h4fc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7420; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13564 = 12'h4fc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10492; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16636 = 12'h4fc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13564; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19708 = 12'h4fc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16636; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22780 = 12'h4fc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19708; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25852 = 12'h4fc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22780; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1276 = io_valid_in ? _GEN_25852 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1276 = 12'h4fc == _T_2[11:0] ? image_1276 : _GEN_1275; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4349 = 12'h4fd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7421 = 12'h4fd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4349; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10493 = 12'h4fd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7421; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13565 = 12'h4fd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10493; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16637 = 12'h4fd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13565; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19709 = 12'h4fd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16637; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22781 = 12'h4fd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19709; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25853 = 12'h4fd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22781; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1277 = io_valid_in ? _GEN_25853 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1277 = 12'h4fd == _T_2[11:0] ? image_1277 : _GEN_1276; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4350 = 12'h4fe == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7422 = 12'h4fe == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4350; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10494 = 12'h4fe == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7422; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13566 = 12'h4fe == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10494; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16638 = 12'h4fe == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13566; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19710 = 12'h4fe == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16638; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22782 = 12'h4fe == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19710; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25854 = 12'h4fe == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22782; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1278 = io_valid_in ? _GEN_25854 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1278 = 12'h4fe == _T_2[11:0] ? image_1278 : _GEN_1277; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4351 = 12'h4ff == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7423 = 12'h4ff == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4351; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10495 = 12'h4ff == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7423; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13567 = 12'h4ff == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10495; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16639 = 12'h4ff == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13567; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19711 = 12'h4ff == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16639; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22783 = 12'h4ff == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19711; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25855 = 12'h4ff == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22783; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1279 = io_valid_in ? _GEN_25855 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1279 = 12'h4ff == _T_2[11:0] ? image_1279 : _GEN_1278; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4352 = 12'h500 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7424 = 12'h500 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4352; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10496 = 12'h500 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7424; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13568 = 12'h500 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10496; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16640 = 12'h500 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13568; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19712 = 12'h500 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16640; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22784 = 12'h500 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19712; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25856 = 12'h500 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22784; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1280 = io_valid_in ? _GEN_25856 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1280 = 12'h500 == _T_2[11:0] ? image_1280 : _GEN_1279; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4353 = 12'h501 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7425 = 12'h501 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4353; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10497 = 12'h501 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7425; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13569 = 12'h501 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10497; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16641 = 12'h501 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13569; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19713 = 12'h501 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16641; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22785 = 12'h501 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19713; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25857 = 12'h501 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22785; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1281 = io_valid_in ? _GEN_25857 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1281 = 12'h501 == _T_2[11:0] ? image_1281 : _GEN_1280; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4354 = 12'h502 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7426 = 12'h502 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4354; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10498 = 12'h502 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7426; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13570 = 12'h502 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10498; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16642 = 12'h502 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13570; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19714 = 12'h502 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16642; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22786 = 12'h502 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19714; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25858 = 12'h502 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22786; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1282 = io_valid_in ? _GEN_25858 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1282 = 12'h502 == _T_2[11:0] ? image_1282 : _GEN_1281; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4355 = 12'h503 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7427 = 12'h503 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4355; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10499 = 12'h503 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7427; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13571 = 12'h503 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10499; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16643 = 12'h503 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13571; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19715 = 12'h503 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16643; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22787 = 12'h503 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19715; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25859 = 12'h503 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22787; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1283 = io_valid_in ? _GEN_25859 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1283 = 12'h503 == _T_2[11:0] ? image_1283 : _GEN_1282; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4356 = 12'h504 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7428 = 12'h504 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4356; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10500 = 12'h504 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7428; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13572 = 12'h504 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10500; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16644 = 12'h504 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13572; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19716 = 12'h504 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16644; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22788 = 12'h504 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19716; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25860 = 12'h504 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22788; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1284 = io_valid_in ? _GEN_25860 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1284 = 12'h504 == _T_2[11:0] ? image_1284 : _GEN_1283; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4357 = 12'h505 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7429 = 12'h505 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4357; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10501 = 12'h505 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7429; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13573 = 12'h505 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10501; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16645 = 12'h505 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13573; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19717 = 12'h505 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16645; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22789 = 12'h505 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19717; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25861 = 12'h505 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22789; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1285 = io_valid_in ? _GEN_25861 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1285 = 12'h505 == _T_2[11:0] ? image_1285 : _GEN_1284; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4358 = 12'h506 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7430 = 12'h506 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4358; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10502 = 12'h506 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7430; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13574 = 12'h506 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10502; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16646 = 12'h506 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13574; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19718 = 12'h506 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16646; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22790 = 12'h506 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19718; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25862 = 12'h506 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22790; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1286 = io_valid_in ? _GEN_25862 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1286 = 12'h506 == _T_2[11:0] ? image_1286 : _GEN_1285; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4359 = 12'h507 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7431 = 12'h507 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4359; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10503 = 12'h507 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7431; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13575 = 12'h507 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10503; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16647 = 12'h507 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13575; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19719 = 12'h507 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16647; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22791 = 12'h507 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19719; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25863 = 12'h507 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22791; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1287 = io_valid_in ? _GEN_25863 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1287 = 12'h507 == _T_2[11:0] ? image_1287 : _GEN_1286; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4360 = 12'h508 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7432 = 12'h508 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4360; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10504 = 12'h508 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7432; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13576 = 12'h508 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10504; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16648 = 12'h508 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13576; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19720 = 12'h508 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16648; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22792 = 12'h508 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19720; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25864 = 12'h508 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22792; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1288 = io_valid_in ? _GEN_25864 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1288 = 12'h508 == _T_2[11:0] ? image_1288 : _GEN_1287; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4361 = 12'h509 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7433 = 12'h509 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4361; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10505 = 12'h509 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7433; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13577 = 12'h509 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10505; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16649 = 12'h509 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13577; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19721 = 12'h509 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16649; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22793 = 12'h509 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19721; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25865 = 12'h509 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22793; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1289 = io_valid_in ? _GEN_25865 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1289 = 12'h509 == _T_2[11:0] ? image_1289 : _GEN_1288; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4362 = 12'h50a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7434 = 12'h50a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4362; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10506 = 12'h50a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7434; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13578 = 12'h50a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10506; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16650 = 12'h50a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13578; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19722 = 12'h50a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16650; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22794 = 12'h50a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19722; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25866 = 12'h50a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22794; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1290 = io_valid_in ? _GEN_25866 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1290 = 12'h50a == _T_2[11:0] ? image_1290 : _GEN_1289; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4363 = 12'h50b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7435 = 12'h50b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4363; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10507 = 12'h50b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7435; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13579 = 12'h50b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10507; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16651 = 12'h50b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13579; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19723 = 12'h50b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16651; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22795 = 12'h50b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19723; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25867 = 12'h50b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22795; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1291 = io_valid_in ? _GEN_25867 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1291 = 12'h50b == _T_2[11:0] ? image_1291 : _GEN_1290; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4364 = 12'h50c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7436 = 12'h50c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4364; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10508 = 12'h50c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7436; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13580 = 12'h50c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10508; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16652 = 12'h50c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13580; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19724 = 12'h50c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16652; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22796 = 12'h50c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19724; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25868 = 12'h50c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22796; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1292 = io_valid_in ? _GEN_25868 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1292 = 12'h50c == _T_2[11:0] ? image_1292 : _GEN_1291; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4365 = 12'h50d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7437 = 12'h50d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4365; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10509 = 12'h50d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7437; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13581 = 12'h50d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10509; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16653 = 12'h50d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13581; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19725 = 12'h50d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16653; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22797 = 12'h50d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19725; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25869 = 12'h50d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22797; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1293 = io_valid_in ? _GEN_25869 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1293 = 12'h50d == _T_2[11:0] ? image_1293 : _GEN_1292; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4366 = 12'h50e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7438 = 12'h50e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4366; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10510 = 12'h50e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7438; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13582 = 12'h50e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10510; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16654 = 12'h50e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13582; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19726 = 12'h50e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16654; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22798 = 12'h50e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19726; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25870 = 12'h50e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22798; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1294 = io_valid_in ? _GEN_25870 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1294 = 12'h50e == _T_2[11:0] ? image_1294 : _GEN_1293; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4367 = 12'h50f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7439 = 12'h50f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4367; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10511 = 12'h50f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7439; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13583 = 12'h50f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10511; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16655 = 12'h50f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13583; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19727 = 12'h50f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16655; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22799 = 12'h50f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19727; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25871 = 12'h50f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22799; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1295 = io_valid_in ? _GEN_25871 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1295 = 12'h50f == _T_2[11:0] ? image_1295 : _GEN_1294; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4368 = 12'h510 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7440 = 12'h510 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4368; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10512 = 12'h510 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7440; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13584 = 12'h510 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10512; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16656 = 12'h510 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13584; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19728 = 12'h510 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16656; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22800 = 12'h510 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19728; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25872 = 12'h510 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22800; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1296 = io_valid_in ? _GEN_25872 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1296 = 12'h510 == _T_2[11:0] ? image_1296 : _GEN_1295; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4369 = 12'h511 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7441 = 12'h511 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4369; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10513 = 12'h511 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7441; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13585 = 12'h511 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10513; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16657 = 12'h511 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13585; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19729 = 12'h511 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16657; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22801 = 12'h511 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19729; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25873 = 12'h511 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22801; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1297 = io_valid_in ? _GEN_25873 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1297 = 12'h511 == _T_2[11:0] ? image_1297 : _GEN_1296; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4370 = 12'h512 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7442 = 12'h512 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4370; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10514 = 12'h512 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7442; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13586 = 12'h512 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10514; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16658 = 12'h512 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13586; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19730 = 12'h512 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16658; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22802 = 12'h512 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19730; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25874 = 12'h512 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22802; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1298 = io_valid_in ? _GEN_25874 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1298 = 12'h512 == _T_2[11:0] ? image_1298 : _GEN_1297; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4371 = 12'h513 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7443 = 12'h513 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4371; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10515 = 12'h513 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7443; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13587 = 12'h513 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10515; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16659 = 12'h513 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13587; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19731 = 12'h513 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16659; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22803 = 12'h513 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19731; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25875 = 12'h513 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22803; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1299 = io_valid_in ? _GEN_25875 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1299 = 12'h513 == _T_2[11:0] ? image_1299 : _GEN_1298; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4372 = 12'h514 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7444 = 12'h514 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4372; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10516 = 12'h514 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7444; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13588 = 12'h514 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10516; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16660 = 12'h514 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13588; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19732 = 12'h514 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16660; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22804 = 12'h514 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19732; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25876 = 12'h514 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22804; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1300 = io_valid_in ? _GEN_25876 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1300 = 12'h514 == _T_2[11:0] ? image_1300 : _GEN_1299; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4373 = 12'h515 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7445 = 12'h515 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4373; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10517 = 12'h515 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7445; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13589 = 12'h515 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10517; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16661 = 12'h515 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13589; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19733 = 12'h515 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16661; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22805 = 12'h515 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19733; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25877 = 12'h515 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22805; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1301 = io_valid_in ? _GEN_25877 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1301 = 12'h515 == _T_2[11:0] ? image_1301 : _GEN_1300; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4374 = 12'h516 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7446 = 12'h516 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4374; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10518 = 12'h516 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7446; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13590 = 12'h516 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10518; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16662 = 12'h516 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13590; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19734 = 12'h516 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16662; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22806 = 12'h516 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19734; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25878 = 12'h516 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22806; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1302 = io_valid_in ? _GEN_25878 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1302 = 12'h516 == _T_2[11:0] ? image_1302 : _GEN_1301; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4375 = 12'h517 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7447 = 12'h517 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4375; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10519 = 12'h517 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7447; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13591 = 12'h517 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10519; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16663 = 12'h517 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13591; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19735 = 12'h517 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16663; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22807 = 12'h517 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19735; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25879 = 12'h517 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22807; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1303 = io_valid_in ? _GEN_25879 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1303 = 12'h517 == _T_2[11:0] ? image_1303 : _GEN_1302; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4376 = 12'h518 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7448 = 12'h518 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4376; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10520 = 12'h518 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7448; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13592 = 12'h518 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10520; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16664 = 12'h518 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13592; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19736 = 12'h518 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16664; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22808 = 12'h518 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19736; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25880 = 12'h518 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22808; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1304 = io_valid_in ? _GEN_25880 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1304 = 12'h518 == _T_2[11:0] ? image_1304 : _GEN_1303; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4377 = 12'h519 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7449 = 12'h519 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4377; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10521 = 12'h519 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7449; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13593 = 12'h519 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10521; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16665 = 12'h519 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13593; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19737 = 12'h519 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16665; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22809 = 12'h519 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19737; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25881 = 12'h519 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22809; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1305 = io_valid_in ? _GEN_25881 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1305 = 12'h519 == _T_2[11:0] ? image_1305 : _GEN_1304; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4378 = 12'h51a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7450 = 12'h51a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4378; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10522 = 12'h51a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7450; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13594 = 12'h51a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10522; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16666 = 12'h51a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13594; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19738 = 12'h51a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16666; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22810 = 12'h51a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19738; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25882 = 12'h51a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22810; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1306 = io_valid_in ? _GEN_25882 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1306 = 12'h51a == _T_2[11:0] ? image_1306 : _GEN_1305; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4379 = 12'h51b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7451 = 12'h51b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4379; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10523 = 12'h51b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7451; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13595 = 12'h51b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10523; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16667 = 12'h51b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13595; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19739 = 12'h51b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16667; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22811 = 12'h51b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19739; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25883 = 12'h51b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22811; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1307 = io_valid_in ? _GEN_25883 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1307 = 12'h51b == _T_2[11:0] ? image_1307 : _GEN_1306; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4380 = 12'h51c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7452 = 12'h51c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4380; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10524 = 12'h51c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7452; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13596 = 12'h51c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10524; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16668 = 12'h51c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13596; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19740 = 12'h51c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16668; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22812 = 12'h51c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19740; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25884 = 12'h51c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22812; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1308 = io_valid_in ? _GEN_25884 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1308 = 12'h51c == _T_2[11:0] ? image_1308 : _GEN_1307; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4381 = 12'h51d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7453 = 12'h51d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4381; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10525 = 12'h51d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7453; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13597 = 12'h51d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10525; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16669 = 12'h51d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13597; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19741 = 12'h51d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16669; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22813 = 12'h51d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19741; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25885 = 12'h51d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22813; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1309 = io_valid_in ? _GEN_25885 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1309 = 12'h51d == _T_2[11:0] ? image_1309 : _GEN_1308; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4382 = 12'h51e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7454 = 12'h51e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4382; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10526 = 12'h51e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7454; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13598 = 12'h51e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10526; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16670 = 12'h51e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13598; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19742 = 12'h51e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16670; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22814 = 12'h51e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19742; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25886 = 12'h51e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22814; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1310 = io_valid_in ? _GEN_25886 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1310 = 12'h51e == _T_2[11:0] ? image_1310 : _GEN_1309; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4383 = 12'h51f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7455 = 12'h51f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4383; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10527 = 12'h51f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7455; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13599 = 12'h51f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10527; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16671 = 12'h51f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13599; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19743 = 12'h51f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16671; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22815 = 12'h51f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19743; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25887 = 12'h51f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22815; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1311 = io_valid_in ? _GEN_25887 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1311 = 12'h51f == _T_2[11:0] ? image_1311 : _GEN_1310; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4384 = 12'h520 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7456 = 12'h520 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4384; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10528 = 12'h520 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7456; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13600 = 12'h520 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10528; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16672 = 12'h520 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13600; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19744 = 12'h520 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16672; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22816 = 12'h520 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19744; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25888 = 12'h520 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22816; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1312 = io_valid_in ? _GEN_25888 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1312 = 12'h520 == _T_2[11:0] ? image_1312 : _GEN_1311; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4385 = 12'h521 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7457 = 12'h521 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4385; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10529 = 12'h521 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7457; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13601 = 12'h521 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10529; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16673 = 12'h521 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13601; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19745 = 12'h521 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16673; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22817 = 12'h521 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19745; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25889 = 12'h521 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22817; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1313 = io_valid_in ? _GEN_25889 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1313 = 12'h521 == _T_2[11:0] ? image_1313 : _GEN_1312; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4386 = 12'h522 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7458 = 12'h522 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4386; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10530 = 12'h522 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7458; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13602 = 12'h522 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10530; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16674 = 12'h522 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13602; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19746 = 12'h522 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16674; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22818 = 12'h522 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19746; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25890 = 12'h522 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22818; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1314 = io_valid_in ? _GEN_25890 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1314 = 12'h522 == _T_2[11:0] ? image_1314 : _GEN_1313; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4387 = 12'h523 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7459 = 12'h523 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4387; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10531 = 12'h523 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7459; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13603 = 12'h523 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10531; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16675 = 12'h523 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13603; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19747 = 12'h523 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16675; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22819 = 12'h523 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19747; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25891 = 12'h523 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22819; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1315 = io_valid_in ? _GEN_25891 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1315 = 12'h523 == _T_2[11:0] ? image_1315 : _GEN_1314; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4388 = 12'h524 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7460 = 12'h524 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4388; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10532 = 12'h524 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7460; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13604 = 12'h524 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10532; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16676 = 12'h524 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13604; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19748 = 12'h524 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16676; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22820 = 12'h524 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19748; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25892 = 12'h524 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22820; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1316 = io_valid_in ? _GEN_25892 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1316 = 12'h524 == _T_2[11:0] ? image_1316 : _GEN_1315; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4389 = 12'h525 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7461 = 12'h525 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4389; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10533 = 12'h525 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7461; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13605 = 12'h525 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10533; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16677 = 12'h525 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13605; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19749 = 12'h525 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16677; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22821 = 12'h525 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19749; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25893 = 12'h525 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22821; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1317 = io_valid_in ? _GEN_25893 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1317 = 12'h525 == _T_2[11:0] ? image_1317 : _GEN_1316; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4390 = 12'h526 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7462 = 12'h526 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4390; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10534 = 12'h526 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7462; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13606 = 12'h526 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10534; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16678 = 12'h526 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13606; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19750 = 12'h526 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16678; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22822 = 12'h526 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19750; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25894 = 12'h526 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22822; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1318 = io_valid_in ? _GEN_25894 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1318 = 12'h526 == _T_2[11:0] ? image_1318 : _GEN_1317; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4391 = 12'h527 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7463 = 12'h527 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4391; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10535 = 12'h527 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7463; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13607 = 12'h527 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10535; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16679 = 12'h527 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13607; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19751 = 12'h527 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16679; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22823 = 12'h527 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19751; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25895 = 12'h527 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22823; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1319 = io_valid_in ? _GEN_25895 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1319 = 12'h527 == _T_2[11:0] ? image_1319 : _GEN_1318; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4392 = 12'h528 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7464 = 12'h528 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4392; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10536 = 12'h528 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7464; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13608 = 12'h528 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10536; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16680 = 12'h528 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13608; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19752 = 12'h528 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16680; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22824 = 12'h528 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19752; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25896 = 12'h528 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22824; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1320 = io_valid_in ? _GEN_25896 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1320 = 12'h528 == _T_2[11:0] ? image_1320 : _GEN_1319; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4393 = 12'h529 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7465 = 12'h529 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4393; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10537 = 12'h529 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7465; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13609 = 12'h529 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10537; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16681 = 12'h529 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13609; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19753 = 12'h529 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16681; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22825 = 12'h529 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19753; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25897 = 12'h529 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22825; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1321 = io_valid_in ? _GEN_25897 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1321 = 12'h529 == _T_2[11:0] ? image_1321 : _GEN_1320; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4394 = 12'h52a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7466 = 12'h52a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4394; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10538 = 12'h52a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7466; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13610 = 12'h52a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10538; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16682 = 12'h52a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13610; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19754 = 12'h52a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16682; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22826 = 12'h52a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19754; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25898 = 12'h52a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22826; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1322 = io_valid_in ? _GEN_25898 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1322 = 12'h52a == _T_2[11:0] ? image_1322 : _GEN_1321; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4395 = 12'h52b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7467 = 12'h52b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4395; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10539 = 12'h52b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7467; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13611 = 12'h52b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10539; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16683 = 12'h52b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13611; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19755 = 12'h52b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16683; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22827 = 12'h52b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19755; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25899 = 12'h52b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22827; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1323 = io_valid_in ? _GEN_25899 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1323 = 12'h52b == _T_2[11:0] ? image_1323 : _GEN_1322; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4396 = 12'h52c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7468 = 12'h52c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4396; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10540 = 12'h52c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7468; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13612 = 12'h52c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10540; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16684 = 12'h52c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13612; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19756 = 12'h52c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16684; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22828 = 12'h52c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19756; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25900 = 12'h52c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22828; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1324 = io_valid_in ? _GEN_25900 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1324 = 12'h52c == _T_2[11:0] ? image_1324 : _GEN_1323; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4397 = 12'h52d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7469 = 12'h52d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4397; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10541 = 12'h52d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7469; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13613 = 12'h52d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10541; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16685 = 12'h52d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13613; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19757 = 12'h52d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16685; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22829 = 12'h52d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19757; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25901 = 12'h52d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22829; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1325 = io_valid_in ? _GEN_25901 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1325 = 12'h52d == _T_2[11:0] ? image_1325 : _GEN_1324; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4398 = 12'h52e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7470 = 12'h52e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4398; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10542 = 12'h52e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7470; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13614 = 12'h52e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10542; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16686 = 12'h52e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13614; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19758 = 12'h52e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16686; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22830 = 12'h52e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19758; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25902 = 12'h52e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22830; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1326 = io_valid_in ? _GEN_25902 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1326 = 12'h52e == _T_2[11:0] ? image_1326 : _GEN_1325; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4399 = 12'h52f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7471 = 12'h52f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4399; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10543 = 12'h52f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7471; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13615 = 12'h52f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10543; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16687 = 12'h52f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13615; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19759 = 12'h52f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16687; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22831 = 12'h52f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19759; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25903 = 12'h52f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22831; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1327 = io_valid_in ? _GEN_25903 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1327 = 12'h52f == _T_2[11:0] ? image_1327 : _GEN_1326; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4400 = 12'h530 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7472 = 12'h530 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4400; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10544 = 12'h530 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7472; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13616 = 12'h530 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10544; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16688 = 12'h530 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13616; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19760 = 12'h530 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16688; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22832 = 12'h530 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19760; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25904 = 12'h530 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22832; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1328 = io_valid_in ? _GEN_25904 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1328 = 12'h530 == _T_2[11:0] ? image_1328 : _GEN_1327; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4401 = 12'h531 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7473 = 12'h531 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4401; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10545 = 12'h531 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7473; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13617 = 12'h531 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10545; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16689 = 12'h531 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13617; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19761 = 12'h531 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16689; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22833 = 12'h531 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19761; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25905 = 12'h531 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22833; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1329 = io_valid_in ? _GEN_25905 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1329 = 12'h531 == _T_2[11:0] ? image_1329 : _GEN_1328; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4402 = 12'h532 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7474 = 12'h532 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4402; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10546 = 12'h532 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7474; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13618 = 12'h532 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10546; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16690 = 12'h532 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13618; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19762 = 12'h532 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16690; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22834 = 12'h532 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19762; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25906 = 12'h532 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22834; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1330 = io_valid_in ? _GEN_25906 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1330 = 12'h532 == _T_2[11:0] ? image_1330 : _GEN_1329; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4403 = 12'h533 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7475 = 12'h533 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4403; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10547 = 12'h533 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7475; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13619 = 12'h533 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10547; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16691 = 12'h533 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13619; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19763 = 12'h533 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16691; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22835 = 12'h533 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19763; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25907 = 12'h533 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22835; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1331 = io_valid_in ? _GEN_25907 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1331 = 12'h533 == _T_2[11:0] ? image_1331 : _GEN_1330; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4404 = 12'h534 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7476 = 12'h534 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4404; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10548 = 12'h534 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7476; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13620 = 12'h534 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10548; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16692 = 12'h534 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13620; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19764 = 12'h534 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16692; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22836 = 12'h534 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19764; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25908 = 12'h534 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22836; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1332 = io_valid_in ? _GEN_25908 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1332 = 12'h534 == _T_2[11:0] ? image_1332 : _GEN_1331; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4405 = 12'h535 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7477 = 12'h535 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4405; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10549 = 12'h535 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7477; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13621 = 12'h535 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10549; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16693 = 12'h535 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13621; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19765 = 12'h535 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16693; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22837 = 12'h535 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19765; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25909 = 12'h535 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22837; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1333 = io_valid_in ? _GEN_25909 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1333 = 12'h535 == _T_2[11:0] ? image_1333 : _GEN_1332; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4406 = 12'h536 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7478 = 12'h536 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4406; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10550 = 12'h536 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7478; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13622 = 12'h536 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10550; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16694 = 12'h536 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13622; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19766 = 12'h536 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16694; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22838 = 12'h536 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19766; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25910 = 12'h536 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22838; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1334 = io_valid_in ? _GEN_25910 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1334 = 12'h536 == _T_2[11:0] ? image_1334 : _GEN_1333; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4407 = 12'h537 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7479 = 12'h537 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4407; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10551 = 12'h537 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7479; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13623 = 12'h537 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10551; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16695 = 12'h537 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13623; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19767 = 12'h537 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16695; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22839 = 12'h537 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19767; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25911 = 12'h537 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22839; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1335 = io_valid_in ? _GEN_25911 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1335 = 12'h537 == _T_2[11:0] ? image_1335 : _GEN_1334; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4408 = 12'h538 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7480 = 12'h538 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4408; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10552 = 12'h538 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7480; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13624 = 12'h538 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10552; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16696 = 12'h538 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13624; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19768 = 12'h538 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16696; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22840 = 12'h538 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19768; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25912 = 12'h538 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22840; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1336 = io_valid_in ? _GEN_25912 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1336 = 12'h538 == _T_2[11:0] ? image_1336 : _GEN_1335; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4409 = 12'h539 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7481 = 12'h539 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4409; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10553 = 12'h539 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7481; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13625 = 12'h539 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10553; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16697 = 12'h539 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13625; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19769 = 12'h539 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16697; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22841 = 12'h539 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19769; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25913 = 12'h539 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22841; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1337 = io_valid_in ? _GEN_25913 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1337 = 12'h539 == _T_2[11:0] ? image_1337 : _GEN_1336; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4410 = 12'h53a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7482 = 12'h53a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4410; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10554 = 12'h53a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7482; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13626 = 12'h53a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10554; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16698 = 12'h53a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13626; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19770 = 12'h53a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16698; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22842 = 12'h53a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19770; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25914 = 12'h53a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22842; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1338 = io_valid_in ? _GEN_25914 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1338 = 12'h53a == _T_2[11:0] ? image_1338 : _GEN_1337; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4411 = 12'h53b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7483 = 12'h53b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4411; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10555 = 12'h53b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7483; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13627 = 12'h53b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10555; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16699 = 12'h53b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13627; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19771 = 12'h53b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16699; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22843 = 12'h53b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19771; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25915 = 12'h53b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22843; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1339 = io_valid_in ? _GEN_25915 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1339 = 12'h53b == _T_2[11:0] ? image_1339 : _GEN_1338; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4412 = 12'h53c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7484 = 12'h53c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4412; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10556 = 12'h53c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7484; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13628 = 12'h53c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10556; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16700 = 12'h53c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13628; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19772 = 12'h53c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16700; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22844 = 12'h53c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19772; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25916 = 12'h53c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22844; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1340 = io_valid_in ? _GEN_25916 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1340 = 12'h53c == _T_2[11:0] ? image_1340 : _GEN_1339; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4413 = 12'h53d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7485 = 12'h53d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4413; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10557 = 12'h53d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7485; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13629 = 12'h53d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10557; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16701 = 12'h53d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13629; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19773 = 12'h53d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16701; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22845 = 12'h53d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19773; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25917 = 12'h53d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22845; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1341 = io_valid_in ? _GEN_25917 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1341 = 12'h53d == _T_2[11:0] ? image_1341 : _GEN_1340; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4414 = 12'h53e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7486 = 12'h53e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4414; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10558 = 12'h53e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7486; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13630 = 12'h53e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10558; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16702 = 12'h53e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13630; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19774 = 12'h53e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16702; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22846 = 12'h53e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19774; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25918 = 12'h53e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22846; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1342 = io_valid_in ? _GEN_25918 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1342 = 12'h53e == _T_2[11:0] ? image_1342 : _GEN_1341; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4415 = 12'h53f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7487 = 12'h53f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4415; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10559 = 12'h53f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7487; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13631 = 12'h53f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10559; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16703 = 12'h53f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13631; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19775 = 12'h53f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16703; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22847 = 12'h53f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19775; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25919 = 12'h53f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22847; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1343 = io_valid_in ? _GEN_25919 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1343 = 12'h53f == _T_2[11:0] ? image_1343 : _GEN_1342; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4416 = 12'h540 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7488 = 12'h540 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4416; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10560 = 12'h540 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7488; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13632 = 12'h540 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10560; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16704 = 12'h540 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13632; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19776 = 12'h540 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16704; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22848 = 12'h540 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19776; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25920 = 12'h540 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22848; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1344 = io_valid_in ? _GEN_25920 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1344 = 12'h540 == _T_2[11:0] ? image_1344 : _GEN_1343; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4417 = 12'h541 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7489 = 12'h541 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4417; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10561 = 12'h541 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7489; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13633 = 12'h541 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10561; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16705 = 12'h541 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13633; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19777 = 12'h541 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16705; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22849 = 12'h541 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19777; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25921 = 12'h541 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22849; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1345 = io_valid_in ? _GEN_25921 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1345 = 12'h541 == _T_2[11:0] ? image_1345 : _GEN_1344; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4418 = 12'h542 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7490 = 12'h542 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4418; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10562 = 12'h542 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7490; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13634 = 12'h542 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10562; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16706 = 12'h542 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13634; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19778 = 12'h542 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16706; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22850 = 12'h542 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19778; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25922 = 12'h542 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22850; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1346 = io_valid_in ? _GEN_25922 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1346 = 12'h542 == _T_2[11:0] ? image_1346 : _GEN_1345; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4419 = 12'h543 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7491 = 12'h543 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4419; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10563 = 12'h543 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7491; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13635 = 12'h543 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10563; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16707 = 12'h543 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13635; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19779 = 12'h543 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16707; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22851 = 12'h543 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19779; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25923 = 12'h543 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22851; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1347 = io_valid_in ? _GEN_25923 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1347 = 12'h543 == _T_2[11:0] ? image_1347 : _GEN_1346; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4420 = 12'h544 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7492 = 12'h544 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4420; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10564 = 12'h544 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7492; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13636 = 12'h544 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10564; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16708 = 12'h544 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13636; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19780 = 12'h544 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16708; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22852 = 12'h544 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19780; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25924 = 12'h544 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22852; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1348 = io_valid_in ? _GEN_25924 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1348 = 12'h544 == _T_2[11:0] ? image_1348 : _GEN_1347; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4421 = 12'h545 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7493 = 12'h545 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4421; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10565 = 12'h545 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7493; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13637 = 12'h545 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10565; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16709 = 12'h545 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13637; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19781 = 12'h545 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16709; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22853 = 12'h545 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19781; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25925 = 12'h545 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22853; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1349 = io_valid_in ? _GEN_25925 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1349 = 12'h545 == _T_2[11:0] ? image_1349 : _GEN_1348; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4422 = 12'h546 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7494 = 12'h546 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4422; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10566 = 12'h546 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7494; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13638 = 12'h546 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10566; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16710 = 12'h546 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13638; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19782 = 12'h546 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16710; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22854 = 12'h546 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19782; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25926 = 12'h546 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22854; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1350 = io_valid_in ? _GEN_25926 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1350 = 12'h546 == _T_2[11:0] ? image_1350 : _GEN_1349; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4423 = 12'h547 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7495 = 12'h547 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4423; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10567 = 12'h547 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7495; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13639 = 12'h547 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10567; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16711 = 12'h547 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13639; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19783 = 12'h547 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16711; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22855 = 12'h547 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19783; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25927 = 12'h547 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22855; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1351 = io_valid_in ? _GEN_25927 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1351 = 12'h547 == _T_2[11:0] ? image_1351 : _GEN_1350; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4424 = 12'h548 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7496 = 12'h548 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4424; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10568 = 12'h548 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7496; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13640 = 12'h548 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10568; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16712 = 12'h548 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13640; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19784 = 12'h548 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16712; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22856 = 12'h548 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19784; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25928 = 12'h548 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22856; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1352 = io_valid_in ? _GEN_25928 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1352 = 12'h548 == _T_2[11:0] ? image_1352 : _GEN_1351; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4425 = 12'h549 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7497 = 12'h549 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4425; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10569 = 12'h549 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7497; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13641 = 12'h549 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10569; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16713 = 12'h549 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13641; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19785 = 12'h549 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16713; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22857 = 12'h549 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19785; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25929 = 12'h549 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22857; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1353 = io_valid_in ? _GEN_25929 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1353 = 12'h549 == _T_2[11:0] ? image_1353 : _GEN_1352; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4426 = 12'h54a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7498 = 12'h54a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4426; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10570 = 12'h54a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7498; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13642 = 12'h54a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10570; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16714 = 12'h54a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13642; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19786 = 12'h54a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16714; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22858 = 12'h54a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19786; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25930 = 12'h54a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22858; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1354 = io_valid_in ? _GEN_25930 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1354 = 12'h54a == _T_2[11:0] ? image_1354 : _GEN_1353; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4427 = 12'h54b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7499 = 12'h54b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4427; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10571 = 12'h54b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7499; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13643 = 12'h54b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10571; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16715 = 12'h54b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13643; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19787 = 12'h54b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16715; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22859 = 12'h54b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19787; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25931 = 12'h54b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22859; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1355 = io_valid_in ? _GEN_25931 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1355 = 12'h54b == _T_2[11:0] ? image_1355 : _GEN_1354; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4428 = 12'h54c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7500 = 12'h54c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4428; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10572 = 12'h54c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7500; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13644 = 12'h54c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10572; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16716 = 12'h54c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13644; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19788 = 12'h54c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16716; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22860 = 12'h54c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19788; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25932 = 12'h54c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22860; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1356 = io_valid_in ? _GEN_25932 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1356 = 12'h54c == _T_2[11:0] ? image_1356 : _GEN_1355; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4429 = 12'h54d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7501 = 12'h54d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4429; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10573 = 12'h54d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7501; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13645 = 12'h54d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10573; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16717 = 12'h54d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13645; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19789 = 12'h54d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16717; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22861 = 12'h54d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19789; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25933 = 12'h54d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22861; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1357 = io_valid_in ? _GEN_25933 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1357 = 12'h54d == _T_2[11:0] ? image_1357 : _GEN_1356; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4430 = 12'h54e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7502 = 12'h54e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4430; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10574 = 12'h54e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7502; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13646 = 12'h54e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10574; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16718 = 12'h54e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13646; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19790 = 12'h54e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16718; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22862 = 12'h54e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19790; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25934 = 12'h54e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22862; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1358 = io_valid_in ? _GEN_25934 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1358 = 12'h54e == _T_2[11:0] ? image_1358 : _GEN_1357; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4431 = 12'h54f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7503 = 12'h54f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4431; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10575 = 12'h54f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7503; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13647 = 12'h54f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10575; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16719 = 12'h54f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13647; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19791 = 12'h54f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16719; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22863 = 12'h54f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19791; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25935 = 12'h54f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22863; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1359 = io_valid_in ? _GEN_25935 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1359 = 12'h54f == _T_2[11:0] ? image_1359 : _GEN_1358; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4432 = 12'h550 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7504 = 12'h550 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4432; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10576 = 12'h550 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7504; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13648 = 12'h550 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10576; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16720 = 12'h550 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13648; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19792 = 12'h550 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16720; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22864 = 12'h550 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19792; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25936 = 12'h550 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22864; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1360 = io_valid_in ? _GEN_25936 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1360 = 12'h550 == _T_2[11:0] ? image_1360 : _GEN_1359; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4433 = 12'h551 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7505 = 12'h551 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4433; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10577 = 12'h551 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7505; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13649 = 12'h551 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10577; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16721 = 12'h551 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13649; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19793 = 12'h551 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16721; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22865 = 12'h551 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19793; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25937 = 12'h551 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22865; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1361 = io_valid_in ? _GEN_25937 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1361 = 12'h551 == _T_2[11:0] ? image_1361 : _GEN_1360; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4434 = 12'h552 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7506 = 12'h552 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4434; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10578 = 12'h552 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7506; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13650 = 12'h552 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10578; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16722 = 12'h552 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13650; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19794 = 12'h552 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16722; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22866 = 12'h552 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19794; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25938 = 12'h552 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22866; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1362 = io_valid_in ? _GEN_25938 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1362 = 12'h552 == _T_2[11:0] ? image_1362 : _GEN_1361; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4435 = 12'h553 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7507 = 12'h553 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4435; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10579 = 12'h553 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7507; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13651 = 12'h553 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10579; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16723 = 12'h553 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13651; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19795 = 12'h553 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16723; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22867 = 12'h553 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19795; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25939 = 12'h553 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22867; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1363 = io_valid_in ? _GEN_25939 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1363 = 12'h553 == _T_2[11:0] ? image_1363 : _GEN_1362; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4436 = 12'h554 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7508 = 12'h554 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4436; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10580 = 12'h554 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7508; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13652 = 12'h554 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10580; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16724 = 12'h554 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13652; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19796 = 12'h554 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16724; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22868 = 12'h554 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19796; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25940 = 12'h554 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22868; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1364 = io_valid_in ? _GEN_25940 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1364 = 12'h554 == _T_2[11:0] ? image_1364 : _GEN_1363; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4437 = 12'h555 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7509 = 12'h555 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4437; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10581 = 12'h555 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7509; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13653 = 12'h555 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10581; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16725 = 12'h555 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13653; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19797 = 12'h555 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16725; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22869 = 12'h555 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19797; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25941 = 12'h555 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22869; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1365 = io_valid_in ? _GEN_25941 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1365 = 12'h555 == _T_2[11:0] ? image_1365 : _GEN_1364; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4438 = 12'h556 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7510 = 12'h556 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4438; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10582 = 12'h556 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7510; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13654 = 12'h556 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10582; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16726 = 12'h556 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13654; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19798 = 12'h556 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16726; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22870 = 12'h556 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19798; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25942 = 12'h556 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22870; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1366 = io_valid_in ? _GEN_25942 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1366 = 12'h556 == _T_2[11:0] ? image_1366 : _GEN_1365; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4439 = 12'h557 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7511 = 12'h557 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4439; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10583 = 12'h557 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7511; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13655 = 12'h557 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10583; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16727 = 12'h557 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13655; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19799 = 12'h557 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16727; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22871 = 12'h557 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19799; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25943 = 12'h557 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22871; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1367 = io_valid_in ? _GEN_25943 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1367 = 12'h557 == _T_2[11:0] ? image_1367 : _GEN_1366; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4440 = 12'h558 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7512 = 12'h558 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4440; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10584 = 12'h558 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7512; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13656 = 12'h558 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10584; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16728 = 12'h558 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13656; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19800 = 12'h558 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16728; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22872 = 12'h558 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19800; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25944 = 12'h558 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22872; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1368 = io_valid_in ? _GEN_25944 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1368 = 12'h558 == _T_2[11:0] ? image_1368 : _GEN_1367; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4441 = 12'h559 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7513 = 12'h559 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4441; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10585 = 12'h559 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7513; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13657 = 12'h559 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10585; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16729 = 12'h559 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13657; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19801 = 12'h559 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16729; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22873 = 12'h559 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19801; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25945 = 12'h559 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22873; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1369 = io_valid_in ? _GEN_25945 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1369 = 12'h559 == _T_2[11:0] ? image_1369 : _GEN_1368; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4442 = 12'h55a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7514 = 12'h55a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4442; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10586 = 12'h55a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7514; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13658 = 12'h55a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10586; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16730 = 12'h55a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13658; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19802 = 12'h55a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16730; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22874 = 12'h55a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19802; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25946 = 12'h55a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22874; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1370 = io_valid_in ? _GEN_25946 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1370 = 12'h55a == _T_2[11:0] ? image_1370 : _GEN_1369; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4443 = 12'h55b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7515 = 12'h55b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4443; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10587 = 12'h55b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7515; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13659 = 12'h55b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10587; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16731 = 12'h55b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13659; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19803 = 12'h55b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16731; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22875 = 12'h55b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19803; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25947 = 12'h55b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22875; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1371 = io_valid_in ? _GEN_25947 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1371 = 12'h55b == _T_2[11:0] ? image_1371 : _GEN_1370; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4444 = 12'h55c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7516 = 12'h55c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4444; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10588 = 12'h55c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7516; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13660 = 12'h55c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10588; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16732 = 12'h55c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13660; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19804 = 12'h55c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16732; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22876 = 12'h55c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19804; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25948 = 12'h55c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22876; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1372 = io_valid_in ? _GEN_25948 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1372 = 12'h55c == _T_2[11:0] ? image_1372 : _GEN_1371; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4445 = 12'h55d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7517 = 12'h55d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4445; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10589 = 12'h55d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7517; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13661 = 12'h55d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10589; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16733 = 12'h55d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13661; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19805 = 12'h55d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16733; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22877 = 12'h55d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19805; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25949 = 12'h55d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22877; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1373 = io_valid_in ? _GEN_25949 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1373 = 12'h55d == _T_2[11:0] ? image_1373 : _GEN_1372; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4446 = 12'h55e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7518 = 12'h55e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4446; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10590 = 12'h55e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7518; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13662 = 12'h55e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10590; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16734 = 12'h55e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13662; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19806 = 12'h55e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16734; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22878 = 12'h55e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19806; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25950 = 12'h55e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22878; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1374 = io_valid_in ? _GEN_25950 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1374 = 12'h55e == _T_2[11:0] ? image_1374 : _GEN_1373; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4447 = 12'h55f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7519 = 12'h55f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4447; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10591 = 12'h55f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7519; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13663 = 12'h55f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10591; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16735 = 12'h55f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13663; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19807 = 12'h55f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16735; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22879 = 12'h55f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19807; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25951 = 12'h55f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22879; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1375 = io_valid_in ? _GEN_25951 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1375 = 12'h55f == _T_2[11:0] ? image_1375 : _GEN_1374; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4448 = 12'h560 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7520 = 12'h560 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4448; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10592 = 12'h560 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7520; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13664 = 12'h560 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10592; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16736 = 12'h560 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13664; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19808 = 12'h560 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16736; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22880 = 12'h560 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19808; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25952 = 12'h560 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22880; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1376 = io_valid_in ? _GEN_25952 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1376 = 12'h560 == _T_2[11:0] ? image_1376 : _GEN_1375; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4449 = 12'h561 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7521 = 12'h561 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4449; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10593 = 12'h561 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7521; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13665 = 12'h561 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10593; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16737 = 12'h561 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13665; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19809 = 12'h561 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16737; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22881 = 12'h561 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19809; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25953 = 12'h561 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22881; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1377 = io_valid_in ? _GEN_25953 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1377 = 12'h561 == _T_2[11:0] ? image_1377 : _GEN_1376; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4450 = 12'h562 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7522 = 12'h562 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4450; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10594 = 12'h562 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7522; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13666 = 12'h562 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10594; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16738 = 12'h562 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13666; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19810 = 12'h562 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16738; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22882 = 12'h562 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19810; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25954 = 12'h562 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22882; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1378 = io_valid_in ? _GEN_25954 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1378 = 12'h562 == _T_2[11:0] ? image_1378 : _GEN_1377; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4451 = 12'h563 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7523 = 12'h563 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4451; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10595 = 12'h563 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7523; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13667 = 12'h563 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10595; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16739 = 12'h563 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13667; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19811 = 12'h563 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16739; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22883 = 12'h563 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19811; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25955 = 12'h563 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22883; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1379 = io_valid_in ? _GEN_25955 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1379 = 12'h563 == _T_2[11:0] ? image_1379 : _GEN_1378; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4452 = 12'h564 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7524 = 12'h564 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4452; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10596 = 12'h564 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7524; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13668 = 12'h564 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10596; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16740 = 12'h564 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13668; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19812 = 12'h564 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16740; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22884 = 12'h564 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19812; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25956 = 12'h564 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22884; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1380 = io_valid_in ? _GEN_25956 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1380 = 12'h564 == _T_2[11:0] ? image_1380 : _GEN_1379; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4453 = 12'h565 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7525 = 12'h565 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4453; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10597 = 12'h565 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7525; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13669 = 12'h565 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10597; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16741 = 12'h565 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13669; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19813 = 12'h565 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16741; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22885 = 12'h565 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19813; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25957 = 12'h565 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22885; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1381 = io_valid_in ? _GEN_25957 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1381 = 12'h565 == _T_2[11:0] ? image_1381 : _GEN_1380; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4454 = 12'h566 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7526 = 12'h566 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4454; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10598 = 12'h566 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7526; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13670 = 12'h566 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10598; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16742 = 12'h566 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13670; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19814 = 12'h566 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16742; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22886 = 12'h566 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19814; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25958 = 12'h566 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22886; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1382 = io_valid_in ? _GEN_25958 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1382 = 12'h566 == _T_2[11:0] ? image_1382 : _GEN_1381; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4455 = 12'h567 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7527 = 12'h567 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4455; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10599 = 12'h567 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7527; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13671 = 12'h567 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10599; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16743 = 12'h567 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13671; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19815 = 12'h567 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16743; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22887 = 12'h567 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19815; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25959 = 12'h567 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22887; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1383 = io_valid_in ? _GEN_25959 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1383 = 12'h567 == _T_2[11:0] ? image_1383 : _GEN_1382; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4456 = 12'h568 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7528 = 12'h568 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4456; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10600 = 12'h568 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7528; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13672 = 12'h568 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10600; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16744 = 12'h568 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13672; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19816 = 12'h568 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16744; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22888 = 12'h568 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19816; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25960 = 12'h568 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22888; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1384 = io_valid_in ? _GEN_25960 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1384 = 12'h568 == _T_2[11:0] ? image_1384 : _GEN_1383; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4457 = 12'h569 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7529 = 12'h569 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4457; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10601 = 12'h569 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7529; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13673 = 12'h569 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10601; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16745 = 12'h569 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13673; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19817 = 12'h569 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16745; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22889 = 12'h569 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19817; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25961 = 12'h569 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22889; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1385 = io_valid_in ? _GEN_25961 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1385 = 12'h569 == _T_2[11:0] ? image_1385 : _GEN_1384; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4458 = 12'h56a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7530 = 12'h56a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4458; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10602 = 12'h56a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7530; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13674 = 12'h56a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10602; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16746 = 12'h56a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13674; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19818 = 12'h56a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16746; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22890 = 12'h56a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19818; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25962 = 12'h56a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22890; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1386 = io_valid_in ? _GEN_25962 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1386 = 12'h56a == _T_2[11:0] ? image_1386 : _GEN_1385; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4459 = 12'h56b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7531 = 12'h56b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4459; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10603 = 12'h56b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7531; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13675 = 12'h56b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10603; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16747 = 12'h56b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13675; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19819 = 12'h56b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16747; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22891 = 12'h56b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19819; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25963 = 12'h56b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22891; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1387 = io_valid_in ? _GEN_25963 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1387 = 12'h56b == _T_2[11:0] ? image_1387 : _GEN_1386; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4460 = 12'h56c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7532 = 12'h56c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4460; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10604 = 12'h56c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7532; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13676 = 12'h56c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10604; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16748 = 12'h56c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13676; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19820 = 12'h56c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16748; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22892 = 12'h56c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19820; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25964 = 12'h56c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22892; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1388 = io_valid_in ? _GEN_25964 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1388 = 12'h56c == _T_2[11:0] ? image_1388 : _GEN_1387; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4461 = 12'h56d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7533 = 12'h56d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4461; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10605 = 12'h56d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7533; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13677 = 12'h56d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10605; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16749 = 12'h56d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13677; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19821 = 12'h56d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16749; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22893 = 12'h56d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19821; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25965 = 12'h56d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22893; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1389 = io_valid_in ? _GEN_25965 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1389 = 12'h56d == _T_2[11:0] ? image_1389 : _GEN_1388; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4462 = 12'h56e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7534 = 12'h56e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4462; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10606 = 12'h56e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7534; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13678 = 12'h56e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10606; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16750 = 12'h56e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13678; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19822 = 12'h56e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16750; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22894 = 12'h56e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19822; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25966 = 12'h56e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22894; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1390 = io_valid_in ? _GEN_25966 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1390 = 12'h56e == _T_2[11:0] ? image_1390 : _GEN_1389; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4463 = 12'h56f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7535 = 12'h56f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4463; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10607 = 12'h56f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7535; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13679 = 12'h56f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10607; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16751 = 12'h56f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13679; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19823 = 12'h56f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16751; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22895 = 12'h56f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19823; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25967 = 12'h56f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22895; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1391 = io_valid_in ? _GEN_25967 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1391 = 12'h56f == _T_2[11:0] ? image_1391 : _GEN_1390; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4464 = 12'h570 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7536 = 12'h570 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4464; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10608 = 12'h570 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7536; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13680 = 12'h570 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10608; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16752 = 12'h570 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13680; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19824 = 12'h570 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16752; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22896 = 12'h570 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19824; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25968 = 12'h570 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22896; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1392 = io_valid_in ? _GEN_25968 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1392 = 12'h570 == _T_2[11:0] ? image_1392 : _GEN_1391; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4465 = 12'h571 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7537 = 12'h571 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4465; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10609 = 12'h571 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7537; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13681 = 12'h571 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10609; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16753 = 12'h571 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13681; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19825 = 12'h571 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16753; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22897 = 12'h571 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19825; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25969 = 12'h571 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22897; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1393 = io_valid_in ? _GEN_25969 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1393 = 12'h571 == _T_2[11:0] ? image_1393 : _GEN_1392; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4466 = 12'h572 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7538 = 12'h572 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4466; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10610 = 12'h572 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7538; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13682 = 12'h572 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10610; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16754 = 12'h572 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13682; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19826 = 12'h572 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16754; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22898 = 12'h572 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19826; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25970 = 12'h572 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22898; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1394 = io_valid_in ? _GEN_25970 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1394 = 12'h572 == _T_2[11:0] ? image_1394 : _GEN_1393; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4467 = 12'h573 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7539 = 12'h573 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4467; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10611 = 12'h573 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7539; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13683 = 12'h573 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10611; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16755 = 12'h573 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13683; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19827 = 12'h573 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16755; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22899 = 12'h573 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19827; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25971 = 12'h573 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22899; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1395 = io_valid_in ? _GEN_25971 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1395 = 12'h573 == _T_2[11:0] ? image_1395 : _GEN_1394; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4468 = 12'h574 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7540 = 12'h574 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4468; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10612 = 12'h574 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7540; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13684 = 12'h574 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10612; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16756 = 12'h574 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13684; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19828 = 12'h574 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16756; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22900 = 12'h574 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19828; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25972 = 12'h574 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22900; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1396 = io_valid_in ? _GEN_25972 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1396 = 12'h574 == _T_2[11:0] ? image_1396 : _GEN_1395; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4469 = 12'h575 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7541 = 12'h575 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4469; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10613 = 12'h575 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7541; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13685 = 12'h575 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10613; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16757 = 12'h575 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13685; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19829 = 12'h575 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16757; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22901 = 12'h575 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19829; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25973 = 12'h575 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22901; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1397 = io_valid_in ? _GEN_25973 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1397 = 12'h575 == _T_2[11:0] ? image_1397 : _GEN_1396; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4470 = 12'h576 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7542 = 12'h576 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4470; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10614 = 12'h576 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7542; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13686 = 12'h576 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10614; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16758 = 12'h576 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13686; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19830 = 12'h576 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16758; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22902 = 12'h576 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19830; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25974 = 12'h576 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22902; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1398 = io_valid_in ? _GEN_25974 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1398 = 12'h576 == _T_2[11:0] ? image_1398 : _GEN_1397; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4471 = 12'h577 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7543 = 12'h577 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4471; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10615 = 12'h577 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7543; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13687 = 12'h577 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10615; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16759 = 12'h577 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13687; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19831 = 12'h577 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16759; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22903 = 12'h577 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19831; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25975 = 12'h577 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22903; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1399 = io_valid_in ? _GEN_25975 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1399 = 12'h577 == _T_2[11:0] ? image_1399 : _GEN_1398; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4472 = 12'h578 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7544 = 12'h578 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4472; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10616 = 12'h578 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7544; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13688 = 12'h578 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10616; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16760 = 12'h578 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13688; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19832 = 12'h578 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16760; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22904 = 12'h578 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19832; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25976 = 12'h578 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22904; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1400 = io_valid_in ? _GEN_25976 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1400 = 12'h578 == _T_2[11:0] ? image_1400 : _GEN_1399; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4473 = 12'h579 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7545 = 12'h579 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4473; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10617 = 12'h579 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7545; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13689 = 12'h579 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10617; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16761 = 12'h579 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13689; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19833 = 12'h579 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16761; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22905 = 12'h579 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19833; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25977 = 12'h579 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22905; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1401 = io_valid_in ? _GEN_25977 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1401 = 12'h579 == _T_2[11:0] ? image_1401 : _GEN_1400; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4474 = 12'h57a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7546 = 12'h57a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4474; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10618 = 12'h57a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7546; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13690 = 12'h57a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10618; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16762 = 12'h57a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13690; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19834 = 12'h57a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16762; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22906 = 12'h57a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19834; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25978 = 12'h57a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22906; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1402 = io_valid_in ? _GEN_25978 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1402 = 12'h57a == _T_2[11:0] ? image_1402 : _GEN_1401; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4475 = 12'h57b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7547 = 12'h57b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4475; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10619 = 12'h57b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7547; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13691 = 12'h57b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10619; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16763 = 12'h57b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13691; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19835 = 12'h57b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16763; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22907 = 12'h57b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19835; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25979 = 12'h57b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22907; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1403 = io_valid_in ? _GEN_25979 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1403 = 12'h57b == _T_2[11:0] ? image_1403 : _GEN_1402; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4476 = 12'h57c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7548 = 12'h57c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4476; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10620 = 12'h57c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7548; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13692 = 12'h57c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10620; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16764 = 12'h57c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13692; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19836 = 12'h57c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16764; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22908 = 12'h57c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19836; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25980 = 12'h57c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22908; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1404 = io_valid_in ? _GEN_25980 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1404 = 12'h57c == _T_2[11:0] ? image_1404 : _GEN_1403; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4477 = 12'h57d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7549 = 12'h57d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4477; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10621 = 12'h57d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7549; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13693 = 12'h57d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10621; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16765 = 12'h57d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13693; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19837 = 12'h57d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16765; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22909 = 12'h57d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19837; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25981 = 12'h57d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22909; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1405 = io_valid_in ? _GEN_25981 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1405 = 12'h57d == _T_2[11:0] ? image_1405 : _GEN_1404; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4478 = 12'h57e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7550 = 12'h57e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4478; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10622 = 12'h57e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7550; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13694 = 12'h57e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10622; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16766 = 12'h57e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13694; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19838 = 12'h57e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16766; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22910 = 12'h57e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19838; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25982 = 12'h57e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22910; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1406 = io_valid_in ? _GEN_25982 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1406 = 12'h57e == _T_2[11:0] ? image_1406 : _GEN_1405; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4479 = 12'h57f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7551 = 12'h57f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4479; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10623 = 12'h57f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7551; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13695 = 12'h57f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10623; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16767 = 12'h57f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13695; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19839 = 12'h57f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16767; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22911 = 12'h57f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19839; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25983 = 12'h57f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22911; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1407 = io_valid_in ? _GEN_25983 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1407 = 12'h57f == _T_2[11:0] ? image_1407 : _GEN_1406; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4480 = 12'h580 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7552 = 12'h580 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4480; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10624 = 12'h580 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7552; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13696 = 12'h580 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10624; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16768 = 12'h580 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13696; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19840 = 12'h580 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16768; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22912 = 12'h580 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19840; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25984 = 12'h580 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22912; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1408 = io_valid_in ? _GEN_25984 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1408 = 12'h580 == _T_2[11:0] ? image_1408 : _GEN_1407; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4481 = 12'h581 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7553 = 12'h581 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4481; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10625 = 12'h581 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7553; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13697 = 12'h581 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10625; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16769 = 12'h581 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13697; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19841 = 12'h581 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16769; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22913 = 12'h581 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19841; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25985 = 12'h581 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22913; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1409 = io_valid_in ? _GEN_25985 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1409 = 12'h581 == _T_2[11:0] ? image_1409 : _GEN_1408; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4482 = 12'h582 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7554 = 12'h582 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4482; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10626 = 12'h582 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7554; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13698 = 12'h582 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10626; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16770 = 12'h582 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13698; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19842 = 12'h582 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16770; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22914 = 12'h582 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19842; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25986 = 12'h582 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22914; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1410 = io_valid_in ? _GEN_25986 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1410 = 12'h582 == _T_2[11:0] ? image_1410 : _GEN_1409; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4483 = 12'h583 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7555 = 12'h583 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4483; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10627 = 12'h583 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7555; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13699 = 12'h583 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10627; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16771 = 12'h583 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13699; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19843 = 12'h583 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16771; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22915 = 12'h583 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19843; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25987 = 12'h583 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22915; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1411 = io_valid_in ? _GEN_25987 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1411 = 12'h583 == _T_2[11:0] ? image_1411 : _GEN_1410; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4484 = 12'h584 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7556 = 12'h584 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4484; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10628 = 12'h584 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7556; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13700 = 12'h584 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10628; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16772 = 12'h584 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13700; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19844 = 12'h584 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16772; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22916 = 12'h584 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19844; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25988 = 12'h584 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22916; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1412 = io_valid_in ? _GEN_25988 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1412 = 12'h584 == _T_2[11:0] ? image_1412 : _GEN_1411; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4485 = 12'h585 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7557 = 12'h585 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4485; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10629 = 12'h585 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7557; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13701 = 12'h585 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10629; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16773 = 12'h585 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13701; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19845 = 12'h585 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16773; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22917 = 12'h585 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19845; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25989 = 12'h585 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22917; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1413 = io_valid_in ? _GEN_25989 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1413 = 12'h585 == _T_2[11:0] ? image_1413 : _GEN_1412; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4486 = 12'h586 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7558 = 12'h586 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4486; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10630 = 12'h586 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7558; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13702 = 12'h586 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10630; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16774 = 12'h586 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13702; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19846 = 12'h586 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16774; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22918 = 12'h586 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19846; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25990 = 12'h586 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22918; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1414 = io_valid_in ? _GEN_25990 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1414 = 12'h586 == _T_2[11:0] ? image_1414 : _GEN_1413; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4487 = 12'h587 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7559 = 12'h587 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4487; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10631 = 12'h587 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7559; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13703 = 12'h587 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10631; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16775 = 12'h587 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13703; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19847 = 12'h587 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16775; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22919 = 12'h587 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19847; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25991 = 12'h587 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22919; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1415 = io_valid_in ? _GEN_25991 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1415 = 12'h587 == _T_2[11:0] ? image_1415 : _GEN_1414; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4488 = 12'h588 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7560 = 12'h588 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4488; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10632 = 12'h588 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7560; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13704 = 12'h588 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10632; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16776 = 12'h588 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13704; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19848 = 12'h588 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16776; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22920 = 12'h588 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19848; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25992 = 12'h588 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22920; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1416 = io_valid_in ? _GEN_25992 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1416 = 12'h588 == _T_2[11:0] ? image_1416 : _GEN_1415; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4489 = 12'h589 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7561 = 12'h589 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4489; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10633 = 12'h589 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7561; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13705 = 12'h589 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10633; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16777 = 12'h589 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13705; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19849 = 12'h589 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16777; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22921 = 12'h589 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19849; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25993 = 12'h589 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22921; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1417 = io_valid_in ? _GEN_25993 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1417 = 12'h589 == _T_2[11:0] ? image_1417 : _GEN_1416; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4490 = 12'h58a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7562 = 12'h58a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4490; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10634 = 12'h58a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7562; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13706 = 12'h58a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10634; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16778 = 12'h58a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13706; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19850 = 12'h58a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16778; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22922 = 12'h58a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19850; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25994 = 12'h58a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22922; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1418 = io_valid_in ? _GEN_25994 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1418 = 12'h58a == _T_2[11:0] ? image_1418 : _GEN_1417; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4491 = 12'h58b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7563 = 12'h58b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4491; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10635 = 12'h58b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7563; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13707 = 12'h58b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10635; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16779 = 12'h58b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13707; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19851 = 12'h58b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16779; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22923 = 12'h58b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19851; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25995 = 12'h58b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22923; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1419 = io_valid_in ? _GEN_25995 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1419 = 12'h58b == _T_2[11:0] ? image_1419 : _GEN_1418; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4492 = 12'h58c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7564 = 12'h58c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4492; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10636 = 12'h58c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7564; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13708 = 12'h58c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10636; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16780 = 12'h58c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13708; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19852 = 12'h58c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16780; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22924 = 12'h58c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19852; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25996 = 12'h58c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22924; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1420 = io_valid_in ? _GEN_25996 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1420 = 12'h58c == _T_2[11:0] ? image_1420 : _GEN_1419; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4493 = 12'h58d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7565 = 12'h58d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4493; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10637 = 12'h58d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7565; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13709 = 12'h58d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10637; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16781 = 12'h58d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13709; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19853 = 12'h58d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16781; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22925 = 12'h58d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19853; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25997 = 12'h58d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22925; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1421 = io_valid_in ? _GEN_25997 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1421 = 12'h58d == _T_2[11:0] ? image_1421 : _GEN_1420; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4494 = 12'h58e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7566 = 12'h58e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4494; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10638 = 12'h58e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7566; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13710 = 12'h58e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10638; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16782 = 12'h58e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13710; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19854 = 12'h58e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16782; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22926 = 12'h58e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19854; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25998 = 12'h58e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22926; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1422 = io_valid_in ? _GEN_25998 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1422 = 12'h58e == _T_2[11:0] ? image_1422 : _GEN_1421; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4495 = 12'h58f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7567 = 12'h58f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4495; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10639 = 12'h58f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7567; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13711 = 12'h58f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10639; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16783 = 12'h58f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13711; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19855 = 12'h58f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16783; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22927 = 12'h58f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19855; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_25999 = 12'h58f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22927; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1423 = io_valid_in ? _GEN_25999 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1423 = 12'h58f == _T_2[11:0] ? image_1423 : _GEN_1422; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4496 = 12'h590 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7568 = 12'h590 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4496; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10640 = 12'h590 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7568; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13712 = 12'h590 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10640; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16784 = 12'h590 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13712; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19856 = 12'h590 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16784; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22928 = 12'h590 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19856; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26000 = 12'h590 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22928; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1424 = io_valid_in ? _GEN_26000 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1424 = 12'h590 == _T_2[11:0] ? image_1424 : _GEN_1423; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4497 = 12'h591 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7569 = 12'h591 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4497; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10641 = 12'h591 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7569; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13713 = 12'h591 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10641; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16785 = 12'h591 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13713; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19857 = 12'h591 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16785; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22929 = 12'h591 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19857; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26001 = 12'h591 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22929; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1425 = io_valid_in ? _GEN_26001 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1425 = 12'h591 == _T_2[11:0] ? image_1425 : _GEN_1424; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4498 = 12'h592 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7570 = 12'h592 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4498; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10642 = 12'h592 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7570; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13714 = 12'h592 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10642; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16786 = 12'h592 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13714; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19858 = 12'h592 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16786; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22930 = 12'h592 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19858; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26002 = 12'h592 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22930; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1426 = io_valid_in ? _GEN_26002 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1426 = 12'h592 == _T_2[11:0] ? image_1426 : _GEN_1425; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4499 = 12'h593 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7571 = 12'h593 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4499; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10643 = 12'h593 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7571; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13715 = 12'h593 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10643; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16787 = 12'h593 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13715; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19859 = 12'h593 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16787; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22931 = 12'h593 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19859; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26003 = 12'h593 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22931; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1427 = io_valid_in ? _GEN_26003 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1427 = 12'h593 == _T_2[11:0] ? image_1427 : _GEN_1426; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4500 = 12'h594 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7572 = 12'h594 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4500; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10644 = 12'h594 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7572; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13716 = 12'h594 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10644; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16788 = 12'h594 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13716; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19860 = 12'h594 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16788; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22932 = 12'h594 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19860; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26004 = 12'h594 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22932; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1428 = io_valid_in ? _GEN_26004 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1428 = 12'h594 == _T_2[11:0] ? image_1428 : _GEN_1427; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4501 = 12'h595 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7573 = 12'h595 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4501; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10645 = 12'h595 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7573; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13717 = 12'h595 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10645; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16789 = 12'h595 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13717; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19861 = 12'h595 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16789; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22933 = 12'h595 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19861; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26005 = 12'h595 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22933; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1429 = io_valid_in ? _GEN_26005 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1429 = 12'h595 == _T_2[11:0] ? image_1429 : _GEN_1428; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4502 = 12'h596 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7574 = 12'h596 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4502; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10646 = 12'h596 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7574; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13718 = 12'h596 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10646; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16790 = 12'h596 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13718; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19862 = 12'h596 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16790; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22934 = 12'h596 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19862; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26006 = 12'h596 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22934; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1430 = io_valid_in ? _GEN_26006 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1430 = 12'h596 == _T_2[11:0] ? image_1430 : _GEN_1429; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4503 = 12'h597 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7575 = 12'h597 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4503; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10647 = 12'h597 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7575; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13719 = 12'h597 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10647; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16791 = 12'h597 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13719; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19863 = 12'h597 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16791; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22935 = 12'h597 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19863; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26007 = 12'h597 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22935; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1431 = io_valid_in ? _GEN_26007 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1431 = 12'h597 == _T_2[11:0] ? image_1431 : _GEN_1430; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4504 = 12'h598 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7576 = 12'h598 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4504; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10648 = 12'h598 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7576; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13720 = 12'h598 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10648; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16792 = 12'h598 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13720; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19864 = 12'h598 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16792; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22936 = 12'h598 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19864; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26008 = 12'h598 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22936; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1432 = io_valid_in ? _GEN_26008 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1432 = 12'h598 == _T_2[11:0] ? image_1432 : _GEN_1431; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4505 = 12'h599 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7577 = 12'h599 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4505; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10649 = 12'h599 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7577; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13721 = 12'h599 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10649; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16793 = 12'h599 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13721; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19865 = 12'h599 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16793; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22937 = 12'h599 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19865; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26009 = 12'h599 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22937; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1433 = io_valid_in ? _GEN_26009 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1433 = 12'h599 == _T_2[11:0] ? image_1433 : _GEN_1432; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4506 = 12'h59a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7578 = 12'h59a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4506; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10650 = 12'h59a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7578; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13722 = 12'h59a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10650; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16794 = 12'h59a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13722; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19866 = 12'h59a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16794; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22938 = 12'h59a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19866; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26010 = 12'h59a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22938; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1434 = io_valid_in ? _GEN_26010 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1434 = 12'h59a == _T_2[11:0] ? image_1434 : _GEN_1433; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4507 = 12'h59b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7579 = 12'h59b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4507; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10651 = 12'h59b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7579; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13723 = 12'h59b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10651; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16795 = 12'h59b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13723; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19867 = 12'h59b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16795; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22939 = 12'h59b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19867; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26011 = 12'h59b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22939; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1435 = io_valid_in ? _GEN_26011 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1435 = 12'h59b == _T_2[11:0] ? image_1435 : _GEN_1434; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4508 = 12'h59c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7580 = 12'h59c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4508; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10652 = 12'h59c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7580; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13724 = 12'h59c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10652; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16796 = 12'h59c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13724; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19868 = 12'h59c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16796; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22940 = 12'h59c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19868; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26012 = 12'h59c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22940; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1436 = io_valid_in ? _GEN_26012 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1436 = 12'h59c == _T_2[11:0] ? image_1436 : _GEN_1435; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4509 = 12'h59d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7581 = 12'h59d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4509; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10653 = 12'h59d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7581; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13725 = 12'h59d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10653; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16797 = 12'h59d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13725; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19869 = 12'h59d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16797; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22941 = 12'h59d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19869; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26013 = 12'h59d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22941; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1437 = io_valid_in ? _GEN_26013 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1437 = 12'h59d == _T_2[11:0] ? image_1437 : _GEN_1436; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4510 = 12'h59e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7582 = 12'h59e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4510; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10654 = 12'h59e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7582; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13726 = 12'h59e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10654; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16798 = 12'h59e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13726; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19870 = 12'h59e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16798; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22942 = 12'h59e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19870; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26014 = 12'h59e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22942; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1438 = io_valid_in ? _GEN_26014 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1438 = 12'h59e == _T_2[11:0] ? image_1438 : _GEN_1437; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4511 = 12'h59f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7583 = 12'h59f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4511; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10655 = 12'h59f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7583; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13727 = 12'h59f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10655; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16799 = 12'h59f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13727; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19871 = 12'h59f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16799; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22943 = 12'h59f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19871; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26015 = 12'h59f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22943; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1439 = io_valid_in ? _GEN_26015 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1439 = 12'h59f == _T_2[11:0] ? image_1439 : _GEN_1438; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4512 = 12'h5a0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7584 = 12'h5a0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4512; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10656 = 12'h5a0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7584; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13728 = 12'h5a0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10656; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16800 = 12'h5a0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13728; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19872 = 12'h5a0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16800; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22944 = 12'h5a0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19872; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26016 = 12'h5a0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22944; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1440 = io_valid_in ? _GEN_26016 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1440 = 12'h5a0 == _T_2[11:0] ? image_1440 : _GEN_1439; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4513 = 12'h5a1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7585 = 12'h5a1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4513; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10657 = 12'h5a1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7585; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13729 = 12'h5a1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10657; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16801 = 12'h5a1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13729; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19873 = 12'h5a1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16801; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22945 = 12'h5a1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19873; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26017 = 12'h5a1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22945; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1441 = io_valid_in ? _GEN_26017 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1441 = 12'h5a1 == _T_2[11:0] ? image_1441 : _GEN_1440; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4514 = 12'h5a2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7586 = 12'h5a2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4514; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10658 = 12'h5a2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7586; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13730 = 12'h5a2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10658; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16802 = 12'h5a2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13730; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19874 = 12'h5a2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16802; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22946 = 12'h5a2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19874; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26018 = 12'h5a2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22946; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1442 = io_valid_in ? _GEN_26018 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1442 = 12'h5a2 == _T_2[11:0] ? image_1442 : _GEN_1441; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4515 = 12'h5a3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7587 = 12'h5a3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4515; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10659 = 12'h5a3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7587; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13731 = 12'h5a3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10659; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16803 = 12'h5a3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13731; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19875 = 12'h5a3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16803; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22947 = 12'h5a3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19875; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26019 = 12'h5a3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22947; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1443 = io_valid_in ? _GEN_26019 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1443 = 12'h5a3 == _T_2[11:0] ? image_1443 : _GEN_1442; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4516 = 12'h5a4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7588 = 12'h5a4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4516; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10660 = 12'h5a4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7588; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13732 = 12'h5a4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10660; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16804 = 12'h5a4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13732; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19876 = 12'h5a4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16804; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22948 = 12'h5a4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19876; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26020 = 12'h5a4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22948; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1444 = io_valid_in ? _GEN_26020 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1444 = 12'h5a4 == _T_2[11:0] ? image_1444 : _GEN_1443; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4517 = 12'h5a5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7589 = 12'h5a5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4517; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10661 = 12'h5a5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7589; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13733 = 12'h5a5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10661; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16805 = 12'h5a5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13733; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19877 = 12'h5a5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16805; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22949 = 12'h5a5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19877; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26021 = 12'h5a5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22949; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1445 = io_valid_in ? _GEN_26021 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1445 = 12'h5a5 == _T_2[11:0] ? image_1445 : _GEN_1444; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4518 = 12'h5a6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7590 = 12'h5a6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4518; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10662 = 12'h5a6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7590; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13734 = 12'h5a6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10662; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16806 = 12'h5a6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13734; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19878 = 12'h5a6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16806; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22950 = 12'h5a6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19878; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26022 = 12'h5a6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22950; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1446 = io_valid_in ? _GEN_26022 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1446 = 12'h5a6 == _T_2[11:0] ? image_1446 : _GEN_1445; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4519 = 12'h5a7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7591 = 12'h5a7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4519; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10663 = 12'h5a7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7591; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13735 = 12'h5a7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10663; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16807 = 12'h5a7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13735; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19879 = 12'h5a7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16807; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22951 = 12'h5a7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19879; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26023 = 12'h5a7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22951; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1447 = io_valid_in ? _GEN_26023 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1447 = 12'h5a7 == _T_2[11:0] ? image_1447 : _GEN_1446; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4520 = 12'h5a8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7592 = 12'h5a8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4520; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10664 = 12'h5a8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7592; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13736 = 12'h5a8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10664; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16808 = 12'h5a8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13736; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19880 = 12'h5a8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16808; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22952 = 12'h5a8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19880; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26024 = 12'h5a8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22952; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1448 = io_valid_in ? _GEN_26024 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1448 = 12'h5a8 == _T_2[11:0] ? image_1448 : _GEN_1447; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4521 = 12'h5a9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7593 = 12'h5a9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4521; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10665 = 12'h5a9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7593; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13737 = 12'h5a9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10665; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16809 = 12'h5a9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13737; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19881 = 12'h5a9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16809; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22953 = 12'h5a9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19881; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26025 = 12'h5a9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22953; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1449 = io_valid_in ? _GEN_26025 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1449 = 12'h5a9 == _T_2[11:0] ? image_1449 : _GEN_1448; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4522 = 12'h5aa == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7594 = 12'h5aa == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4522; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10666 = 12'h5aa == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7594; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13738 = 12'h5aa == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10666; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16810 = 12'h5aa == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13738; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19882 = 12'h5aa == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16810; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22954 = 12'h5aa == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19882; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26026 = 12'h5aa == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22954; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1450 = io_valid_in ? _GEN_26026 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1450 = 12'h5aa == _T_2[11:0] ? image_1450 : _GEN_1449; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4523 = 12'h5ab == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7595 = 12'h5ab == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4523; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10667 = 12'h5ab == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7595; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13739 = 12'h5ab == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10667; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16811 = 12'h5ab == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13739; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19883 = 12'h5ab == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16811; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22955 = 12'h5ab == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19883; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26027 = 12'h5ab == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22955; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1451 = io_valid_in ? _GEN_26027 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1451 = 12'h5ab == _T_2[11:0] ? image_1451 : _GEN_1450; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4524 = 12'h5ac == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7596 = 12'h5ac == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4524; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10668 = 12'h5ac == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7596; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13740 = 12'h5ac == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10668; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16812 = 12'h5ac == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13740; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19884 = 12'h5ac == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16812; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22956 = 12'h5ac == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19884; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26028 = 12'h5ac == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22956; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1452 = io_valid_in ? _GEN_26028 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1452 = 12'h5ac == _T_2[11:0] ? image_1452 : _GEN_1451; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4525 = 12'h5ad == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7597 = 12'h5ad == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4525; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10669 = 12'h5ad == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7597; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13741 = 12'h5ad == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10669; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16813 = 12'h5ad == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13741; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19885 = 12'h5ad == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16813; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22957 = 12'h5ad == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19885; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26029 = 12'h5ad == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22957; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1453 = io_valid_in ? _GEN_26029 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1453 = 12'h5ad == _T_2[11:0] ? image_1453 : _GEN_1452; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4526 = 12'h5ae == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7598 = 12'h5ae == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4526; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10670 = 12'h5ae == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7598; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13742 = 12'h5ae == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10670; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16814 = 12'h5ae == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13742; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19886 = 12'h5ae == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16814; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22958 = 12'h5ae == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19886; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26030 = 12'h5ae == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22958; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1454 = io_valid_in ? _GEN_26030 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1454 = 12'h5ae == _T_2[11:0] ? image_1454 : _GEN_1453; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4527 = 12'h5af == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7599 = 12'h5af == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4527; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10671 = 12'h5af == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7599; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13743 = 12'h5af == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10671; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16815 = 12'h5af == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13743; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19887 = 12'h5af == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16815; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22959 = 12'h5af == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19887; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26031 = 12'h5af == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22959; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1455 = io_valid_in ? _GEN_26031 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1455 = 12'h5af == _T_2[11:0] ? image_1455 : _GEN_1454; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4528 = 12'h5b0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7600 = 12'h5b0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4528; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10672 = 12'h5b0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7600; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13744 = 12'h5b0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10672; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16816 = 12'h5b0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13744; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19888 = 12'h5b0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16816; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22960 = 12'h5b0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19888; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26032 = 12'h5b0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22960; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1456 = io_valid_in ? _GEN_26032 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1456 = 12'h5b0 == _T_2[11:0] ? image_1456 : _GEN_1455; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4529 = 12'h5b1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7601 = 12'h5b1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4529; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10673 = 12'h5b1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7601; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13745 = 12'h5b1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10673; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16817 = 12'h5b1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13745; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19889 = 12'h5b1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16817; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22961 = 12'h5b1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19889; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26033 = 12'h5b1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22961; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1457 = io_valid_in ? _GEN_26033 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1457 = 12'h5b1 == _T_2[11:0] ? image_1457 : _GEN_1456; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4530 = 12'h5b2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7602 = 12'h5b2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4530; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10674 = 12'h5b2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7602; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13746 = 12'h5b2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10674; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16818 = 12'h5b2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13746; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19890 = 12'h5b2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16818; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22962 = 12'h5b2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19890; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26034 = 12'h5b2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22962; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1458 = io_valid_in ? _GEN_26034 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1458 = 12'h5b2 == _T_2[11:0] ? image_1458 : _GEN_1457; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4531 = 12'h5b3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7603 = 12'h5b3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4531; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10675 = 12'h5b3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7603; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13747 = 12'h5b3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10675; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16819 = 12'h5b3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13747; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19891 = 12'h5b3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16819; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22963 = 12'h5b3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19891; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26035 = 12'h5b3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22963; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1459 = io_valid_in ? _GEN_26035 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1459 = 12'h5b3 == _T_2[11:0] ? image_1459 : _GEN_1458; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4532 = 12'h5b4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7604 = 12'h5b4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4532; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10676 = 12'h5b4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7604; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13748 = 12'h5b4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10676; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16820 = 12'h5b4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13748; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19892 = 12'h5b4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16820; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22964 = 12'h5b4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19892; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26036 = 12'h5b4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22964; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1460 = io_valid_in ? _GEN_26036 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1460 = 12'h5b4 == _T_2[11:0] ? image_1460 : _GEN_1459; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4533 = 12'h5b5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7605 = 12'h5b5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4533; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10677 = 12'h5b5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7605; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13749 = 12'h5b5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10677; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16821 = 12'h5b5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13749; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19893 = 12'h5b5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16821; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22965 = 12'h5b5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19893; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26037 = 12'h5b5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22965; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1461 = io_valid_in ? _GEN_26037 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1461 = 12'h5b5 == _T_2[11:0] ? image_1461 : _GEN_1460; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4534 = 12'h5b6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7606 = 12'h5b6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4534; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10678 = 12'h5b6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7606; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13750 = 12'h5b6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10678; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16822 = 12'h5b6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13750; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19894 = 12'h5b6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16822; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22966 = 12'h5b6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19894; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26038 = 12'h5b6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22966; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1462 = io_valid_in ? _GEN_26038 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1462 = 12'h5b6 == _T_2[11:0] ? image_1462 : _GEN_1461; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4535 = 12'h5b7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7607 = 12'h5b7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4535; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10679 = 12'h5b7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7607; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13751 = 12'h5b7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10679; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16823 = 12'h5b7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13751; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19895 = 12'h5b7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16823; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22967 = 12'h5b7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19895; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26039 = 12'h5b7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22967; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1463 = io_valid_in ? _GEN_26039 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1463 = 12'h5b7 == _T_2[11:0] ? image_1463 : _GEN_1462; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4536 = 12'h5b8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7608 = 12'h5b8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4536; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10680 = 12'h5b8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7608; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13752 = 12'h5b8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10680; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16824 = 12'h5b8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13752; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19896 = 12'h5b8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16824; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22968 = 12'h5b8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19896; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26040 = 12'h5b8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22968; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1464 = io_valid_in ? _GEN_26040 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1464 = 12'h5b8 == _T_2[11:0] ? image_1464 : _GEN_1463; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4537 = 12'h5b9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7609 = 12'h5b9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4537; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10681 = 12'h5b9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7609; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13753 = 12'h5b9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10681; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16825 = 12'h5b9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13753; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19897 = 12'h5b9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16825; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22969 = 12'h5b9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19897; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26041 = 12'h5b9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22969; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1465 = io_valid_in ? _GEN_26041 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1465 = 12'h5b9 == _T_2[11:0] ? image_1465 : _GEN_1464; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4538 = 12'h5ba == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7610 = 12'h5ba == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4538; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10682 = 12'h5ba == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7610; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13754 = 12'h5ba == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10682; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16826 = 12'h5ba == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13754; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19898 = 12'h5ba == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16826; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22970 = 12'h5ba == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19898; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26042 = 12'h5ba == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22970; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1466 = io_valid_in ? _GEN_26042 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1466 = 12'h5ba == _T_2[11:0] ? image_1466 : _GEN_1465; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4539 = 12'h5bb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7611 = 12'h5bb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4539; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10683 = 12'h5bb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7611; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13755 = 12'h5bb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10683; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16827 = 12'h5bb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13755; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19899 = 12'h5bb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16827; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22971 = 12'h5bb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19899; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26043 = 12'h5bb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22971; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1467 = io_valid_in ? _GEN_26043 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1467 = 12'h5bb == _T_2[11:0] ? image_1467 : _GEN_1466; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4540 = 12'h5bc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7612 = 12'h5bc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4540; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10684 = 12'h5bc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7612; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13756 = 12'h5bc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10684; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16828 = 12'h5bc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13756; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19900 = 12'h5bc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16828; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22972 = 12'h5bc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19900; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26044 = 12'h5bc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22972; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1468 = io_valid_in ? _GEN_26044 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1468 = 12'h5bc == _T_2[11:0] ? image_1468 : _GEN_1467; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4541 = 12'h5bd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7613 = 12'h5bd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4541; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10685 = 12'h5bd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7613; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13757 = 12'h5bd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10685; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16829 = 12'h5bd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13757; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19901 = 12'h5bd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16829; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22973 = 12'h5bd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19901; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26045 = 12'h5bd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22973; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1469 = io_valid_in ? _GEN_26045 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1469 = 12'h5bd == _T_2[11:0] ? image_1469 : _GEN_1468; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4542 = 12'h5be == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7614 = 12'h5be == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4542; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10686 = 12'h5be == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7614; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13758 = 12'h5be == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10686; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16830 = 12'h5be == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13758; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19902 = 12'h5be == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16830; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22974 = 12'h5be == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19902; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26046 = 12'h5be == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22974; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1470 = io_valid_in ? _GEN_26046 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1470 = 12'h5be == _T_2[11:0] ? image_1470 : _GEN_1469; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4543 = 12'h5bf == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7615 = 12'h5bf == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4543; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10687 = 12'h5bf == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7615; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13759 = 12'h5bf == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10687; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16831 = 12'h5bf == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13759; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19903 = 12'h5bf == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16831; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22975 = 12'h5bf == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19903; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26047 = 12'h5bf == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22975; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1471 = io_valid_in ? _GEN_26047 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1471 = 12'h5bf == _T_2[11:0] ? image_1471 : _GEN_1470; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4544 = 12'h5c0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7616 = 12'h5c0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4544; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10688 = 12'h5c0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7616; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13760 = 12'h5c0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10688; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16832 = 12'h5c0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13760; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19904 = 12'h5c0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16832; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22976 = 12'h5c0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19904; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26048 = 12'h5c0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22976; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1472 = io_valid_in ? _GEN_26048 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1472 = 12'h5c0 == _T_2[11:0] ? image_1472 : _GEN_1471; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4545 = 12'h5c1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7617 = 12'h5c1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4545; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10689 = 12'h5c1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7617; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13761 = 12'h5c1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10689; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16833 = 12'h5c1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13761; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19905 = 12'h5c1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16833; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22977 = 12'h5c1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19905; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26049 = 12'h5c1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22977; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1473 = io_valid_in ? _GEN_26049 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1473 = 12'h5c1 == _T_2[11:0] ? image_1473 : _GEN_1472; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4546 = 12'h5c2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7618 = 12'h5c2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4546; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10690 = 12'h5c2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7618; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13762 = 12'h5c2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10690; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16834 = 12'h5c2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13762; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19906 = 12'h5c2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16834; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22978 = 12'h5c2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19906; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26050 = 12'h5c2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22978; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1474 = io_valid_in ? _GEN_26050 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1474 = 12'h5c2 == _T_2[11:0] ? image_1474 : _GEN_1473; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4547 = 12'h5c3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7619 = 12'h5c3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4547; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10691 = 12'h5c3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7619; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13763 = 12'h5c3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10691; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16835 = 12'h5c3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13763; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19907 = 12'h5c3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16835; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22979 = 12'h5c3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19907; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26051 = 12'h5c3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22979; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1475 = io_valid_in ? _GEN_26051 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1475 = 12'h5c3 == _T_2[11:0] ? image_1475 : _GEN_1474; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4548 = 12'h5c4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7620 = 12'h5c4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4548; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10692 = 12'h5c4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7620; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13764 = 12'h5c4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10692; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16836 = 12'h5c4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13764; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19908 = 12'h5c4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16836; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22980 = 12'h5c4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19908; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26052 = 12'h5c4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22980; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1476 = io_valid_in ? _GEN_26052 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1476 = 12'h5c4 == _T_2[11:0] ? image_1476 : _GEN_1475; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4549 = 12'h5c5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7621 = 12'h5c5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4549; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10693 = 12'h5c5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7621; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13765 = 12'h5c5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10693; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16837 = 12'h5c5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13765; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19909 = 12'h5c5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16837; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22981 = 12'h5c5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19909; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26053 = 12'h5c5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22981; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1477 = io_valid_in ? _GEN_26053 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1477 = 12'h5c5 == _T_2[11:0] ? image_1477 : _GEN_1476; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4550 = 12'h5c6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7622 = 12'h5c6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4550; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10694 = 12'h5c6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7622; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13766 = 12'h5c6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10694; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16838 = 12'h5c6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13766; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19910 = 12'h5c6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16838; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22982 = 12'h5c6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19910; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26054 = 12'h5c6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22982; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1478 = io_valid_in ? _GEN_26054 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1478 = 12'h5c6 == _T_2[11:0] ? image_1478 : _GEN_1477; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4551 = 12'h5c7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7623 = 12'h5c7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4551; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10695 = 12'h5c7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7623; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13767 = 12'h5c7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10695; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16839 = 12'h5c7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13767; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19911 = 12'h5c7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16839; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22983 = 12'h5c7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19911; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26055 = 12'h5c7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22983; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1479 = io_valid_in ? _GEN_26055 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1479 = 12'h5c7 == _T_2[11:0] ? image_1479 : _GEN_1478; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4552 = 12'h5c8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7624 = 12'h5c8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4552; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10696 = 12'h5c8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7624; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13768 = 12'h5c8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10696; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16840 = 12'h5c8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13768; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19912 = 12'h5c8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16840; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22984 = 12'h5c8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19912; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26056 = 12'h5c8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22984; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1480 = io_valid_in ? _GEN_26056 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1480 = 12'h5c8 == _T_2[11:0] ? image_1480 : _GEN_1479; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4553 = 12'h5c9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7625 = 12'h5c9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4553; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10697 = 12'h5c9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7625; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13769 = 12'h5c9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10697; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16841 = 12'h5c9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13769; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19913 = 12'h5c9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16841; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22985 = 12'h5c9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19913; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26057 = 12'h5c9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22985; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1481 = io_valid_in ? _GEN_26057 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1481 = 12'h5c9 == _T_2[11:0] ? image_1481 : _GEN_1480; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4554 = 12'h5ca == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7626 = 12'h5ca == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4554; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10698 = 12'h5ca == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7626; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13770 = 12'h5ca == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10698; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16842 = 12'h5ca == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13770; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19914 = 12'h5ca == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16842; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22986 = 12'h5ca == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19914; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26058 = 12'h5ca == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22986; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1482 = io_valid_in ? _GEN_26058 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1482 = 12'h5ca == _T_2[11:0] ? image_1482 : _GEN_1481; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4555 = 12'h5cb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7627 = 12'h5cb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4555; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10699 = 12'h5cb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7627; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13771 = 12'h5cb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10699; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16843 = 12'h5cb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13771; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19915 = 12'h5cb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16843; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22987 = 12'h5cb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19915; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26059 = 12'h5cb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22987; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1483 = io_valid_in ? _GEN_26059 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1483 = 12'h5cb == _T_2[11:0] ? image_1483 : _GEN_1482; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4556 = 12'h5cc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7628 = 12'h5cc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4556; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10700 = 12'h5cc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7628; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13772 = 12'h5cc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10700; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16844 = 12'h5cc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13772; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19916 = 12'h5cc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16844; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22988 = 12'h5cc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19916; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26060 = 12'h5cc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22988; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1484 = io_valid_in ? _GEN_26060 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1484 = 12'h5cc == _T_2[11:0] ? image_1484 : _GEN_1483; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4557 = 12'h5cd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7629 = 12'h5cd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4557; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10701 = 12'h5cd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7629; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13773 = 12'h5cd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10701; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16845 = 12'h5cd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13773; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19917 = 12'h5cd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16845; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22989 = 12'h5cd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19917; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26061 = 12'h5cd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22989; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1485 = io_valid_in ? _GEN_26061 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1485 = 12'h5cd == _T_2[11:0] ? image_1485 : _GEN_1484; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4558 = 12'h5ce == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7630 = 12'h5ce == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4558; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10702 = 12'h5ce == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7630; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13774 = 12'h5ce == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10702; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16846 = 12'h5ce == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13774; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19918 = 12'h5ce == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16846; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22990 = 12'h5ce == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19918; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26062 = 12'h5ce == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22990; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1486 = io_valid_in ? _GEN_26062 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1486 = 12'h5ce == _T_2[11:0] ? image_1486 : _GEN_1485; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4559 = 12'h5cf == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7631 = 12'h5cf == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4559; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10703 = 12'h5cf == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7631; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13775 = 12'h5cf == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10703; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16847 = 12'h5cf == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13775; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19919 = 12'h5cf == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16847; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22991 = 12'h5cf == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19919; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26063 = 12'h5cf == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22991; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1487 = io_valid_in ? _GEN_26063 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1487 = 12'h5cf == _T_2[11:0] ? image_1487 : _GEN_1486; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4560 = 12'h5d0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7632 = 12'h5d0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4560; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10704 = 12'h5d0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7632; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13776 = 12'h5d0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10704; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16848 = 12'h5d0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13776; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19920 = 12'h5d0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16848; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22992 = 12'h5d0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19920; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26064 = 12'h5d0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22992; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1488 = io_valid_in ? _GEN_26064 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1488 = 12'h5d0 == _T_2[11:0] ? image_1488 : _GEN_1487; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4561 = 12'h5d1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7633 = 12'h5d1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4561; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10705 = 12'h5d1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7633; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13777 = 12'h5d1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10705; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16849 = 12'h5d1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13777; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19921 = 12'h5d1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16849; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22993 = 12'h5d1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19921; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26065 = 12'h5d1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22993; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1489 = io_valid_in ? _GEN_26065 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1489 = 12'h5d1 == _T_2[11:0] ? image_1489 : _GEN_1488; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4562 = 12'h5d2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7634 = 12'h5d2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4562; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10706 = 12'h5d2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7634; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13778 = 12'h5d2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10706; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16850 = 12'h5d2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13778; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19922 = 12'h5d2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16850; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22994 = 12'h5d2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19922; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26066 = 12'h5d2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22994; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1490 = io_valid_in ? _GEN_26066 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1490 = 12'h5d2 == _T_2[11:0] ? image_1490 : _GEN_1489; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4563 = 12'h5d3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7635 = 12'h5d3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4563; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10707 = 12'h5d3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7635; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13779 = 12'h5d3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10707; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16851 = 12'h5d3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13779; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19923 = 12'h5d3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16851; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22995 = 12'h5d3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19923; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26067 = 12'h5d3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22995; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1491 = io_valid_in ? _GEN_26067 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1491 = 12'h5d3 == _T_2[11:0] ? image_1491 : _GEN_1490; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4564 = 12'h5d4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7636 = 12'h5d4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4564; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10708 = 12'h5d4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7636; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13780 = 12'h5d4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10708; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16852 = 12'h5d4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13780; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19924 = 12'h5d4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16852; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22996 = 12'h5d4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19924; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26068 = 12'h5d4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22996; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1492 = io_valid_in ? _GEN_26068 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1492 = 12'h5d4 == _T_2[11:0] ? image_1492 : _GEN_1491; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4565 = 12'h5d5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7637 = 12'h5d5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4565; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10709 = 12'h5d5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7637; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13781 = 12'h5d5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10709; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16853 = 12'h5d5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13781; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19925 = 12'h5d5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16853; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22997 = 12'h5d5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19925; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26069 = 12'h5d5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22997; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1493 = io_valid_in ? _GEN_26069 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1493 = 12'h5d5 == _T_2[11:0] ? image_1493 : _GEN_1492; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4566 = 12'h5d6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7638 = 12'h5d6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4566; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10710 = 12'h5d6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7638; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13782 = 12'h5d6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10710; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16854 = 12'h5d6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13782; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19926 = 12'h5d6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16854; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22998 = 12'h5d6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19926; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26070 = 12'h5d6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22998; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1494 = io_valid_in ? _GEN_26070 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1494 = 12'h5d6 == _T_2[11:0] ? image_1494 : _GEN_1493; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4567 = 12'h5d7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7639 = 12'h5d7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4567; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10711 = 12'h5d7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7639; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13783 = 12'h5d7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10711; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16855 = 12'h5d7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13783; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19927 = 12'h5d7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16855; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_22999 = 12'h5d7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19927; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26071 = 12'h5d7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_22999; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1495 = io_valid_in ? _GEN_26071 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1495 = 12'h5d7 == _T_2[11:0] ? image_1495 : _GEN_1494; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4568 = 12'h5d8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7640 = 12'h5d8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4568; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10712 = 12'h5d8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7640; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13784 = 12'h5d8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10712; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16856 = 12'h5d8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13784; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19928 = 12'h5d8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16856; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23000 = 12'h5d8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19928; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26072 = 12'h5d8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23000; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1496 = io_valid_in ? _GEN_26072 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1496 = 12'h5d8 == _T_2[11:0] ? image_1496 : _GEN_1495; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4569 = 12'h5d9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7641 = 12'h5d9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4569; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10713 = 12'h5d9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7641; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13785 = 12'h5d9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10713; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16857 = 12'h5d9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13785; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19929 = 12'h5d9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16857; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23001 = 12'h5d9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19929; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26073 = 12'h5d9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23001; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1497 = io_valid_in ? _GEN_26073 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1497 = 12'h5d9 == _T_2[11:0] ? image_1497 : _GEN_1496; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4570 = 12'h5da == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7642 = 12'h5da == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4570; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10714 = 12'h5da == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7642; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13786 = 12'h5da == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10714; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16858 = 12'h5da == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13786; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19930 = 12'h5da == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16858; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23002 = 12'h5da == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19930; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26074 = 12'h5da == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23002; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1498 = io_valid_in ? _GEN_26074 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1498 = 12'h5da == _T_2[11:0] ? image_1498 : _GEN_1497; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4571 = 12'h5db == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7643 = 12'h5db == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4571; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10715 = 12'h5db == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7643; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13787 = 12'h5db == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10715; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16859 = 12'h5db == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13787; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19931 = 12'h5db == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16859; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23003 = 12'h5db == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19931; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26075 = 12'h5db == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23003; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1499 = io_valid_in ? _GEN_26075 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1499 = 12'h5db == _T_2[11:0] ? image_1499 : _GEN_1498; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4572 = 12'h5dc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7644 = 12'h5dc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4572; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10716 = 12'h5dc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7644; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13788 = 12'h5dc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10716; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16860 = 12'h5dc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13788; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19932 = 12'h5dc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16860; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23004 = 12'h5dc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19932; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26076 = 12'h5dc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23004; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1500 = io_valid_in ? _GEN_26076 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1500 = 12'h5dc == _T_2[11:0] ? image_1500 : _GEN_1499; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4573 = 12'h5dd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7645 = 12'h5dd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4573; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10717 = 12'h5dd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7645; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13789 = 12'h5dd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10717; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16861 = 12'h5dd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13789; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19933 = 12'h5dd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16861; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23005 = 12'h5dd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19933; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26077 = 12'h5dd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23005; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1501 = io_valid_in ? _GEN_26077 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1501 = 12'h5dd == _T_2[11:0] ? image_1501 : _GEN_1500; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4574 = 12'h5de == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7646 = 12'h5de == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4574; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10718 = 12'h5de == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7646; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13790 = 12'h5de == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10718; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16862 = 12'h5de == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13790; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19934 = 12'h5de == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16862; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23006 = 12'h5de == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19934; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26078 = 12'h5de == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23006; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1502 = io_valid_in ? _GEN_26078 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1502 = 12'h5de == _T_2[11:0] ? image_1502 : _GEN_1501; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4575 = 12'h5df == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7647 = 12'h5df == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4575; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10719 = 12'h5df == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7647; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13791 = 12'h5df == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10719; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16863 = 12'h5df == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13791; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19935 = 12'h5df == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16863; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23007 = 12'h5df == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19935; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26079 = 12'h5df == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23007; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1503 = io_valid_in ? _GEN_26079 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1503 = 12'h5df == _T_2[11:0] ? image_1503 : _GEN_1502; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4576 = 12'h5e0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7648 = 12'h5e0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4576; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10720 = 12'h5e0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7648; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13792 = 12'h5e0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10720; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16864 = 12'h5e0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13792; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19936 = 12'h5e0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16864; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23008 = 12'h5e0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19936; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26080 = 12'h5e0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23008; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1504 = io_valid_in ? _GEN_26080 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1504 = 12'h5e0 == _T_2[11:0] ? image_1504 : _GEN_1503; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4577 = 12'h5e1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7649 = 12'h5e1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4577; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10721 = 12'h5e1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7649; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13793 = 12'h5e1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10721; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16865 = 12'h5e1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13793; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19937 = 12'h5e1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16865; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23009 = 12'h5e1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19937; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26081 = 12'h5e1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23009; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1505 = io_valid_in ? _GEN_26081 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1505 = 12'h5e1 == _T_2[11:0] ? image_1505 : _GEN_1504; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4578 = 12'h5e2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7650 = 12'h5e2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4578; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10722 = 12'h5e2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7650; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13794 = 12'h5e2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10722; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16866 = 12'h5e2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13794; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19938 = 12'h5e2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16866; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23010 = 12'h5e2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19938; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26082 = 12'h5e2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23010; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1506 = io_valid_in ? _GEN_26082 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1506 = 12'h5e2 == _T_2[11:0] ? image_1506 : _GEN_1505; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4579 = 12'h5e3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7651 = 12'h5e3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4579; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10723 = 12'h5e3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7651; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13795 = 12'h5e3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10723; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16867 = 12'h5e3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13795; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19939 = 12'h5e3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16867; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23011 = 12'h5e3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19939; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26083 = 12'h5e3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23011; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1507 = io_valid_in ? _GEN_26083 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1507 = 12'h5e3 == _T_2[11:0] ? image_1507 : _GEN_1506; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4580 = 12'h5e4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7652 = 12'h5e4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4580; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10724 = 12'h5e4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7652; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13796 = 12'h5e4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10724; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16868 = 12'h5e4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13796; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19940 = 12'h5e4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16868; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23012 = 12'h5e4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19940; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26084 = 12'h5e4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23012; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1508 = io_valid_in ? _GEN_26084 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1508 = 12'h5e4 == _T_2[11:0] ? image_1508 : _GEN_1507; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4581 = 12'h5e5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7653 = 12'h5e5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4581; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10725 = 12'h5e5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7653; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13797 = 12'h5e5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10725; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16869 = 12'h5e5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13797; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19941 = 12'h5e5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16869; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23013 = 12'h5e5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19941; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26085 = 12'h5e5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23013; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1509 = io_valid_in ? _GEN_26085 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1509 = 12'h5e5 == _T_2[11:0] ? image_1509 : _GEN_1508; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4582 = 12'h5e6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7654 = 12'h5e6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4582; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10726 = 12'h5e6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7654; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13798 = 12'h5e6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10726; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16870 = 12'h5e6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13798; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19942 = 12'h5e6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16870; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23014 = 12'h5e6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19942; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26086 = 12'h5e6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23014; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1510 = io_valid_in ? _GEN_26086 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1510 = 12'h5e6 == _T_2[11:0] ? image_1510 : _GEN_1509; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4583 = 12'h5e7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7655 = 12'h5e7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4583; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10727 = 12'h5e7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7655; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13799 = 12'h5e7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10727; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16871 = 12'h5e7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13799; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19943 = 12'h5e7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16871; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23015 = 12'h5e7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19943; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26087 = 12'h5e7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23015; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1511 = io_valid_in ? _GEN_26087 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1511 = 12'h5e7 == _T_2[11:0] ? image_1511 : _GEN_1510; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4584 = 12'h5e8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7656 = 12'h5e8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4584; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10728 = 12'h5e8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7656; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13800 = 12'h5e8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10728; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16872 = 12'h5e8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13800; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19944 = 12'h5e8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16872; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23016 = 12'h5e8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19944; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26088 = 12'h5e8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23016; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1512 = io_valid_in ? _GEN_26088 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1512 = 12'h5e8 == _T_2[11:0] ? image_1512 : _GEN_1511; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4585 = 12'h5e9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7657 = 12'h5e9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4585; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10729 = 12'h5e9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7657; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13801 = 12'h5e9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10729; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16873 = 12'h5e9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13801; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19945 = 12'h5e9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16873; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23017 = 12'h5e9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19945; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26089 = 12'h5e9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23017; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1513 = io_valid_in ? _GEN_26089 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1513 = 12'h5e9 == _T_2[11:0] ? image_1513 : _GEN_1512; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4586 = 12'h5ea == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7658 = 12'h5ea == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4586; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10730 = 12'h5ea == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7658; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13802 = 12'h5ea == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10730; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16874 = 12'h5ea == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13802; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19946 = 12'h5ea == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16874; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23018 = 12'h5ea == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19946; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26090 = 12'h5ea == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23018; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1514 = io_valid_in ? _GEN_26090 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1514 = 12'h5ea == _T_2[11:0] ? image_1514 : _GEN_1513; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4587 = 12'h5eb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7659 = 12'h5eb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4587; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10731 = 12'h5eb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7659; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13803 = 12'h5eb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10731; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16875 = 12'h5eb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13803; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19947 = 12'h5eb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16875; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23019 = 12'h5eb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19947; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26091 = 12'h5eb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23019; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1515 = io_valid_in ? _GEN_26091 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1515 = 12'h5eb == _T_2[11:0] ? image_1515 : _GEN_1514; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4588 = 12'h5ec == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7660 = 12'h5ec == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4588; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10732 = 12'h5ec == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7660; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13804 = 12'h5ec == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10732; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16876 = 12'h5ec == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13804; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19948 = 12'h5ec == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16876; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23020 = 12'h5ec == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19948; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26092 = 12'h5ec == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23020; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1516 = io_valid_in ? _GEN_26092 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1516 = 12'h5ec == _T_2[11:0] ? image_1516 : _GEN_1515; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4589 = 12'h5ed == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7661 = 12'h5ed == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4589; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10733 = 12'h5ed == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7661; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13805 = 12'h5ed == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10733; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16877 = 12'h5ed == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13805; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19949 = 12'h5ed == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16877; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23021 = 12'h5ed == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19949; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26093 = 12'h5ed == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23021; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1517 = io_valid_in ? _GEN_26093 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1517 = 12'h5ed == _T_2[11:0] ? image_1517 : _GEN_1516; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4590 = 12'h5ee == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7662 = 12'h5ee == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4590; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10734 = 12'h5ee == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7662; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13806 = 12'h5ee == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10734; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16878 = 12'h5ee == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13806; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19950 = 12'h5ee == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16878; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23022 = 12'h5ee == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19950; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26094 = 12'h5ee == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23022; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1518 = io_valid_in ? _GEN_26094 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1518 = 12'h5ee == _T_2[11:0] ? image_1518 : _GEN_1517; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4591 = 12'h5ef == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7663 = 12'h5ef == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4591; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10735 = 12'h5ef == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7663; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13807 = 12'h5ef == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10735; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16879 = 12'h5ef == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13807; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19951 = 12'h5ef == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16879; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23023 = 12'h5ef == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19951; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26095 = 12'h5ef == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23023; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1519 = io_valid_in ? _GEN_26095 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1519 = 12'h5ef == _T_2[11:0] ? image_1519 : _GEN_1518; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4592 = 12'h5f0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7664 = 12'h5f0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4592; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10736 = 12'h5f0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7664; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13808 = 12'h5f0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10736; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16880 = 12'h5f0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13808; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19952 = 12'h5f0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16880; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23024 = 12'h5f0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19952; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26096 = 12'h5f0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23024; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1520 = io_valid_in ? _GEN_26096 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1520 = 12'h5f0 == _T_2[11:0] ? image_1520 : _GEN_1519; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4593 = 12'h5f1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7665 = 12'h5f1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4593; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10737 = 12'h5f1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7665; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13809 = 12'h5f1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10737; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16881 = 12'h5f1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13809; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19953 = 12'h5f1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16881; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23025 = 12'h5f1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19953; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26097 = 12'h5f1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23025; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1521 = io_valid_in ? _GEN_26097 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1521 = 12'h5f1 == _T_2[11:0] ? image_1521 : _GEN_1520; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4594 = 12'h5f2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7666 = 12'h5f2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4594; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10738 = 12'h5f2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7666; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13810 = 12'h5f2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10738; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16882 = 12'h5f2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13810; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19954 = 12'h5f2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16882; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23026 = 12'h5f2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19954; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26098 = 12'h5f2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23026; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1522 = io_valid_in ? _GEN_26098 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1522 = 12'h5f2 == _T_2[11:0] ? image_1522 : _GEN_1521; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4595 = 12'h5f3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7667 = 12'h5f3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4595; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10739 = 12'h5f3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7667; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13811 = 12'h5f3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10739; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16883 = 12'h5f3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13811; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19955 = 12'h5f3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16883; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23027 = 12'h5f3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19955; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26099 = 12'h5f3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23027; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1523 = io_valid_in ? _GEN_26099 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1523 = 12'h5f3 == _T_2[11:0] ? image_1523 : _GEN_1522; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4596 = 12'h5f4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7668 = 12'h5f4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4596; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10740 = 12'h5f4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7668; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13812 = 12'h5f4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10740; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16884 = 12'h5f4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13812; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19956 = 12'h5f4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16884; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23028 = 12'h5f4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19956; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26100 = 12'h5f4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23028; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1524 = io_valid_in ? _GEN_26100 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1524 = 12'h5f4 == _T_2[11:0] ? image_1524 : _GEN_1523; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4597 = 12'h5f5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7669 = 12'h5f5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4597; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10741 = 12'h5f5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7669; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13813 = 12'h5f5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10741; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16885 = 12'h5f5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13813; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19957 = 12'h5f5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16885; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23029 = 12'h5f5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19957; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26101 = 12'h5f5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23029; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1525 = io_valid_in ? _GEN_26101 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1525 = 12'h5f5 == _T_2[11:0] ? image_1525 : _GEN_1524; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4598 = 12'h5f6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7670 = 12'h5f6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4598; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10742 = 12'h5f6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7670; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13814 = 12'h5f6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10742; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16886 = 12'h5f6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13814; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19958 = 12'h5f6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16886; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23030 = 12'h5f6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19958; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26102 = 12'h5f6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23030; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1526 = io_valid_in ? _GEN_26102 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1526 = 12'h5f6 == _T_2[11:0] ? image_1526 : _GEN_1525; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4599 = 12'h5f7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7671 = 12'h5f7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4599; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10743 = 12'h5f7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7671; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13815 = 12'h5f7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10743; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16887 = 12'h5f7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13815; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19959 = 12'h5f7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16887; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23031 = 12'h5f7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19959; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26103 = 12'h5f7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23031; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1527 = io_valid_in ? _GEN_26103 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1527 = 12'h5f7 == _T_2[11:0] ? image_1527 : _GEN_1526; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4600 = 12'h5f8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7672 = 12'h5f8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4600; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10744 = 12'h5f8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7672; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13816 = 12'h5f8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10744; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16888 = 12'h5f8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13816; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19960 = 12'h5f8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16888; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23032 = 12'h5f8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19960; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26104 = 12'h5f8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23032; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1528 = io_valid_in ? _GEN_26104 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1528 = 12'h5f8 == _T_2[11:0] ? image_1528 : _GEN_1527; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4601 = 12'h5f9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7673 = 12'h5f9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4601; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10745 = 12'h5f9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7673; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13817 = 12'h5f9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10745; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16889 = 12'h5f9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13817; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19961 = 12'h5f9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16889; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23033 = 12'h5f9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19961; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26105 = 12'h5f9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23033; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1529 = io_valid_in ? _GEN_26105 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1529 = 12'h5f9 == _T_2[11:0] ? image_1529 : _GEN_1528; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4602 = 12'h5fa == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7674 = 12'h5fa == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4602; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10746 = 12'h5fa == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7674; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13818 = 12'h5fa == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10746; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16890 = 12'h5fa == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13818; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19962 = 12'h5fa == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16890; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23034 = 12'h5fa == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19962; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26106 = 12'h5fa == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23034; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1530 = io_valid_in ? _GEN_26106 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1530 = 12'h5fa == _T_2[11:0] ? image_1530 : _GEN_1529; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4603 = 12'h5fb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7675 = 12'h5fb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4603; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10747 = 12'h5fb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7675; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13819 = 12'h5fb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10747; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16891 = 12'h5fb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13819; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19963 = 12'h5fb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16891; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23035 = 12'h5fb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19963; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26107 = 12'h5fb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23035; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1531 = io_valid_in ? _GEN_26107 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1531 = 12'h5fb == _T_2[11:0] ? image_1531 : _GEN_1530; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4604 = 12'h5fc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7676 = 12'h5fc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4604; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10748 = 12'h5fc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7676; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13820 = 12'h5fc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10748; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16892 = 12'h5fc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13820; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19964 = 12'h5fc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16892; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23036 = 12'h5fc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19964; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26108 = 12'h5fc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23036; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1532 = io_valid_in ? _GEN_26108 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1532 = 12'h5fc == _T_2[11:0] ? image_1532 : _GEN_1531; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4605 = 12'h5fd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7677 = 12'h5fd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4605; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10749 = 12'h5fd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7677; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13821 = 12'h5fd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10749; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16893 = 12'h5fd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13821; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19965 = 12'h5fd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16893; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23037 = 12'h5fd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19965; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26109 = 12'h5fd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23037; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1533 = io_valid_in ? _GEN_26109 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1533 = 12'h5fd == _T_2[11:0] ? image_1533 : _GEN_1532; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4606 = 12'h5fe == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7678 = 12'h5fe == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4606; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10750 = 12'h5fe == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7678; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13822 = 12'h5fe == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10750; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16894 = 12'h5fe == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13822; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19966 = 12'h5fe == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16894; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23038 = 12'h5fe == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19966; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26110 = 12'h5fe == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23038; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1534 = io_valid_in ? _GEN_26110 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1534 = 12'h5fe == _T_2[11:0] ? image_1534 : _GEN_1533; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4607 = 12'h5ff == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7679 = 12'h5ff == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4607; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10751 = 12'h5ff == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7679; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13823 = 12'h5ff == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10751; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16895 = 12'h5ff == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13823; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19967 = 12'h5ff == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16895; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23039 = 12'h5ff == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19967; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26111 = 12'h5ff == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23039; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1535 = io_valid_in ? _GEN_26111 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1535 = 12'h5ff == _T_2[11:0] ? image_1535 : _GEN_1534; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4608 = 12'h600 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7680 = 12'h600 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4608; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10752 = 12'h600 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7680; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13824 = 12'h600 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10752; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16896 = 12'h600 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13824; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19968 = 12'h600 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16896; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23040 = 12'h600 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19968; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26112 = 12'h600 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23040; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1536 = io_valid_in ? _GEN_26112 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1536 = 12'h600 == _T_2[11:0] ? image_1536 : _GEN_1535; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4609 = 12'h601 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7681 = 12'h601 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4609; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10753 = 12'h601 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7681; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13825 = 12'h601 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10753; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16897 = 12'h601 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13825; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19969 = 12'h601 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16897; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23041 = 12'h601 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19969; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26113 = 12'h601 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23041; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1537 = io_valid_in ? _GEN_26113 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1537 = 12'h601 == _T_2[11:0] ? image_1537 : _GEN_1536; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4610 = 12'h602 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7682 = 12'h602 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4610; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10754 = 12'h602 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7682; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13826 = 12'h602 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10754; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16898 = 12'h602 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13826; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19970 = 12'h602 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16898; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23042 = 12'h602 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19970; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26114 = 12'h602 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23042; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1538 = io_valid_in ? _GEN_26114 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1538 = 12'h602 == _T_2[11:0] ? image_1538 : _GEN_1537; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4611 = 12'h603 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7683 = 12'h603 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4611; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10755 = 12'h603 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7683; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13827 = 12'h603 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10755; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16899 = 12'h603 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13827; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19971 = 12'h603 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16899; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23043 = 12'h603 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19971; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26115 = 12'h603 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23043; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1539 = io_valid_in ? _GEN_26115 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1539 = 12'h603 == _T_2[11:0] ? image_1539 : _GEN_1538; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4612 = 12'h604 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7684 = 12'h604 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4612; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10756 = 12'h604 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7684; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13828 = 12'h604 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10756; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16900 = 12'h604 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13828; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19972 = 12'h604 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16900; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23044 = 12'h604 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19972; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26116 = 12'h604 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23044; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1540 = io_valid_in ? _GEN_26116 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1540 = 12'h604 == _T_2[11:0] ? image_1540 : _GEN_1539; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4613 = 12'h605 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7685 = 12'h605 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4613; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10757 = 12'h605 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7685; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13829 = 12'h605 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10757; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16901 = 12'h605 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13829; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19973 = 12'h605 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16901; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23045 = 12'h605 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19973; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26117 = 12'h605 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23045; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1541 = io_valid_in ? _GEN_26117 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1541 = 12'h605 == _T_2[11:0] ? image_1541 : _GEN_1540; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4614 = 12'h606 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7686 = 12'h606 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4614; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10758 = 12'h606 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7686; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13830 = 12'h606 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10758; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16902 = 12'h606 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13830; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19974 = 12'h606 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16902; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23046 = 12'h606 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19974; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26118 = 12'h606 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23046; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1542 = io_valid_in ? _GEN_26118 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1542 = 12'h606 == _T_2[11:0] ? image_1542 : _GEN_1541; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4615 = 12'h607 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7687 = 12'h607 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4615; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10759 = 12'h607 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7687; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13831 = 12'h607 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10759; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16903 = 12'h607 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13831; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19975 = 12'h607 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16903; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23047 = 12'h607 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19975; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26119 = 12'h607 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23047; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1543 = io_valid_in ? _GEN_26119 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1543 = 12'h607 == _T_2[11:0] ? image_1543 : _GEN_1542; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4616 = 12'h608 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7688 = 12'h608 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4616; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10760 = 12'h608 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7688; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13832 = 12'h608 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10760; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16904 = 12'h608 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13832; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19976 = 12'h608 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16904; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23048 = 12'h608 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19976; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26120 = 12'h608 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23048; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1544 = io_valid_in ? _GEN_26120 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1544 = 12'h608 == _T_2[11:0] ? image_1544 : _GEN_1543; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4617 = 12'h609 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7689 = 12'h609 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4617; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10761 = 12'h609 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7689; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13833 = 12'h609 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10761; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16905 = 12'h609 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13833; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19977 = 12'h609 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16905; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23049 = 12'h609 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19977; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26121 = 12'h609 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23049; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1545 = io_valid_in ? _GEN_26121 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1545 = 12'h609 == _T_2[11:0] ? image_1545 : _GEN_1544; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4618 = 12'h60a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7690 = 12'h60a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4618; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10762 = 12'h60a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7690; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13834 = 12'h60a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10762; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16906 = 12'h60a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13834; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19978 = 12'h60a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16906; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23050 = 12'h60a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19978; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26122 = 12'h60a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23050; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1546 = io_valid_in ? _GEN_26122 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1546 = 12'h60a == _T_2[11:0] ? image_1546 : _GEN_1545; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4619 = 12'h60b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7691 = 12'h60b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4619; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10763 = 12'h60b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7691; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13835 = 12'h60b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10763; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16907 = 12'h60b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13835; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19979 = 12'h60b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16907; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23051 = 12'h60b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19979; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26123 = 12'h60b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23051; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1547 = io_valid_in ? _GEN_26123 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1547 = 12'h60b == _T_2[11:0] ? image_1547 : _GEN_1546; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4620 = 12'h60c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7692 = 12'h60c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4620; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10764 = 12'h60c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7692; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13836 = 12'h60c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10764; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16908 = 12'h60c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13836; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19980 = 12'h60c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16908; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23052 = 12'h60c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19980; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26124 = 12'h60c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23052; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1548 = io_valid_in ? _GEN_26124 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1548 = 12'h60c == _T_2[11:0] ? image_1548 : _GEN_1547; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4621 = 12'h60d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7693 = 12'h60d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4621; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10765 = 12'h60d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7693; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13837 = 12'h60d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10765; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16909 = 12'h60d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13837; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19981 = 12'h60d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16909; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23053 = 12'h60d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19981; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26125 = 12'h60d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23053; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1549 = io_valid_in ? _GEN_26125 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1549 = 12'h60d == _T_2[11:0] ? image_1549 : _GEN_1548; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4622 = 12'h60e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7694 = 12'h60e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4622; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10766 = 12'h60e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7694; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13838 = 12'h60e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10766; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16910 = 12'h60e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13838; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19982 = 12'h60e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16910; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23054 = 12'h60e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19982; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26126 = 12'h60e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23054; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1550 = io_valid_in ? _GEN_26126 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1550 = 12'h60e == _T_2[11:0] ? image_1550 : _GEN_1549; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4623 = 12'h60f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7695 = 12'h60f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4623; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10767 = 12'h60f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7695; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13839 = 12'h60f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10767; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16911 = 12'h60f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13839; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19983 = 12'h60f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16911; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23055 = 12'h60f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19983; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26127 = 12'h60f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23055; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1551 = io_valid_in ? _GEN_26127 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1551 = 12'h60f == _T_2[11:0] ? image_1551 : _GEN_1550; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4624 = 12'h610 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7696 = 12'h610 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4624; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10768 = 12'h610 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7696; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13840 = 12'h610 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10768; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16912 = 12'h610 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13840; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19984 = 12'h610 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16912; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23056 = 12'h610 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19984; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26128 = 12'h610 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23056; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1552 = io_valid_in ? _GEN_26128 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1552 = 12'h610 == _T_2[11:0] ? image_1552 : _GEN_1551; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4625 = 12'h611 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7697 = 12'h611 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4625; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10769 = 12'h611 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7697; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13841 = 12'h611 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10769; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16913 = 12'h611 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13841; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19985 = 12'h611 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16913; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23057 = 12'h611 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19985; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26129 = 12'h611 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23057; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1553 = io_valid_in ? _GEN_26129 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1553 = 12'h611 == _T_2[11:0] ? image_1553 : _GEN_1552; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4626 = 12'h612 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7698 = 12'h612 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4626; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10770 = 12'h612 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7698; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13842 = 12'h612 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10770; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16914 = 12'h612 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13842; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19986 = 12'h612 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16914; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23058 = 12'h612 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19986; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26130 = 12'h612 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23058; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1554 = io_valid_in ? _GEN_26130 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1554 = 12'h612 == _T_2[11:0] ? image_1554 : _GEN_1553; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4627 = 12'h613 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7699 = 12'h613 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4627; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10771 = 12'h613 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7699; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13843 = 12'h613 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10771; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16915 = 12'h613 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13843; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19987 = 12'h613 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16915; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23059 = 12'h613 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19987; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26131 = 12'h613 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23059; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1555 = io_valid_in ? _GEN_26131 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1555 = 12'h613 == _T_2[11:0] ? image_1555 : _GEN_1554; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4628 = 12'h614 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7700 = 12'h614 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4628; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10772 = 12'h614 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7700; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13844 = 12'h614 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10772; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16916 = 12'h614 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13844; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19988 = 12'h614 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16916; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23060 = 12'h614 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19988; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26132 = 12'h614 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23060; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1556 = io_valid_in ? _GEN_26132 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1556 = 12'h614 == _T_2[11:0] ? image_1556 : _GEN_1555; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4629 = 12'h615 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7701 = 12'h615 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4629; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10773 = 12'h615 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7701; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13845 = 12'h615 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10773; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16917 = 12'h615 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13845; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19989 = 12'h615 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16917; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23061 = 12'h615 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19989; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26133 = 12'h615 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23061; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1557 = io_valid_in ? _GEN_26133 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1557 = 12'h615 == _T_2[11:0] ? image_1557 : _GEN_1556; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4630 = 12'h616 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7702 = 12'h616 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4630; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10774 = 12'h616 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7702; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13846 = 12'h616 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10774; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16918 = 12'h616 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13846; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19990 = 12'h616 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16918; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23062 = 12'h616 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19990; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26134 = 12'h616 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23062; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1558 = io_valid_in ? _GEN_26134 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1558 = 12'h616 == _T_2[11:0] ? image_1558 : _GEN_1557; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4631 = 12'h617 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7703 = 12'h617 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4631; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10775 = 12'h617 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7703; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13847 = 12'h617 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10775; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16919 = 12'h617 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13847; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19991 = 12'h617 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16919; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23063 = 12'h617 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19991; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26135 = 12'h617 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23063; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1559 = io_valid_in ? _GEN_26135 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1559 = 12'h617 == _T_2[11:0] ? image_1559 : _GEN_1558; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4632 = 12'h618 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7704 = 12'h618 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4632; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10776 = 12'h618 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7704; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13848 = 12'h618 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10776; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16920 = 12'h618 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13848; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19992 = 12'h618 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16920; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23064 = 12'h618 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19992; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26136 = 12'h618 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23064; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1560 = io_valid_in ? _GEN_26136 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1560 = 12'h618 == _T_2[11:0] ? image_1560 : _GEN_1559; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4633 = 12'h619 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7705 = 12'h619 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4633; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10777 = 12'h619 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7705; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13849 = 12'h619 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10777; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16921 = 12'h619 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13849; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19993 = 12'h619 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16921; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23065 = 12'h619 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19993; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26137 = 12'h619 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23065; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1561 = io_valid_in ? _GEN_26137 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1561 = 12'h619 == _T_2[11:0] ? image_1561 : _GEN_1560; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4634 = 12'h61a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7706 = 12'h61a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4634; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10778 = 12'h61a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7706; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13850 = 12'h61a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10778; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16922 = 12'h61a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13850; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19994 = 12'h61a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16922; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23066 = 12'h61a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19994; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26138 = 12'h61a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23066; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1562 = io_valid_in ? _GEN_26138 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1562 = 12'h61a == _T_2[11:0] ? image_1562 : _GEN_1561; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4635 = 12'h61b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7707 = 12'h61b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4635; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10779 = 12'h61b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7707; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13851 = 12'h61b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10779; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16923 = 12'h61b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13851; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19995 = 12'h61b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16923; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23067 = 12'h61b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19995; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26139 = 12'h61b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23067; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1563 = io_valid_in ? _GEN_26139 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1563 = 12'h61b == _T_2[11:0] ? image_1563 : _GEN_1562; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4636 = 12'h61c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7708 = 12'h61c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4636; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10780 = 12'h61c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7708; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13852 = 12'h61c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10780; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16924 = 12'h61c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13852; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19996 = 12'h61c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16924; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23068 = 12'h61c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19996; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26140 = 12'h61c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23068; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1564 = io_valid_in ? _GEN_26140 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1564 = 12'h61c == _T_2[11:0] ? image_1564 : _GEN_1563; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4637 = 12'h61d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7709 = 12'h61d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4637; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10781 = 12'h61d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7709; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13853 = 12'h61d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10781; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16925 = 12'h61d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13853; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19997 = 12'h61d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16925; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23069 = 12'h61d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19997; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26141 = 12'h61d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23069; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1565 = io_valid_in ? _GEN_26141 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1565 = 12'h61d == _T_2[11:0] ? image_1565 : _GEN_1564; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4638 = 12'h61e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7710 = 12'h61e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4638; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10782 = 12'h61e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7710; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13854 = 12'h61e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10782; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16926 = 12'h61e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13854; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19998 = 12'h61e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16926; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23070 = 12'h61e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19998; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26142 = 12'h61e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23070; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1566 = io_valid_in ? _GEN_26142 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1566 = 12'h61e == _T_2[11:0] ? image_1566 : _GEN_1565; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4639 = 12'h61f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7711 = 12'h61f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4639; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10783 = 12'h61f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7711; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13855 = 12'h61f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10783; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16927 = 12'h61f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13855; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_19999 = 12'h61f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16927; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23071 = 12'h61f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_19999; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26143 = 12'h61f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23071; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1567 = io_valid_in ? _GEN_26143 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1567 = 12'h61f == _T_2[11:0] ? image_1567 : _GEN_1566; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4640 = 12'h620 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7712 = 12'h620 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4640; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10784 = 12'h620 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7712; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13856 = 12'h620 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10784; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16928 = 12'h620 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13856; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20000 = 12'h620 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16928; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23072 = 12'h620 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20000; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26144 = 12'h620 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23072; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1568 = io_valid_in ? _GEN_26144 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1568 = 12'h620 == _T_2[11:0] ? image_1568 : _GEN_1567; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4641 = 12'h621 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7713 = 12'h621 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4641; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10785 = 12'h621 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7713; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13857 = 12'h621 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10785; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16929 = 12'h621 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13857; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20001 = 12'h621 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16929; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23073 = 12'h621 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20001; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26145 = 12'h621 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23073; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1569 = io_valid_in ? _GEN_26145 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1569 = 12'h621 == _T_2[11:0] ? image_1569 : _GEN_1568; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4642 = 12'h622 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7714 = 12'h622 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4642; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10786 = 12'h622 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7714; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13858 = 12'h622 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10786; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16930 = 12'h622 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13858; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20002 = 12'h622 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16930; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23074 = 12'h622 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20002; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26146 = 12'h622 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23074; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1570 = io_valid_in ? _GEN_26146 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1570 = 12'h622 == _T_2[11:0] ? image_1570 : _GEN_1569; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4643 = 12'h623 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7715 = 12'h623 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4643; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10787 = 12'h623 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7715; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13859 = 12'h623 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10787; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16931 = 12'h623 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13859; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20003 = 12'h623 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16931; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23075 = 12'h623 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20003; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26147 = 12'h623 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23075; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1571 = io_valid_in ? _GEN_26147 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1571 = 12'h623 == _T_2[11:0] ? image_1571 : _GEN_1570; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4644 = 12'h624 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7716 = 12'h624 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4644; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10788 = 12'h624 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7716; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13860 = 12'h624 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10788; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16932 = 12'h624 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13860; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20004 = 12'h624 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16932; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23076 = 12'h624 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20004; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26148 = 12'h624 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23076; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1572 = io_valid_in ? _GEN_26148 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1572 = 12'h624 == _T_2[11:0] ? image_1572 : _GEN_1571; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4645 = 12'h625 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7717 = 12'h625 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4645; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10789 = 12'h625 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7717; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13861 = 12'h625 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10789; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16933 = 12'h625 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13861; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20005 = 12'h625 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16933; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23077 = 12'h625 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20005; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26149 = 12'h625 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23077; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1573 = io_valid_in ? _GEN_26149 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1573 = 12'h625 == _T_2[11:0] ? image_1573 : _GEN_1572; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4646 = 12'h626 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7718 = 12'h626 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4646; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10790 = 12'h626 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7718; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13862 = 12'h626 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10790; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16934 = 12'h626 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13862; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20006 = 12'h626 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16934; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23078 = 12'h626 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20006; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26150 = 12'h626 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23078; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1574 = io_valid_in ? _GEN_26150 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1574 = 12'h626 == _T_2[11:0] ? image_1574 : _GEN_1573; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4647 = 12'h627 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7719 = 12'h627 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4647; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10791 = 12'h627 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7719; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13863 = 12'h627 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10791; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16935 = 12'h627 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13863; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20007 = 12'h627 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16935; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23079 = 12'h627 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20007; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26151 = 12'h627 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23079; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1575 = io_valid_in ? _GEN_26151 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1575 = 12'h627 == _T_2[11:0] ? image_1575 : _GEN_1574; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4648 = 12'h628 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7720 = 12'h628 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4648; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10792 = 12'h628 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7720; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13864 = 12'h628 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10792; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16936 = 12'h628 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13864; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20008 = 12'h628 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16936; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23080 = 12'h628 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20008; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26152 = 12'h628 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23080; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1576 = io_valid_in ? _GEN_26152 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1576 = 12'h628 == _T_2[11:0] ? image_1576 : _GEN_1575; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4649 = 12'h629 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7721 = 12'h629 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4649; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10793 = 12'h629 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7721; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13865 = 12'h629 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10793; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16937 = 12'h629 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13865; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20009 = 12'h629 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16937; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23081 = 12'h629 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20009; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26153 = 12'h629 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23081; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1577 = io_valid_in ? _GEN_26153 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1577 = 12'h629 == _T_2[11:0] ? image_1577 : _GEN_1576; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4650 = 12'h62a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7722 = 12'h62a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4650; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10794 = 12'h62a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7722; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13866 = 12'h62a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10794; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16938 = 12'h62a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13866; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20010 = 12'h62a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16938; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23082 = 12'h62a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20010; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26154 = 12'h62a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23082; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1578 = io_valid_in ? _GEN_26154 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1578 = 12'h62a == _T_2[11:0] ? image_1578 : _GEN_1577; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4651 = 12'h62b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7723 = 12'h62b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4651; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10795 = 12'h62b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7723; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13867 = 12'h62b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10795; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16939 = 12'h62b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13867; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20011 = 12'h62b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16939; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23083 = 12'h62b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20011; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26155 = 12'h62b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23083; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1579 = io_valid_in ? _GEN_26155 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1579 = 12'h62b == _T_2[11:0] ? image_1579 : _GEN_1578; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4652 = 12'h62c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7724 = 12'h62c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4652; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10796 = 12'h62c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7724; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13868 = 12'h62c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10796; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16940 = 12'h62c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13868; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20012 = 12'h62c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16940; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23084 = 12'h62c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20012; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26156 = 12'h62c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23084; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1580 = io_valid_in ? _GEN_26156 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1580 = 12'h62c == _T_2[11:0] ? image_1580 : _GEN_1579; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4653 = 12'h62d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7725 = 12'h62d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4653; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10797 = 12'h62d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7725; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13869 = 12'h62d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10797; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16941 = 12'h62d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13869; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20013 = 12'h62d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16941; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23085 = 12'h62d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20013; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26157 = 12'h62d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23085; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1581 = io_valid_in ? _GEN_26157 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1581 = 12'h62d == _T_2[11:0] ? image_1581 : _GEN_1580; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4654 = 12'h62e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7726 = 12'h62e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4654; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10798 = 12'h62e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7726; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13870 = 12'h62e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10798; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16942 = 12'h62e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13870; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20014 = 12'h62e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16942; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23086 = 12'h62e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20014; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26158 = 12'h62e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23086; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1582 = io_valid_in ? _GEN_26158 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1582 = 12'h62e == _T_2[11:0] ? image_1582 : _GEN_1581; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4655 = 12'h62f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7727 = 12'h62f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4655; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10799 = 12'h62f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7727; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13871 = 12'h62f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10799; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16943 = 12'h62f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13871; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20015 = 12'h62f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16943; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23087 = 12'h62f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20015; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26159 = 12'h62f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23087; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1583 = io_valid_in ? _GEN_26159 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1583 = 12'h62f == _T_2[11:0] ? image_1583 : _GEN_1582; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4656 = 12'h630 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7728 = 12'h630 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4656; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10800 = 12'h630 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7728; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13872 = 12'h630 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10800; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16944 = 12'h630 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13872; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20016 = 12'h630 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16944; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23088 = 12'h630 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20016; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26160 = 12'h630 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23088; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1584 = io_valid_in ? _GEN_26160 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1584 = 12'h630 == _T_2[11:0] ? image_1584 : _GEN_1583; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4657 = 12'h631 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7729 = 12'h631 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4657; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10801 = 12'h631 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7729; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13873 = 12'h631 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10801; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16945 = 12'h631 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13873; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20017 = 12'h631 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16945; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23089 = 12'h631 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20017; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26161 = 12'h631 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23089; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1585 = io_valid_in ? _GEN_26161 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1585 = 12'h631 == _T_2[11:0] ? image_1585 : _GEN_1584; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4658 = 12'h632 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7730 = 12'h632 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4658; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10802 = 12'h632 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7730; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13874 = 12'h632 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10802; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16946 = 12'h632 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13874; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20018 = 12'h632 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16946; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23090 = 12'h632 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20018; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26162 = 12'h632 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23090; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1586 = io_valid_in ? _GEN_26162 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1586 = 12'h632 == _T_2[11:0] ? image_1586 : _GEN_1585; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4659 = 12'h633 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7731 = 12'h633 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4659; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10803 = 12'h633 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7731; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13875 = 12'h633 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10803; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16947 = 12'h633 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13875; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20019 = 12'h633 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16947; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23091 = 12'h633 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20019; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26163 = 12'h633 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23091; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1587 = io_valid_in ? _GEN_26163 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1587 = 12'h633 == _T_2[11:0] ? image_1587 : _GEN_1586; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4660 = 12'h634 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7732 = 12'h634 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4660; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10804 = 12'h634 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7732; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13876 = 12'h634 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10804; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16948 = 12'h634 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13876; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20020 = 12'h634 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16948; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23092 = 12'h634 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20020; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26164 = 12'h634 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23092; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1588 = io_valid_in ? _GEN_26164 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1588 = 12'h634 == _T_2[11:0] ? image_1588 : _GEN_1587; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4661 = 12'h635 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7733 = 12'h635 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4661; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10805 = 12'h635 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7733; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13877 = 12'h635 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10805; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16949 = 12'h635 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13877; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20021 = 12'h635 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16949; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23093 = 12'h635 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20021; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26165 = 12'h635 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23093; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1589 = io_valid_in ? _GEN_26165 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1589 = 12'h635 == _T_2[11:0] ? image_1589 : _GEN_1588; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4662 = 12'h636 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7734 = 12'h636 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4662; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10806 = 12'h636 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7734; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13878 = 12'h636 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10806; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16950 = 12'h636 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13878; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20022 = 12'h636 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16950; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23094 = 12'h636 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20022; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26166 = 12'h636 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23094; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1590 = io_valid_in ? _GEN_26166 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1590 = 12'h636 == _T_2[11:0] ? image_1590 : _GEN_1589; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4663 = 12'h637 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7735 = 12'h637 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4663; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10807 = 12'h637 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7735; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13879 = 12'h637 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10807; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16951 = 12'h637 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13879; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20023 = 12'h637 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16951; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23095 = 12'h637 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20023; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26167 = 12'h637 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23095; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1591 = io_valid_in ? _GEN_26167 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1591 = 12'h637 == _T_2[11:0] ? image_1591 : _GEN_1590; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4664 = 12'h638 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7736 = 12'h638 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4664; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10808 = 12'h638 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7736; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13880 = 12'h638 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10808; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16952 = 12'h638 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13880; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20024 = 12'h638 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16952; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23096 = 12'h638 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20024; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26168 = 12'h638 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23096; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1592 = io_valid_in ? _GEN_26168 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1592 = 12'h638 == _T_2[11:0] ? image_1592 : _GEN_1591; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4665 = 12'h639 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7737 = 12'h639 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4665; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10809 = 12'h639 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7737; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13881 = 12'h639 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10809; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16953 = 12'h639 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13881; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20025 = 12'h639 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16953; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23097 = 12'h639 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20025; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26169 = 12'h639 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23097; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1593 = io_valid_in ? _GEN_26169 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1593 = 12'h639 == _T_2[11:0] ? image_1593 : _GEN_1592; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4666 = 12'h63a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7738 = 12'h63a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4666; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10810 = 12'h63a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7738; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13882 = 12'h63a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10810; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16954 = 12'h63a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13882; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20026 = 12'h63a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16954; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23098 = 12'h63a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20026; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26170 = 12'h63a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23098; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1594 = io_valid_in ? _GEN_26170 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1594 = 12'h63a == _T_2[11:0] ? image_1594 : _GEN_1593; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4667 = 12'h63b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7739 = 12'h63b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4667; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10811 = 12'h63b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7739; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13883 = 12'h63b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10811; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16955 = 12'h63b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13883; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20027 = 12'h63b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16955; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23099 = 12'h63b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20027; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26171 = 12'h63b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23099; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1595 = io_valid_in ? _GEN_26171 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1595 = 12'h63b == _T_2[11:0] ? image_1595 : _GEN_1594; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4668 = 12'h63c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7740 = 12'h63c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4668; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10812 = 12'h63c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7740; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13884 = 12'h63c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10812; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16956 = 12'h63c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13884; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20028 = 12'h63c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16956; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23100 = 12'h63c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20028; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26172 = 12'h63c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23100; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1596 = io_valid_in ? _GEN_26172 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1596 = 12'h63c == _T_2[11:0] ? image_1596 : _GEN_1595; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4669 = 12'h63d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7741 = 12'h63d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4669; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10813 = 12'h63d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7741; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13885 = 12'h63d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10813; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16957 = 12'h63d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13885; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20029 = 12'h63d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16957; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23101 = 12'h63d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20029; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26173 = 12'h63d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23101; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1597 = io_valid_in ? _GEN_26173 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1597 = 12'h63d == _T_2[11:0] ? image_1597 : _GEN_1596; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4670 = 12'h63e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7742 = 12'h63e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4670; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10814 = 12'h63e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7742; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13886 = 12'h63e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10814; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16958 = 12'h63e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13886; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20030 = 12'h63e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16958; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23102 = 12'h63e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20030; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26174 = 12'h63e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23102; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1598 = io_valid_in ? _GEN_26174 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1598 = 12'h63e == _T_2[11:0] ? image_1598 : _GEN_1597; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4671 = 12'h63f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7743 = 12'h63f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4671; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10815 = 12'h63f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7743; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13887 = 12'h63f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10815; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16959 = 12'h63f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13887; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20031 = 12'h63f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16959; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23103 = 12'h63f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20031; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26175 = 12'h63f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23103; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1599 = io_valid_in ? _GEN_26175 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1599 = 12'h63f == _T_2[11:0] ? image_1599 : _GEN_1598; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4672 = 12'h640 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7744 = 12'h640 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4672; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10816 = 12'h640 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7744; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13888 = 12'h640 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10816; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16960 = 12'h640 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13888; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20032 = 12'h640 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16960; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23104 = 12'h640 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20032; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26176 = 12'h640 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23104; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1600 = io_valid_in ? _GEN_26176 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1600 = 12'h640 == _T_2[11:0] ? image_1600 : _GEN_1599; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4673 = 12'h641 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7745 = 12'h641 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4673; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10817 = 12'h641 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7745; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13889 = 12'h641 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10817; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16961 = 12'h641 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13889; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20033 = 12'h641 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16961; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23105 = 12'h641 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20033; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26177 = 12'h641 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23105; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1601 = io_valid_in ? _GEN_26177 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1601 = 12'h641 == _T_2[11:0] ? image_1601 : _GEN_1600; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4674 = 12'h642 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7746 = 12'h642 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4674; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10818 = 12'h642 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7746; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13890 = 12'h642 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10818; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16962 = 12'h642 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13890; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20034 = 12'h642 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16962; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23106 = 12'h642 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20034; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26178 = 12'h642 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23106; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1602 = io_valid_in ? _GEN_26178 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1602 = 12'h642 == _T_2[11:0] ? image_1602 : _GEN_1601; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4675 = 12'h643 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7747 = 12'h643 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4675; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10819 = 12'h643 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7747; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13891 = 12'h643 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10819; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16963 = 12'h643 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13891; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20035 = 12'h643 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16963; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23107 = 12'h643 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20035; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26179 = 12'h643 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23107; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1603 = io_valid_in ? _GEN_26179 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1603 = 12'h643 == _T_2[11:0] ? image_1603 : _GEN_1602; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4676 = 12'h644 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7748 = 12'h644 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4676; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10820 = 12'h644 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7748; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13892 = 12'h644 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10820; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16964 = 12'h644 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13892; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20036 = 12'h644 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16964; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23108 = 12'h644 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20036; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26180 = 12'h644 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23108; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1604 = io_valid_in ? _GEN_26180 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1604 = 12'h644 == _T_2[11:0] ? image_1604 : _GEN_1603; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4677 = 12'h645 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7749 = 12'h645 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4677; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10821 = 12'h645 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7749; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13893 = 12'h645 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10821; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16965 = 12'h645 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13893; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20037 = 12'h645 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16965; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23109 = 12'h645 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20037; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26181 = 12'h645 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23109; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1605 = io_valid_in ? _GEN_26181 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1605 = 12'h645 == _T_2[11:0] ? image_1605 : _GEN_1604; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4678 = 12'h646 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7750 = 12'h646 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4678; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10822 = 12'h646 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7750; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13894 = 12'h646 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10822; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16966 = 12'h646 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13894; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20038 = 12'h646 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16966; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23110 = 12'h646 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20038; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26182 = 12'h646 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23110; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1606 = io_valid_in ? _GEN_26182 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1606 = 12'h646 == _T_2[11:0] ? image_1606 : _GEN_1605; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4679 = 12'h647 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7751 = 12'h647 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4679; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10823 = 12'h647 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7751; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13895 = 12'h647 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10823; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16967 = 12'h647 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13895; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20039 = 12'h647 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16967; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23111 = 12'h647 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20039; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26183 = 12'h647 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23111; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1607 = io_valid_in ? _GEN_26183 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1607 = 12'h647 == _T_2[11:0] ? image_1607 : _GEN_1606; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4680 = 12'h648 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7752 = 12'h648 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4680; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10824 = 12'h648 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7752; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13896 = 12'h648 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10824; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16968 = 12'h648 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13896; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20040 = 12'h648 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16968; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23112 = 12'h648 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20040; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26184 = 12'h648 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23112; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1608 = io_valid_in ? _GEN_26184 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1608 = 12'h648 == _T_2[11:0] ? image_1608 : _GEN_1607; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4681 = 12'h649 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7753 = 12'h649 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4681; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10825 = 12'h649 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7753; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13897 = 12'h649 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10825; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16969 = 12'h649 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13897; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20041 = 12'h649 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16969; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23113 = 12'h649 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20041; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26185 = 12'h649 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23113; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1609 = io_valid_in ? _GEN_26185 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1609 = 12'h649 == _T_2[11:0] ? image_1609 : _GEN_1608; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4682 = 12'h64a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7754 = 12'h64a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4682; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10826 = 12'h64a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7754; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13898 = 12'h64a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10826; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16970 = 12'h64a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13898; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20042 = 12'h64a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16970; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23114 = 12'h64a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20042; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26186 = 12'h64a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23114; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1610 = io_valid_in ? _GEN_26186 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1610 = 12'h64a == _T_2[11:0] ? image_1610 : _GEN_1609; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4683 = 12'h64b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7755 = 12'h64b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4683; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10827 = 12'h64b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7755; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13899 = 12'h64b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10827; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16971 = 12'h64b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13899; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20043 = 12'h64b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16971; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23115 = 12'h64b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20043; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26187 = 12'h64b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23115; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1611 = io_valid_in ? _GEN_26187 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1611 = 12'h64b == _T_2[11:0] ? image_1611 : _GEN_1610; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4684 = 12'h64c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7756 = 12'h64c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4684; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10828 = 12'h64c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7756; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13900 = 12'h64c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10828; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16972 = 12'h64c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13900; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20044 = 12'h64c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16972; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23116 = 12'h64c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20044; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26188 = 12'h64c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23116; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1612 = io_valid_in ? _GEN_26188 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1612 = 12'h64c == _T_2[11:0] ? image_1612 : _GEN_1611; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4685 = 12'h64d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7757 = 12'h64d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4685; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10829 = 12'h64d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7757; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13901 = 12'h64d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10829; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16973 = 12'h64d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13901; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20045 = 12'h64d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16973; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23117 = 12'h64d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20045; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26189 = 12'h64d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23117; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1613 = io_valid_in ? _GEN_26189 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1613 = 12'h64d == _T_2[11:0] ? image_1613 : _GEN_1612; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4686 = 12'h64e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7758 = 12'h64e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4686; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10830 = 12'h64e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7758; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13902 = 12'h64e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10830; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16974 = 12'h64e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13902; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20046 = 12'h64e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16974; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23118 = 12'h64e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20046; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26190 = 12'h64e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23118; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1614 = io_valid_in ? _GEN_26190 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1614 = 12'h64e == _T_2[11:0] ? image_1614 : _GEN_1613; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4687 = 12'h64f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7759 = 12'h64f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4687; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10831 = 12'h64f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7759; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13903 = 12'h64f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10831; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16975 = 12'h64f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13903; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20047 = 12'h64f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16975; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23119 = 12'h64f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20047; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26191 = 12'h64f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23119; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1615 = io_valid_in ? _GEN_26191 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1615 = 12'h64f == _T_2[11:0] ? image_1615 : _GEN_1614; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4688 = 12'h650 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7760 = 12'h650 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4688; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10832 = 12'h650 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7760; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13904 = 12'h650 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10832; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16976 = 12'h650 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13904; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20048 = 12'h650 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16976; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23120 = 12'h650 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20048; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26192 = 12'h650 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23120; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1616 = io_valid_in ? _GEN_26192 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1616 = 12'h650 == _T_2[11:0] ? image_1616 : _GEN_1615; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4689 = 12'h651 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7761 = 12'h651 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4689; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10833 = 12'h651 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7761; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13905 = 12'h651 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10833; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16977 = 12'h651 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13905; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20049 = 12'h651 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16977; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23121 = 12'h651 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20049; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26193 = 12'h651 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23121; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1617 = io_valid_in ? _GEN_26193 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1617 = 12'h651 == _T_2[11:0] ? image_1617 : _GEN_1616; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4690 = 12'h652 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7762 = 12'h652 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4690; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10834 = 12'h652 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7762; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13906 = 12'h652 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10834; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16978 = 12'h652 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13906; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20050 = 12'h652 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16978; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23122 = 12'h652 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20050; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26194 = 12'h652 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23122; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1618 = io_valid_in ? _GEN_26194 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1618 = 12'h652 == _T_2[11:0] ? image_1618 : _GEN_1617; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4691 = 12'h653 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7763 = 12'h653 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4691; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10835 = 12'h653 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7763; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13907 = 12'h653 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10835; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16979 = 12'h653 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13907; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20051 = 12'h653 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16979; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23123 = 12'h653 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20051; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26195 = 12'h653 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23123; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1619 = io_valid_in ? _GEN_26195 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1619 = 12'h653 == _T_2[11:0] ? image_1619 : _GEN_1618; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4692 = 12'h654 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7764 = 12'h654 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4692; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10836 = 12'h654 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7764; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13908 = 12'h654 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10836; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16980 = 12'h654 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13908; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20052 = 12'h654 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16980; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23124 = 12'h654 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20052; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26196 = 12'h654 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23124; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1620 = io_valid_in ? _GEN_26196 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1620 = 12'h654 == _T_2[11:0] ? image_1620 : _GEN_1619; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4693 = 12'h655 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7765 = 12'h655 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4693; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10837 = 12'h655 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7765; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13909 = 12'h655 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10837; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16981 = 12'h655 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13909; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20053 = 12'h655 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16981; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23125 = 12'h655 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20053; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26197 = 12'h655 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23125; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1621 = io_valid_in ? _GEN_26197 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1621 = 12'h655 == _T_2[11:0] ? image_1621 : _GEN_1620; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4694 = 12'h656 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7766 = 12'h656 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4694; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10838 = 12'h656 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7766; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13910 = 12'h656 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10838; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16982 = 12'h656 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13910; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20054 = 12'h656 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16982; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23126 = 12'h656 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20054; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26198 = 12'h656 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23126; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1622 = io_valid_in ? _GEN_26198 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1622 = 12'h656 == _T_2[11:0] ? image_1622 : _GEN_1621; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4695 = 12'h657 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7767 = 12'h657 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4695; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10839 = 12'h657 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7767; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13911 = 12'h657 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10839; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16983 = 12'h657 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13911; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20055 = 12'h657 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16983; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23127 = 12'h657 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20055; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26199 = 12'h657 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23127; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1623 = io_valid_in ? _GEN_26199 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1623 = 12'h657 == _T_2[11:0] ? image_1623 : _GEN_1622; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4696 = 12'h658 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7768 = 12'h658 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4696; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10840 = 12'h658 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7768; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13912 = 12'h658 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10840; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16984 = 12'h658 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13912; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20056 = 12'h658 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16984; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23128 = 12'h658 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20056; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26200 = 12'h658 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23128; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1624 = io_valid_in ? _GEN_26200 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1624 = 12'h658 == _T_2[11:0] ? image_1624 : _GEN_1623; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4697 = 12'h659 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7769 = 12'h659 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4697; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10841 = 12'h659 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7769; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13913 = 12'h659 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10841; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16985 = 12'h659 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13913; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20057 = 12'h659 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16985; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23129 = 12'h659 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20057; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26201 = 12'h659 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23129; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1625 = io_valid_in ? _GEN_26201 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1625 = 12'h659 == _T_2[11:0] ? image_1625 : _GEN_1624; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4698 = 12'h65a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7770 = 12'h65a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4698; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10842 = 12'h65a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7770; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13914 = 12'h65a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10842; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16986 = 12'h65a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13914; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20058 = 12'h65a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16986; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23130 = 12'h65a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20058; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26202 = 12'h65a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23130; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1626 = io_valid_in ? _GEN_26202 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1626 = 12'h65a == _T_2[11:0] ? image_1626 : _GEN_1625; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4699 = 12'h65b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7771 = 12'h65b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4699; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10843 = 12'h65b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7771; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13915 = 12'h65b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10843; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16987 = 12'h65b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13915; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20059 = 12'h65b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16987; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23131 = 12'h65b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20059; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26203 = 12'h65b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23131; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1627 = io_valid_in ? _GEN_26203 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1627 = 12'h65b == _T_2[11:0] ? image_1627 : _GEN_1626; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4700 = 12'h65c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7772 = 12'h65c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4700; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10844 = 12'h65c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7772; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13916 = 12'h65c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10844; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16988 = 12'h65c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13916; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20060 = 12'h65c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16988; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23132 = 12'h65c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20060; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26204 = 12'h65c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23132; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1628 = io_valid_in ? _GEN_26204 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1628 = 12'h65c == _T_2[11:0] ? image_1628 : _GEN_1627; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4701 = 12'h65d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7773 = 12'h65d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4701; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10845 = 12'h65d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7773; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13917 = 12'h65d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10845; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16989 = 12'h65d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13917; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20061 = 12'h65d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16989; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23133 = 12'h65d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20061; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26205 = 12'h65d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23133; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1629 = io_valid_in ? _GEN_26205 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1629 = 12'h65d == _T_2[11:0] ? image_1629 : _GEN_1628; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4702 = 12'h65e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7774 = 12'h65e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4702; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10846 = 12'h65e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7774; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13918 = 12'h65e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10846; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16990 = 12'h65e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13918; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20062 = 12'h65e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16990; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23134 = 12'h65e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20062; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26206 = 12'h65e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23134; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1630 = io_valid_in ? _GEN_26206 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1630 = 12'h65e == _T_2[11:0] ? image_1630 : _GEN_1629; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4703 = 12'h65f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7775 = 12'h65f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4703; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10847 = 12'h65f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7775; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13919 = 12'h65f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10847; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16991 = 12'h65f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13919; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20063 = 12'h65f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16991; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23135 = 12'h65f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20063; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26207 = 12'h65f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23135; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1631 = io_valid_in ? _GEN_26207 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1631 = 12'h65f == _T_2[11:0] ? image_1631 : _GEN_1630; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4704 = 12'h660 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7776 = 12'h660 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4704; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10848 = 12'h660 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7776; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13920 = 12'h660 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10848; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16992 = 12'h660 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13920; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20064 = 12'h660 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16992; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23136 = 12'h660 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20064; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26208 = 12'h660 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23136; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1632 = io_valid_in ? _GEN_26208 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1632 = 12'h660 == _T_2[11:0] ? image_1632 : _GEN_1631; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4705 = 12'h661 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7777 = 12'h661 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4705; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10849 = 12'h661 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7777; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13921 = 12'h661 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10849; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16993 = 12'h661 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13921; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20065 = 12'h661 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16993; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23137 = 12'h661 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20065; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26209 = 12'h661 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23137; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1633 = io_valid_in ? _GEN_26209 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1633 = 12'h661 == _T_2[11:0] ? image_1633 : _GEN_1632; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4706 = 12'h662 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7778 = 12'h662 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4706; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10850 = 12'h662 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7778; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13922 = 12'h662 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10850; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16994 = 12'h662 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13922; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20066 = 12'h662 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16994; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23138 = 12'h662 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20066; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26210 = 12'h662 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23138; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1634 = io_valid_in ? _GEN_26210 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1634 = 12'h662 == _T_2[11:0] ? image_1634 : _GEN_1633; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4707 = 12'h663 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7779 = 12'h663 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4707; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10851 = 12'h663 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7779; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13923 = 12'h663 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10851; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16995 = 12'h663 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13923; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20067 = 12'h663 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16995; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23139 = 12'h663 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20067; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26211 = 12'h663 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23139; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1635 = io_valid_in ? _GEN_26211 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1635 = 12'h663 == _T_2[11:0] ? image_1635 : _GEN_1634; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4708 = 12'h664 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7780 = 12'h664 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4708; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10852 = 12'h664 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7780; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13924 = 12'h664 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10852; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16996 = 12'h664 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13924; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20068 = 12'h664 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16996; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23140 = 12'h664 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20068; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26212 = 12'h664 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23140; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1636 = io_valid_in ? _GEN_26212 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1636 = 12'h664 == _T_2[11:0] ? image_1636 : _GEN_1635; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4709 = 12'h665 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7781 = 12'h665 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4709; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10853 = 12'h665 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7781; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13925 = 12'h665 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10853; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16997 = 12'h665 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13925; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20069 = 12'h665 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16997; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23141 = 12'h665 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20069; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26213 = 12'h665 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23141; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1637 = io_valid_in ? _GEN_26213 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1637 = 12'h665 == _T_2[11:0] ? image_1637 : _GEN_1636; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4710 = 12'h666 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7782 = 12'h666 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4710; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10854 = 12'h666 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7782; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13926 = 12'h666 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10854; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16998 = 12'h666 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13926; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20070 = 12'h666 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16998; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23142 = 12'h666 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20070; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26214 = 12'h666 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23142; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1638 = io_valid_in ? _GEN_26214 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1638 = 12'h666 == _T_2[11:0] ? image_1638 : _GEN_1637; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4711 = 12'h667 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7783 = 12'h667 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4711; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10855 = 12'h667 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7783; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13927 = 12'h667 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10855; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_16999 = 12'h667 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13927; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20071 = 12'h667 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_16999; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23143 = 12'h667 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20071; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26215 = 12'h667 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23143; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1639 = io_valid_in ? _GEN_26215 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1639 = 12'h667 == _T_2[11:0] ? image_1639 : _GEN_1638; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4712 = 12'h668 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7784 = 12'h668 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4712; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10856 = 12'h668 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7784; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13928 = 12'h668 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10856; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17000 = 12'h668 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13928; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20072 = 12'h668 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17000; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23144 = 12'h668 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20072; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26216 = 12'h668 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23144; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1640 = io_valid_in ? _GEN_26216 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1640 = 12'h668 == _T_2[11:0] ? image_1640 : _GEN_1639; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4713 = 12'h669 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7785 = 12'h669 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4713; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10857 = 12'h669 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7785; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13929 = 12'h669 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10857; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17001 = 12'h669 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13929; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20073 = 12'h669 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17001; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23145 = 12'h669 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20073; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26217 = 12'h669 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23145; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1641 = io_valid_in ? _GEN_26217 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1641 = 12'h669 == _T_2[11:0] ? image_1641 : _GEN_1640; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4714 = 12'h66a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7786 = 12'h66a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4714; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10858 = 12'h66a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7786; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13930 = 12'h66a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10858; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17002 = 12'h66a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13930; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20074 = 12'h66a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17002; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23146 = 12'h66a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20074; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26218 = 12'h66a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23146; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1642 = io_valid_in ? _GEN_26218 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1642 = 12'h66a == _T_2[11:0] ? image_1642 : _GEN_1641; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4715 = 12'h66b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7787 = 12'h66b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4715; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10859 = 12'h66b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7787; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13931 = 12'h66b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10859; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17003 = 12'h66b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13931; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20075 = 12'h66b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17003; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23147 = 12'h66b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20075; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26219 = 12'h66b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23147; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1643 = io_valid_in ? _GEN_26219 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1643 = 12'h66b == _T_2[11:0] ? image_1643 : _GEN_1642; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4716 = 12'h66c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7788 = 12'h66c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4716; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10860 = 12'h66c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7788; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13932 = 12'h66c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10860; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17004 = 12'h66c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13932; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20076 = 12'h66c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17004; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23148 = 12'h66c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20076; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26220 = 12'h66c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23148; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1644 = io_valid_in ? _GEN_26220 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1644 = 12'h66c == _T_2[11:0] ? image_1644 : _GEN_1643; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4717 = 12'h66d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7789 = 12'h66d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4717; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10861 = 12'h66d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7789; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13933 = 12'h66d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10861; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17005 = 12'h66d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13933; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20077 = 12'h66d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17005; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23149 = 12'h66d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20077; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26221 = 12'h66d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23149; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1645 = io_valid_in ? _GEN_26221 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1645 = 12'h66d == _T_2[11:0] ? image_1645 : _GEN_1644; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4718 = 12'h66e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7790 = 12'h66e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4718; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10862 = 12'h66e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7790; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13934 = 12'h66e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10862; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17006 = 12'h66e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13934; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20078 = 12'h66e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17006; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23150 = 12'h66e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20078; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26222 = 12'h66e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23150; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1646 = io_valid_in ? _GEN_26222 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1646 = 12'h66e == _T_2[11:0] ? image_1646 : _GEN_1645; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4719 = 12'h66f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7791 = 12'h66f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4719; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10863 = 12'h66f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7791; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13935 = 12'h66f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10863; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17007 = 12'h66f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13935; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20079 = 12'h66f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17007; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23151 = 12'h66f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20079; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26223 = 12'h66f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23151; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1647 = io_valid_in ? _GEN_26223 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1647 = 12'h66f == _T_2[11:0] ? image_1647 : _GEN_1646; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4720 = 12'h670 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7792 = 12'h670 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4720; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10864 = 12'h670 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7792; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13936 = 12'h670 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10864; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17008 = 12'h670 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13936; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20080 = 12'h670 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17008; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23152 = 12'h670 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20080; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26224 = 12'h670 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23152; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1648 = io_valid_in ? _GEN_26224 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1648 = 12'h670 == _T_2[11:0] ? image_1648 : _GEN_1647; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4721 = 12'h671 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7793 = 12'h671 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4721; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10865 = 12'h671 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7793; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13937 = 12'h671 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10865; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17009 = 12'h671 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13937; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20081 = 12'h671 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17009; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23153 = 12'h671 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20081; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26225 = 12'h671 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23153; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1649 = io_valid_in ? _GEN_26225 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1649 = 12'h671 == _T_2[11:0] ? image_1649 : _GEN_1648; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4722 = 12'h672 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7794 = 12'h672 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4722; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10866 = 12'h672 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7794; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13938 = 12'h672 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10866; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17010 = 12'h672 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13938; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20082 = 12'h672 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17010; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23154 = 12'h672 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20082; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26226 = 12'h672 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23154; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1650 = io_valid_in ? _GEN_26226 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1650 = 12'h672 == _T_2[11:0] ? image_1650 : _GEN_1649; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4723 = 12'h673 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7795 = 12'h673 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4723; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10867 = 12'h673 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7795; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13939 = 12'h673 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10867; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17011 = 12'h673 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13939; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20083 = 12'h673 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17011; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23155 = 12'h673 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20083; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26227 = 12'h673 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23155; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1651 = io_valid_in ? _GEN_26227 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1651 = 12'h673 == _T_2[11:0] ? image_1651 : _GEN_1650; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4724 = 12'h674 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7796 = 12'h674 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4724; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10868 = 12'h674 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7796; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13940 = 12'h674 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10868; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17012 = 12'h674 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13940; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20084 = 12'h674 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17012; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23156 = 12'h674 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20084; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26228 = 12'h674 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23156; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1652 = io_valid_in ? _GEN_26228 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1652 = 12'h674 == _T_2[11:0] ? image_1652 : _GEN_1651; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4725 = 12'h675 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7797 = 12'h675 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4725; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10869 = 12'h675 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7797; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13941 = 12'h675 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10869; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17013 = 12'h675 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13941; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20085 = 12'h675 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17013; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23157 = 12'h675 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20085; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26229 = 12'h675 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23157; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1653 = io_valid_in ? _GEN_26229 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1653 = 12'h675 == _T_2[11:0] ? image_1653 : _GEN_1652; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4726 = 12'h676 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7798 = 12'h676 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4726; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10870 = 12'h676 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7798; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13942 = 12'h676 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10870; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17014 = 12'h676 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13942; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20086 = 12'h676 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17014; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23158 = 12'h676 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20086; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26230 = 12'h676 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23158; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1654 = io_valid_in ? _GEN_26230 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1654 = 12'h676 == _T_2[11:0] ? image_1654 : _GEN_1653; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4727 = 12'h677 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7799 = 12'h677 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4727; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10871 = 12'h677 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7799; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13943 = 12'h677 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10871; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17015 = 12'h677 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13943; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20087 = 12'h677 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17015; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23159 = 12'h677 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20087; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26231 = 12'h677 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23159; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1655 = io_valid_in ? _GEN_26231 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1655 = 12'h677 == _T_2[11:0] ? image_1655 : _GEN_1654; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4728 = 12'h678 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7800 = 12'h678 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4728; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10872 = 12'h678 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7800; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13944 = 12'h678 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10872; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17016 = 12'h678 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13944; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20088 = 12'h678 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17016; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23160 = 12'h678 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20088; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26232 = 12'h678 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23160; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1656 = io_valid_in ? _GEN_26232 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1656 = 12'h678 == _T_2[11:0] ? image_1656 : _GEN_1655; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4729 = 12'h679 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7801 = 12'h679 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4729; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10873 = 12'h679 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7801; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13945 = 12'h679 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10873; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17017 = 12'h679 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13945; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20089 = 12'h679 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17017; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23161 = 12'h679 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20089; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26233 = 12'h679 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23161; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1657 = io_valid_in ? _GEN_26233 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1657 = 12'h679 == _T_2[11:0] ? image_1657 : _GEN_1656; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4730 = 12'h67a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7802 = 12'h67a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4730; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10874 = 12'h67a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7802; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13946 = 12'h67a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10874; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17018 = 12'h67a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13946; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20090 = 12'h67a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17018; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23162 = 12'h67a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20090; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26234 = 12'h67a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23162; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1658 = io_valid_in ? _GEN_26234 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1658 = 12'h67a == _T_2[11:0] ? image_1658 : _GEN_1657; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4731 = 12'h67b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7803 = 12'h67b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4731; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10875 = 12'h67b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7803; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13947 = 12'h67b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10875; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17019 = 12'h67b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13947; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20091 = 12'h67b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17019; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23163 = 12'h67b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20091; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26235 = 12'h67b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23163; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1659 = io_valid_in ? _GEN_26235 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1659 = 12'h67b == _T_2[11:0] ? image_1659 : _GEN_1658; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4732 = 12'h67c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7804 = 12'h67c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4732; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10876 = 12'h67c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7804; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13948 = 12'h67c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10876; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17020 = 12'h67c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13948; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20092 = 12'h67c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17020; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23164 = 12'h67c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20092; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26236 = 12'h67c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23164; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1660 = io_valid_in ? _GEN_26236 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1660 = 12'h67c == _T_2[11:0] ? image_1660 : _GEN_1659; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4733 = 12'h67d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7805 = 12'h67d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4733; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10877 = 12'h67d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7805; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13949 = 12'h67d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10877; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17021 = 12'h67d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13949; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20093 = 12'h67d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17021; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23165 = 12'h67d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20093; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26237 = 12'h67d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23165; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1661 = io_valid_in ? _GEN_26237 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1661 = 12'h67d == _T_2[11:0] ? image_1661 : _GEN_1660; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4734 = 12'h67e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7806 = 12'h67e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4734; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10878 = 12'h67e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7806; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13950 = 12'h67e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10878; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17022 = 12'h67e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13950; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20094 = 12'h67e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17022; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23166 = 12'h67e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20094; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26238 = 12'h67e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23166; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1662 = io_valid_in ? _GEN_26238 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1662 = 12'h67e == _T_2[11:0] ? image_1662 : _GEN_1661; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4735 = 12'h67f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7807 = 12'h67f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4735; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10879 = 12'h67f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7807; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13951 = 12'h67f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10879; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17023 = 12'h67f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13951; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20095 = 12'h67f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17023; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23167 = 12'h67f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20095; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26239 = 12'h67f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23167; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1663 = io_valid_in ? _GEN_26239 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1663 = 12'h67f == _T_2[11:0] ? image_1663 : _GEN_1662; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4736 = 12'h680 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7808 = 12'h680 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4736; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10880 = 12'h680 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7808; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13952 = 12'h680 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10880; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17024 = 12'h680 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13952; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20096 = 12'h680 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17024; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23168 = 12'h680 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20096; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26240 = 12'h680 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23168; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1664 = io_valid_in ? _GEN_26240 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1664 = 12'h680 == _T_2[11:0] ? image_1664 : _GEN_1663; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4737 = 12'h681 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7809 = 12'h681 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4737; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10881 = 12'h681 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7809; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13953 = 12'h681 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10881; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17025 = 12'h681 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13953; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20097 = 12'h681 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17025; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23169 = 12'h681 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20097; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26241 = 12'h681 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23169; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1665 = io_valid_in ? _GEN_26241 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1665 = 12'h681 == _T_2[11:0] ? image_1665 : _GEN_1664; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4738 = 12'h682 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7810 = 12'h682 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4738; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10882 = 12'h682 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7810; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13954 = 12'h682 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10882; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17026 = 12'h682 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13954; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20098 = 12'h682 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17026; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23170 = 12'h682 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20098; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26242 = 12'h682 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23170; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1666 = io_valid_in ? _GEN_26242 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1666 = 12'h682 == _T_2[11:0] ? image_1666 : _GEN_1665; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4739 = 12'h683 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7811 = 12'h683 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4739; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10883 = 12'h683 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7811; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13955 = 12'h683 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10883; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17027 = 12'h683 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13955; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20099 = 12'h683 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17027; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23171 = 12'h683 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20099; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26243 = 12'h683 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23171; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1667 = io_valid_in ? _GEN_26243 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1667 = 12'h683 == _T_2[11:0] ? image_1667 : _GEN_1666; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4740 = 12'h684 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7812 = 12'h684 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4740; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10884 = 12'h684 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7812; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13956 = 12'h684 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10884; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17028 = 12'h684 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13956; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20100 = 12'h684 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17028; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23172 = 12'h684 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20100; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26244 = 12'h684 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23172; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1668 = io_valid_in ? _GEN_26244 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1668 = 12'h684 == _T_2[11:0] ? image_1668 : _GEN_1667; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4741 = 12'h685 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7813 = 12'h685 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4741; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10885 = 12'h685 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7813; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13957 = 12'h685 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10885; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17029 = 12'h685 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13957; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20101 = 12'h685 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17029; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23173 = 12'h685 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20101; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26245 = 12'h685 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23173; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1669 = io_valid_in ? _GEN_26245 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1669 = 12'h685 == _T_2[11:0] ? image_1669 : _GEN_1668; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4742 = 12'h686 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7814 = 12'h686 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4742; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10886 = 12'h686 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7814; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13958 = 12'h686 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10886; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17030 = 12'h686 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13958; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20102 = 12'h686 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17030; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23174 = 12'h686 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20102; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26246 = 12'h686 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23174; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1670 = io_valid_in ? _GEN_26246 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1670 = 12'h686 == _T_2[11:0] ? image_1670 : _GEN_1669; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4743 = 12'h687 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7815 = 12'h687 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4743; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10887 = 12'h687 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7815; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13959 = 12'h687 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10887; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17031 = 12'h687 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13959; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20103 = 12'h687 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17031; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23175 = 12'h687 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20103; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26247 = 12'h687 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23175; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1671 = io_valid_in ? _GEN_26247 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1671 = 12'h687 == _T_2[11:0] ? image_1671 : _GEN_1670; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4744 = 12'h688 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7816 = 12'h688 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4744; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10888 = 12'h688 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7816; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13960 = 12'h688 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10888; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17032 = 12'h688 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13960; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20104 = 12'h688 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17032; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23176 = 12'h688 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20104; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26248 = 12'h688 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23176; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1672 = io_valid_in ? _GEN_26248 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1672 = 12'h688 == _T_2[11:0] ? image_1672 : _GEN_1671; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4745 = 12'h689 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7817 = 12'h689 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4745; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10889 = 12'h689 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7817; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13961 = 12'h689 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10889; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17033 = 12'h689 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13961; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20105 = 12'h689 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17033; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23177 = 12'h689 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20105; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26249 = 12'h689 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23177; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1673 = io_valid_in ? _GEN_26249 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1673 = 12'h689 == _T_2[11:0] ? image_1673 : _GEN_1672; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4746 = 12'h68a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7818 = 12'h68a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4746; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10890 = 12'h68a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7818; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13962 = 12'h68a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10890; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17034 = 12'h68a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13962; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20106 = 12'h68a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17034; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23178 = 12'h68a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20106; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26250 = 12'h68a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23178; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1674 = io_valid_in ? _GEN_26250 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1674 = 12'h68a == _T_2[11:0] ? image_1674 : _GEN_1673; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4747 = 12'h68b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7819 = 12'h68b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4747; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10891 = 12'h68b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7819; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13963 = 12'h68b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10891; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17035 = 12'h68b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13963; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20107 = 12'h68b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17035; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23179 = 12'h68b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20107; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26251 = 12'h68b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23179; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1675 = io_valid_in ? _GEN_26251 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1675 = 12'h68b == _T_2[11:0] ? image_1675 : _GEN_1674; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4748 = 12'h68c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7820 = 12'h68c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4748; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10892 = 12'h68c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7820; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13964 = 12'h68c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10892; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17036 = 12'h68c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13964; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20108 = 12'h68c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17036; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23180 = 12'h68c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20108; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26252 = 12'h68c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23180; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1676 = io_valid_in ? _GEN_26252 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1676 = 12'h68c == _T_2[11:0] ? image_1676 : _GEN_1675; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4749 = 12'h68d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7821 = 12'h68d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4749; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10893 = 12'h68d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7821; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13965 = 12'h68d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10893; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17037 = 12'h68d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13965; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20109 = 12'h68d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17037; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23181 = 12'h68d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20109; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26253 = 12'h68d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23181; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1677 = io_valid_in ? _GEN_26253 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1677 = 12'h68d == _T_2[11:0] ? image_1677 : _GEN_1676; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4750 = 12'h68e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7822 = 12'h68e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4750; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10894 = 12'h68e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7822; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13966 = 12'h68e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10894; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17038 = 12'h68e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13966; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20110 = 12'h68e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17038; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23182 = 12'h68e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20110; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26254 = 12'h68e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23182; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1678 = io_valid_in ? _GEN_26254 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1678 = 12'h68e == _T_2[11:0] ? image_1678 : _GEN_1677; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4751 = 12'h68f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7823 = 12'h68f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4751; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10895 = 12'h68f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7823; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13967 = 12'h68f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10895; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17039 = 12'h68f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13967; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20111 = 12'h68f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17039; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23183 = 12'h68f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20111; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26255 = 12'h68f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23183; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1679 = io_valid_in ? _GEN_26255 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1679 = 12'h68f == _T_2[11:0] ? image_1679 : _GEN_1678; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4752 = 12'h690 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7824 = 12'h690 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4752; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10896 = 12'h690 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7824; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13968 = 12'h690 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10896; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17040 = 12'h690 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13968; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20112 = 12'h690 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17040; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23184 = 12'h690 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20112; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26256 = 12'h690 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23184; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1680 = io_valid_in ? _GEN_26256 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1680 = 12'h690 == _T_2[11:0] ? image_1680 : _GEN_1679; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4753 = 12'h691 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7825 = 12'h691 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4753; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10897 = 12'h691 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7825; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13969 = 12'h691 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10897; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17041 = 12'h691 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13969; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20113 = 12'h691 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17041; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23185 = 12'h691 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20113; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26257 = 12'h691 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23185; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1681 = io_valid_in ? _GEN_26257 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1681 = 12'h691 == _T_2[11:0] ? image_1681 : _GEN_1680; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4754 = 12'h692 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7826 = 12'h692 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4754; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10898 = 12'h692 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7826; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13970 = 12'h692 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10898; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17042 = 12'h692 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13970; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20114 = 12'h692 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17042; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23186 = 12'h692 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20114; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26258 = 12'h692 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23186; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1682 = io_valid_in ? _GEN_26258 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1682 = 12'h692 == _T_2[11:0] ? image_1682 : _GEN_1681; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4755 = 12'h693 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7827 = 12'h693 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4755; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10899 = 12'h693 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7827; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13971 = 12'h693 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10899; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17043 = 12'h693 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13971; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20115 = 12'h693 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17043; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23187 = 12'h693 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20115; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26259 = 12'h693 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23187; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1683 = io_valid_in ? _GEN_26259 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1683 = 12'h693 == _T_2[11:0] ? image_1683 : _GEN_1682; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4756 = 12'h694 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7828 = 12'h694 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4756; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10900 = 12'h694 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7828; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13972 = 12'h694 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10900; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17044 = 12'h694 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13972; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20116 = 12'h694 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17044; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23188 = 12'h694 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20116; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26260 = 12'h694 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23188; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1684 = io_valid_in ? _GEN_26260 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1684 = 12'h694 == _T_2[11:0] ? image_1684 : _GEN_1683; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4757 = 12'h695 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7829 = 12'h695 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4757; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10901 = 12'h695 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7829; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13973 = 12'h695 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10901; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17045 = 12'h695 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13973; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20117 = 12'h695 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17045; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23189 = 12'h695 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20117; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26261 = 12'h695 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23189; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1685 = io_valid_in ? _GEN_26261 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1685 = 12'h695 == _T_2[11:0] ? image_1685 : _GEN_1684; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4758 = 12'h696 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7830 = 12'h696 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4758; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10902 = 12'h696 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7830; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13974 = 12'h696 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10902; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17046 = 12'h696 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13974; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20118 = 12'h696 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17046; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23190 = 12'h696 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20118; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26262 = 12'h696 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23190; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1686 = io_valid_in ? _GEN_26262 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1686 = 12'h696 == _T_2[11:0] ? image_1686 : _GEN_1685; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4759 = 12'h697 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7831 = 12'h697 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4759; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10903 = 12'h697 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7831; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13975 = 12'h697 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10903; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17047 = 12'h697 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13975; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20119 = 12'h697 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17047; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23191 = 12'h697 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20119; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26263 = 12'h697 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23191; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1687 = io_valid_in ? _GEN_26263 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1687 = 12'h697 == _T_2[11:0] ? image_1687 : _GEN_1686; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4760 = 12'h698 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7832 = 12'h698 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4760; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10904 = 12'h698 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7832; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13976 = 12'h698 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10904; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17048 = 12'h698 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13976; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20120 = 12'h698 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17048; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23192 = 12'h698 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20120; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26264 = 12'h698 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23192; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1688 = io_valid_in ? _GEN_26264 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1688 = 12'h698 == _T_2[11:0] ? image_1688 : _GEN_1687; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4761 = 12'h699 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7833 = 12'h699 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4761; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10905 = 12'h699 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7833; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13977 = 12'h699 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10905; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17049 = 12'h699 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13977; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20121 = 12'h699 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17049; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23193 = 12'h699 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20121; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26265 = 12'h699 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23193; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1689 = io_valid_in ? _GEN_26265 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1689 = 12'h699 == _T_2[11:0] ? image_1689 : _GEN_1688; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4762 = 12'h69a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7834 = 12'h69a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4762; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10906 = 12'h69a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7834; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13978 = 12'h69a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10906; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17050 = 12'h69a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13978; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20122 = 12'h69a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17050; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23194 = 12'h69a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20122; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26266 = 12'h69a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23194; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1690 = io_valid_in ? _GEN_26266 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1690 = 12'h69a == _T_2[11:0] ? image_1690 : _GEN_1689; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4763 = 12'h69b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7835 = 12'h69b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4763; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10907 = 12'h69b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7835; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13979 = 12'h69b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10907; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17051 = 12'h69b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13979; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20123 = 12'h69b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17051; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23195 = 12'h69b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20123; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26267 = 12'h69b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23195; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1691 = io_valid_in ? _GEN_26267 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1691 = 12'h69b == _T_2[11:0] ? image_1691 : _GEN_1690; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4764 = 12'h69c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7836 = 12'h69c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4764; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10908 = 12'h69c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7836; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13980 = 12'h69c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10908; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17052 = 12'h69c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13980; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20124 = 12'h69c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17052; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23196 = 12'h69c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20124; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26268 = 12'h69c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23196; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1692 = io_valid_in ? _GEN_26268 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1692 = 12'h69c == _T_2[11:0] ? image_1692 : _GEN_1691; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4765 = 12'h69d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7837 = 12'h69d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4765; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10909 = 12'h69d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7837; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13981 = 12'h69d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10909; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17053 = 12'h69d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13981; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20125 = 12'h69d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17053; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23197 = 12'h69d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20125; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26269 = 12'h69d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23197; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1693 = io_valid_in ? _GEN_26269 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1693 = 12'h69d == _T_2[11:0] ? image_1693 : _GEN_1692; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4766 = 12'h69e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7838 = 12'h69e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4766; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10910 = 12'h69e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7838; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13982 = 12'h69e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10910; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17054 = 12'h69e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13982; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20126 = 12'h69e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17054; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23198 = 12'h69e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20126; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26270 = 12'h69e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23198; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1694 = io_valid_in ? _GEN_26270 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1694 = 12'h69e == _T_2[11:0] ? image_1694 : _GEN_1693; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4767 = 12'h69f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7839 = 12'h69f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4767; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10911 = 12'h69f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7839; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13983 = 12'h69f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10911; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17055 = 12'h69f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13983; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20127 = 12'h69f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17055; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23199 = 12'h69f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20127; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26271 = 12'h69f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23199; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1695 = io_valid_in ? _GEN_26271 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1695 = 12'h69f == _T_2[11:0] ? image_1695 : _GEN_1694; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4768 = 12'h6a0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7840 = 12'h6a0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4768; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10912 = 12'h6a0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7840; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13984 = 12'h6a0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10912; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17056 = 12'h6a0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13984; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20128 = 12'h6a0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17056; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23200 = 12'h6a0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20128; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26272 = 12'h6a0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23200; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1696 = io_valid_in ? _GEN_26272 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1696 = 12'h6a0 == _T_2[11:0] ? image_1696 : _GEN_1695; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4769 = 12'h6a1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7841 = 12'h6a1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4769; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10913 = 12'h6a1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7841; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13985 = 12'h6a1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10913; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17057 = 12'h6a1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13985; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20129 = 12'h6a1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17057; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23201 = 12'h6a1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20129; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26273 = 12'h6a1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23201; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1697 = io_valid_in ? _GEN_26273 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1697 = 12'h6a1 == _T_2[11:0] ? image_1697 : _GEN_1696; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4770 = 12'h6a2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7842 = 12'h6a2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4770; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10914 = 12'h6a2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7842; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13986 = 12'h6a2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10914; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17058 = 12'h6a2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13986; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20130 = 12'h6a2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17058; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23202 = 12'h6a2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20130; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26274 = 12'h6a2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23202; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1698 = io_valid_in ? _GEN_26274 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1698 = 12'h6a2 == _T_2[11:0] ? image_1698 : _GEN_1697; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4771 = 12'h6a3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7843 = 12'h6a3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4771; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10915 = 12'h6a3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7843; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13987 = 12'h6a3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10915; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17059 = 12'h6a3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13987; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20131 = 12'h6a3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17059; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23203 = 12'h6a3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20131; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26275 = 12'h6a3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23203; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1699 = io_valid_in ? _GEN_26275 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1699 = 12'h6a3 == _T_2[11:0] ? image_1699 : _GEN_1698; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4772 = 12'h6a4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7844 = 12'h6a4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4772; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10916 = 12'h6a4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7844; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13988 = 12'h6a4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10916; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17060 = 12'h6a4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13988; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20132 = 12'h6a4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17060; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23204 = 12'h6a4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20132; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26276 = 12'h6a4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23204; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1700 = io_valid_in ? _GEN_26276 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1700 = 12'h6a4 == _T_2[11:0] ? image_1700 : _GEN_1699; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4773 = 12'h6a5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7845 = 12'h6a5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4773; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10917 = 12'h6a5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7845; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13989 = 12'h6a5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10917; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17061 = 12'h6a5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13989; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20133 = 12'h6a5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17061; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23205 = 12'h6a5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20133; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26277 = 12'h6a5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23205; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1701 = io_valid_in ? _GEN_26277 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1701 = 12'h6a5 == _T_2[11:0] ? image_1701 : _GEN_1700; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4774 = 12'h6a6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7846 = 12'h6a6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4774; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10918 = 12'h6a6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7846; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13990 = 12'h6a6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10918; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17062 = 12'h6a6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13990; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20134 = 12'h6a6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17062; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23206 = 12'h6a6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20134; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26278 = 12'h6a6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23206; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1702 = io_valid_in ? _GEN_26278 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1702 = 12'h6a6 == _T_2[11:0] ? image_1702 : _GEN_1701; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4775 = 12'h6a7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7847 = 12'h6a7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4775; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10919 = 12'h6a7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7847; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13991 = 12'h6a7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10919; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17063 = 12'h6a7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13991; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20135 = 12'h6a7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17063; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23207 = 12'h6a7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20135; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26279 = 12'h6a7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23207; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1703 = io_valid_in ? _GEN_26279 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1703 = 12'h6a7 == _T_2[11:0] ? image_1703 : _GEN_1702; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4776 = 12'h6a8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7848 = 12'h6a8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4776; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10920 = 12'h6a8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7848; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13992 = 12'h6a8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10920; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17064 = 12'h6a8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13992; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20136 = 12'h6a8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17064; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23208 = 12'h6a8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20136; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26280 = 12'h6a8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23208; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1704 = io_valid_in ? _GEN_26280 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1704 = 12'h6a8 == _T_2[11:0] ? image_1704 : _GEN_1703; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4777 = 12'h6a9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7849 = 12'h6a9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4777; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10921 = 12'h6a9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7849; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13993 = 12'h6a9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10921; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17065 = 12'h6a9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13993; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20137 = 12'h6a9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17065; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23209 = 12'h6a9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20137; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26281 = 12'h6a9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23209; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1705 = io_valid_in ? _GEN_26281 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1705 = 12'h6a9 == _T_2[11:0] ? image_1705 : _GEN_1704; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4778 = 12'h6aa == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7850 = 12'h6aa == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4778; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10922 = 12'h6aa == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7850; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13994 = 12'h6aa == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10922; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17066 = 12'h6aa == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13994; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20138 = 12'h6aa == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17066; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23210 = 12'h6aa == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20138; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26282 = 12'h6aa == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23210; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1706 = io_valid_in ? _GEN_26282 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1706 = 12'h6aa == _T_2[11:0] ? image_1706 : _GEN_1705; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4779 = 12'h6ab == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7851 = 12'h6ab == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4779; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10923 = 12'h6ab == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7851; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13995 = 12'h6ab == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10923; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17067 = 12'h6ab == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13995; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20139 = 12'h6ab == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17067; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23211 = 12'h6ab == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20139; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26283 = 12'h6ab == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23211; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1707 = io_valid_in ? _GEN_26283 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1707 = 12'h6ab == _T_2[11:0] ? image_1707 : _GEN_1706; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4780 = 12'h6ac == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7852 = 12'h6ac == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4780; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10924 = 12'h6ac == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7852; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13996 = 12'h6ac == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10924; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17068 = 12'h6ac == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13996; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20140 = 12'h6ac == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17068; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23212 = 12'h6ac == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20140; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26284 = 12'h6ac == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23212; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1708 = io_valid_in ? _GEN_26284 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1708 = 12'h6ac == _T_2[11:0] ? image_1708 : _GEN_1707; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4781 = 12'h6ad == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7853 = 12'h6ad == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4781; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10925 = 12'h6ad == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7853; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13997 = 12'h6ad == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10925; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17069 = 12'h6ad == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13997; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20141 = 12'h6ad == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17069; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23213 = 12'h6ad == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20141; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26285 = 12'h6ad == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23213; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1709 = io_valid_in ? _GEN_26285 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1709 = 12'h6ad == _T_2[11:0] ? image_1709 : _GEN_1708; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4782 = 12'h6ae == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7854 = 12'h6ae == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4782; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10926 = 12'h6ae == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7854; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13998 = 12'h6ae == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10926; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17070 = 12'h6ae == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13998; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20142 = 12'h6ae == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17070; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23214 = 12'h6ae == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20142; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26286 = 12'h6ae == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23214; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1710 = io_valid_in ? _GEN_26286 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1710 = 12'h6ae == _T_2[11:0] ? image_1710 : _GEN_1709; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4783 = 12'h6af == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7855 = 12'h6af == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4783; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10927 = 12'h6af == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7855; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_13999 = 12'h6af == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10927; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17071 = 12'h6af == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_13999; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20143 = 12'h6af == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17071; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23215 = 12'h6af == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20143; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26287 = 12'h6af == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23215; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1711 = io_valid_in ? _GEN_26287 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1711 = 12'h6af == _T_2[11:0] ? image_1711 : _GEN_1710; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4784 = 12'h6b0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7856 = 12'h6b0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4784; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10928 = 12'h6b0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7856; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14000 = 12'h6b0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10928; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17072 = 12'h6b0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14000; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20144 = 12'h6b0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17072; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23216 = 12'h6b0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20144; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26288 = 12'h6b0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23216; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1712 = io_valid_in ? _GEN_26288 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1712 = 12'h6b0 == _T_2[11:0] ? image_1712 : _GEN_1711; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4785 = 12'h6b1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7857 = 12'h6b1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4785; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10929 = 12'h6b1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7857; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14001 = 12'h6b1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10929; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17073 = 12'h6b1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14001; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20145 = 12'h6b1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17073; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23217 = 12'h6b1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20145; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26289 = 12'h6b1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23217; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1713 = io_valid_in ? _GEN_26289 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1713 = 12'h6b1 == _T_2[11:0] ? image_1713 : _GEN_1712; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4786 = 12'h6b2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7858 = 12'h6b2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4786; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10930 = 12'h6b2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7858; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14002 = 12'h6b2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10930; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17074 = 12'h6b2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14002; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20146 = 12'h6b2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17074; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23218 = 12'h6b2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20146; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26290 = 12'h6b2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23218; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1714 = io_valid_in ? _GEN_26290 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1714 = 12'h6b2 == _T_2[11:0] ? image_1714 : _GEN_1713; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4787 = 12'h6b3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7859 = 12'h6b3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4787; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10931 = 12'h6b3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7859; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14003 = 12'h6b3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10931; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17075 = 12'h6b3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14003; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20147 = 12'h6b3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17075; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23219 = 12'h6b3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20147; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26291 = 12'h6b3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23219; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1715 = io_valid_in ? _GEN_26291 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1715 = 12'h6b3 == _T_2[11:0] ? image_1715 : _GEN_1714; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4788 = 12'h6b4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7860 = 12'h6b4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4788; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10932 = 12'h6b4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7860; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14004 = 12'h6b4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10932; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17076 = 12'h6b4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14004; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20148 = 12'h6b4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17076; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23220 = 12'h6b4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20148; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26292 = 12'h6b4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23220; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1716 = io_valid_in ? _GEN_26292 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1716 = 12'h6b4 == _T_2[11:0] ? image_1716 : _GEN_1715; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4789 = 12'h6b5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7861 = 12'h6b5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4789; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10933 = 12'h6b5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7861; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14005 = 12'h6b5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10933; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17077 = 12'h6b5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14005; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20149 = 12'h6b5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17077; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23221 = 12'h6b5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20149; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26293 = 12'h6b5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23221; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1717 = io_valid_in ? _GEN_26293 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1717 = 12'h6b5 == _T_2[11:0] ? image_1717 : _GEN_1716; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4790 = 12'h6b6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7862 = 12'h6b6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4790; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10934 = 12'h6b6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7862; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14006 = 12'h6b6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10934; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17078 = 12'h6b6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14006; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20150 = 12'h6b6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17078; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23222 = 12'h6b6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20150; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26294 = 12'h6b6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23222; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1718 = io_valid_in ? _GEN_26294 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1718 = 12'h6b6 == _T_2[11:0] ? image_1718 : _GEN_1717; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4791 = 12'h6b7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7863 = 12'h6b7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4791; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10935 = 12'h6b7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7863; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14007 = 12'h6b7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10935; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17079 = 12'h6b7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14007; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20151 = 12'h6b7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17079; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23223 = 12'h6b7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20151; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26295 = 12'h6b7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23223; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1719 = io_valid_in ? _GEN_26295 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1719 = 12'h6b7 == _T_2[11:0] ? image_1719 : _GEN_1718; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4792 = 12'h6b8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7864 = 12'h6b8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4792; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10936 = 12'h6b8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7864; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14008 = 12'h6b8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10936; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17080 = 12'h6b8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14008; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20152 = 12'h6b8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17080; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23224 = 12'h6b8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20152; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26296 = 12'h6b8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23224; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1720 = io_valid_in ? _GEN_26296 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1720 = 12'h6b8 == _T_2[11:0] ? image_1720 : _GEN_1719; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4793 = 12'h6b9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7865 = 12'h6b9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4793; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10937 = 12'h6b9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7865; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14009 = 12'h6b9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10937; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17081 = 12'h6b9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14009; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20153 = 12'h6b9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17081; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23225 = 12'h6b9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20153; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26297 = 12'h6b9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23225; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1721 = io_valid_in ? _GEN_26297 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1721 = 12'h6b9 == _T_2[11:0] ? image_1721 : _GEN_1720; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4794 = 12'h6ba == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7866 = 12'h6ba == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4794; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10938 = 12'h6ba == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7866; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14010 = 12'h6ba == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10938; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17082 = 12'h6ba == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14010; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20154 = 12'h6ba == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17082; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23226 = 12'h6ba == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20154; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26298 = 12'h6ba == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23226; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1722 = io_valid_in ? _GEN_26298 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1722 = 12'h6ba == _T_2[11:0] ? image_1722 : _GEN_1721; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4795 = 12'h6bb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7867 = 12'h6bb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4795; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10939 = 12'h6bb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7867; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14011 = 12'h6bb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10939; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17083 = 12'h6bb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14011; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20155 = 12'h6bb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17083; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23227 = 12'h6bb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20155; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26299 = 12'h6bb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23227; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1723 = io_valid_in ? _GEN_26299 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1723 = 12'h6bb == _T_2[11:0] ? image_1723 : _GEN_1722; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4796 = 12'h6bc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7868 = 12'h6bc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4796; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10940 = 12'h6bc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7868; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14012 = 12'h6bc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10940; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17084 = 12'h6bc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14012; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20156 = 12'h6bc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17084; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23228 = 12'h6bc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20156; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26300 = 12'h6bc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23228; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1724 = io_valid_in ? _GEN_26300 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1724 = 12'h6bc == _T_2[11:0] ? image_1724 : _GEN_1723; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4797 = 12'h6bd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7869 = 12'h6bd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4797; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10941 = 12'h6bd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7869; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14013 = 12'h6bd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10941; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17085 = 12'h6bd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14013; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20157 = 12'h6bd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17085; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23229 = 12'h6bd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20157; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26301 = 12'h6bd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23229; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1725 = io_valid_in ? _GEN_26301 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1725 = 12'h6bd == _T_2[11:0] ? image_1725 : _GEN_1724; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4798 = 12'h6be == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7870 = 12'h6be == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4798; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10942 = 12'h6be == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7870; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14014 = 12'h6be == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10942; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17086 = 12'h6be == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14014; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20158 = 12'h6be == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17086; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23230 = 12'h6be == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20158; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26302 = 12'h6be == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23230; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1726 = io_valid_in ? _GEN_26302 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1726 = 12'h6be == _T_2[11:0] ? image_1726 : _GEN_1725; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4799 = 12'h6bf == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7871 = 12'h6bf == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4799; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10943 = 12'h6bf == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7871; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14015 = 12'h6bf == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10943; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17087 = 12'h6bf == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14015; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20159 = 12'h6bf == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17087; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23231 = 12'h6bf == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20159; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26303 = 12'h6bf == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23231; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1727 = io_valid_in ? _GEN_26303 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1727 = 12'h6bf == _T_2[11:0] ? image_1727 : _GEN_1726; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4800 = 12'h6c0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7872 = 12'h6c0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4800; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10944 = 12'h6c0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7872; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14016 = 12'h6c0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10944; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17088 = 12'h6c0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14016; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20160 = 12'h6c0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17088; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23232 = 12'h6c0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20160; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26304 = 12'h6c0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23232; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1728 = io_valid_in ? _GEN_26304 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1728 = 12'h6c0 == _T_2[11:0] ? image_1728 : _GEN_1727; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4801 = 12'h6c1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7873 = 12'h6c1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4801; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10945 = 12'h6c1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7873; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14017 = 12'h6c1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10945; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17089 = 12'h6c1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14017; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20161 = 12'h6c1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17089; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23233 = 12'h6c1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20161; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26305 = 12'h6c1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23233; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1729 = io_valid_in ? _GEN_26305 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1729 = 12'h6c1 == _T_2[11:0] ? image_1729 : _GEN_1728; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4802 = 12'h6c2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7874 = 12'h6c2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4802; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10946 = 12'h6c2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7874; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14018 = 12'h6c2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10946; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17090 = 12'h6c2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14018; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20162 = 12'h6c2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17090; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23234 = 12'h6c2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20162; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26306 = 12'h6c2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23234; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1730 = io_valid_in ? _GEN_26306 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1730 = 12'h6c2 == _T_2[11:0] ? image_1730 : _GEN_1729; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4803 = 12'h6c3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7875 = 12'h6c3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4803; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10947 = 12'h6c3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7875; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14019 = 12'h6c3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10947; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17091 = 12'h6c3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14019; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20163 = 12'h6c3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17091; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23235 = 12'h6c3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20163; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26307 = 12'h6c3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23235; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1731 = io_valid_in ? _GEN_26307 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1731 = 12'h6c3 == _T_2[11:0] ? image_1731 : _GEN_1730; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4804 = 12'h6c4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7876 = 12'h6c4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4804; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10948 = 12'h6c4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7876; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14020 = 12'h6c4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10948; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17092 = 12'h6c4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14020; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20164 = 12'h6c4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17092; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23236 = 12'h6c4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20164; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26308 = 12'h6c4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23236; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1732 = io_valid_in ? _GEN_26308 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1732 = 12'h6c4 == _T_2[11:0] ? image_1732 : _GEN_1731; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4805 = 12'h6c5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7877 = 12'h6c5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4805; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10949 = 12'h6c5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7877; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14021 = 12'h6c5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10949; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17093 = 12'h6c5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14021; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20165 = 12'h6c5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17093; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23237 = 12'h6c5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20165; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26309 = 12'h6c5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23237; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1733 = io_valid_in ? _GEN_26309 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1733 = 12'h6c5 == _T_2[11:0] ? image_1733 : _GEN_1732; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4806 = 12'h6c6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7878 = 12'h6c6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4806; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10950 = 12'h6c6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7878; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14022 = 12'h6c6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10950; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17094 = 12'h6c6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14022; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20166 = 12'h6c6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17094; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23238 = 12'h6c6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20166; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26310 = 12'h6c6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23238; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1734 = io_valid_in ? _GEN_26310 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1734 = 12'h6c6 == _T_2[11:0] ? image_1734 : _GEN_1733; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4807 = 12'h6c7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7879 = 12'h6c7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4807; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10951 = 12'h6c7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7879; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14023 = 12'h6c7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10951; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17095 = 12'h6c7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14023; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20167 = 12'h6c7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17095; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23239 = 12'h6c7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20167; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26311 = 12'h6c7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23239; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1735 = io_valid_in ? _GEN_26311 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1735 = 12'h6c7 == _T_2[11:0] ? image_1735 : _GEN_1734; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4808 = 12'h6c8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7880 = 12'h6c8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4808; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10952 = 12'h6c8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7880; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14024 = 12'h6c8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10952; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17096 = 12'h6c8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14024; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20168 = 12'h6c8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17096; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23240 = 12'h6c8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20168; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26312 = 12'h6c8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23240; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1736 = io_valid_in ? _GEN_26312 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1736 = 12'h6c8 == _T_2[11:0] ? image_1736 : _GEN_1735; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4809 = 12'h6c9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7881 = 12'h6c9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4809; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10953 = 12'h6c9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7881; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14025 = 12'h6c9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10953; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17097 = 12'h6c9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14025; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20169 = 12'h6c9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17097; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23241 = 12'h6c9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20169; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26313 = 12'h6c9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23241; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1737 = io_valid_in ? _GEN_26313 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1737 = 12'h6c9 == _T_2[11:0] ? image_1737 : _GEN_1736; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4810 = 12'h6ca == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7882 = 12'h6ca == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4810; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10954 = 12'h6ca == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7882; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14026 = 12'h6ca == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10954; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17098 = 12'h6ca == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14026; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20170 = 12'h6ca == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17098; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23242 = 12'h6ca == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20170; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26314 = 12'h6ca == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23242; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1738 = io_valid_in ? _GEN_26314 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1738 = 12'h6ca == _T_2[11:0] ? image_1738 : _GEN_1737; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4811 = 12'h6cb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7883 = 12'h6cb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4811; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10955 = 12'h6cb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7883; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14027 = 12'h6cb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10955; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17099 = 12'h6cb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14027; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20171 = 12'h6cb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17099; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23243 = 12'h6cb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20171; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26315 = 12'h6cb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23243; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1739 = io_valid_in ? _GEN_26315 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1739 = 12'h6cb == _T_2[11:0] ? image_1739 : _GEN_1738; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4812 = 12'h6cc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7884 = 12'h6cc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4812; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10956 = 12'h6cc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7884; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14028 = 12'h6cc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10956; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17100 = 12'h6cc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14028; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20172 = 12'h6cc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17100; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23244 = 12'h6cc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20172; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26316 = 12'h6cc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23244; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1740 = io_valid_in ? _GEN_26316 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1740 = 12'h6cc == _T_2[11:0] ? image_1740 : _GEN_1739; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4813 = 12'h6cd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7885 = 12'h6cd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4813; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10957 = 12'h6cd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7885; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14029 = 12'h6cd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10957; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17101 = 12'h6cd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14029; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20173 = 12'h6cd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17101; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23245 = 12'h6cd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20173; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26317 = 12'h6cd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23245; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1741 = io_valid_in ? _GEN_26317 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1741 = 12'h6cd == _T_2[11:0] ? image_1741 : _GEN_1740; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4814 = 12'h6ce == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7886 = 12'h6ce == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4814; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10958 = 12'h6ce == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7886; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14030 = 12'h6ce == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10958; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17102 = 12'h6ce == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14030; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20174 = 12'h6ce == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17102; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23246 = 12'h6ce == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20174; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26318 = 12'h6ce == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23246; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1742 = io_valid_in ? _GEN_26318 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1742 = 12'h6ce == _T_2[11:0] ? image_1742 : _GEN_1741; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4815 = 12'h6cf == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7887 = 12'h6cf == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4815; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10959 = 12'h6cf == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7887; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14031 = 12'h6cf == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10959; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17103 = 12'h6cf == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14031; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20175 = 12'h6cf == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17103; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23247 = 12'h6cf == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20175; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26319 = 12'h6cf == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23247; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1743 = io_valid_in ? _GEN_26319 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1743 = 12'h6cf == _T_2[11:0] ? image_1743 : _GEN_1742; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4816 = 12'h6d0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7888 = 12'h6d0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4816; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10960 = 12'h6d0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7888; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14032 = 12'h6d0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10960; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17104 = 12'h6d0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14032; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20176 = 12'h6d0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17104; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23248 = 12'h6d0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20176; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26320 = 12'h6d0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23248; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1744 = io_valid_in ? _GEN_26320 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1744 = 12'h6d0 == _T_2[11:0] ? image_1744 : _GEN_1743; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4817 = 12'h6d1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7889 = 12'h6d1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4817; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10961 = 12'h6d1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7889; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14033 = 12'h6d1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10961; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17105 = 12'h6d1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14033; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20177 = 12'h6d1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17105; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23249 = 12'h6d1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20177; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26321 = 12'h6d1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23249; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1745 = io_valid_in ? _GEN_26321 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1745 = 12'h6d1 == _T_2[11:0] ? image_1745 : _GEN_1744; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4818 = 12'h6d2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7890 = 12'h6d2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4818; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10962 = 12'h6d2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7890; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14034 = 12'h6d2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10962; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17106 = 12'h6d2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14034; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20178 = 12'h6d2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17106; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23250 = 12'h6d2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20178; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26322 = 12'h6d2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23250; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1746 = io_valid_in ? _GEN_26322 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1746 = 12'h6d2 == _T_2[11:0] ? image_1746 : _GEN_1745; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4819 = 12'h6d3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7891 = 12'h6d3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4819; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10963 = 12'h6d3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7891; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14035 = 12'h6d3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10963; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17107 = 12'h6d3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14035; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20179 = 12'h6d3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17107; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23251 = 12'h6d3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20179; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26323 = 12'h6d3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23251; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1747 = io_valid_in ? _GEN_26323 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1747 = 12'h6d3 == _T_2[11:0] ? image_1747 : _GEN_1746; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4820 = 12'h6d4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7892 = 12'h6d4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4820; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10964 = 12'h6d4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7892; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14036 = 12'h6d4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10964; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17108 = 12'h6d4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14036; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20180 = 12'h6d4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17108; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23252 = 12'h6d4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20180; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26324 = 12'h6d4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23252; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1748 = io_valid_in ? _GEN_26324 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1748 = 12'h6d4 == _T_2[11:0] ? image_1748 : _GEN_1747; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4821 = 12'h6d5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7893 = 12'h6d5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4821; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10965 = 12'h6d5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7893; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14037 = 12'h6d5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10965; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17109 = 12'h6d5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14037; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20181 = 12'h6d5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17109; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23253 = 12'h6d5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20181; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26325 = 12'h6d5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23253; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1749 = io_valid_in ? _GEN_26325 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1749 = 12'h6d5 == _T_2[11:0] ? image_1749 : _GEN_1748; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4822 = 12'h6d6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7894 = 12'h6d6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4822; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10966 = 12'h6d6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7894; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14038 = 12'h6d6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10966; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17110 = 12'h6d6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14038; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20182 = 12'h6d6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17110; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23254 = 12'h6d6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20182; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26326 = 12'h6d6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23254; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1750 = io_valid_in ? _GEN_26326 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1750 = 12'h6d6 == _T_2[11:0] ? image_1750 : _GEN_1749; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4823 = 12'h6d7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7895 = 12'h6d7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4823; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10967 = 12'h6d7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7895; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14039 = 12'h6d7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10967; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17111 = 12'h6d7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14039; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20183 = 12'h6d7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17111; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23255 = 12'h6d7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20183; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26327 = 12'h6d7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23255; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1751 = io_valid_in ? _GEN_26327 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1751 = 12'h6d7 == _T_2[11:0] ? image_1751 : _GEN_1750; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4824 = 12'h6d8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7896 = 12'h6d8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4824; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10968 = 12'h6d8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7896; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14040 = 12'h6d8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10968; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17112 = 12'h6d8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14040; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20184 = 12'h6d8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17112; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23256 = 12'h6d8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20184; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26328 = 12'h6d8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23256; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1752 = io_valid_in ? _GEN_26328 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1752 = 12'h6d8 == _T_2[11:0] ? image_1752 : _GEN_1751; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4825 = 12'h6d9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7897 = 12'h6d9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4825; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10969 = 12'h6d9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7897; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14041 = 12'h6d9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10969; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17113 = 12'h6d9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14041; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20185 = 12'h6d9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17113; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23257 = 12'h6d9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20185; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26329 = 12'h6d9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23257; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1753 = io_valid_in ? _GEN_26329 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1753 = 12'h6d9 == _T_2[11:0] ? image_1753 : _GEN_1752; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4826 = 12'h6da == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7898 = 12'h6da == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4826; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10970 = 12'h6da == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7898; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14042 = 12'h6da == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10970; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17114 = 12'h6da == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14042; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20186 = 12'h6da == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17114; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23258 = 12'h6da == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20186; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26330 = 12'h6da == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23258; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1754 = io_valid_in ? _GEN_26330 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1754 = 12'h6da == _T_2[11:0] ? image_1754 : _GEN_1753; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4827 = 12'h6db == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7899 = 12'h6db == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4827; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10971 = 12'h6db == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7899; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14043 = 12'h6db == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10971; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17115 = 12'h6db == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14043; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20187 = 12'h6db == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17115; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23259 = 12'h6db == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20187; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26331 = 12'h6db == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23259; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1755 = io_valid_in ? _GEN_26331 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1755 = 12'h6db == _T_2[11:0] ? image_1755 : _GEN_1754; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4828 = 12'h6dc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7900 = 12'h6dc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4828; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10972 = 12'h6dc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7900; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14044 = 12'h6dc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10972; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17116 = 12'h6dc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14044; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20188 = 12'h6dc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17116; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23260 = 12'h6dc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20188; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26332 = 12'h6dc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23260; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1756 = io_valid_in ? _GEN_26332 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1756 = 12'h6dc == _T_2[11:0] ? image_1756 : _GEN_1755; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4829 = 12'h6dd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7901 = 12'h6dd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4829; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10973 = 12'h6dd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7901; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14045 = 12'h6dd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10973; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17117 = 12'h6dd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14045; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20189 = 12'h6dd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17117; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23261 = 12'h6dd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20189; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26333 = 12'h6dd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23261; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1757 = io_valid_in ? _GEN_26333 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1757 = 12'h6dd == _T_2[11:0] ? image_1757 : _GEN_1756; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4830 = 12'h6de == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7902 = 12'h6de == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4830; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10974 = 12'h6de == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7902; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14046 = 12'h6de == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10974; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17118 = 12'h6de == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14046; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20190 = 12'h6de == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17118; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23262 = 12'h6de == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20190; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26334 = 12'h6de == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23262; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1758 = io_valid_in ? _GEN_26334 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1758 = 12'h6de == _T_2[11:0] ? image_1758 : _GEN_1757; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4831 = 12'h6df == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7903 = 12'h6df == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4831; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10975 = 12'h6df == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7903; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14047 = 12'h6df == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10975; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17119 = 12'h6df == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14047; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20191 = 12'h6df == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17119; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23263 = 12'h6df == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20191; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26335 = 12'h6df == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23263; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1759 = io_valid_in ? _GEN_26335 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1759 = 12'h6df == _T_2[11:0] ? image_1759 : _GEN_1758; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4832 = 12'h6e0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7904 = 12'h6e0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4832; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10976 = 12'h6e0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7904; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14048 = 12'h6e0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10976; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17120 = 12'h6e0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14048; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20192 = 12'h6e0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17120; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23264 = 12'h6e0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20192; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26336 = 12'h6e0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23264; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1760 = io_valid_in ? _GEN_26336 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1760 = 12'h6e0 == _T_2[11:0] ? image_1760 : _GEN_1759; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4833 = 12'h6e1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7905 = 12'h6e1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4833; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10977 = 12'h6e1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7905; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14049 = 12'h6e1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10977; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17121 = 12'h6e1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14049; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20193 = 12'h6e1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17121; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23265 = 12'h6e1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20193; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26337 = 12'h6e1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23265; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1761 = io_valid_in ? _GEN_26337 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1761 = 12'h6e1 == _T_2[11:0] ? image_1761 : _GEN_1760; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4834 = 12'h6e2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7906 = 12'h6e2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4834; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10978 = 12'h6e2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7906; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14050 = 12'h6e2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10978; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17122 = 12'h6e2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14050; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20194 = 12'h6e2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17122; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23266 = 12'h6e2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20194; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26338 = 12'h6e2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23266; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1762 = io_valid_in ? _GEN_26338 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1762 = 12'h6e2 == _T_2[11:0] ? image_1762 : _GEN_1761; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4835 = 12'h6e3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7907 = 12'h6e3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4835; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10979 = 12'h6e3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7907; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14051 = 12'h6e3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10979; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17123 = 12'h6e3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14051; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20195 = 12'h6e3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17123; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23267 = 12'h6e3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20195; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26339 = 12'h6e3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23267; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1763 = io_valid_in ? _GEN_26339 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1763 = 12'h6e3 == _T_2[11:0] ? image_1763 : _GEN_1762; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4836 = 12'h6e4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7908 = 12'h6e4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4836; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10980 = 12'h6e4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7908; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14052 = 12'h6e4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10980; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17124 = 12'h6e4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14052; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20196 = 12'h6e4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17124; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23268 = 12'h6e4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20196; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26340 = 12'h6e4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23268; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1764 = io_valid_in ? _GEN_26340 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1764 = 12'h6e4 == _T_2[11:0] ? image_1764 : _GEN_1763; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4837 = 12'h6e5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7909 = 12'h6e5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4837; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10981 = 12'h6e5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7909; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14053 = 12'h6e5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10981; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17125 = 12'h6e5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14053; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20197 = 12'h6e5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17125; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23269 = 12'h6e5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20197; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26341 = 12'h6e5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23269; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1765 = io_valid_in ? _GEN_26341 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1765 = 12'h6e5 == _T_2[11:0] ? image_1765 : _GEN_1764; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4838 = 12'h6e6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7910 = 12'h6e6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4838; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10982 = 12'h6e6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7910; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14054 = 12'h6e6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10982; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17126 = 12'h6e6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14054; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20198 = 12'h6e6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17126; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23270 = 12'h6e6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20198; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26342 = 12'h6e6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23270; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1766 = io_valid_in ? _GEN_26342 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1766 = 12'h6e6 == _T_2[11:0] ? image_1766 : _GEN_1765; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4839 = 12'h6e7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7911 = 12'h6e7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4839; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10983 = 12'h6e7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7911; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14055 = 12'h6e7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10983; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17127 = 12'h6e7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14055; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20199 = 12'h6e7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17127; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23271 = 12'h6e7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20199; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26343 = 12'h6e7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23271; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1767 = io_valid_in ? _GEN_26343 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1767 = 12'h6e7 == _T_2[11:0] ? image_1767 : _GEN_1766; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4840 = 12'h6e8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7912 = 12'h6e8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4840; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10984 = 12'h6e8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7912; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14056 = 12'h6e8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10984; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17128 = 12'h6e8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14056; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20200 = 12'h6e8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17128; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23272 = 12'h6e8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20200; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26344 = 12'h6e8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23272; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1768 = io_valid_in ? _GEN_26344 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1768 = 12'h6e8 == _T_2[11:0] ? image_1768 : _GEN_1767; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4841 = 12'h6e9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7913 = 12'h6e9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4841; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10985 = 12'h6e9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7913; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14057 = 12'h6e9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10985; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17129 = 12'h6e9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14057; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20201 = 12'h6e9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17129; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23273 = 12'h6e9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20201; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26345 = 12'h6e9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23273; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1769 = io_valid_in ? _GEN_26345 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1769 = 12'h6e9 == _T_2[11:0] ? image_1769 : _GEN_1768; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4842 = 12'h6ea == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7914 = 12'h6ea == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4842; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10986 = 12'h6ea == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7914; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14058 = 12'h6ea == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10986; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17130 = 12'h6ea == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14058; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20202 = 12'h6ea == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17130; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23274 = 12'h6ea == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20202; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26346 = 12'h6ea == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23274; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1770 = io_valid_in ? _GEN_26346 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1770 = 12'h6ea == _T_2[11:0] ? image_1770 : _GEN_1769; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4843 = 12'h6eb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7915 = 12'h6eb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4843; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10987 = 12'h6eb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7915; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14059 = 12'h6eb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10987; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17131 = 12'h6eb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14059; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20203 = 12'h6eb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17131; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23275 = 12'h6eb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20203; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26347 = 12'h6eb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23275; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1771 = io_valid_in ? _GEN_26347 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1771 = 12'h6eb == _T_2[11:0] ? image_1771 : _GEN_1770; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4844 = 12'h6ec == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7916 = 12'h6ec == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4844; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10988 = 12'h6ec == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7916; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14060 = 12'h6ec == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10988; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17132 = 12'h6ec == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14060; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20204 = 12'h6ec == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17132; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23276 = 12'h6ec == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20204; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26348 = 12'h6ec == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23276; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1772 = io_valid_in ? _GEN_26348 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1772 = 12'h6ec == _T_2[11:0] ? image_1772 : _GEN_1771; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4845 = 12'h6ed == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7917 = 12'h6ed == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4845; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10989 = 12'h6ed == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7917; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14061 = 12'h6ed == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10989; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17133 = 12'h6ed == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14061; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20205 = 12'h6ed == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17133; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23277 = 12'h6ed == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20205; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26349 = 12'h6ed == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23277; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1773 = io_valid_in ? _GEN_26349 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1773 = 12'h6ed == _T_2[11:0] ? image_1773 : _GEN_1772; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4846 = 12'h6ee == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7918 = 12'h6ee == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4846; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10990 = 12'h6ee == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7918; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14062 = 12'h6ee == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10990; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17134 = 12'h6ee == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14062; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20206 = 12'h6ee == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17134; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23278 = 12'h6ee == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20206; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26350 = 12'h6ee == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23278; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1774 = io_valid_in ? _GEN_26350 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1774 = 12'h6ee == _T_2[11:0] ? image_1774 : _GEN_1773; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4847 = 12'h6ef == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7919 = 12'h6ef == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4847; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10991 = 12'h6ef == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7919; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14063 = 12'h6ef == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10991; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17135 = 12'h6ef == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14063; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20207 = 12'h6ef == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17135; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23279 = 12'h6ef == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20207; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26351 = 12'h6ef == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23279; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1775 = io_valid_in ? _GEN_26351 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1775 = 12'h6ef == _T_2[11:0] ? image_1775 : _GEN_1774; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4848 = 12'h6f0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7920 = 12'h6f0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4848; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10992 = 12'h6f0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7920; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14064 = 12'h6f0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10992; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17136 = 12'h6f0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14064; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20208 = 12'h6f0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17136; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23280 = 12'h6f0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20208; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26352 = 12'h6f0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23280; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1776 = io_valid_in ? _GEN_26352 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1776 = 12'h6f0 == _T_2[11:0] ? image_1776 : _GEN_1775; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4849 = 12'h6f1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7921 = 12'h6f1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4849; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10993 = 12'h6f1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7921; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14065 = 12'h6f1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10993; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17137 = 12'h6f1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14065; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20209 = 12'h6f1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17137; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23281 = 12'h6f1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20209; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26353 = 12'h6f1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23281; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1777 = io_valid_in ? _GEN_26353 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1777 = 12'h6f1 == _T_2[11:0] ? image_1777 : _GEN_1776; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4850 = 12'h6f2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7922 = 12'h6f2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4850; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10994 = 12'h6f2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7922; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14066 = 12'h6f2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10994; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17138 = 12'h6f2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14066; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20210 = 12'h6f2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17138; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23282 = 12'h6f2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20210; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26354 = 12'h6f2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23282; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1778 = io_valid_in ? _GEN_26354 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1778 = 12'h6f2 == _T_2[11:0] ? image_1778 : _GEN_1777; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4851 = 12'h6f3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7923 = 12'h6f3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4851; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10995 = 12'h6f3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7923; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14067 = 12'h6f3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10995; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17139 = 12'h6f3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14067; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20211 = 12'h6f3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17139; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23283 = 12'h6f3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20211; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26355 = 12'h6f3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23283; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1779 = io_valid_in ? _GEN_26355 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1779 = 12'h6f3 == _T_2[11:0] ? image_1779 : _GEN_1778; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4852 = 12'h6f4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7924 = 12'h6f4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4852; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10996 = 12'h6f4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7924; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14068 = 12'h6f4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10996; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17140 = 12'h6f4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14068; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20212 = 12'h6f4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17140; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23284 = 12'h6f4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20212; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26356 = 12'h6f4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23284; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1780 = io_valid_in ? _GEN_26356 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1780 = 12'h6f4 == _T_2[11:0] ? image_1780 : _GEN_1779; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4853 = 12'h6f5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7925 = 12'h6f5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4853; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10997 = 12'h6f5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7925; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14069 = 12'h6f5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10997; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17141 = 12'h6f5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14069; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20213 = 12'h6f5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17141; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23285 = 12'h6f5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20213; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26357 = 12'h6f5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23285; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1781 = io_valid_in ? _GEN_26357 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1781 = 12'h6f5 == _T_2[11:0] ? image_1781 : _GEN_1780; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4854 = 12'h6f6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7926 = 12'h6f6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4854; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10998 = 12'h6f6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7926; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14070 = 12'h6f6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10998; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17142 = 12'h6f6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14070; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20214 = 12'h6f6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17142; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23286 = 12'h6f6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20214; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26358 = 12'h6f6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23286; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1782 = io_valid_in ? _GEN_26358 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1782 = 12'h6f6 == _T_2[11:0] ? image_1782 : _GEN_1781; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4855 = 12'h6f7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7927 = 12'h6f7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4855; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_10999 = 12'h6f7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7927; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14071 = 12'h6f7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_10999; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17143 = 12'h6f7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14071; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20215 = 12'h6f7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17143; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23287 = 12'h6f7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20215; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26359 = 12'h6f7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23287; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1783 = io_valid_in ? _GEN_26359 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1783 = 12'h6f7 == _T_2[11:0] ? image_1783 : _GEN_1782; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4856 = 12'h6f8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7928 = 12'h6f8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4856; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11000 = 12'h6f8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7928; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14072 = 12'h6f8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11000; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17144 = 12'h6f8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14072; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20216 = 12'h6f8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17144; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23288 = 12'h6f8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20216; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26360 = 12'h6f8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23288; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1784 = io_valid_in ? _GEN_26360 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1784 = 12'h6f8 == _T_2[11:0] ? image_1784 : _GEN_1783; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4857 = 12'h6f9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7929 = 12'h6f9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4857; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11001 = 12'h6f9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7929; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14073 = 12'h6f9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11001; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17145 = 12'h6f9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14073; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20217 = 12'h6f9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17145; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23289 = 12'h6f9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20217; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26361 = 12'h6f9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23289; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1785 = io_valid_in ? _GEN_26361 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1785 = 12'h6f9 == _T_2[11:0] ? image_1785 : _GEN_1784; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4858 = 12'h6fa == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7930 = 12'h6fa == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4858; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11002 = 12'h6fa == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7930; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14074 = 12'h6fa == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11002; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17146 = 12'h6fa == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14074; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20218 = 12'h6fa == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17146; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23290 = 12'h6fa == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20218; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26362 = 12'h6fa == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23290; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1786 = io_valid_in ? _GEN_26362 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1786 = 12'h6fa == _T_2[11:0] ? image_1786 : _GEN_1785; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4859 = 12'h6fb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7931 = 12'h6fb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4859; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11003 = 12'h6fb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7931; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14075 = 12'h6fb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11003; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17147 = 12'h6fb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14075; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20219 = 12'h6fb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17147; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23291 = 12'h6fb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20219; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26363 = 12'h6fb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23291; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1787 = io_valid_in ? _GEN_26363 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1787 = 12'h6fb == _T_2[11:0] ? image_1787 : _GEN_1786; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4860 = 12'h6fc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7932 = 12'h6fc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4860; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11004 = 12'h6fc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7932; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14076 = 12'h6fc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11004; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17148 = 12'h6fc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14076; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20220 = 12'h6fc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17148; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23292 = 12'h6fc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20220; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26364 = 12'h6fc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23292; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1788 = io_valid_in ? _GEN_26364 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1788 = 12'h6fc == _T_2[11:0] ? image_1788 : _GEN_1787; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4861 = 12'h6fd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7933 = 12'h6fd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4861; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11005 = 12'h6fd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7933; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14077 = 12'h6fd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11005; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17149 = 12'h6fd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14077; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20221 = 12'h6fd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17149; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23293 = 12'h6fd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20221; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26365 = 12'h6fd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23293; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1789 = io_valid_in ? _GEN_26365 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1789 = 12'h6fd == _T_2[11:0] ? image_1789 : _GEN_1788; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4862 = 12'h6fe == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7934 = 12'h6fe == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4862; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11006 = 12'h6fe == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7934; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14078 = 12'h6fe == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11006; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17150 = 12'h6fe == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14078; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20222 = 12'h6fe == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17150; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23294 = 12'h6fe == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20222; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26366 = 12'h6fe == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23294; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1790 = io_valid_in ? _GEN_26366 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1790 = 12'h6fe == _T_2[11:0] ? image_1790 : _GEN_1789; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4863 = 12'h6ff == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7935 = 12'h6ff == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4863; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11007 = 12'h6ff == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7935; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14079 = 12'h6ff == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11007; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17151 = 12'h6ff == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14079; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20223 = 12'h6ff == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17151; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23295 = 12'h6ff == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20223; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26367 = 12'h6ff == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23295; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1791 = io_valid_in ? _GEN_26367 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1791 = 12'h6ff == _T_2[11:0] ? image_1791 : _GEN_1790; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4864 = 12'h700 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7936 = 12'h700 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4864; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11008 = 12'h700 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7936; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14080 = 12'h700 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11008; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17152 = 12'h700 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14080; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20224 = 12'h700 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17152; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23296 = 12'h700 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20224; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26368 = 12'h700 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23296; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1792 = io_valid_in ? _GEN_26368 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1792 = 12'h700 == _T_2[11:0] ? image_1792 : _GEN_1791; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4865 = 12'h701 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7937 = 12'h701 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4865; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11009 = 12'h701 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7937; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14081 = 12'h701 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11009; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17153 = 12'h701 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14081; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20225 = 12'h701 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17153; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23297 = 12'h701 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20225; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26369 = 12'h701 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23297; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1793 = io_valid_in ? _GEN_26369 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1793 = 12'h701 == _T_2[11:0] ? image_1793 : _GEN_1792; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4866 = 12'h702 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7938 = 12'h702 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4866; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11010 = 12'h702 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7938; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14082 = 12'h702 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11010; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17154 = 12'h702 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14082; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20226 = 12'h702 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17154; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23298 = 12'h702 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20226; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26370 = 12'h702 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23298; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1794 = io_valid_in ? _GEN_26370 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1794 = 12'h702 == _T_2[11:0] ? image_1794 : _GEN_1793; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4867 = 12'h703 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7939 = 12'h703 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4867; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11011 = 12'h703 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7939; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14083 = 12'h703 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11011; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17155 = 12'h703 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14083; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20227 = 12'h703 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17155; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23299 = 12'h703 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20227; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26371 = 12'h703 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23299; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1795 = io_valid_in ? _GEN_26371 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1795 = 12'h703 == _T_2[11:0] ? image_1795 : _GEN_1794; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4868 = 12'h704 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7940 = 12'h704 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4868; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11012 = 12'h704 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7940; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14084 = 12'h704 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11012; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17156 = 12'h704 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14084; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20228 = 12'h704 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17156; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23300 = 12'h704 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20228; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26372 = 12'h704 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23300; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1796 = io_valid_in ? _GEN_26372 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1796 = 12'h704 == _T_2[11:0] ? image_1796 : _GEN_1795; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4869 = 12'h705 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7941 = 12'h705 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4869; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11013 = 12'h705 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7941; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14085 = 12'h705 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11013; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17157 = 12'h705 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14085; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20229 = 12'h705 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17157; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23301 = 12'h705 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20229; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26373 = 12'h705 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23301; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1797 = io_valid_in ? _GEN_26373 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1797 = 12'h705 == _T_2[11:0] ? image_1797 : _GEN_1796; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4870 = 12'h706 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7942 = 12'h706 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4870; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11014 = 12'h706 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7942; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14086 = 12'h706 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11014; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17158 = 12'h706 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14086; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20230 = 12'h706 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17158; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23302 = 12'h706 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20230; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26374 = 12'h706 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23302; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1798 = io_valid_in ? _GEN_26374 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1798 = 12'h706 == _T_2[11:0] ? image_1798 : _GEN_1797; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4871 = 12'h707 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7943 = 12'h707 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4871; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11015 = 12'h707 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7943; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14087 = 12'h707 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11015; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17159 = 12'h707 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14087; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20231 = 12'h707 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17159; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23303 = 12'h707 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20231; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26375 = 12'h707 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23303; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1799 = io_valid_in ? _GEN_26375 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1799 = 12'h707 == _T_2[11:0] ? image_1799 : _GEN_1798; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4872 = 12'h708 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7944 = 12'h708 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4872; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11016 = 12'h708 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7944; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14088 = 12'h708 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11016; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17160 = 12'h708 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14088; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20232 = 12'h708 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17160; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23304 = 12'h708 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20232; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26376 = 12'h708 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23304; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1800 = io_valid_in ? _GEN_26376 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1800 = 12'h708 == _T_2[11:0] ? image_1800 : _GEN_1799; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4873 = 12'h709 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7945 = 12'h709 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4873; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11017 = 12'h709 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7945; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14089 = 12'h709 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11017; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17161 = 12'h709 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14089; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20233 = 12'h709 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17161; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23305 = 12'h709 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20233; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26377 = 12'h709 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23305; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1801 = io_valid_in ? _GEN_26377 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1801 = 12'h709 == _T_2[11:0] ? image_1801 : _GEN_1800; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4874 = 12'h70a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7946 = 12'h70a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4874; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11018 = 12'h70a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7946; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14090 = 12'h70a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11018; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17162 = 12'h70a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14090; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20234 = 12'h70a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17162; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23306 = 12'h70a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20234; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26378 = 12'h70a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23306; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1802 = io_valid_in ? _GEN_26378 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1802 = 12'h70a == _T_2[11:0] ? image_1802 : _GEN_1801; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4875 = 12'h70b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7947 = 12'h70b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4875; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11019 = 12'h70b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7947; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14091 = 12'h70b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11019; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17163 = 12'h70b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14091; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20235 = 12'h70b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17163; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23307 = 12'h70b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20235; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26379 = 12'h70b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23307; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1803 = io_valid_in ? _GEN_26379 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1803 = 12'h70b == _T_2[11:0] ? image_1803 : _GEN_1802; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4876 = 12'h70c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7948 = 12'h70c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4876; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11020 = 12'h70c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7948; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14092 = 12'h70c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11020; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17164 = 12'h70c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14092; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20236 = 12'h70c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17164; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23308 = 12'h70c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20236; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26380 = 12'h70c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23308; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1804 = io_valid_in ? _GEN_26380 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1804 = 12'h70c == _T_2[11:0] ? image_1804 : _GEN_1803; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4877 = 12'h70d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7949 = 12'h70d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4877; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11021 = 12'h70d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7949; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14093 = 12'h70d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11021; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17165 = 12'h70d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14093; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20237 = 12'h70d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17165; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23309 = 12'h70d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20237; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26381 = 12'h70d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23309; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1805 = io_valid_in ? _GEN_26381 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1805 = 12'h70d == _T_2[11:0] ? image_1805 : _GEN_1804; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4878 = 12'h70e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7950 = 12'h70e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4878; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11022 = 12'h70e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7950; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14094 = 12'h70e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11022; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17166 = 12'h70e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14094; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20238 = 12'h70e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17166; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23310 = 12'h70e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20238; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26382 = 12'h70e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23310; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1806 = io_valid_in ? _GEN_26382 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1806 = 12'h70e == _T_2[11:0] ? image_1806 : _GEN_1805; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4879 = 12'h70f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7951 = 12'h70f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4879; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11023 = 12'h70f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7951; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14095 = 12'h70f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11023; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17167 = 12'h70f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14095; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20239 = 12'h70f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17167; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23311 = 12'h70f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20239; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26383 = 12'h70f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23311; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1807 = io_valid_in ? _GEN_26383 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1807 = 12'h70f == _T_2[11:0] ? image_1807 : _GEN_1806; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4880 = 12'h710 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7952 = 12'h710 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4880; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11024 = 12'h710 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7952; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14096 = 12'h710 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11024; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17168 = 12'h710 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14096; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20240 = 12'h710 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17168; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23312 = 12'h710 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20240; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26384 = 12'h710 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23312; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1808 = io_valid_in ? _GEN_26384 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1808 = 12'h710 == _T_2[11:0] ? image_1808 : _GEN_1807; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4881 = 12'h711 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7953 = 12'h711 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4881; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11025 = 12'h711 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7953; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14097 = 12'h711 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11025; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17169 = 12'h711 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14097; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20241 = 12'h711 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17169; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23313 = 12'h711 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20241; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26385 = 12'h711 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23313; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1809 = io_valid_in ? _GEN_26385 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1809 = 12'h711 == _T_2[11:0] ? image_1809 : _GEN_1808; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4882 = 12'h712 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7954 = 12'h712 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4882; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11026 = 12'h712 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7954; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14098 = 12'h712 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11026; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17170 = 12'h712 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14098; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20242 = 12'h712 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17170; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23314 = 12'h712 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20242; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26386 = 12'h712 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23314; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1810 = io_valid_in ? _GEN_26386 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1810 = 12'h712 == _T_2[11:0] ? image_1810 : _GEN_1809; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4883 = 12'h713 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7955 = 12'h713 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4883; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11027 = 12'h713 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7955; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14099 = 12'h713 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11027; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17171 = 12'h713 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14099; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20243 = 12'h713 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17171; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23315 = 12'h713 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20243; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26387 = 12'h713 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23315; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1811 = io_valid_in ? _GEN_26387 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1811 = 12'h713 == _T_2[11:0] ? image_1811 : _GEN_1810; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4884 = 12'h714 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7956 = 12'h714 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4884; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11028 = 12'h714 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7956; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14100 = 12'h714 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11028; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17172 = 12'h714 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14100; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20244 = 12'h714 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17172; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23316 = 12'h714 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20244; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26388 = 12'h714 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23316; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1812 = io_valid_in ? _GEN_26388 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1812 = 12'h714 == _T_2[11:0] ? image_1812 : _GEN_1811; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4885 = 12'h715 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7957 = 12'h715 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4885; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11029 = 12'h715 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7957; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14101 = 12'h715 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11029; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17173 = 12'h715 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14101; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20245 = 12'h715 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17173; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23317 = 12'h715 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20245; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26389 = 12'h715 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23317; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1813 = io_valid_in ? _GEN_26389 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1813 = 12'h715 == _T_2[11:0] ? image_1813 : _GEN_1812; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4886 = 12'h716 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7958 = 12'h716 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4886; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11030 = 12'h716 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7958; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14102 = 12'h716 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11030; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17174 = 12'h716 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14102; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20246 = 12'h716 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17174; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23318 = 12'h716 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20246; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26390 = 12'h716 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23318; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1814 = io_valid_in ? _GEN_26390 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1814 = 12'h716 == _T_2[11:0] ? image_1814 : _GEN_1813; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4887 = 12'h717 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7959 = 12'h717 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4887; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11031 = 12'h717 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7959; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14103 = 12'h717 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11031; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17175 = 12'h717 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14103; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20247 = 12'h717 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17175; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23319 = 12'h717 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20247; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26391 = 12'h717 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23319; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1815 = io_valid_in ? _GEN_26391 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1815 = 12'h717 == _T_2[11:0] ? image_1815 : _GEN_1814; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4888 = 12'h718 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7960 = 12'h718 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4888; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11032 = 12'h718 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7960; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14104 = 12'h718 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11032; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17176 = 12'h718 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14104; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20248 = 12'h718 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17176; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23320 = 12'h718 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20248; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26392 = 12'h718 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23320; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1816 = io_valid_in ? _GEN_26392 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1816 = 12'h718 == _T_2[11:0] ? image_1816 : _GEN_1815; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4889 = 12'h719 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7961 = 12'h719 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4889; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11033 = 12'h719 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7961; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14105 = 12'h719 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11033; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17177 = 12'h719 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14105; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20249 = 12'h719 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17177; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23321 = 12'h719 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20249; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26393 = 12'h719 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23321; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1817 = io_valid_in ? _GEN_26393 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1817 = 12'h719 == _T_2[11:0] ? image_1817 : _GEN_1816; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4890 = 12'h71a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7962 = 12'h71a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4890; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11034 = 12'h71a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7962; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14106 = 12'h71a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11034; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17178 = 12'h71a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14106; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20250 = 12'h71a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17178; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23322 = 12'h71a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20250; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26394 = 12'h71a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23322; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1818 = io_valid_in ? _GEN_26394 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1818 = 12'h71a == _T_2[11:0] ? image_1818 : _GEN_1817; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4891 = 12'h71b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7963 = 12'h71b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4891; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11035 = 12'h71b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7963; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14107 = 12'h71b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11035; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17179 = 12'h71b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14107; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20251 = 12'h71b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17179; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23323 = 12'h71b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20251; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26395 = 12'h71b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23323; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1819 = io_valid_in ? _GEN_26395 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1819 = 12'h71b == _T_2[11:0] ? image_1819 : _GEN_1818; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4892 = 12'h71c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7964 = 12'h71c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4892; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11036 = 12'h71c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7964; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14108 = 12'h71c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11036; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17180 = 12'h71c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14108; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20252 = 12'h71c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17180; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23324 = 12'h71c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20252; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26396 = 12'h71c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23324; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1820 = io_valid_in ? _GEN_26396 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1820 = 12'h71c == _T_2[11:0] ? image_1820 : _GEN_1819; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4893 = 12'h71d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7965 = 12'h71d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4893; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11037 = 12'h71d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7965; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14109 = 12'h71d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11037; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17181 = 12'h71d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14109; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20253 = 12'h71d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17181; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23325 = 12'h71d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20253; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26397 = 12'h71d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23325; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1821 = io_valid_in ? _GEN_26397 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1821 = 12'h71d == _T_2[11:0] ? image_1821 : _GEN_1820; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4894 = 12'h71e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7966 = 12'h71e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4894; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11038 = 12'h71e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7966; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14110 = 12'h71e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11038; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17182 = 12'h71e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14110; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20254 = 12'h71e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17182; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23326 = 12'h71e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20254; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26398 = 12'h71e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23326; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1822 = io_valid_in ? _GEN_26398 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1822 = 12'h71e == _T_2[11:0] ? image_1822 : _GEN_1821; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4895 = 12'h71f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7967 = 12'h71f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4895; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11039 = 12'h71f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7967; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14111 = 12'h71f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11039; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17183 = 12'h71f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14111; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20255 = 12'h71f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17183; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23327 = 12'h71f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20255; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26399 = 12'h71f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23327; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1823 = io_valid_in ? _GEN_26399 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1823 = 12'h71f == _T_2[11:0] ? image_1823 : _GEN_1822; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4896 = 12'h720 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7968 = 12'h720 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4896; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11040 = 12'h720 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7968; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14112 = 12'h720 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11040; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17184 = 12'h720 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14112; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20256 = 12'h720 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17184; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23328 = 12'h720 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20256; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26400 = 12'h720 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23328; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1824 = io_valid_in ? _GEN_26400 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1824 = 12'h720 == _T_2[11:0] ? image_1824 : _GEN_1823; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4897 = 12'h721 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7969 = 12'h721 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4897; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11041 = 12'h721 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7969; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14113 = 12'h721 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11041; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17185 = 12'h721 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14113; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20257 = 12'h721 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17185; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23329 = 12'h721 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20257; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26401 = 12'h721 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23329; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1825 = io_valid_in ? _GEN_26401 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1825 = 12'h721 == _T_2[11:0] ? image_1825 : _GEN_1824; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4898 = 12'h722 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7970 = 12'h722 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4898; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11042 = 12'h722 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7970; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14114 = 12'h722 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11042; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17186 = 12'h722 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14114; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20258 = 12'h722 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17186; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23330 = 12'h722 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20258; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26402 = 12'h722 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23330; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1826 = io_valid_in ? _GEN_26402 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1826 = 12'h722 == _T_2[11:0] ? image_1826 : _GEN_1825; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4899 = 12'h723 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7971 = 12'h723 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4899; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11043 = 12'h723 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7971; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14115 = 12'h723 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11043; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17187 = 12'h723 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14115; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20259 = 12'h723 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17187; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23331 = 12'h723 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20259; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26403 = 12'h723 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23331; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1827 = io_valid_in ? _GEN_26403 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1827 = 12'h723 == _T_2[11:0] ? image_1827 : _GEN_1826; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4900 = 12'h724 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7972 = 12'h724 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4900; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11044 = 12'h724 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7972; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14116 = 12'h724 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11044; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17188 = 12'h724 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14116; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20260 = 12'h724 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17188; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23332 = 12'h724 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20260; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26404 = 12'h724 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23332; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1828 = io_valid_in ? _GEN_26404 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1828 = 12'h724 == _T_2[11:0] ? image_1828 : _GEN_1827; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4901 = 12'h725 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7973 = 12'h725 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4901; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11045 = 12'h725 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7973; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14117 = 12'h725 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11045; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17189 = 12'h725 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14117; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20261 = 12'h725 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17189; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23333 = 12'h725 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20261; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26405 = 12'h725 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23333; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1829 = io_valid_in ? _GEN_26405 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1829 = 12'h725 == _T_2[11:0] ? image_1829 : _GEN_1828; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4902 = 12'h726 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7974 = 12'h726 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4902; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11046 = 12'h726 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7974; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14118 = 12'h726 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11046; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17190 = 12'h726 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14118; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20262 = 12'h726 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17190; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23334 = 12'h726 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20262; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26406 = 12'h726 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23334; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1830 = io_valid_in ? _GEN_26406 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1830 = 12'h726 == _T_2[11:0] ? image_1830 : _GEN_1829; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4903 = 12'h727 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7975 = 12'h727 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4903; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11047 = 12'h727 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7975; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14119 = 12'h727 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11047; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17191 = 12'h727 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14119; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20263 = 12'h727 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17191; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23335 = 12'h727 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20263; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26407 = 12'h727 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23335; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1831 = io_valid_in ? _GEN_26407 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1831 = 12'h727 == _T_2[11:0] ? image_1831 : _GEN_1830; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4904 = 12'h728 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7976 = 12'h728 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4904; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11048 = 12'h728 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7976; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14120 = 12'h728 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11048; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17192 = 12'h728 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14120; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20264 = 12'h728 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17192; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23336 = 12'h728 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20264; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26408 = 12'h728 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23336; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1832 = io_valid_in ? _GEN_26408 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1832 = 12'h728 == _T_2[11:0] ? image_1832 : _GEN_1831; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4905 = 12'h729 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7977 = 12'h729 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4905; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11049 = 12'h729 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7977; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14121 = 12'h729 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11049; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17193 = 12'h729 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14121; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20265 = 12'h729 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17193; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23337 = 12'h729 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20265; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26409 = 12'h729 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23337; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1833 = io_valid_in ? _GEN_26409 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1833 = 12'h729 == _T_2[11:0] ? image_1833 : _GEN_1832; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4906 = 12'h72a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7978 = 12'h72a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4906; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11050 = 12'h72a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7978; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14122 = 12'h72a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11050; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17194 = 12'h72a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14122; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20266 = 12'h72a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17194; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23338 = 12'h72a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20266; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26410 = 12'h72a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23338; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1834 = io_valid_in ? _GEN_26410 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1834 = 12'h72a == _T_2[11:0] ? image_1834 : _GEN_1833; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4907 = 12'h72b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7979 = 12'h72b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4907; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11051 = 12'h72b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7979; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14123 = 12'h72b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11051; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17195 = 12'h72b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14123; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20267 = 12'h72b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17195; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23339 = 12'h72b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20267; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26411 = 12'h72b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23339; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1835 = io_valid_in ? _GEN_26411 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1835 = 12'h72b == _T_2[11:0] ? image_1835 : _GEN_1834; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4908 = 12'h72c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7980 = 12'h72c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4908; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11052 = 12'h72c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7980; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14124 = 12'h72c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11052; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17196 = 12'h72c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14124; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20268 = 12'h72c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17196; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23340 = 12'h72c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20268; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26412 = 12'h72c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23340; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1836 = io_valid_in ? _GEN_26412 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1836 = 12'h72c == _T_2[11:0] ? image_1836 : _GEN_1835; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4909 = 12'h72d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7981 = 12'h72d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4909; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11053 = 12'h72d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7981; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14125 = 12'h72d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11053; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17197 = 12'h72d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14125; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20269 = 12'h72d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17197; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23341 = 12'h72d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20269; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26413 = 12'h72d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23341; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1837 = io_valid_in ? _GEN_26413 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1837 = 12'h72d == _T_2[11:0] ? image_1837 : _GEN_1836; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4910 = 12'h72e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7982 = 12'h72e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4910; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11054 = 12'h72e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7982; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14126 = 12'h72e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11054; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17198 = 12'h72e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14126; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20270 = 12'h72e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17198; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23342 = 12'h72e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20270; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26414 = 12'h72e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23342; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1838 = io_valid_in ? _GEN_26414 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1838 = 12'h72e == _T_2[11:0] ? image_1838 : _GEN_1837; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4911 = 12'h72f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7983 = 12'h72f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4911; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11055 = 12'h72f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7983; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14127 = 12'h72f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11055; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17199 = 12'h72f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14127; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20271 = 12'h72f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17199; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23343 = 12'h72f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20271; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26415 = 12'h72f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23343; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1839 = io_valid_in ? _GEN_26415 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1839 = 12'h72f == _T_2[11:0] ? image_1839 : _GEN_1838; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4912 = 12'h730 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7984 = 12'h730 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4912; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11056 = 12'h730 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7984; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14128 = 12'h730 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11056; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17200 = 12'h730 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14128; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20272 = 12'h730 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17200; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23344 = 12'h730 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20272; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26416 = 12'h730 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23344; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1840 = io_valid_in ? _GEN_26416 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1840 = 12'h730 == _T_2[11:0] ? image_1840 : _GEN_1839; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4913 = 12'h731 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7985 = 12'h731 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4913; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11057 = 12'h731 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7985; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14129 = 12'h731 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11057; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17201 = 12'h731 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14129; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20273 = 12'h731 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17201; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23345 = 12'h731 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20273; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26417 = 12'h731 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23345; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1841 = io_valid_in ? _GEN_26417 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1841 = 12'h731 == _T_2[11:0] ? image_1841 : _GEN_1840; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4914 = 12'h732 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7986 = 12'h732 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4914; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11058 = 12'h732 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7986; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14130 = 12'h732 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11058; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17202 = 12'h732 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14130; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20274 = 12'h732 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17202; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23346 = 12'h732 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20274; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26418 = 12'h732 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23346; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1842 = io_valid_in ? _GEN_26418 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1842 = 12'h732 == _T_2[11:0] ? image_1842 : _GEN_1841; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4915 = 12'h733 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7987 = 12'h733 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4915; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11059 = 12'h733 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7987; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14131 = 12'h733 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11059; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17203 = 12'h733 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14131; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20275 = 12'h733 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17203; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23347 = 12'h733 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20275; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26419 = 12'h733 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23347; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1843 = io_valid_in ? _GEN_26419 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1843 = 12'h733 == _T_2[11:0] ? image_1843 : _GEN_1842; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4916 = 12'h734 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7988 = 12'h734 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4916; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11060 = 12'h734 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7988; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14132 = 12'h734 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11060; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17204 = 12'h734 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14132; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20276 = 12'h734 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17204; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23348 = 12'h734 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20276; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26420 = 12'h734 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23348; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1844 = io_valid_in ? _GEN_26420 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1844 = 12'h734 == _T_2[11:0] ? image_1844 : _GEN_1843; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4917 = 12'h735 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7989 = 12'h735 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4917; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11061 = 12'h735 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7989; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14133 = 12'h735 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11061; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17205 = 12'h735 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14133; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20277 = 12'h735 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17205; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23349 = 12'h735 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20277; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26421 = 12'h735 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23349; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1845 = io_valid_in ? _GEN_26421 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1845 = 12'h735 == _T_2[11:0] ? image_1845 : _GEN_1844; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4918 = 12'h736 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7990 = 12'h736 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4918; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11062 = 12'h736 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7990; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14134 = 12'h736 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11062; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17206 = 12'h736 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14134; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20278 = 12'h736 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17206; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23350 = 12'h736 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20278; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26422 = 12'h736 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23350; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1846 = io_valid_in ? _GEN_26422 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1846 = 12'h736 == _T_2[11:0] ? image_1846 : _GEN_1845; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4919 = 12'h737 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7991 = 12'h737 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4919; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11063 = 12'h737 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7991; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14135 = 12'h737 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11063; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17207 = 12'h737 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14135; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20279 = 12'h737 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17207; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23351 = 12'h737 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20279; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26423 = 12'h737 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23351; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1847 = io_valid_in ? _GEN_26423 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1847 = 12'h737 == _T_2[11:0] ? image_1847 : _GEN_1846; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4920 = 12'h738 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7992 = 12'h738 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4920; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11064 = 12'h738 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7992; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14136 = 12'h738 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11064; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17208 = 12'h738 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14136; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20280 = 12'h738 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17208; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23352 = 12'h738 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20280; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26424 = 12'h738 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23352; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1848 = io_valid_in ? _GEN_26424 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1848 = 12'h738 == _T_2[11:0] ? image_1848 : _GEN_1847; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4921 = 12'h739 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7993 = 12'h739 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4921; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11065 = 12'h739 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7993; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14137 = 12'h739 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11065; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17209 = 12'h739 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14137; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20281 = 12'h739 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17209; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23353 = 12'h739 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20281; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26425 = 12'h739 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23353; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1849 = io_valid_in ? _GEN_26425 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1849 = 12'h739 == _T_2[11:0] ? image_1849 : _GEN_1848; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4922 = 12'h73a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7994 = 12'h73a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4922; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11066 = 12'h73a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7994; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14138 = 12'h73a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11066; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17210 = 12'h73a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14138; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20282 = 12'h73a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17210; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23354 = 12'h73a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20282; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26426 = 12'h73a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23354; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1850 = io_valid_in ? _GEN_26426 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1850 = 12'h73a == _T_2[11:0] ? image_1850 : _GEN_1849; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4923 = 12'h73b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7995 = 12'h73b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4923; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11067 = 12'h73b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7995; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14139 = 12'h73b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11067; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17211 = 12'h73b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14139; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20283 = 12'h73b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17211; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23355 = 12'h73b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20283; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26427 = 12'h73b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23355; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1851 = io_valid_in ? _GEN_26427 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1851 = 12'h73b == _T_2[11:0] ? image_1851 : _GEN_1850; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4924 = 12'h73c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7996 = 12'h73c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4924; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11068 = 12'h73c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7996; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14140 = 12'h73c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11068; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17212 = 12'h73c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14140; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20284 = 12'h73c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17212; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23356 = 12'h73c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20284; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26428 = 12'h73c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23356; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1852 = io_valid_in ? _GEN_26428 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1852 = 12'h73c == _T_2[11:0] ? image_1852 : _GEN_1851; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4925 = 12'h73d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7997 = 12'h73d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4925; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11069 = 12'h73d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7997; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14141 = 12'h73d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11069; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17213 = 12'h73d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14141; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20285 = 12'h73d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17213; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23357 = 12'h73d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20285; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26429 = 12'h73d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23357; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1853 = io_valid_in ? _GEN_26429 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1853 = 12'h73d == _T_2[11:0] ? image_1853 : _GEN_1852; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4926 = 12'h73e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7998 = 12'h73e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4926; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11070 = 12'h73e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7998; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14142 = 12'h73e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11070; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17214 = 12'h73e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14142; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20286 = 12'h73e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17214; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23358 = 12'h73e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20286; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26430 = 12'h73e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23358; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1854 = io_valid_in ? _GEN_26430 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1854 = 12'h73e == _T_2[11:0] ? image_1854 : _GEN_1853; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4927 = 12'h73f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_7999 = 12'h73f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4927; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11071 = 12'h73f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_7999; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14143 = 12'h73f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11071; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17215 = 12'h73f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14143; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20287 = 12'h73f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17215; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23359 = 12'h73f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20287; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26431 = 12'h73f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23359; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1855 = io_valid_in ? _GEN_26431 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1855 = 12'h73f == _T_2[11:0] ? image_1855 : _GEN_1854; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4928 = 12'h740 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8000 = 12'h740 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4928; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11072 = 12'h740 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8000; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14144 = 12'h740 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11072; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17216 = 12'h740 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14144; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20288 = 12'h740 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17216; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23360 = 12'h740 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20288; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26432 = 12'h740 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23360; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1856 = io_valid_in ? _GEN_26432 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1856 = 12'h740 == _T_2[11:0] ? image_1856 : _GEN_1855; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4929 = 12'h741 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8001 = 12'h741 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4929; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11073 = 12'h741 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8001; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14145 = 12'h741 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11073; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17217 = 12'h741 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14145; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20289 = 12'h741 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17217; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23361 = 12'h741 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20289; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26433 = 12'h741 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23361; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1857 = io_valid_in ? _GEN_26433 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1857 = 12'h741 == _T_2[11:0] ? image_1857 : _GEN_1856; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4930 = 12'h742 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8002 = 12'h742 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4930; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11074 = 12'h742 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8002; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14146 = 12'h742 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11074; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17218 = 12'h742 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14146; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20290 = 12'h742 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17218; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23362 = 12'h742 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20290; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26434 = 12'h742 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23362; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1858 = io_valid_in ? _GEN_26434 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1858 = 12'h742 == _T_2[11:0] ? image_1858 : _GEN_1857; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4931 = 12'h743 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8003 = 12'h743 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4931; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11075 = 12'h743 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8003; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14147 = 12'h743 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11075; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17219 = 12'h743 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14147; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20291 = 12'h743 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17219; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23363 = 12'h743 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20291; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26435 = 12'h743 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23363; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1859 = io_valid_in ? _GEN_26435 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1859 = 12'h743 == _T_2[11:0] ? image_1859 : _GEN_1858; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4932 = 12'h744 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8004 = 12'h744 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4932; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11076 = 12'h744 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8004; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14148 = 12'h744 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11076; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17220 = 12'h744 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14148; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20292 = 12'h744 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17220; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23364 = 12'h744 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20292; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26436 = 12'h744 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23364; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1860 = io_valid_in ? _GEN_26436 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1860 = 12'h744 == _T_2[11:0] ? image_1860 : _GEN_1859; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4933 = 12'h745 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8005 = 12'h745 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4933; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11077 = 12'h745 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8005; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14149 = 12'h745 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11077; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17221 = 12'h745 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14149; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20293 = 12'h745 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17221; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23365 = 12'h745 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20293; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26437 = 12'h745 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23365; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1861 = io_valid_in ? _GEN_26437 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1861 = 12'h745 == _T_2[11:0] ? image_1861 : _GEN_1860; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4934 = 12'h746 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8006 = 12'h746 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4934; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11078 = 12'h746 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8006; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14150 = 12'h746 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11078; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17222 = 12'h746 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14150; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20294 = 12'h746 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17222; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23366 = 12'h746 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20294; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26438 = 12'h746 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23366; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1862 = io_valid_in ? _GEN_26438 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1862 = 12'h746 == _T_2[11:0] ? image_1862 : _GEN_1861; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4935 = 12'h747 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8007 = 12'h747 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4935; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11079 = 12'h747 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8007; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14151 = 12'h747 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11079; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17223 = 12'h747 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14151; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20295 = 12'h747 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17223; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23367 = 12'h747 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20295; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26439 = 12'h747 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23367; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1863 = io_valid_in ? _GEN_26439 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1863 = 12'h747 == _T_2[11:0] ? image_1863 : _GEN_1862; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4936 = 12'h748 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8008 = 12'h748 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4936; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11080 = 12'h748 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8008; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14152 = 12'h748 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11080; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17224 = 12'h748 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14152; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20296 = 12'h748 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17224; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23368 = 12'h748 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20296; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26440 = 12'h748 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23368; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1864 = io_valid_in ? _GEN_26440 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1864 = 12'h748 == _T_2[11:0] ? image_1864 : _GEN_1863; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4937 = 12'h749 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8009 = 12'h749 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4937; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11081 = 12'h749 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8009; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14153 = 12'h749 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11081; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17225 = 12'h749 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14153; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20297 = 12'h749 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17225; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23369 = 12'h749 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20297; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26441 = 12'h749 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23369; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1865 = io_valid_in ? _GEN_26441 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1865 = 12'h749 == _T_2[11:0] ? image_1865 : _GEN_1864; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4938 = 12'h74a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8010 = 12'h74a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4938; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11082 = 12'h74a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8010; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14154 = 12'h74a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11082; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17226 = 12'h74a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14154; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20298 = 12'h74a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17226; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23370 = 12'h74a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20298; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26442 = 12'h74a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23370; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1866 = io_valid_in ? _GEN_26442 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1866 = 12'h74a == _T_2[11:0] ? image_1866 : _GEN_1865; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4939 = 12'h74b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8011 = 12'h74b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4939; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11083 = 12'h74b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8011; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14155 = 12'h74b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11083; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17227 = 12'h74b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14155; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20299 = 12'h74b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17227; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23371 = 12'h74b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20299; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26443 = 12'h74b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23371; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1867 = io_valid_in ? _GEN_26443 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1867 = 12'h74b == _T_2[11:0] ? image_1867 : _GEN_1866; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4940 = 12'h74c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8012 = 12'h74c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4940; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11084 = 12'h74c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8012; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14156 = 12'h74c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11084; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17228 = 12'h74c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14156; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20300 = 12'h74c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17228; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23372 = 12'h74c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20300; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26444 = 12'h74c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23372; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1868 = io_valid_in ? _GEN_26444 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1868 = 12'h74c == _T_2[11:0] ? image_1868 : _GEN_1867; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4941 = 12'h74d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8013 = 12'h74d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4941; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11085 = 12'h74d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8013; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14157 = 12'h74d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11085; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17229 = 12'h74d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14157; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20301 = 12'h74d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17229; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23373 = 12'h74d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20301; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26445 = 12'h74d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23373; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1869 = io_valid_in ? _GEN_26445 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1869 = 12'h74d == _T_2[11:0] ? image_1869 : _GEN_1868; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4942 = 12'h74e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8014 = 12'h74e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4942; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11086 = 12'h74e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8014; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14158 = 12'h74e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11086; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17230 = 12'h74e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14158; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20302 = 12'h74e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17230; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23374 = 12'h74e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20302; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26446 = 12'h74e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23374; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1870 = io_valid_in ? _GEN_26446 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1870 = 12'h74e == _T_2[11:0] ? image_1870 : _GEN_1869; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4943 = 12'h74f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8015 = 12'h74f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4943; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11087 = 12'h74f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8015; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14159 = 12'h74f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11087; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17231 = 12'h74f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14159; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20303 = 12'h74f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17231; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23375 = 12'h74f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20303; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26447 = 12'h74f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23375; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1871 = io_valid_in ? _GEN_26447 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1871 = 12'h74f == _T_2[11:0] ? image_1871 : _GEN_1870; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4944 = 12'h750 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8016 = 12'h750 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4944; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11088 = 12'h750 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8016; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14160 = 12'h750 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11088; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17232 = 12'h750 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14160; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20304 = 12'h750 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17232; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23376 = 12'h750 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20304; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26448 = 12'h750 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23376; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1872 = io_valid_in ? _GEN_26448 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1872 = 12'h750 == _T_2[11:0] ? image_1872 : _GEN_1871; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4945 = 12'h751 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8017 = 12'h751 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4945; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11089 = 12'h751 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8017; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14161 = 12'h751 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11089; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17233 = 12'h751 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14161; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20305 = 12'h751 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17233; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23377 = 12'h751 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20305; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26449 = 12'h751 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23377; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1873 = io_valid_in ? _GEN_26449 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1873 = 12'h751 == _T_2[11:0] ? image_1873 : _GEN_1872; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4946 = 12'h752 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8018 = 12'h752 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4946; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11090 = 12'h752 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8018; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14162 = 12'h752 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11090; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17234 = 12'h752 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14162; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20306 = 12'h752 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17234; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23378 = 12'h752 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20306; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26450 = 12'h752 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23378; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1874 = io_valid_in ? _GEN_26450 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1874 = 12'h752 == _T_2[11:0] ? image_1874 : _GEN_1873; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4947 = 12'h753 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8019 = 12'h753 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4947; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11091 = 12'h753 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8019; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14163 = 12'h753 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11091; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17235 = 12'h753 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14163; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20307 = 12'h753 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17235; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23379 = 12'h753 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20307; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26451 = 12'h753 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23379; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1875 = io_valid_in ? _GEN_26451 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1875 = 12'h753 == _T_2[11:0] ? image_1875 : _GEN_1874; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4948 = 12'h754 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8020 = 12'h754 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4948; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11092 = 12'h754 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8020; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14164 = 12'h754 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11092; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17236 = 12'h754 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14164; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20308 = 12'h754 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17236; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23380 = 12'h754 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20308; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26452 = 12'h754 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23380; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1876 = io_valid_in ? _GEN_26452 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1876 = 12'h754 == _T_2[11:0] ? image_1876 : _GEN_1875; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4949 = 12'h755 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8021 = 12'h755 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4949; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11093 = 12'h755 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8021; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14165 = 12'h755 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11093; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17237 = 12'h755 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14165; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20309 = 12'h755 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17237; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23381 = 12'h755 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20309; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26453 = 12'h755 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23381; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1877 = io_valid_in ? _GEN_26453 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1877 = 12'h755 == _T_2[11:0] ? image_1877 : _GEN_1876; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4950 = 12'h756 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8022 = 12'h756 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4950; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11094 = 12'h756 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8022; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14166 = 12'h756 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11094; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17238 = 12'h756 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14166; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20310 = 12'h756 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17238; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23382 = 12'h756 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20310; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26454 = 12'h756 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23382; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1878 = io_valid_in ? _GEN_26454 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1878 = 12'h756 == _T_2[11:0] ? image_1878 : _GEN_1877; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4951 = 12'h757 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8023 = 12'h757 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4951; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11095 = 12'h757 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8023; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14167 = 12'h757 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11095; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17239 = 12'h757 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14167; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20311 = 12'h757 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17239; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23383 = 12'h757 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20311; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26455 = 12'h757 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23383; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1879 = io_valid_in ? _GEN_26455 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1879 = 12'h757 == _T_2[11:0] ? image_1879 : _GEN_1878; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4952 = 12'h758 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8024 = 12'h758 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4952; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11096 = 12'h758 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8024; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14168 = 12'h758 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11096; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17240 = 12'h758 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14168; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20312 = 12'h758 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17240; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23384 = 12'h758 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20312; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26456 = 12'h758 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23384; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1880 = io_valid_in ? _GEN_26456 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1880 = 12'h758 == _T_2[11:0] ? image_1880 : _GEN_1879; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4953 = 12'h759 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8025 = 12'h759 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4953; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11097 = 12'h759 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8025; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14169 = 12'h759 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11097; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17241 = 12'h759 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14169; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20313 = 12'h759 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17241; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23385 = 12'h759 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20313; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26457 = 12'h759 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23385; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1881 = io_valid_in ? _GEN_26457 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1881 = 12'h759 == _T_2[11:0] ? image_1881 : _GEN_1880; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4954 = 12'h75a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8026 = 12'h75a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4954; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11098 = 12'h75a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8026; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14170 = 12'h75a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11098; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17242 = 12'h75a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14170; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20314 = 12'h75a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17242; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23386 = 12'h75a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20314; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26458 = 12'h75a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23386; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1882 = io_valid_in ? _GEN_26458 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1882 = 12'h75a == _T_2[11:0] ? image_1882 : _GEN_1881; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4955 = 12'h75b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8027 = 12'h75b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4955; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11099 = 12'h75b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8027; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14171 = 12'h75b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11099; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17243 = 12'h75b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14171; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20315 = 12'h75b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17243; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23387 = 12'h75b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20315; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26459 = 12'h75b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23387; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1883 = io_valid_in ? _GEN_26459 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1883 = 12'h75b == _T_2[11:0] ? image_1883 : _GEN_1882; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4956 = 12'h75c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8028 = 12'h75c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4956; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11100 = 12'h75c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8028; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14172 = 12'h75c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11100; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17244 = 12'h75c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14172; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20316 = 12'h75c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17244; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23388 = 12'h75c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20316; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26460 = 12'h75c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23388; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1884 = io_valid_in ? _GEN_26460 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1884 = 12'h75c == _T_2[11:0] ? image_1884 : _GEN_1883; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4957 = 12'h75d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8029 = 12'h75d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4957; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11101 = 12'h75d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8029; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14173 = 12'h75d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11101; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17245 = 12'h75d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14173; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20317 = 12'h75d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17245; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23389 = 12'h75d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20317; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26461 = 12'h75d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23389; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1885 = io_valid_in ? _GEN_26461 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1885 = 12'h75d == _T_2[11:0] ? image_1885 : _GEN_1884; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4958 = 12'h75e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8030 = 12'h75e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4958; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11102 = 12'h75e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8030; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14174 = 12'h75e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11102; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17246 = 12'h75e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14174; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20318 = 12'h75e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17246; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23390 = 12'h75e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20318; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26462 = 12'h75e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23390; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1886 = io_valid_in ? _GEN_26462 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1886 = 12'h75e == _T_2[11:0] ? image_1886 : _GEN_1885; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4959 = 12'h75f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8031 = 12'h75f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4959; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11103 = 12'h75f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8031; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14175 = 12'h75f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11103; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17247 = 12'h75f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14175; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20319 = 12'h75f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17247; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23391 = 12'h75f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20319; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26463 = 12'h75f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23391; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1887 = io_valid_in ? _GEN_26463 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1887 = 12'h75f == _T_2[11:0] ? image_1887 : _GEN_1886; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4960 = 12'h760 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8032 = 12'h760 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4960; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11104 = 12'h760 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8032; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14176 = 12'h760 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11104; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17248 = 12'h760 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14176; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20320 = 12'h760 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17248; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23392 = 12'h760 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20320; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26464 = 12'h760 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23392; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1888 = io_valid_in ? _GEN_26464 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1888 = 12'h760 == _T_2[11:0] ? image_1888 : _GEN_1887; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4961 = 12'h761 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8033 = 12'h761 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4961; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11105 = 12'h761 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8033; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14177 = 12'h761 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11105; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17249 = 12'h761 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14177; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20321 = 12'h761 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17249; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23393 = 12'h761 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20321; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26465 = 12'h761 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23393; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1889 = io_valid_in ? _GEN_26465 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1889 = 12'h761 == _T_2[11:0] ? image_1889 : _GEN_1888; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4962 = 12'h762 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8034 = 12'h762 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4962; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11106 = 12'h762 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8034; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14178 = 12'h762 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11106; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17250 = 12'h762 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14178; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20322 = 12'h762 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17250; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23394 = 12'h762 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20322; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26466 = 12'h762 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23394; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1890 = io_valid_in ? _GEN_26466 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1890 = 12'h762 == _T_2[11:0] ? image_1890 : _GEN_1889; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4963 = 12'h763 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8035 = 12'h763 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4963; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11107 = 12'h763 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8035; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14179 = 12'h763 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11107; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17251 = 12'h763 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14179; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20323 = 12'h763 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17251; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23395 = 12'h763 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20323; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26467 = 12'h763 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23395; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1891 = io_valid_in ? _GEN_26467 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1891 = 12'h763 == _T_2[11:0] ? image_1891 : _GEN_1890; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4964 = 12'h764 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8036 = 12'h764 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4964; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11108 = 12'h764 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8036; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14180 = 12'h764 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11108; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17252 = 12'h764 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14180; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20324 = 12'h764 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17252; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23396 = 12'h764 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20324; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26468 = 12'h764 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23396; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1892 = io_valid_in ? _GEN_26468 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1892 = 12'h764 == _T_2[11:0] ? image_1892 : _GEN_1891; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4965 = 12'h765 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8037 = 12'h765 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4965; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11109 = 12'h765 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8037; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14181 = 12'h765 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11109; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17253 = 12'h765 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14181; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20325 = 12'h765 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17253; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23397 = 12'h765 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20325; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26469 = 12'h765 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23397; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1893 = io_valid_in ? _GEN_26469 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1893 = 12'h765 == _T_2[11:0] ? image_1893 : _GEN_1892; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4966 = 12'h766 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8038 = 12'h766 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4966; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11110 = 12'h766 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8038; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14182 = 12'h766 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11110; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17254 = 12'h766 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14182; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20326 = 12'h766 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17254; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23398 = 12'h766 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20326; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26470 = 12'h766 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23398; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1894 = io_valid_in ? _GEN_26470 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1894 = 12'h766 == _T_2[11:0] ? image_1894 : _GEN_1893; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4967 = 12'h767 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8039 = 12'h767 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4967; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11111 = 12'h767 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8039; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14183 = 12'h767 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11111; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17255 = 12'h767 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14183; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20327 = 12'h767 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17255; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23399 = 12'h767 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20327; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26471 = 12'h767 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23399; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1895 = io_valid_in ? _GEN_26471 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1895 = 12'h767 == _T_2[11:0] ? image_1895 : _GEN_1894; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4968 = 12'h768 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8040 = 12'h768 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4968; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11112 = 12'h768 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8040; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14184 = 12'h768 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11112; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17256 = 12'h768 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14184; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20328 = 12'h768 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17256; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23400 = 12'h768 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20328; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26472 = 12'h768 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23400; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1896 = io_valid_in ? _GEN_26472 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1896 = 12'h768 == _T_2[11:0] ? image_1896 : _GEN_1895; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4969 = 12'h769 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8041 = 12'h769 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4969; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11113 = 12'h769 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8041; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14185 = 12'h769 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11113; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17257 = 12'h769 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14185; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20329 = 12'h769 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17257; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23401 = 12'h769 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20329; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26473 = 12'h769 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23401; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1897 = io_valid_in ? _GEN_26473 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1897 = 12'h769 == _T_2[11:0] ? image_1897 : _GEN_1896; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4970 = 12'h76a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8042 = 12'h76a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4970; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11114 = 12'h76a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8042; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14186 = 12'h76a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11114; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17258 = 12'h76a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14186; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20330 = 12'h76a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17258; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23402 = 12'h76a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20330; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26474 = 12'h76a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23402; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1898 = io_valid_in ? _GEN_26474 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1898 = 12'h76a == _T_2[11:0] ? image_1898 : _GEN_1897; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4971 = 12'h76b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8043 = 12'h76b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4971; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11115 = 12'h76b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8043; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14187 = 12'h76b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11115; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17259 = 12'h76b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14187; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20331 = 12'h76b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17259; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23403 = 12'h76b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20331; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26475 = 12'h76b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23403; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1899 = io_valid_in ? _GEN_26475 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1899 = 12'h76b == _T_2[11:0] ? image_1899 : _GEN_1898; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4972 = 12'h76c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8044 = 12'h76c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4972; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11116 = 12'h76c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8044; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14188 = 12'h76c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11116; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17260 = 12'h76c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14188; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20332 = 12'h76c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17260; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23404 = 12'h76c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20332; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26476 = 12'h76c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23404; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1900 = io_valid_in ? _GEN_26476 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1900 = 12'h76c == _T_2[11:0] ? image_1900 : _GEN_1899; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4973 = 12'h76d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8045 = 12'h76d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4973; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11117 = 12'h76d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8045; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14189 = 12'h76d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11117; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17261 = 12'h76d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14189; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20333 = 12'h76d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17261; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23405 = 12'h76d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20333; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26477 = 12'h76d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23405; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1901 = io_valid_in ? _GEN_26477 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1901 = 12'h76d == _T_2[11:0] ? image_1901 : _GEN_1900; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4974 = 12'h76e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8046 = 12'h76e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4974; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11118 = 12'h76e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8046; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14190 = 12'h76e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11118; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17262 = 12'h76e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14190; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20334 = 12'h76e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17262; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23406 = 12'h76e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20334; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26478 = 12'h76e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23406; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1902 = io_valid_in ? _GEN_26478 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1902 = 12'h76e == _T_2[11:0] ? image_1902 : _GEN_1901; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4975 = 12'h76f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8047 = 12'h76f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4975; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11119 = 12'h76f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8047; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14191 = 12'h76f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11119; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17263 = 12'h76f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14191; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20335 = 12'h76f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17263; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23407 = 12'h76f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20335; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26479 = 12'h76f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23407; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1903 = io_valid_in ? _GEN_26479 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1903 = 12'h76f == _T_2[11:0] ? image_1903 : _GEN_1902; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4976 = 12'h770 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8048 = 12'h770 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4976; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11120 = 12'h770 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8048; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14192 = 12'h770 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11120; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17264 = 12'h770 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14192; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20336 = 12'h770 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17264; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23408 = 12'h770 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20336; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26480 = 12'h770 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23408; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1904 = io_valid_in ? _GEN_26480 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1904 = 12'h770 == _T_2[11:0] ? image_1904 : _GEN_1903; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4977 = 12'h771 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8049 = 12'h771 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4977; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11121 = 12'h771 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8049; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14193 = 12'h771 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11121; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17265 = 12'h771 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14193; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20337 = 12'h771 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17265; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23409 = 12'h771 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20337; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26481 = 12'h771 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23409; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1905 = io_valid_in ? _GEN_26481 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1905 = 12'h771 == _T_2[11:0] ? image_1905 : _GEN_1904; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4978 = 12'h772 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8050 = 12'h772 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4978; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11122 = 12'h772 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8050; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14194 = 12'h772 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11122; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17266 = 12'h772 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14194; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20338 = 12'h772 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17266; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23410 = 12'h772 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20338; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26482 = 12'h772 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23410; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1906 = io_valid_in ? _GEN_26482 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1906 = 12'h772 == _T_2[11:0] ? image_1906 : _GEN_1905; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4979 = 12'h773 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8051 = 12'h773 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4979; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11123 = 12'h773 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8051; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14195 = 12'h773 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11123; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17267 = 12'h773 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14195; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20339 = 12'h773 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17267; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23411 = 12'h773 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20339; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26483 = 12'h773 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23411; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1907 = io_valid_in ? _GEN_26483 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1907 = 12'h773 == _T_2[11:0] ? image_1907 : _GEN_1906; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4980 = 12'h774 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8052 = 12'h774 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4980; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11124 = 12'h774 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8052; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14196 = 12'h774 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11124; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17268 = 12'h774 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14196; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20340 = 12'h774 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17268; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23412 = 12'h774 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20340; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26484 = 12'h774 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23412; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1908 = io_valid_in ? _GEN_26484 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1908 = 12'h774 == _T_2[11:0] ? image_1908 : _GEN_1907; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4981 = 12'h775 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8053 = 12'h775 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4981; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11125 = 12'h775 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8053; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14197 = 12'h775 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11125; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17269 = 12'h775 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14197; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20341 = 12'h775 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17269; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23413 = 12'h775 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20341; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26485 = 12'h775 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23413; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1909 = io_valid_in ? _GEN_26485 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1909 = 12'h775 == _T_2[11:0] ? image_1909 : _GEN_1908; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4982 = 12'h776 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8054 = 12'h776 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4982; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11126 = 12'h776 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8054; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14198 = 12'h776 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11126; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17270 = 12'h776 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14198; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20342 = 12'h776 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17270; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23414 = 12'h776 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20342; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26486 = 12'h776 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23414; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1910 = io_valid_in ? _GEN_26486 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1910 = 12'h776 == _T_2[11:0] ? image_1910 : _GEN_1909; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4983 = 12'h777 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8055 = 12'h777 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4983; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11127 = 12'h777 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8055; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14199 = 12'h777 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11127; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17271 = 12'h777 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14199; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20343 = 12'h777 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17271; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23415 = 12'h777 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20343; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26487 = 12'h777 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23415; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1911 = io_valid_in ? _GEN_26487 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1911 = 12'h777 == _T_2[11:0] ? image_1911 : _GEN_1910; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4984 = 12'h778 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8056 = 12'h778 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4984; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11128 = 12'h778 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8056; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14200 = 12'h778 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11128; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17272 = 12'h778 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14200; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20344 = 12'h778 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17272; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23416 = 12'h778 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20344; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26488 = 12'h778 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23416; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1912 = io_valid_in ? _GEN_26488 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1912 = 12'h778 == _T_2[11:0] ? image_1912 : _GEN_1911; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4985 = 12'h779 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8057 = 12'h779 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4985; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11129 = 12'h779 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8057; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14201 = 12'h779 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11129; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17273 = 12'h779 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14201; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20345 = 12'h779 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17273; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23417 = 12'h779 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20345; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26489 = 12'h779 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23417; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1913 = io_valid_in ? _GEN_26489 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1913 = 12'h779 == _T_2[11:0] ? image_1913 : _GEN_1912; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4986 = 12'h77a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8058 = 12'h77a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4986; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11130 = 12'h77a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8058; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14202 = 12'h77a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11130; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17274 = 12'h77a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14202; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20346 = 12'h77a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17274; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23418 = 12'h77a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20346; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26490 = 12'h77a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23418; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1914 = io_valid_in ? _GEN_26490 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1914 = 12'h77a == _T_2[11:0] ? image_1914 : _GEN_1913; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4987 = 12'h77b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8059 = 12'h77b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4987; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11131 = 12'h77b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8059; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14203 = 12'h77b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11131; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17275 = 12'h77b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14203; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20347 = 12'h77b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17275; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23419 = 12'h77b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20347; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26491 = 12'h77b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23419; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1915 = io_valid_in ? _GEN_26491 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1915 = 12'h77b == _T_2[11:0] ? image_1915 : _GEN_1914; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4988 = 12'h77c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8060 = 12'h77c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4988; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11132 = 12'h77c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8060; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14204 = 12'h77c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11132; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17276 = 12'h77c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14204; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20348 = 12'h77c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17276; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23420 = 12'h77c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20348; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26492 = 12'h77c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23420; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1916 = io_valid_in ? _GEN_26492 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1916 = 12'h77c == _T_2[11:0] ? image_1916 : _GEN_1915; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4989 = 12'h77d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8061 = 12'h77d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4989; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11133 = 12'h77d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8061; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14205 = 12'h77d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11133; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17277 = 12'h77d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14205; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20349 = 12'h77d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17277; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23421 = 12'h77d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20349; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26493 = 12'h77d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23421; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1917 = io_valid_in ? _GEN_26493 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1917 = 12'h77d == _T_2[11:0] ? image_1917 : _GEN_1916; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4990 = 12'h77e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8062 = 12'h77e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4990; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11134 = 12'h77e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8062; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14206 = 12'h77e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11134; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17278 = 12'h77e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14206; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20350 = 12'h77e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17278; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23422 = 12'h77e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20350; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26494 = 12'h77e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23422; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1918 = io_valid_in ? _GEN_26494 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1918 = 12'h77e == _T_2[11:0] ? image_1918 : _GEN_1917; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4991 = 12'h77f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8063 = 12'h77f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4991; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11135 = 12'h77f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8063; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14207 = 12'h77f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11135; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17279 = 12'h77f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14207; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20351 = 12'h77f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17279; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23423 = 12'h77f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20351; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26495 = 12'h77f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23423; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1919 = io_valid_in ? _GEN_26495 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1919 = 12'h77f == _T_2[11:0] ? image_1919 : _GEN_1918; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4992 = 12'h780 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8064 = 12'h780 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4992; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11136 = 12'h780 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8064; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14208 = 12'h780 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11136; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17280 = 12'h780 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14208; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20352 = 12'h780 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17280; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23424 = 12'h780 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20352; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26496 = 12'h780 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23424; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1920 = io_valid_in ? _GEN_26496 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1920 = 12'h780 == _T_2[11:0] ? image_1920 : _GEN_1919; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4993 = 12'h781 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8065 = 12'h781 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4993; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11137 = 12'h781 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8065; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14209 = 12'h781 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11137; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17281 = 12'h781 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14209; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20353 = 12'h781 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17281; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23425 = 12'h781 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20353; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26497 = 12'h781 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23425; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1921 = io_valid_in ? _GEN_26497 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1921 = 12'h781 == _T_2[11:0] ? image_1921 : _GEN_1920; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4994 = 12'h782 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8066 = 12'h782 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4994; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11138 = 12'h782 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8066; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14210 = 12'h782 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11138; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17282 = 12'h782 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14210; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20354 = 12'h782 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17282; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23426 = 12'h782 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20354; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26498 = 12'h782 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23426; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1922 = io_valid_in ? _GEN_26498 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1922 = 12'h782 == _T_2[11:0] ? image_1922 : _GEN_1921; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4995 = 12'h783 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8067 = 12'h783 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4995; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11139 = 12'h783 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8067; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14211 = 12'h783 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11139; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17283 = 12'h783 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14211; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20355 = 12'h783 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17283; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23427 = 12'h783 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20355; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26499 = 12'h783 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23427; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1923 = io_valid_in ? _GEN_26499 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1923 = 12'h783 == _T_2[11:0] ? image_1923 : _GEN_1922; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4996 = 12'h784 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8068 = 12'h784 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4996; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11140 = 12'h784 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8068; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14212 = 12'h784 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11140; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17284 = 12'h784 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14212; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20356 = 12'h784 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17284; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23428 = 12'h784 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20356; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26500 = 12'h784 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23428; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1924 = io_valid_in ? _GEN_26500 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1924 = 12'h784 == _T_2[11:0] ? image_1924 : _GEN_1923; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4997 = 12'h785 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8069 = 12'h785 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4997; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11141 = 12'h785 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8069; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14213 = 12'h785 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11141; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17285 = 12'h785 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14213; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20357 = 12'h785 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17285; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23429 = 12'h785 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20357; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26501 = 12'h785 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23429; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1925 = io_valid_in ? _GEN_26501 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1925 = 12'h785 == _T_2[11:0] ? image_1925 : _GEN_1924; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4998 = 12'h786 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8070 = 12'h786 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4998; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11142 = 12'h786 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8070; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14214 = 12'h786 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11142; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17286 = 12'h786 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14214; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20358 = 12'h786 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17286; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23430 = 12'h786 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20358; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26502 = 12'h786 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23430; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1926 = io_valid_in ? _GEN_26502 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1926 = 12'h786 == _T_2[11:0] ? image_1926 : _GEN_1925; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_4999 = 12'h787 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8071 = 12'h787 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_4999; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11143 = 12'h787 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8071; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14215 = 12'h787 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11143; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17287 = 12'h787 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14215; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20359 = 12'h787 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17287; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23431 = 12'h787 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20359; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26503 = 12'h787 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23431; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1927 = io_valid_in ? _GEN_26503 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1927 = 12'h787 == _T_2[11:0] ? image_1927 : _GEN_1926; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5000 = 12'h788 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8072 = 12'h788 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5000; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11144 = 12'h788 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8072; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14216 = 12'h788 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11144; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17288 = 12'h788 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14216; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20360 = 12'h788 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17288; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23432 = 12'h788 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20360; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26504 = 12'h788 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23432; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1928 = io_valid_in ? _GEN_26504 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1928 = 12'h788 == _T_2[11:0] ? image_1928 : _GEN_1927; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5001 = 12'h789 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8073 = 12'h789 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5001; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11145 = 12'h789 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8073; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14217 = 12'h789 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11145; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17289 = 12'h789 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14217; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20361 = 12'h789 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17289; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23433 = 12'h789 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20361; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26505 = 12'h789 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23433; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1929 = io_valid_in ? _GEN_26505 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1929 = 12'h789 == _T_2[11:0] ? image_1929 : _GEN_1928; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5002 = 12'h78a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8074 = 12'h78a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5002; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11146 = 12'h78a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8074; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14218 = 12'h78a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11146; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17290 = 12'h78a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14218; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20362 = 12'h78a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17290; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23434 = 12'h78a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20362; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26506 = 12'h78a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23434; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1930 = io_valid_in ? _GEN_26506 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1930 = 12'h78a == _T_2[11:0] ? image_1930 : _GEN_1929; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5003 = 12'h78b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8075 = 12'h78b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5003; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11147 = 12'h78b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8075; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14219 = 12'h78b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11147; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17291 = 12'h78b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14219; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20363 = 12'h78b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17291; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23435 = 12'h78b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20363; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26507 = 12'h78b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23435; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1931 = io_valid_in ? _GEN_26507 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1931 = 12'h78b == _T_2[11:0] ? image_1931 : _GEN_1930; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5004 = 12'h78c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8076 = 12'h78c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5004; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11148 = 12'h78c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8076; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14220 = 12'h78c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11148; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17292 = 12'h78c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14220; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20364 = 12'h78c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17292; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23436 = 12'h78c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20364; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26508 = 12'h78c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23436; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1932 = io_valid_in ? _GEN_26508 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1932 = 12'h78c == _T_2[11:0] ? image_1932 : _GEN_1931; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5005 = 12'h78d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8077 = 12'h78d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5005; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11149 = 12'h78d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8077; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14221 = 12'h78d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11149; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17293 = 12'h78d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14221; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20365 = 12'h78d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17293; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23437 = 12'h78d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20365; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26509 = 12'h78d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23437; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1933 = io_valid_in ? _GEN_26509 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1933 = 12'h78d == _T_2[11:0] ? image_1933 : _GEN_1932; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5006 = 12'h78e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8078 = 12'h78e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5006; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11150 = 12'h78e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8078; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14222 = 12'h78e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11150; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17294 = 12'h78e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14222; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20366 = 12'h78e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17294; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23438 = 12'h78e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20366; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26510 = 12'h78e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23438; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1934 = io_valid_in ? _GEN_26510 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1934 = 12'h78e == _T_2[11:0] ? image_1934 : _GEN_1933; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5007 = 12'h78f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8079 = 12'h78f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5007; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11151 = 12'h78f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8079; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14223 = 12'h78f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11151; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17295 = 12'h78f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14223; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20367 = 12'h78f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17295; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23439 = 12'h78f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20367; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26511 = 12'h78f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23439; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1935 = io_valid_in ? _GEN_26511 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1935 = 12'h78f == _T_2[11:0] ? image_1935 : _GEN_1934; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5008 = 12'h790 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8080 = 12'h790 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5008; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11152 = 12'h790 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8080; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14224 = 12'h790 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11152; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17296 = 12'h790 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14224; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20368 = 12'h790 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17296; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23440 = 12'h790 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20368; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26512 = 12'h790 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23440; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1936 = io_valid_in ? _GEN_26512 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1936 = 12'h790 == _T_2[11:0] ? image_1936 : _GEN_1935; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5009 = 12'h791 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8081 = 12'h791 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5009; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11153 = 12'h791 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8081; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14225 = 12'h791 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11153; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17297 = 12'h791 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14225; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20369 = 12'h791 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17297; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23441 = 12'h791 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20369; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26513 = 12'h791 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23441; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1937 = io_valid_in ? _GEN_26513 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1937 = 12'h791 == _T_2[11:0] ? image_1937 : _GEN_1936; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5010 = 12'h792 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8082 = 12'h792 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5010; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11154 = 12'h792 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8082; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14226 = 12'h792 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11154; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17298 = 12'h792 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14226; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20370 = 12'h792 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17298; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23442 = 12'h792 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20370; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26514 = 12'h792 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23442; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1938 = io_valid_in ? _GEN_26514 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1938 = 12'h792 == _T_2[11:0] ? image_1938 : _GEN_1937; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5011 = 12'h793 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8083 = 12'h793 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5011; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11155 = 12'h793 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8083; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14227 = 12'h793 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11155; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17299 = 12'h793 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14227; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20371 = 12'h793 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17299; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23443 = 12'h793 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20371; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26515 = 12'h793 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23443; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1939 = io_valid_in ? _GEN_26515 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1939 = 12'h793 == _T_2[11:0] ? image_1939 : _GEN_1938; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5012 = 12'h794 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8084 = 12'h794 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5012; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11156 = 12'h794 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8084; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14228 = 12'h794 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11156; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17300 = 12'h794 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14228; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20372 = 12'h794 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17300; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23444 = 12'h794 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20372; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26516 = 12'h794 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23444; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1940 = io_valid_in ? _GEN_26516 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1940 = 12'h794 == _T_2[11:0] ? image_1940 : _GEN_1939; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5013 = 12'h795 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8085 = 12'h795 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5013; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11157 = 12'h795 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8085; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14229 = 12'h795 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11157; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17301 = 12'h795 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14229; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20373 = 12'h795 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17301; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23445 = 12'h795 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20373; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26517 = 12'h795 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23445; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1941 = io_valid_in ? _GEN_26517 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1941 = 12'h795 == _T_2[11:0] ? image_1941 : _GEN_1940; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5014 = 12'h796 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8086 = 12'h796 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5014; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11158 = 12'h796 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8086; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14230 = 12'h796 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11158; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17302 = 12'h796 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14230; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20374 = 12'h796 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17302; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23446 = 12'h796 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20374; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26518 = 12'h796 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23446; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1942 = io_valid_in ? _GEN_26518 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1942 = 12'h796 == _T_2[11:0] ? image_1942 : _GEN_1941; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5015 = 12'h797 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8087 = 12'h797 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5015; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11159 = 12'h797 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8087; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14231 = 12'h797 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11159; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17303 = 12'h797 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14231; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20375 = 12'h797 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17303; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23447 = 12'h797 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20375; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26519 = 12'h797 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23447; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1943 = io_valid_in ? _GEN_26519 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1943 = 12'h797 == _T_2[11:0] ? image_1943 : _GEN_1942; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5016 = 12'h798 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8088 = 12'h798 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5016; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11160 = 12'h798 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8088; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14232 = 12'h798 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11160; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17304 = 12'h798 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14232; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20376 = 12'h798 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17304; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23448 = 12'h798 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20376; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26520 = 12'h798 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23448; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1944 = io_valid_in ? _GEN_26520 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1944 = 12'h798 == _T_2[11:0] ? image_1944 : _GEN_1943; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5017 = 12'h799 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8089 = 12'h799 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5017; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11161 = 12'h799 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8089; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14233 = 12'h799 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11161; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17305 = 12'h799 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14233; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20377 = 12'h799 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17305; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23449 = 12'h799 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20377; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26521 = 12'h799 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23449; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1945 = io_valid_in ? _GEN_26521 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1945 = 12'h799 == _T_2[11:0] ? image_1945 : _GEN_1944; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5018 = 12'h79a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8090 = 12'h79a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5018; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11162 = 12'h79a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8090; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14234 = 12'h79a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11162; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17306 = 12'h79a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14234; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20378 = 12'h79a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17306; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23450 = 12'h79a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20378; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26522 = 12'h79a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23450; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1946 = io_valid_in ? _GEN_26522 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1946 = 12'h79a == _T_2[11:0] ? image_1946 : _GEN_1945; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5019 = 12'h79b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8091 = 12'h79b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5019; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11163 = 12'h79b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8091; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14235 = 12'h79b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11163; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17307 = 12'h79b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14235; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20379 = 12'h79b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17307; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23451 = 12'h79b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20379; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26523 = 12'h79b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23451; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1947 = io_valid_in ? _GEN_26523 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1947 = 12'h79b == _T_2[11:0] ? image_1947 : _GEN_1946; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5020 = 12'h79c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8092 = 12'h79c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5020; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11164 = 12'h79c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8092; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14236 = 12'h79c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11164; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17308 = 12'h79c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14236; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20380 = 12'h79c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17308; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23452 = 12'h79c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20380; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26524 = 12'h79c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23452; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1948 = io_valid_in ? _GEN_26524 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1948 = 12'h79c == _T_2[11:0] ? image_1948 : _GEN_1947; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5021 = 12'h79d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8093 = 12'h79d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5021; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11165 = 12'h79d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8093; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14237 = 12'h79d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11165; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17309 = 12'h79d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14237; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20381 = 12'h79d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17309; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23453 = 12'h79d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20381; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26525 = 12'h79d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23453; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1949 = io_valid_in ? _GEN_26525 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1949 = 12'h79d == _T_2[11:0] ? image_1949 : _GEN_1948; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5022 = 12'h79e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8094 = 12'h79e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5022; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11166 = 12'h79e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8094; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14238 = 12'h79e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11166; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17310 = 12'h79e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14238; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20382 = 12'h79e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17310; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23454 = 12'h79e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20382; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26526 = 12'h79e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23454; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1950 = io_valid_in ? _GEN_26526 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1950 = 12'h79e == _T_2[11:0] ? image_1950 : _GEN_1949; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5023 = 12'h79f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8095 = 12'h79f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5023; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11167 = 12'h79f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8095; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14239 = 12'h79f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11167; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17311 = 12'h79f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14239; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20383 = 12'h79f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17311; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23455 = 12'h79f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20383; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26527 = 12'h79f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23455; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1951 = io_valid_in ? _GEN_26527 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1951 = 12'h79f == _T_2[11:0] ? image_1951 : _GEN_1950; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5024 = 12'h7a0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8096 = 12'h7a0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5024; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11168 = 12'h7a0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8096; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14240 = 12'h7a0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11168; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17312 = 12'h7a0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14240; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20384 = 12'h7a0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17312; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23456 = 12'h7a0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20384; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26528 = 12'h7a0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23456; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1952 = io_valid_in ? _GEN_26528 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1952 = 12'h7a0 == _T_2[11:0] ? image_1952 : _GEN_1951; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5025 = 12'h7a1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8097 = 12'h7a1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5025; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11169 = 12'h7a1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8097; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14241 = 12'h7a1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11169; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17313 = 12'h7a1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14241; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20385 = 12'h7a1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17313; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23457 = 12'h7a1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20385; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26529 = 12'h7a1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23457; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1953 = io_valid_in ? _GEN_26529 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1953 = 12'h7a1 == _T_2[11:0] ? image_1953 : _GEN_1952; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5026 = 12'h7a2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8098 = 12'h7a2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5026; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11170 = 12'h7a2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8098; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14242 = 12'h7a2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11170; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17314 = 12'h7a2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14242; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20386 = 12'h7a2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17314; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23458 = 12'h7a2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20386; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26530 = 12'h7a2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23458; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1954 = io_valid_in ? _GEN_26530 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1954 = 12'h7a2 == _T_2[11:0] ? image_1954 : _GEN_1953; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5027 = 12'h7a3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8099 = 12'h7a3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5027; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11171 = 12'h7a3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8099; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14243 = 12'h7a3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11171; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17315 = 12'h7a3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14243; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20387 = 12'h7a3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17315; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23459 = 12'h7a3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20387; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26531 = 12'h7a3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23459; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1955 = io_valid_in ? _GEN_26531 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1955 = 12'h7a3 == _T_2[11:0] ? image_1955 : _GEN_1954; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5028 = 12'h7a4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8100 = 12'h7a4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5028; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11172 = 12'h7a4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8100; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14244 = 12'h7a4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11172; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17316 = 12'h7a4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14244; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20388 = 12'h7a4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17316; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23460 = 12'h7a4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20388; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26532 = 12'h7a4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23460; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1956 = io_valid_in ? _GEN_26532 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1956 = 12'h7a4 == _T_2[11:0] ? image_1956 : _GEN_1955; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5029 = 12'h7a5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8101 = 12'h7a5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5029; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11173 = 12'h7a5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8101; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14245 = 12'h7a5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11173; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17317 = 12'h7a5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14245; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20389 = 12'h7a5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17317; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23461 = 12'h7a5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20389; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26533 = 12'h7a5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23461; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1957 = io_valid_in ? _GEN_26533 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1957 = 12'h7a5 == _T_2[11:0] ? image_1957 : _GEN_1956; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5030 = 12'h7a6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8102 = 12'h7a6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5030; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11174 = 12'h7a6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8102; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14246 = 12'h7a6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11174; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17318 = 12'h7a6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14246; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20390 = 12'h7a6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17318; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23462 = 12'h7a6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20390; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26534 = 12'h7a6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23462; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1958 = io_valid_in ? _GEN_26534 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1958 = 12'h7a6 == _T_2[11:0] ? image_1958 : _GEN_1957; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5031 = 12'h7a7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8103 = 12'h7a7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5031; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11175 = 12'h7a7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8103; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14247 = 12'h7a7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11175; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17319 = 12'h7a7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14247; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20391 = 12'h7a7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17319; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23463 = 12'h7a7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20391; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26535 = 12'h7a7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23463; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1959 = io_valid_in ? _GEN_26535 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1959 = 12'h7a7 == _T_2[11:0] ? image_1959 : _GEN_1958; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5032 = 12'h7a8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8104 = 12'h7a8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5032; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11176 = 12'h7a8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8104; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14248 = 12'h7a8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11176; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17320 = 12'h7a8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14248; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20392 = 12'h7a8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17320; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23464 = 12'h7a8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20392; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26536 = 12'h7a8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23464; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1960 = io_valid_in ? _GEN_26536 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1960 = 12'h7a8 == _T_2[11:0] ? image_1960 : _GEN_1959; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5033 = 12'h7a9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8105 = 12'h7a9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5033; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11177 = 12'h7a9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8105; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14249 = 12'h7a9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11177; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17321 = 12'h7a9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14249; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20393 = 12'h7a9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17321; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23465 = 12'h7a9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20393; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26537 = 12'h7a9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23465; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1961 = io_valid_in ? _GEN_26537 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1961 = 12'h7a9 == _T_2[11:0] ? image_1961 : _GEN_1960; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5034 = 12'h7aa == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8106 = 12'h7aa == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5034; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11178 = 12'h7aa == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8106; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14250 = 12'h7aa == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11178; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17322 = 12'h7aa == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14250; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20394 = 12'h7aa == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17322; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23466 = 12'h7aa == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20394; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26538 = 12'h7aa == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23466; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1962 = io_valid_in ? _GEN_26538 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1962 = 12'h7aa == _T_2[11:0] ? image_1962 : _GEN_1961; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5035 = 12'h7ab == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8107 = 12'h7ab == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5035; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11179 = 12'h7ab == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8107; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14251 = 12'h7ab == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11179; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17323 = 12'h7ab == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14251; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20395 = 12'h7ab == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17323; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23467 = 12'h7ab == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20395; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26539 = 12'h7ab == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23467; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1963 = io_valid_in ? _GEN_26539 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1963 = 12'h7ab == _T_2[11:0] ? image_1963 : _GEN_1962; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5036 = 12'h7ac == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8108 = 12'h7ac == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5036; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11180 = 12'h7ac == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8108; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14252 = 12'h7ac == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11180; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17324 = 12'h7ac == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14252; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20396 = 12'h7ac == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17324; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23468 = 12'h7ac == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20396; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26540 = 12'h7ac == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23468; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1964 = io_valid_in ? _GEN_26540 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1964 = 12'h7ac == _T_2[11:0] ? image_1964 : _GEN_1963; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5037 = 12'h7ad == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8109 = 12'h7ad == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5037; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11181 = 12'h7ad == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8109; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14253 = 12'h7ad == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11181; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17325 = 12'h7ad == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14253; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20397 = 12'h7ad == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17325; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23469 = 12'h7ad == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20397; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26541 = 12'h7ad == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23469; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1965 = io_valid_in ? _GEN_26541 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1965 = 12'h7ad == _T_2[11:0] ? image_1965 : _GEN_1964; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5038 = 12'h7ae == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8110 = 12'h7ae == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5038; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11182 = 12'h7ae == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8110; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14254 = 12'h7ae == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11182; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17326 = 12'h7ae == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14254; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20398 = 12'h7ae == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17326; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23470 = 12'h7ae == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20398; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26542 = 12'h7ae == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23470; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1966 = io_valid_in ? _GEN_26542 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1966 = 12'h7ae == _T_2[11:0] ? image_1966 : _GEN_1965; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5039 = 12'h7af == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8111 = 12'h7af == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5039; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11183 = 12'h7af == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8111; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14255 = 12'h7af == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11183; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17327 = 12'h7af == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14255; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20399 = 12'h7af == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17327; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23471 = 12'h7af == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20399; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26543 = 12'h7af == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23471; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1967 = io_valid_in ? _GEN_26543 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1967 = 12'h7af == _T_2[11:0] ? image_1967 : _GEN_1966; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5040 = 12'h7b0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8112 = 12'h7b0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5040; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11184 = 12'h7b0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8112; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14256 = 12'h7b0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11184; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17328 = 12'h7b0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14256; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20400 = 12'h7b0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17328; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23472 = 12'h7b0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20400; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26544 = 12'h7b0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23472; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1968 = io_valid_in ? _GEN_26544 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1968 = 12'h7b0 == _T_2[11:0] ? image_1968 : _GEN_1967; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5041 = 12'h7b1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8113 = 12'h7b1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5041; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11185 = 12'h7b1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8113; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14257 = 12'h7b1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11185; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17329 = 12'h7b1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14257; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20401 = 12'h7b1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17329; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23473 = 12'h7b1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20401; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26545 = 12'h7b1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23473; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1969 = io_valid_in ? _GEN_26545 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1969 = 12'h7b1 == _T_2[11:0] ? image_1969 : _GEN_1968; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5042 = 12'h7b2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8114 = 12'h7b2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5042; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11186 = 12'h7b2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8114; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14258 = 12'h7b2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11186; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17330 = 12'h7b2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14258; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20402 = 12'h7b2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17330; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23474 = 12'h7b2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20402; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26546 = 12'h7b2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23474; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1970 = io_valid_in ? _GEN_26546 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1970 = 12'h7b2 == _T_2[11:0] ? image_1970 : _GEN_1969; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5043 = 12'h7b3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8115 = 12'h7b3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5043; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11187 = 12'h7b3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8115; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14259 = 12'h7b3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11187; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17331 = 12'h7b3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14259; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20403 = 12'h7b3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17331; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23475 = 12'h7b3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20403; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26547 = 12'h7b3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23475; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1971 = io_valid_in ? _GEN_26547 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1971 = 12'h7b3 == _T_2[11:0] ? image_1971 : _GEN_1970; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5044 = 12'h7b4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8116 = 12'h7b4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5044; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11188 = 12'h7b4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8116; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14260 = 12'h7b4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11188; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17332 = 12'h7b4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14260; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20404 = 12'h7b4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17332; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23476 = 12'h7b4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20404; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26548 = 12'h7b4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23476; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1972 = io_valid_in ? _GEN_26548 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1972 = 12'h7b4 == _T_2[11:0] ? image_1972 : _GEN_1971; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5045 = 12'h7b5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8117 = 12'h7b5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5045; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11189 = 12'h7b5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8117; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14261 = 12'h7b5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11189; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17333 = 12'h7b5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14261; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20405 = 12'h7b5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17333; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23477 = 12'h7b5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20405; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26549 = 12'h7b5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23477; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1973 = io_valid_in ? _GEN_26549 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1973 = 12'h7b5 == _T_2[11:0] ? image_1973 : _GEN_1972; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5046 = 12'h7b6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8118 = 12'h7b6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5046; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11190 = 12'h7b6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8118; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14262 = 12'h7b6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11190; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17334 = 12'h7b6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14262; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20406 = 12'h7b6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17334; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23478 = 12'h7b6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20406; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26550 = 12'h7b6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23478; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1974 = io_valid_in ? _GEN_26550 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1974 = 12'h7b6 == _T_2[11:0] ? image_1974 : _GEN_1973; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5047 = 12'h7b7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8119 = 12'h7b7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5047; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11191 = 12'h7b7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8119; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14263 = 12'h7b7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11191; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17335 = 12'h7b7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14263; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20407 = 12'h7b7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17335; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23479 = 12'h7b7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20407; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26551 = 12'h7b7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23479; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1975 = io_valid_in ? _GEN_26551 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1975 = 12'h7b7 == _T_2[11:0] ? image_1975 : _GEN_1974; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5048 = 12'h7b8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8120 = 12'h7b8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5048; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11192 = 12'h7b8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8120; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14264 = 12'h7b8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11192; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17336 = 12'h7b8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14264; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20408 = 12'h7b8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17336; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23480 = 12'h7b8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20408; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26552 = 12'h7b8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23480; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1976 = io_valid_in ? _GEN_26552 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1976 = 12'h7b8 == _T_2[11:0] ? image_1976 : _GEN_1975; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5049 = 12'h7b9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8121 = 12'h7b9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5049; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11193 = 12'h7b9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8121; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14265 = 12'h7b9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11193; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17337 = 12'h7b9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14265; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20409 = 12'h7b9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17337; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23481 = 12'h7b9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20409; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26553 = 12'h7b9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23481; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1977 = io_valid_in ? _GEN_26553 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1977 = 12'h7b9 == _T_2[11:0] ? image_1977 : _GEN_1976; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5050 = 12'h7ba == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8122 = 12'h7ba == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5050; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11194 = 12'h7ba == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8122; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14266 = 12'h7ba == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11194; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17338 = 12'h7ba == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14266; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20410 = 12'h7ba == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17338; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23482 = 12'h7ba == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20410; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26554 = 12'h7ba == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23482; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1978 = io_valid_in ? _GEN_26554 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1978 = 12'h7ba == _T_2[11:0] ? image_1978 : _GEN_1977; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5051 = 12'h7bb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8123 = 12'h7bb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5051; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11195 = 12'h7bb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8123; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14267 = 12'h7bb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11195; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17339 = 12'h7bb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14267; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20411 = 12'h7bb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17339; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23483 = 12'h7bb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20411; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26555 = 12'h7bb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23483; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1979 = io_valid_in ? _GEN_26555 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1979 = 12'h7bb == _T_2[11:0] ? image_1979 : _GEN_1978; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5052 = 12'h7bc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8124 = 12'h7bc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5052; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11196 = 12'h7bc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8124; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14268 = 12'h7bc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11196; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17340 = 12'h7bc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14268; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20412 = 12'h7bc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17340; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23484 = 12'h7bc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20412; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26556 = 12'h7bc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23484; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1980 = io_valid_in ? _GEN_26556 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1980 = 12'h7bc == _T_2[11:0] ? image_1980 : _GEN_1979; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5053 = 12'h7bd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8125 = 12'h7bd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5053; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11197 = 12'h7bd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8125; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14269 = 12'h7bd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11197; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17341 = 12'h7bd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14269; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20413 = 12'h7bd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17341; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23485 = 12'h7bd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20413; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26557 = 12'h7bd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23485; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1981 = io_valid_in ? _GEN_26557 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1981 = 12'h7bd == _T_2[11:0] ? image_1981 : _GEN_1980; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5054 = 12'h7be == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8126 = 12'h7be == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5054; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11198 = 12'h7be == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8126; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14270 = 12'h7be == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11198; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17342 = 12'h7be == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14270; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20414 = 12'h7be == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17342; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23486 = 12'h7be == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20414; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26558 = 12'h7be == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23486; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1982 = io_valid_in ? _GEN_26558 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1982 = 12'h7be == _T_2[11:0] ? image_1982 : _GEN_1981; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5055 = 12'h7bf == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8127 = 12'h7bf == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5055; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11199 = 12'h7bf == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8127; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14271 = 12'h7bf == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11199; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17343 = 12'h7bf == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14271; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20415 = 12'h7bf == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17343; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23487 = 12'h7bf == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20415; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26559 = 12'h7bf == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23487; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1983 = io_valid_in ? _GEN_26559 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1983 = 12'h7bf == _T_2[11:0] ? image_1983 : _GEN_1982; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5056 = 12'h7c0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8128 = 12'h7c0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5056; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11200 = 12'h7c0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8128; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14272 = 12'h7c0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11200; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17344 = 12'h7c0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14272; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20416 = 12'h7c0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17344; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23488 = 12'h7c0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20416; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26560 = 12'h7c0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23488; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1984 = io_valid_in ? _GEN_26560 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1984 = 12'h7c0 == _T_2[11:0] ? image_1984 : _GEN_1983; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5057 = 12'h7c1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8129 = 12'h7c1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5057; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11201 = 12'h7c1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8129; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14273 = 12'h7c1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11201; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17345 = 12'h7c1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14273; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20417 = 12'h7c1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17345; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23489 = 12'h7c1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20417; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26561 = 12'h7c1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23489; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1985 = io_valid_in ? _GEN_26561 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1985 = 12'h7c1 == _T_2[11:0] ? image_1985 : _GEN_1984; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5058 = 12'h7c2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8130 = 12'h7c2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5058; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11202 = 12'h7c2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8130; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14274 = 12'h7c2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11202; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17346 = 12'h7c2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14274; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20418 = 12'h7c2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17346; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23490 = 12'h7c2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20418; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26562 = 12'h7c2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23490; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1986 = io_valid_in ? _GEN_26562 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1986 = 12'h7c2 == _T_2[11:0] ? image_1986 : _GEN_1985; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5059 = 12'h7c3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8131 = 12'h7c3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5059; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11203 = 12'h7c3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8131; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14275 = 12'h7c3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11203; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17347 = 12'h7c3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14275; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20419 = 12'h7c3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17347; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23491 = 12'h7c3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20419; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26563 = 12'h7c3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23491; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1987 = io_valid_in ? _GEN_26563 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1987 = 12'h7c3 == _T_2[11:0] ? image_1987 : _GEN_1986; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5060 = 12'h7c4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8132 = 12'h7c4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5060; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11204 = 12'h7c4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8132; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14276 = 12'h7c4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11204; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17348 = 12'h7c4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14276; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20420 = 12'h7c4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17348; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23492 = 12'h7c4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20420; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26564 = 12'h7c4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23492; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1988 = io_valid_in ? _GEN_26564 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1988 = 12'h7c4 == _T_2[11:0] ? image_1988 : _GEN_1987; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5061 = 12'h7c5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8133 = 12'h7c5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5061; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11205 = 12'h7c5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8133; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14277 = 12'h7c5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11205; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17349 = 12'h7c5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14277; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20421 = 12'h7c5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17349; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23493 = 12'h7c5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20421; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26565 = 12'h7c5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23493; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1989 = io_valid_in ? _GEN_26565 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1989 = 12'h7c5 == _T_2[11:0] ? image_1989 : _GEN_1988; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5062 = 12'h7c6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8134 = 12'h7c6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5062; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11206 = 12'h7c6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8134; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14278 = 12'h7c6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11206; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17350 = 12'h7c6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14278; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20422 = 12'h7c6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17350; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23494 = 12'h7c6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20422; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26566 = 12'h7c6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23494; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1990 = io_valid_in ? _GEN_26566 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1990 = 12'h7c6 == _T_2[11:0] ? image_1990 : _GEN_1989; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5063 = 12'h7c7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8135 = 12'h7c7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5063; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11207 = 12'h7c7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8135; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14279 = 12'h7c7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11207; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17351 = 12'h7c7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14279; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20423 = 12'h7c7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17351; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23495 = 12'h7c7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20423; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26567 = 12'h7c7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23495; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1991 = io_valid_in ? _GEN_26567 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1991 = 12'h7c7 == _T_2[11:0] ? image_1991 : _GEN_1990; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5064 = 12'h7c8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8136 = 12'h7c8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5064; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11208 = 12'h7c8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8136; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14280 = 12'h7c8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11208; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17352 = 12'h7c8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14280; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20424 = 12'h7c8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17352; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23496 = 12'h7c8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20424; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26568 = 12'h7c8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23496; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1992 = io_valid_in ? _GEN_26568 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1992 = 12'h7c8 == _T_2[11:0] ? image_1992 : _GEN_1991; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5065 = 12'h7c9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8137 = 12'h7c9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5065; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11209 = 12'h7c9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8137; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14281 = 12'h7c9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11209; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17353 = 12'h7c9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14281; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20425 = 12'h7c9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17353; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23497 = 12'h7c9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20425; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26569 = 12'h7c9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23497; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1993 = io_valid_in ? _GEN_26569 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1993 = 12'h7c9 == _T_2[11:0] ? image_1993 : _GEN_1992; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5066 = 12'h7ca == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8138 = 12'h7ca == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5066; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11210 = 12'h7ca == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8138; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14282 = 12'h7ca == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11210; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17354 = 12'h7ca == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14282; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20426 = 12'h7ca == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17354; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23498 = 12'h7ca == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20426; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26570 = 12'h7ca == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23498; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1994 = io_valid_in ? _GEN_26570 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1994 = 12'h7ca == _T_2[11:0] ? image_1994 : _GEN_1993; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5067 = 12'h7cb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8139 = 12'h7cb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5067; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11211 = 12'h7cb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8139; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14283 = 12'h7cb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11211; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17355 = 12'h7cb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14283; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20427 = 12'h7cb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17355; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23499 = 12'h7cb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20427; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26571 = 12'h7cb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23499; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1995 = io_valid_in ? _GEN_26571 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1995 = 12'h7cb == _T_2[11:0] ? image_1995 : _GEN_1994; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5068 = 12'h7cc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8140 = 12'h7cc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5068; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11212 = 12'h7cc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8140; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14284 = 12'h7cc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11212; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17356 = 12'h7cc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14284; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20428 = 12'h7cc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17356; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23500 = 12'h7cc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20428; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26572 = 12'h7cc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23500; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1996 = io_valid_in ? _GEN_26572 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1996 = 12'h7cc == _T_2[11:0] ? image_1996 : _GEN_1995; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5069 = 12'h7cd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8141 = 12'h7cd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5069; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11213 = 12'h7cd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8141; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14285 = 12'h7cd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11213; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17357 = 12'h7cd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14285; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20429 = 12'h7cd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17357; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23501 = 12'h7cd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20429; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26573 = 12'h7cd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23501; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1997 = io_valid_in ? _GEN_26573 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1997 = 12'h7cd == _T_2[11:0] ? image_1997 : _GEN_1996; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5070 = 12'h7ce == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8142 = 12'h7ce == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5070; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11214 = 12'h7ce == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8142; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14286 = 12'h7ce == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11214; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17358 = 12'h7ce == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14286; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20430 = 12'h7ce == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17358; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23502 = 12'h7ce == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20430; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26574 = 12'h7ce == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23502; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1998 = io_valid_in ? _GEN_26574 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1998 = 12'h7ce == _T_2[11:0] ? image_1998 : _GEN_1997; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5071 = 12'h7cf == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8143 = 12'h7cf == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5071; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11215 = 12'h7cf == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8143; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14287 = 12'h7cf == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11215; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17359 = 12'h7cf == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14287; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20431 = 12'h7cf == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17359; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23503 = 12'h7cf == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20431; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26575 = 12'h7cf == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23503; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1999 = io_valid_in ? _GEN_26575 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1999 = 12'h7cf == _T_2[11:0] ? image_1999 : _GEN_1998; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5072 = 12'h7d0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8144 = 12'h7d0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5072; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11216 = 12'h7d0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8144; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14288 = 12'h7d0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11216; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17360 = 12'h7d0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14288; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20432 = 12'h7d0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17360; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23504 = 12'h7d0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20432; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26576 = 12'h7d0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23504; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2000 = io_valid_in ? _GEN_26576 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2000 = 12'h7d0 == _T_2[11:0] ? image_2000 : _GEN_1999; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5073 = 12'h7d1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8145 = 12'h7d1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5073; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11217 = 12'h7d1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8145; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14289 = 12'h7d1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11217; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17361 = 12'h7d1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14289; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20433 = 12'h7d1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17361; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23505 = 12'h7d1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20433; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26577 = 12'h7d1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23505; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2001 = io_valid_in ? _GEN_26577 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2001 = 12'h7d1 == _T_2[11:0] ? image_2001 : _GEN_2000; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5074 = 12'h7d2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8146 = 12'h7d2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5074; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11218 = 12'h7d2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8146; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14290 = 12'h7d2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11218; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17362 = 12'h7d2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14290; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20434 = 12'h7d2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17362; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23506 = 12'h7d2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20434; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26578 = 12'h7d2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23506; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2002 = io_valid_in ? _GEN_26578 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2002 = 12'h7d2 == _T_2[11:0] ? image_2002 : _GEN_2001; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5075 = 12'h7d3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8147 = 12'h7d3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5075; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11219 = 12'h7d3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8147; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14291 = 12'h7d3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11219; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17363 = 12'h7d3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14291; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20435 = 12'h7d3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17363; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23507 = 12'h7d3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20435; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26579 = 12'h7d3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23507; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2003 = io_valid_in ? _GEN_26579 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2003 = 12'h7d3 == _T_2[11:0] ? image_2003 : _GEN_2002; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5076 = 12'h7d4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8148 = 12'h7d4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5076; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11220 = 12'h7d4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8148; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14292 = 12'h7d4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11220; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17364 = 12'h7d4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14292; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20436 = 12'h7d4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17364; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23508 = 12'h7d4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20436; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26580 = 12'h7d4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23508; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2004 = io_valid_in ? _GEN_26580 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2004 = 12'h7d4 == _T_2[11:0] ? image_2004 : _GEN_2003; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5077 = 12'h7d5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8149 = 12'h7d5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5077; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11221 = 12'h7d5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8149; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14293 = 12'h7d5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11221; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17365 = 12'h7d5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14293; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20437 = 12'h7d5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17365; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23509 = 12'h7d5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20437; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26581 = 12'h7d5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23509; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2005 = io_valid_in ? _GEN_26581 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2005 = 12'h7d5 == _T_2[11:0] ? image_2005 : _GEN_2004; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5078 = 12'h7d6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8150 = 12'h7d6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5078; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11222 = 12'h7d6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8150; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14294 = 12'h7d6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11222; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17366 = 12'h7d6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14294; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20438 = 12'h7d6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17366; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23510 = 12'h7d6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20438; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26582 = 12'h7d6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23510; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2006 = io_valid_in ? _GEN_26582 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2006 = 12'h7d6 == _T_2[11:0] ? image_2006 : _GEN_2005; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5079 = 12'h7d7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8151 = 12'h7d7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5079; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11223 = 12'h7d7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8151; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14295 = 12'h7d7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11223; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17367 = 12'h7d7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14295; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20439 = 12'h7d7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17367; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23511 = 12'h7d7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20439; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26583 = 12'h7d7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23511; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2007 = io_valid_in ? _GEN_26583 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2007 = 12'h7d7 == _T_2[11:0] ? image_2007 : _GEN_2006; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5080 = 12'h7d8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8152 = 12'h7d8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5080; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11224 = 12'h7d8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8152; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14296 = 12'h7d8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11224; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17368 = 12'h7d8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14296; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20440 = 12'h7d8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17368; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23512 = 12'h7d8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20440; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26584 = 12'h7d8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23512; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2008 = io_valid_in ? _GEN_26584 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2008 = 12'h7d8 == _T_2[11:0] ? image_2008 : _GEN_2007; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5081 = 12'h7d9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8153 = 12'h7d9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5081; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11225 = 12'h7d9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8153; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14297 = 12'h7d9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11225; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17369 = 12'h7d9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14297; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20441 = 12'h7d9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17369; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23513 = 12'h7d9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20441; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26585 = 12'h7d9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23513; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2009 = io_valid_in ? _GEN_26585 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2009 = 12'h7d9 == _T_2[11:0] ? image_2009 : _GEN_2008; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5082 = 12'h7da == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8154 = 12'h7da == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5082; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11226 = 12'h7da == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8154; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14298 = 12'h7da == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11226; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17370 = 12'h7da == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14298; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20442 = 12'h7da == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17370; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23514 = 12'h7da == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20442; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26586 = 12'h7da == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23514; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2010 = io_valid_in ? _GEN_26586 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2010 = 12'h7da == _T_2[11:0] ? image_2010 : _GEN_2009; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5083 = 12'h7db == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8155 = 12'h7db == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5083; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11227 = 12'h7db == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8155; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14299 = 12'h7db == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11227; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17371 = 12'h7db == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14299; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20443 = 12'h7db == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17371; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23515 = 12'h7db == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20443; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26587 = 12'h7db == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23515; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2011 = io_valid_in ? _GEN_26587 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2011 = 12'h7db == _T_2[11:0] ? image_2011 : _GEN_2010; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5084 = 12'h7dc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8156 = 12'h7dc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5084; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11228 = 12'h7dc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8156; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14300 = 12'h7dc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11228; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17372 = 12'h7dc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14300; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20444 = 12'h7dc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17372; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23516 = 12'h7dc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20444; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26588 = 12'h7dc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23516; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2012 = io_valid_in ? _GEN_26588 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2012 = 12'h7dc == _T_2[11:0] ? image_2012 : _GEN_2011; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5085 = 12'h7dd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8157 = 12'h7dd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5085; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11229 = 12'h7dd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8157; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14301 = 12'h7dd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11229; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17373 = 12'h7dd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14301; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20445 = 12'h7dd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17373; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23517 = 12'h7dd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20445; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26589 = 12'h7dd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23517; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2013 = io_valid_in ? _GEN_26589 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2013 = 12'h7dd == _T_2[11:0] ? image_2013 : _GEN_2012; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5086 = 12'h7de == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8158 = 12'h7de == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5086; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11230 = 12'h7de == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8158; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14302 = 12'h7de == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11230; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17374 = 12'h7de == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14302; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20446 = 12'h7de == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17374; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23518 = 12'h7de == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20446; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26590 = 12'h7de == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23518; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2014 = io_valid_in ? _GEN_26590 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2014 = 12'h7de == _T_2[11:0] ? image_2014 : _GEN_2013; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5087 = 12'h7df == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8159 = 12'h7df == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5087; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11231 = 12'h7df == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8159; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14303 = 12'h7df == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11231; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17375 = 12'h7df == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14303; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20447 = 12'h7df == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17375; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23519 = 12'h7df == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20447; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26591 = 12'h7df == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23519; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2015 = io_valid_in ? _GEN_26591 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2015 = 12'h7df == _T_2[11:0] ? image_2015 : _GEN_2014; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5088 = 12'h7e0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8160 = 12'h7e0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5088; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11232 = 12'h7e0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8160; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14304 = 12'h7e0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11232; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17376 = 12'h7e0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14304; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20448 = 12'h7e0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17376; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23520 = 12'h7e0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20448; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26592 = 12'h7e0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23520; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2016 = io_valid_in ? _GEN_26592 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2016 = 12'h7e0 == _T_2[11:0] ? image_2016 : _GEN_2015; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5089 = 12'h7e1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8161 = 12'h7e1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5089; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11233 = 12'h7e1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8161; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14305 = 12'h7e1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11233; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17377 = 12'h7e1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14305; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20449 = 12'h7e1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17377; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23521 = 12'h7e1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20449; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26593 = 12'h7e1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23521; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2017 = io_valid_in ? _GEN_26593 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2017 = 12'h7e1 == _T_2[11:0] ? image_2017 : _GEN_2016; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5090 = 12'h7e2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8162 = 12'h7e2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5090; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11234 = 12'h7e2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8162; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14306 = 12'h7e2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11234; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17378 = 12'h7e2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14306; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20450 = 12'h7e2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17378; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23522 = 12'h7e2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20450; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26594 = 12'h7e2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23522; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2018 = io_valid_in ? _GEN_26594 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2018 = 12'h7e2 == _T_2[11:0] ? image_2018 : _GEN_2017; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5091 = 12'h7e3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8163 = 12'h7e3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5091; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11235 = 12'h7e3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8163; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14307 = 12'h7e3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11235; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17379 = 12'h7e3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14307; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20451 = 12'h7e3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17379; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23523 = 12'h7e3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20451; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26595 = 12'h7e3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23523; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2019 = io_valid_in ? _GEN_26595 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2019 = 12'h7e3 == _T_2[11:0] ? image_2019 : _GEN_2018; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5092 = 12'h7e4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8164 = 12'h7e4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5092; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11236 = 12'h7e4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8164; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14308 = 12'h7e4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11236; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17380 = 12'h7e4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14308; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20452 = 12'h7e4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17380; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23524 = 12'h7e4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20452; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26596 = 12'h7e4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23524; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2020 = io_valid_in ? _GEN_26596 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2020 = 12'h7e4 == _T_2[11:0] ? image_2020 : _GEN_2019; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5093 = 12'h7e5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8165 = 12'h7e5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5093; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11237 = 12'h7e5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8165; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14309 = 12'h7e5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11237; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17381 = 12'h7e5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14309; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20453 = 12'h7e5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17381; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23525 = 12'h7e5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20453; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26597 = 12'h7e5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23525; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2021 = io_valid_in ? _GEN_26597 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2021 = 12'h7e5 == _T_2[11:0] ? image_2021 : _GEN_2020; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5094 = 12'h7e6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8166 = 12'h7e6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5094; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11238 = 12'h7e6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8166; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14310 = 12'h7e6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11238; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17382 = 12'h7e6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14310; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20454 = 12'h7e6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17382; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23526 = 12'h7e6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20454; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26598 = 12'h7e6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23526; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2022 = io_valid_in ? _GEN_26598 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2022 = 12'h7e6 == _T_2[11:0] ? image_2022 : _GEN_2021; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5095 = 12'h7e7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8167 = 12'h7e7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5095; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11239 = 12'h7e7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8167; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14311 = 12'h7e7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11239; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17383 = 12'h7e7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14311; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20455 = 12'h7e7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17383; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23527 = 12'h7e7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20455; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26599 = 12'h7e7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23527; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2023 = io_valid_in ? _GEN_26599 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2023 = 12'h7e7 == _T_2[11:0] ? image_2023 : _GEN_2022; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5096 = 12'h7e8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8168 = 12'h7e8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5096; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11240 = 12'h7e8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8168; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14312 = 12'h7e8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11240; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17384 = 12'h7e8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14312; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20456 = 12'h7e8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17384; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23528 = 12'h7e8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20456; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26600 = 12'h7e8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23528; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2024 = io_valid_in ? _GEN_26600 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2024 = 12'h7e8 == _T_2[11:0] ? image_2024 : _GEN_2023; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5097 = 12'h7e9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8169 = 12'h7e9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5097; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11241 = 12'h7e9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8169; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14313 = 12'h7e9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11241; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17385 = 12'h7e9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14313; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20457 = 12'h7e9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17385; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23529 = 12'h7e9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20457; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26601 = 12'h7e9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23529; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2025 = io_valid_in ? _GEN_26601 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2025 = 12'h7e9 == _T_2[11:0] ? image_2025 : _GEN_2024; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5098 = 12'h7ea == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8170 = 12'h7ea == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5098; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11242 = 12'h7ea == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8170; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14314 = 12'h7ea == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11242; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17386 = 12'h7ea == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14314; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20458 = 12'h7ea == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17386; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23530 = 12'h7ea == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20458; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26602 = 12'h7ea == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23530; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2026 = io_valid_in ? _GEN_26602 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2026 = 12'h7ea == _T_2[11:0] ? image_2026 : _GEN_2025; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5099 = 12'h7eb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8171 = 12'h7eb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5099; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11243 = 12'h7eb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8171; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14315 = 12'h7eb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11243; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17387 = 12'h7eb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14315; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20459 = 12'h7eb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17387; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23531 = 12'h7eb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20459; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26603 = 12'h7eb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23531; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2027 = io_valid_in ? _GEN_26603 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2027 = 12'h7eb == _T_2[11:0] ? image_2027 : _GEN_2026; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5100 = 12'h7ec == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8172 = 12'h7ec == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5100; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11244 = 12'h7ec == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8172; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14316 = 12'h7ec == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11244; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17388 = 12'h7ec == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14316; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20460 = 12'h7ec == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17388; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23532 = 12'h7ec == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20460; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26604 = 12'h7ec == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23532; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2028 = io_valid_in ? _GEN_26604 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2028 = 12'h7ec == _T_2[11:0] ? image_2028 : _GEN_2027; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5101 = 12'h7ed == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8173 = 12'h7ed == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5101; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11245 = 12'h7ed == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8173; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14317 = 12'h7ed == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11245; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17389 = 12'h7ed == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14317; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20461 = 12'h7ed == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17389; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23533 = 12'h7ed == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20461; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26605 = 12'h7ed == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23533; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2029 = io_valid_in ? _GEN_26605 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2029 = 12'h7ed == _T_2[11:0] ? image_2029 : _GEN_2028; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5102 = 12'h7ee == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8174 = 12'h7ee == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5102; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11246 = 12'h7ee == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8174; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14318 = 12'h7ee == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11246; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17390 = 12'h7ee == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14318; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20462 = 12'h7ee == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17390; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23534 = 12'h7ee == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20462; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26606 = 12'h7ee == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23534; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2030 = io_valid_in ? _GEN_26606 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2030 = 12'h7ee == _T_2[11:0] ? image_2030 : _GEN_2029; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5103 = 12'h7ef == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8175 = 12'h7ef == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5103; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11247 = 12'h7ef == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8175; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14319 = 12'h7ef == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11247; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17391 = 12'h7ef == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14319; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20463 = 12'h7ef == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17391; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23535 = 12'h7ef == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20463; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26607 = 12'h7ef == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23535; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2031 = io_valid_in ? _GEN_26607 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2031 = 12'h7ef == _T_2[11:0] ? image_2031 : _GEN_2030; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5104 = 12'h7f0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8176 = 12'h7f0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5104; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11248 = 12'h7f0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8176; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14320 = 12'h7f0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11248; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17392 = 12'h7f0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14320; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20464 = 12'h7f0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17392; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23536 = 12'h7f0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20464; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26608 = 12'h7f0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23536; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2032 = io_valid_in ? _GEN_26608 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2032 = 12'h7f0 == _T_2[11:0] ? image_2032 : _GEN_2031; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5105 = 12'h7f1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8177 = 12'h7f1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5105; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11249 = 12'h7f1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8177; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14321 = 12'h7f1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11249; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17393 = 12'h7f1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14321; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20465 = 12'h7f1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17393; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23537 = 12'h7f1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20465; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26609 = 12'h7f1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23537; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2033 = io_valid_in ? _GEN_26609 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2033 = 12'h7f1 == _T_2[11:0] ? image_2033 : _GEN_2032; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5106 = 12'h7f2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8178 = 12'h7f2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5106; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11250 = 12'h7f2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8178; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14322 = 12'h7f2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11250; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17394 = 12'h7f2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14322; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20466 = 12'h7f2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17394; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23538 = 12'h7f2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20466; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26610 = 12'h7f2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23538; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2034 = io_valid_in ? _GEN_26610 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2034 = 12'h7f2 == _T_2[11:0] ? image_2034 : _GEN_2033; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5107 = 12'h7f3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8179 = 12'h7f3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5107; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11251 = 12'h7f3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8179; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14323 = 12'h7f3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11251; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17395 = 12'h7f3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14323; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20467 = 12'h7f3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17395; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23539 = 12'h7f3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20467; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26611 = 12'h7f3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23539; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2035 = io_valid_in ? _GEN_26611 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2035 = 12'h7f3 == _T_2[11:0] ? image_2035 : _GEN_2034; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5108 = 12'h7f4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8180 = 12'h7f4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5108; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11252 = 12'h7f4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8180; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14324 = 12'h7f4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11252; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17396 = 12'h7f4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14324; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20468 = 12'h7f4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17396; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23540 = 12'h7f4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20468; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26612 = 12'h7f4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23540; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2036 = io_valid_in ? _GEN_26612 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2036 = 12'h7f4 == _T_2[11:0] ? image_2036 : _GEN_2035; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5109 = 12'h7f5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8181 = 12'h7f5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5109; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11253 = 12'h7f5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8181; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14325 = 12'h7f5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11253; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17397 = 12'h7f5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14325; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20469 = 12'h7f5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17397; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23541 = 12'h7f5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20469; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26613 = 12'h7f5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23541; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2037 = io_valid_in ? _GEN_26613 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2037 = 12'h7f5 == _T_2[11:0] ? image_2037 : _GEN_2036; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5110 = 12'h7f6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8182 = 12'h7f6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5110; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11254 = 12'h7f6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8182; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14326 = 12'h7f6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11254; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17398 = 12'h7f6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14326; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20470 = 12'h7f6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17398; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23542 = 12'h7f6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20470; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26614 = 12'h7f6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23542; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2038 = io_valid_in ? _GEN_26614 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2038 = 12'h7f6 == _T_2[11:0] ? image_2038 : _GEN_2037; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5111 = 12'h7f7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8183 = 12'h7f7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5111; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11255 = 12'h7f7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8183; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14327 = 12'h7f7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11255; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17399 = 12'h7f7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14327; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20471 = 12'h7f7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17399; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23543 = 12'h7f7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20471; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26615 = 12'h7f7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23543; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2039 = io_valid_in ? _GEN_26615 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2039 = 12'h7f7 == _T_2[11:0] ? image_2039 : _GEN_2038; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5112 = 12'h7f8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8184 = 12'h7f8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5112; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11256 = 12'h7f8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8184; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14328 = 12'h7f8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11256; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17400 = 12'h7f8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14328; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20472 = 12'h7f8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17400; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23544 = 12'h7f8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20472; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26616 = 12'h7f8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23544; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2040 = io_valid_in ? _GEN_26616 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2040 = 12'h7f8 == _T_2[11:0] ? image_2040 : _GEN_2039; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5113 = 12'h7f9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8185 = 12'h7f9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5113; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11257 = 12'h7f9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8185; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14329 = 12'h7f9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11257; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17401 = 12'h7f9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14329; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20473 = 12'h7f9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17401; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23545 = 12'h7f9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20473; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26617 = 12'h7f9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23545; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2041 = io_valid_in ? _GEN_26617 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2041 = 12'h7f9 == _T_2[11:0] ? image_2041 : _GEN_2040; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5114 = 12'h7fa == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8186 = 12'h7fa == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5114; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11258 = 12'h7fa == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8186; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14330 = 12'h7fa == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11258; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17402 = 12'h7fa == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14330; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20474 = 12'h7fa == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17402; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23546 = 12'h7fa == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20474; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26618 = 12'h7fa == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23546; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2042 = io_valid_in ? _GEN_26618 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2042 = 12'h7fa == _T_2[11:0] ? image_2042 : _GEN_2041; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5115 = 12'h7fb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8187 = 12'h7fb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5115; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11259 = 12'h7fb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8187; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14331 = 12'h7fb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11259; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17403 = 12'h7fb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14331; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20475 = 12'h7fb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17403; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23547 = 12'h7fb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20475; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26619 = 12'h7fb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23547; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2043 = io_valid_in ? _GEN_26619 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2043 = 12'h7fb == _T_2[11:0] ? image_2043 : _GEN_2042; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5116 = 12'h7fc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8188 = 12'h7fc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5116; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11260 = 12'h7fc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8188; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14332 = 12'h7fc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11260; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17404 = 12'h7fc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14332; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20476 = 12'h7fc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17404; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23548 = 12'h7fc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20476; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26620 = 12'h7fc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23548; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2044 = io_valid_in ? _GEN_26620 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2044 = 12'h7fc == _T_2[11:0] ? image_2044 : _GEN_2043; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5117 = 12'h7fd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8189 = 12'h7fd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5117; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11261 = 12'h7fd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8189; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14333 = 12'h7fd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11261; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17405 = 12'h7fd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14333; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20477 = 12'h7fd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17405; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23549 = 12'h7fd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20477; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26621 = 12'h7fd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23549; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2045 = io_valid_in ? _GEN_26621 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2045 = 12'h7fd == _T_2[11:0] ? image_2045 : _GEN_2044; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5118 = 12'h7fe == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8190 = 12'h7fe == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5118; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11262 = 12'h7fe == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8190; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14334 = 12'h7fe == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11262; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17406 = 12'h7fe == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14334; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20478 = 12'h7fe == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17406; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23550 = 12'h7fe == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20478; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26622 = 12'h7fe == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23550; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2046 = io_valid_in ? _GEN_26622 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2046 = 12'h7fe == _T_2[11:0] ? image_2046 : _GEN_2045; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5119 = 12'h7ff == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8191 = 12'h7ff == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5119; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11263 = 12'h7ff == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8191; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14335 = 12'h7ff == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11263; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17407 = 12'h7ff == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14335; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20479 = 12'h7ff == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17407; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23551 = 12'h7ff == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20479; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26623 = 12'h7ff == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23551; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2047 = io_valid_in ? _GEN_26623 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2047 = 12'h7ff == _T_2[11:0] ? image_2047 : _GEN_2046; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5120 = 12'h800 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8192 = 12'h800 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5120; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11264 = 12'h800 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8192; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14336 = 12'h800 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11264; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17408 = 12'h800 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14336; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20480 = 12'h800 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17408; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23552 = 12'h800 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20480; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26624 = 12'h800 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23552; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2048 = io_valid_in ? _GEN_26624 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2048 = 12'h800 == _T_2[11:0] ? image_2048 : _GEN_2047; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5121 = 12'h801 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8193 = 12'h801 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5121; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11265 = 12'h801 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8193; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14337 = 12'h801 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11265; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17409 = 12'h801 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14337; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20481 = 12'h801 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17409; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23553 = 12'h801 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20481; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26625 = 12'h801 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23553; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2049 = io_valid_in ? _GEN_26625 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2049 = 12'h801 == _T_2[11:0] ? image_2049 : _GEN_2048; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5122 = 12'h802 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8194 = 12'h802 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5122; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11266 = 12'h802 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8194; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14338 = 12'h802 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11266; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17410 = 12'h802 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14338; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20482 = 12'h802 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17410; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23554 = 12'h802 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20482; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26626 = 12'h802 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23554; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2050 = io_valid_in ? _GEN_26626 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2050 = 12'h802 == _T_2[11:0] ? image_2050 : _GEN_2049; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5123 = 12'h803 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8195 = 12'h803 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5123; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11267 = 12'h803 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8195; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14339 = 12'h803 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11267; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17411 = 12'h803 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14339; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20483 = 12'h803 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17411; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23555 = 12'h803 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20483; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26627 = 12'h803 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23555; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2051 = io_valid_in ? _GEN_26627 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2051 = 12'h803 == _T_2[11:0] ? image_2051 : _GEN_2050; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5124 = 12'h804 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8196 = 12'h804 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5124; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11268 = 12'h804 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8196; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14340 = 12'h804 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11268; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17412 = 12'h804 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14340; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20484 = 12'h804 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17412; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23556 = 12'h804 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20484; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26628 = 12'h804 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23556; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2052 = io_valid_in ? _GEN_26628 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2052 = 12'h804 == _T_2[11:0] ? image_2052 : _GEN_2051; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5125 = 12'h805 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8197 = 12'h805 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5125; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11269 = 12'h805 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8197; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14341 = 12'h805 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11269; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17413 = 12'h805 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14341; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20485 = 12'h805 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17413; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23557 = 12'h805 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20485; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26629 = 12'h805 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23557; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2053 = io_valid_in ? _GEN_26629 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2053 = 12'h805 == _T_2[11:0] ? image_2053 : _GEN_2052; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5126 = 12'h806 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8198 = 12'h806 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5126; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11270 = 12'h806 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8198; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14342 = 12'h806 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11270; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17414 = 12'h806 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14342; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20486 = 12'h806 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17414; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23558 = 12'h806 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20486; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26630 = 12'h806 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23558; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2054 = io_valid_in ? _GEN_26630 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2054 = 12'h806 == _T_2[11:0] ? image_2054 : _GEN_2053; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5127 = 12'h807 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8199 = 12'h807 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5127; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11271 = 12'h807 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8199; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14343 = 12'h807 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11271; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17415 = 12'h807 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14343; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20487 = 12'h807 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17415; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23559 = 12'h807 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20487; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26631 = 12'h807 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23559; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2055 = io_valid_in ? _GEN_26631 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2055 = 12'h807 == _T_2[11:0] ? image_2055 : _GEN_2054; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5128 = 12'h808 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8200 = 12'h808 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5128; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11272 = 12'h808 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8200; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14344 = 12'h808 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11272; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17416 = 12'h808 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14344; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20488 = 12'h808 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17416; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23560 = 12'h808 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20488; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26632 = 12'h808 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23560; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2056 = io_valid_in ? _GEN_26632 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2056 = 12'h808 == _T_2[11:0] ? image_2056 : _GEN_2055; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5129 = 12'h809 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8201 = 12'h809 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5129; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11273 = 12'h809 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8201; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14345 = 12'h809 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11273; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17417 = 12'h809 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14345; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20489 = 12'h809 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17417; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23561 = 12'h809 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20489; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26633 = 12'h809 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23561; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2057 = io_valid_in ? _GEN_26633 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2057 = 12'h809 == _T_2[11:0] ? image_2057 : _GEN_2056; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5130 = 12'h80a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8202 = 12'h80a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5130; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11274 = 12'h80a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8202; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14346 = 12'h80a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11274; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17418 = 12'h80a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14346; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20490 = 12'h80a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17418; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23562 = 12'h80a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20490; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26634 = 12'h80a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23562; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2058 = io_valid_in ? _GEN_26634 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2058 = 12'h80a == _T_2[11:0] ? image_2058 : _GEN_2057; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5131 = 12'h80b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8203 = 12'h80b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5131; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11275 = 12'h80b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8203; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14347 = 12'h80b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11275; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17419 = 12'h80b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14347; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20491 = 12'h80b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17419; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23563 = 12'h80b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20491; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26635 = 12'h80b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23563; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2059 = io_valid_in ? _GEN_26635 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2059 = 12'h80b == _T_2[11:0] ? image_2059 : _GEN_2058; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5132 = 12'h80c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8204 = 12'h80c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5132; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11276 = 12'h80c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8204; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14348 = 12'h80c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11276; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17420 = 12'h80c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14348; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20492 = 12'h80c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17420; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23564 = 12'h80c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20492; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26636 = 12'h80c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23564; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2060 = io_valid_in ? _GEN_26636 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2060 = 12'h80c == _T_2[11:0] ? image_2060 : _GEN_2059; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5133 = 12'h80d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8205 = 12'h80d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5133; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11277 = 12'h80d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8205; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14349 = 12'h80d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11277; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17421 = 12'h80d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14349; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20493 = 12'h80d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17421; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23565 = 12'h80d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20493; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26637 = 12'h80d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23565; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2061 = io_valid_in ? _GEN_26637 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2061 = 12'h80d == _T_2[11:0] ? image_2061 : _GEN_2060; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5134 = 12'h80e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8206 = 12'h80e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5134; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11278 = 12'h80e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8206; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14350 = 12'h80e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11278; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17422 = 12'h80e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14350; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20494 = 12'h80e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17422; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23566 = 12'h80e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20494; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26638 = 12'h80e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23566; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2062 = io_valid_in ? _GEN_26638 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2062 = 12'h80e == _T_2[11:0] ? image_2062 : _GEN_2061; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5135 = 12'h80f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8207 = 12'h80f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5135; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11279 = 12'h80f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8207; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14351 = 12'h80f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11279; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17423 = 12'h80f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14351; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20495 = 12'h80f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17423; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23567 = 12'h80f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20495; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26639 = 12'h80f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23567; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2063 = io_valid_in ? _GEN_26639 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2063 = 12'h80f == _T_2[11:0] ? image_2063 : _GEN_2062; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5136 = 12'h810 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8208 = 12'h810 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5136; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11280 = 12'h810 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8208; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14352 = 12'h810 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11280; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17424 = 12'h810 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14352; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20496 = 12'h810 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17424; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23568 = 12'h810 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20496; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26640 = 12'h810 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23568; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2064 = io_valid_in ? _GEN_26640 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2064 = 12'h810 == _T_2[11:0] ? image_2064 : _GEN_2063; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5137 = 12'h811 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8209 = 12'h811 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5137; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11281 = 12'h811 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8209; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14353 = 12'h811 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11281; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17425 = 12'h811 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14353; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20497 = 12'h811 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17425; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23569 = 12'h811 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20497; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26641 = 12'h811 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23569; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2065 = io_valid_in ? _GEN_26641 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2065 = 12'h811 == _T_2[11:0] ? image_2065 : _GEN_2064; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5138 = 12'h812 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8210 = 12'h812 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5138; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11282 = 12'h812 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8210; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14354 = 12'h812 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11282; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17426 = 12'h812 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14354; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20498 = 12'h812 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17426; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23570 = 12'h812 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20498; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26642 = 12'h812 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23570; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2066 = io_valid_in ? _GEN_26642 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2066 = 12'h812 == _T_2[11:0] ? image_2066 : _GEN_2065; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5139 = 12'h813 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8211 = 12'h813 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5139; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11283 = 12'h813 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8211; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14355 = 12'h813 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11283; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17427 = 12'h813 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14355; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20499 = 12'h813 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17427; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23571 = 12'h813 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20499; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26643 = 12'h813 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23571; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2067 = io_valid_in ? _GEN_26643 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2067 = 12'h813 == _T_2[11:0] ? image_2067 : _GEN_2066; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5140 = 12'h814 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8212 = 12'h814 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5140; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11284 = 12'h814 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8212; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14356 = 12'h814 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11284; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17428 = 12'h814 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14356; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20500 = 12'h814 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17428; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23572 = 12'h814 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20500; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26644 = 12'h814 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23572; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2068 = io_valid_in ? _GEN_26644 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2068 = 12'h814 == _T_2[11:0] ? image_2068 : _GEN_2067; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5141 = 12'h815 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8213 = 12'h815 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5141; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11285 = 12'h815 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8213; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14357 = 12'h815 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11285; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17429 = 12'h815 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14357; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20501 = 12'h815 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17429; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23573 = 12'h815 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20501; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26645 = 12'h815 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23573; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2069 = io_valid_in ? _GEN_26645 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2069 = 12'h815 == _T_2[11:0] ? image_2069 : _GEN_2068; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5142 = 12'h816 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8214 = 12'h816 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5142; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11286 = 12'h816 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8214; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14358 = 12'h816 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11286; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17430 = 12'h816 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14358; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20502 = 12'h816 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17430; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23574 = 12'h816 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20502; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26646 = 12'h816 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23574; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2070 = io_valid_in ? _GEN_26646 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2070 = 12'h816 == _T_2[11:0] ? image_2070 : _GEN_2069; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5143 = 12'h817 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8215 = 12'h817 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5143; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11287 = 12'h817 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8215; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14359 = 12'h817 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11287; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17431 = 12'h817 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14359; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20503 = 12'h817 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17431; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23575 = 12'h817 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20503; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26647 = 12'h817 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23575; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2071 = io_valid_in ? _GEN_26647 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2071 = 12'h817 == _T_2[11:0] ? image_2071 : _GEN_2070; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5144 = 12'h818 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8216 = 12'h818 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5144; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11288 = 12'h818 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8216; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14360 = 12'h818 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11288; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17432 = 12'h818 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14360; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20504 = 12'h818 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17432; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23576 = 12'h818 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20504; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26648 = 12'h818 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23576; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2072 = io_valid_in ? _GEN_26648 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2072 = 12'h818 == _T_2[11:0] ? image_2072 : _GEN_2071; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5145 = 12'h819 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8217 = 12'h819 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5145; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11289 = 12'h819 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8217; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14361 = 12'h819 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11289; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17433 = 12'h819 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14361; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20505 = 12'h819 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17433; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23577 = 12'h819 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20505; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26649 = 12'h819 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23577; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2073 = io_valid_in ? _GEN_26649 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2073 = 12'h819 == _T_2[11:0] ? image_2073 : _GEN_2072; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5146 = 12'h81a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8218 = 12'h81a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5146; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11290 = 12'h81a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8218; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14362 = 12'h81a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11290; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17434 = 12'h81a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14362; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20506 = 12'h81a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17434; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23578 = 12'h81a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20506; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26650 = 12'h81a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23578; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2074 = io_valid_in ? _GEN_26650 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2074 = 12'h81a == _T_2[11:0] ? image_2074 : _GEN_2073; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5147 = 12'h81b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8219 = 12'h81b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5147; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11291 = 12'h81b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8219; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14363 = 12'h81b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11291; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17435 = 12'h81b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14363; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20507 = 12'h81b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17435; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23579 = 12'h81b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20507; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26651 = 12'h81b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23579; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2075 = io_valid_in ? _GEN_26651 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2075 = 12'h81b == _T_2[11:0] ? image_2075 : _GEN_2074; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5148 = 12'h81c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8220 = 12'h81c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5148; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11292 = 12'h81c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8220; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14364 = 12'h81c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11292; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17436 = 12'h81c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14364; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20508 = 12'h81c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17436; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23580 = 12'h81c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20508; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26652 = 12'h81c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23580; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2076 = io_valid_in ? _GEN_26652 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2076 = 12'h81c == _T_2[11:0] ? image_2076 : _GEN_2075; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5149 = 12'h81d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8221 = 12'h81d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5149; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11293 = 12'h81d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8221; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14365 = 12'h81d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11293; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17437 = 12'h81d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14365; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20509 = 12'h81d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17437; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23581 = 12'h81d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20509; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26653 = 12'h81d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23581; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2077 = io_valid_in ? _GEN_26653 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2077 = 12'h81d == _T_2[11:0] ? image_2077 : _GEN_2076; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5150 = 12'h81e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8222 = 12'h81e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5150; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11294 = 12'h81e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8222; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14366 = 12'h81e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11294; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17438 = 12'h81e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14366; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20510 = 12'h81e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17438; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23582 = 12'h81e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20510; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26654 = 12'h81e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23582; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2078 = io_valid_in ? _GEN_26654 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2078 = 12'h81e == _T_2[11:0] ? image_2078 : _GEN_2077; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5151 = 12'h81f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8223 = 12'h81f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5151; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11295 = 12'h81f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8223; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14367 = 12'h81f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11295; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17439 = 12'h81f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14367; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20511 = 12'h81f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17439; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23583 = 12'h81f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20511; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26655 = 12'h81f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23583; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2079 = io_valid_in ? _GEN_26655 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2079 = 12'h81f == _T_2[11:0] ? image_2079 : _GEN_2078; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5152 = 12'h820 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8224 = 12'h820 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5152; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11296 = 12'h820 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8224; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14368 = 12'h820 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11296; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17440 = 12'h820 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14368; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20512 = 12'h820 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17440; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23584 = 12'h820 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20512; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26656 = 12'h820 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23584; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2080 = io_valid_in ? _GEN_26656 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2080 = 12'h820 == _T_2[11:0] ? image_2080 : _GEN_2079; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5153 = 12'h821 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8225 = 12'h821 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5153; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11297 = 12'h821 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8225; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14369 = 12'h821 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11297; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17441 = 12'h821 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14369; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20513 = 12'h821 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17441; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23585 = 12'h821 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20513; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26657 = 12'h821 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23585; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2081 = io_valid_in ? _GEN_26657 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2081 = 12'h821 == _T_2[11:0] ? image_2081 : _GEN_2080; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5154 = 12'h822 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8226 = 12'h822 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5154; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11298 = 12'h822 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8226; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14370 = 12'h822 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11298; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17442 = 12'h822 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14370; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20514 = 12'h822 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17442; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23586 = 12'h822 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20514; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26658 = 12'h822 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23586; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2082 = io_valid_in ? _GEN_26658 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2082 = 12'h822 == _T_2[11:0] ? image_2082 : _GEN_2081; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5155 = 12'h823 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8227 = 12'h823 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5155; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11299 = 12'h823 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8227; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14371 = 12'h823 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11299; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17443 = 12'h823 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14371; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20515 = 12'h823 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17443; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23587 = 12'h823 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20515; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26659 = 12'h823 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23587; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2083 = io_valid_in ? _GEN_26659 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2083 = 12'h823 == _T_2[11:0] ? image_2083 : _GEN_2082; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5156 = 12'h824 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8228 = 12'h824 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5156; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11300 = 12'h824 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8228; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14372 = 12'h824 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11300; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17444 = 12'h824 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14372; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20516 = 12'h824 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17444; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23588 = 12'h824 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20516; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26660 = 12'h824 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23588; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2084 = io_valid_in ? _GEN_26660 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2084 = 12'h824 == _T_2[11:0] ? image_2084 : _GEN_2083; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5157 = 12'h825 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8229 = 12'h825 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5157; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11301 = 12'h825 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8229; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14373 = 12'h825 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11301; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17445 = 12'h825 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14373; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20517 = 12'h825 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17445; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23589 = 12'h825 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20517; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26661 = 12'h825 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23589; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2085 = io_valid_in ? _GEN_26661 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2085 = 12'h825 == _T_2[11:0] ? image_2085 : _GEN_2084; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5158 = 12'h826 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8230 = 12'h826 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5158; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11302 = 12'h826 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8230; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14374 = 12'h826 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11302; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17446 = 12'h826 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14374; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20518 = 12'h826 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17446; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23590 = 12'h826 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20518; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26662 = 12'h826 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23590; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2086 = io_valid_in ? _GEN_26662 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2086 = 12'h826 == _T_2[11:0] ? image_2086 : _GEN_2085; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5159 = 12'h827 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8231 = 12'h827 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5159; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11303 = 12'h827 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8231; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14375 = 12'h827 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11303; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17447 = 12'h827 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14375; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20519 = 12'h827 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17447; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23591 = 12'h827 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20519; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26663 = 12'h827 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23591; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2087 = io_valid_in ? _GEN_26663 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2087 = 12'h827 == _T_2[11:0] ? image_2087 : _GEN_2086; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5160 = 12'h828 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8232 = 12'h828 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5160; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11304 = 12'h828 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8232; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14376 = 12'h828 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11304; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17448 = 12'h828 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14376; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20520 = 12'h828 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17448; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23592 = 12'h828 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20520; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26664 = 12'h828 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23592; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2088 = io_valid_in ? _GEN_26664 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2088 = 12'h828 == _T_2[11:0] ? image_2088 : _GEN_2087; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5161 = 12'h829 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8233 = 12'h829 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5161; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11305 = 12'h829 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8233; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14377 = 12'h829 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11305; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17449 = 12'h829 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14377; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20521 = 12'h829 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17449; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23593 = 12'h829 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20521; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26665 = 12'h829 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23593; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2089 = io_valid_in ? _GEN_26665 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2089 = 12'h829 == _T_2[11:0] ? image_2089 : _GEN_2088; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5162 = 12'h82a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8234 = 12'h82a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5162; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11306 = 12'h82a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8234; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14378 = 12'h82a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11306; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17450 = 12'h82a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14378; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20522 = 12'h82a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17450; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23594 = 12'h82a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20522; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26666 = 12'h82a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23594; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2090 = io_valid_in ? _GEN_26666 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2090 = 12'h82a == _T_2[11:0] ? image_2090 : _GEN_2089; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5163 = 12'h82b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8235 = 12'h82b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5163; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11307 = 12'h82b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8235; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14379 = 12'h82b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11307; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17451 = 12'h82b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14379; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20523 = 12'h82b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17451; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23595 = 12'h82b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20523; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26667 = 12'h82b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23595; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2091 = io_valid_in ? _GEN_26667 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2091 = 12'h82b == _T_2[11:0] ? image_2091 : _GEN_2090; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5164 = 12'h82c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8236 = 12'h82c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5164; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11308 = 12'h82c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8236; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14380 = 12'h82c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11308; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17452 = 12'h82c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14380; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20524 = 12'h82c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17452; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23596 = 12'h82c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20524; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26668 = 12'h82c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23596; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2092 = io_valid_in ? _GEN_26668 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2092 = 12'h82c == _T_2[11:0] ? image_2092 : _GEN_2091; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5165 = 12'h82d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8237 = 12'h82d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5165; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11309 = 12'h82d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8237; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14381 = 12'h82d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11309; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17453 = 12'h82d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14381; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20525 = 12'h82d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17453; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23597 = 12'h82d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20525; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26669 = 12'h82d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23597; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2093 = io_valid_in ? _GEN_26669 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2093 = 12'h82d == _T_2[11:0] ? image_2093 : _GEN_2092; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5166 = 12'h82e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8238 = 12'h82e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5166; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11310 = 12'h82e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8238; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14382 = 12'h82e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11310; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17454 = 12'h82e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14382; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20526 = 12'h82e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17454; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23598 = 12'h82e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20526; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26670 = 12'h82e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23598; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2094 = io_valid_in ? _GEN_26670 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2094 = 12'h82e == _T_2[11:0] ? image_2094 : _GEN_2093; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5167 = 12'h82f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8239 = 12'h82f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5167; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11311 = 12'h82f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8239; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14383 = 12'h82f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11311; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17455 = 12'h82f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14383; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20527 = 12'h82f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17455; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23599 = 12'h82f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20527; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26671 = 12'h82f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23599; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2095 = io_valid_in ? _GEN_26671 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2095 = 12'h82f == _T_2[11:0] ? image_2095 : _GEN_2094; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5168 = 12'h830 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8240 = 12'h830 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5168; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11312 = 12'h830 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8240; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14384 = 12'h830 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11312; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17456 = 12'h830 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14384; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20528 = 12'h830 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17456; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23600 = 12'h830 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20528; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26672 = 12'h830 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23600; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2096 = io_valid_in ? _GEN_26672 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2096 = 12'h830 == _T_2[11:0] ? image_2096 : _GEN_2095; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5169 = 12'h831 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8241 = 12'h831 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5169; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11313 = 12'h831 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8241; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14385 = 12'h831 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11313; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17457 = 12'h831 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14385; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20529 = 12'h831 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17457; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23601 = 12'h831 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20529; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26673 = 12'h831 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23601; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2097 = io_valid_in ? _GEN_26673 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2097 = 12'h831 == _T_2[11:0] ? image_2097 : _GEN_2096; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5170 = 12'h832 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8242 = 12'h832 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5170; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11314 = 12'h832 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8242; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14386 = 12'h832 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11314; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17458 = 12'h832 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14386; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20530 = 12'h832 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17458; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23602 = 12'h832 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20530; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26674 = 12'h832 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23602; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2098 = io_valid_in ? _GEN_26674 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2098 = 12'h832 == _T_2[11:0] ? image_2098 : _GEN_2097; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5171 = 12'h833 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8243 = 12'h833 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5171; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11315 = 12'h833 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8243; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14387 = 12'h833 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11315; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17459 = 12'h833 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14387; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20531 = 12'h833 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17459; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23603 = 12'h833 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20531; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26675 = 12'h833 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23603; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2099 = io_valid_in ? _GEN_26675 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2099 = 12'h833 == _T_2[11:0] ? image_2099 : _GEN_2098; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5172 = 12'h834 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8244 = 12'h834 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5172; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11316 = 12'h834 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8244; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14388 = 12'h834 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11316; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17460 = 12'h834 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14388; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20532 = 12'h834 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17460; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23604 = 12'h834 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20532; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26676 = 12'h834 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23604; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2100 = io_valid_in ? _GEN_26676 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2100 = 12'h834 == _T_2[11:0] ? image_2100 : _GEN_2099; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5173 = 12'h835 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8245 = 12'h835 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5173; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11317 = 12'h835 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8245; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14389 = 12'h835 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11317; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17461 = 12'h835 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14389; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20533 = 12'h835 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17461; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23605 = 12'h835 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20533; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26677 = 12'h835 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23605; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2101 = io_valid_in ? _GEN_26677 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2101 = 12'h835 == _T_2[11:0] ? image_2101 : _GEN_2100; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5174 = 12'h836 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8246 = 12'h836 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5174; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11318 = 12'h836 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8246; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14390 = 12'h836 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11318; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17462 = 12'h836 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14390; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20534 = 12'h836 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17462; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23606 = 12'h836 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20534; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26678 = 12'h836 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23606; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2102 = io_valid_in ? _GEN_26678 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2102 = 12'h836 == _T_2[11:0] ? image_2102 : _GEN_2101; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5175 = 12'h837 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8247 = 12'h837 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5175; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11319 = 12'h837 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8247; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14391 = 12'h837 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11319; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17463 = 12'h837 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14391; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20535 = 12'h837 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17463; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23607 = 12'h837 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20535; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26679 = 12'h837 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23607; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2103 = io_valid_in ? _GEN_26679 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2103 = 12'h837 == _T_2[11:0] ? image_2103 : _GEN_2102; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5176 = 12'h838 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8248 = 12'h838 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5176; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11320 = 12'h838 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8248; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14392 = 12'h838 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11320; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17464 = 12'h838 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14392; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20536 = 12'h838 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17464; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23608 = 12'h838 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20536; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26680 = 12'h838 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23608; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2104 = io_valid_in ? _GEN_26680 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2104 = 12'h838 == _T_2[11:0] ? image_2104 : _GEN_2103; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5177 = 12'h839 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8249 = 12'h839 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5177; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11321 = 12'h839 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8249; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14393 = 12'h839 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11321; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17465 = 12'h839 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14393; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20537 = 12'h839 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17465; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23609 = 12'h839 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20537; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26681 = 12'h839 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23609; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2105 = io_valid_in ? _GEN_26681 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2105 = 12'h839 == _T_2[11:0] ? image_2105 : _GEN_2104; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5178 = 12'h83a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8250 = 12'h83a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5178; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11322 = 12'h83a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8250; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14394 = 12'h83a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11322; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17466 = 12'h83a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14394; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20538 = 12'h83a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17466; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23610 = 12'h83a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20538; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26682 = 12'h83a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23610; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2106 = io_valid_in ? _GEN_26682 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2106 = 12'h83a == _T_2[11:0] ? image_2106 : _GEN_2105; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5179 = 12'h83b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8251 = 12'h83b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5179; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11323 = 12'h83b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8251; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14395 = 12'h83b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11323; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17467 = 12'h83b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14395; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20539 = 12'h83b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17467; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23611 = 12'h83b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20539; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26683 = 12'h83b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23611; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2107 = io_valid_in ? _GEN_26683 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2107 = 12'h83b == _T_2[11:0] ? image_2107 : _GEN_2106; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5180 = 12'h83c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8252 = 12'h83c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5180; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11324 = 12'h83c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8252; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14396 = 12'h83c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11324; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17468 = 12'h83c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14396; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20540 = 12'h83c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17468; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23612 = 12'h83c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20540; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26684 = 12'h83c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23612; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2108 = io_valid_in ? _GEN_26684 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2108 = 12'h83c == _T_2[11:0] ? image_2108 : _GEN_2107; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5181 = 12'h83d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8253 = 12'h83d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5181; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11325 = 12'h83d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8253; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14397 = 12'h83d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11325; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17469 = 12'h83d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14397; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20541 = 12'h83d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17469; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23613 = 12'h83d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20541; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26685 = 12'h83d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23613; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2109 = io_valid_in ? _GEN_26685 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2109 = 12'h83d == _T_2[11:0] ? image_2109 : _GEN_2108; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5182 = 12'h83e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8254 = 12'h83e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5182; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11326 = 12'h83e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8254; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14398 = 12'h83e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11326; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17470 = 12'h83e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14398; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20542 = 12'h83e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17470; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23614 = 12'h83e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20542; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26686 = 12'h83e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23614; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2110 = io_valid_in ? _GEN_26686 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2110 = 12'h83e == _T_2[11:0] ? image_2110 : _GEN_2109; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5183 = 12'h83f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8255 = 12'h83f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5183; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11327 = 12'h83f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8255; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14399 = 12'h83f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11327; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17471 = 12'h83f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14399; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20543 = 12'h83f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17471; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23615 = 12'h83f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20543; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26687 = 12'h83f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23615; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2111 = io_valid_in ? _GEN_26687 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2111 = 12'h83f == _T_2[11:0] ? image_2111 : _GEN_2110; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5184 = 12'h840 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8256 = 12'h840 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5184; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11328 = 12'h840 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8256; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14400 = 12'h840 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11328; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17472 = 12'h840 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14400; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20544 = 12'h840 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17472; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23616 = 12'h840 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20544; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26688 = 12'h840 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23616; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2112 = io_valid_in ? _GEN_26688 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2112 = 12'h840 == _T_2[11:0] ? image_2112 : _GEN_2111; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5185 = 12'h841 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8257 = 12'h841 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5185; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11329 = 12'h841 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8257; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14401 = 12'h841 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11329; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17473 = 12'h841 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14401; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20545 = 12'h841 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17473; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23617 = 12'h841 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20545; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26689 = 12'h841 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23617; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2113 = io_valid_in ? _GEN_26689 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2113 = 12'h841 == _T_2[11:0] ? image_2113 : _GEN_2112; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5186 = 12'h842 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8258 = 12'h842 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5186; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11330 = 12'h842 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8258; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14402 = 12'h842 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11330; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17474 = 12'h842 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14402; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20546 = 12'h842 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17474; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23618 = 12'h842 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20546; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26690 = 12'h842 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23618; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2114 = io_valid_in ? _GEN_26690 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2114 = 12'h842 == _T_2[11:0] ? image_2114 : _GEN_2113; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5187 = 12'h843 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8259 = 12'h843 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5187; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11331 = 12'h843 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8259; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14403 = 12'h843 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11331; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17475 = 12'h843 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14403; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20547 = 12'h843 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17475; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23619 = 12'h843 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20547; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26691 = 12'h843 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23619; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2115 = io_valid_in ? _GEN_26691 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2115 = 12'h843 == _T_2[11:0] ? image_2115 : _GEN_2114; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5188 = 12'h844 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8260 = 12'h844 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5188; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11332 = 12'h844 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8260; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14404 = 12'h844 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11332; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17476 = 12'h844 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14404; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20548 = 12'h844 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17476; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23620 = 12'h844 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20548; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26692 = 12'h844 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23620; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2116 = io_valid_in ? _GEN_26692 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2116 = 12'h844 == _T_2[11:0] ? image_2116 : _GEN_2115; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5189 = 12'h845 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8261 = 12'h845 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5189; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11333 = 12'h845 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8261; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14405 = 12'h845 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11333; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17477 = 12'h845 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14405; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20549 = 12'h845 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17477; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23621 = 12'h845 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20549; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26693 = 12'h845 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23621; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2117 = io_valid_in ? _GEN_26693 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2117 = 12'h845 == _T_2[11:0] ? image_2117 : _GEN_2116; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5190 = 12'h846 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8262 = 12'h846 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5190; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11334 = 12'h846 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8262; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14406 = 12'h846 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11334; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17478 = 12'h846 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14406; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20550 = 12'h846 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17478; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23622 = 12'h846 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20550; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26694 = 12'h846 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23622; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2118 = io_valid_in ? _GEN_26694 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2118 = 12'h846 == _T_2[11:0] ? image_2118 : _GEN_2117; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5191 = 12'h847 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8263 = 12'h847 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5191; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11335 = 12'h847 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8263; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14407 = 12'h847 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11335; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17479 = 12'h847 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14407; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20551 = 12'h847 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17479; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23623 = 12'h847 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20551; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26695 = 12'h847 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23623; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2119 = io_valid_in ? _GEN_26695 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2119 = 12'h847 == _T_2[11:0] ? image_2119 : _GEN_2118; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5192 = 12'h848 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8264 = 12'h848 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5192; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11336 = 12'h848 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8264; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14408 = 12'h848 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11336; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17480 = 12'h848 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14408; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20552 = 12'h848 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17480; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23624 = 12'h848 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20552; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26696 = 12'h848 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23624; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2120 = io_valid_in ? _GEN_26696 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2120 = 12'h848 == _T_2[11:0] ? image_2120 : _GEN_2119; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5193 = 12'h849 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8265 = 12'h849 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5193; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11337 = 12'h849 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8265; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14409 = 12'h849 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11337; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17481 = 12'h849 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14409; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20553 = 12'h849 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17481; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23625 = 12'h849 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20553; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26697 = 12'h849 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23625; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2121 = io_valid_in ? _GEN_26697 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2121 = 12'h849 == _T_2[11:0] ? image_2121 : _GEN_2120; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5194 = 12'h84a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8266 = 12'h84a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5194; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11338 = 12'h84a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8266; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14410 = 12'h84a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11338; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17482 = 12'h84a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14410; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20554 = 12'h84a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17482; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23626 = 12'h84a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20554; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26698 = 12'h84a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23626; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2122 = io_valid_in ? _GEN_26698 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2122 = 12'h84a == _T_2[11:0] ? image_2122 : _GEN_2121; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5195 = 12'h84b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8267 = 12'h84b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5195; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11339 = 12'h84b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8267; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14411 = 12'h84b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11339; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17483 = 12'h84b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14411; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20555 = 12'h84b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17483; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23627 = 12'h84b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20555; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26699 = 12'h84b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23627; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2123 = io_valid_in ? _GEN_26699 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2123 = 12'h84b == _T_2[11:0] ? image_2123 : _GEN_2122; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5196 = 12'h84c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8268 = 12'h84c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5196; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11340 = 12'h84c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8268; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14412 = 12'h84c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11340; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17484 = 12'h84c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14412; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20556 = 12'h84c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17484; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23628 = 12'h84c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20556; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26700 = 12'h84c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23628; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2124 = io_valid_in ? _GEN_26700 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2124 = 12'h84c == _T_2[11:0] ? image_2124 : _GEN_2123; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5197 = 12'h84d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8269 = 12'h84d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5197; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11341 = 12'h84d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8269; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14413 = 12'h84d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11341; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17485 = 12'h84d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14413; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20557 = 12'h84d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17485; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23629 = 12'h84d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20557; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26701 = 12'h84d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23629; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2125 = io_valid_in ? _GEN_26701 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2125 = 12'h84d == _T_2[11:0] ? image_2125 : _GEN_2124; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5198 = 12'h84e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8270 = 12'h84e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5198; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11342 = 12'h84e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8270; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14414 = 12'h84e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11342; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17486 = 12'h84e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14414; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20558 = 12'h84e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17486; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23630 = 12'h84e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20558; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26702 = 12'h84e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23630; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2126 = io_valid_in ? _GEN_26702 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2126 = 12'h84e == _T_2[11:0] ? image_2126 : _GEN_2125; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5199 = 12'h84f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8271 = 12'h84f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5199; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11343 = 12'h84f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8271; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14415 = 12'h84f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11343; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17487 = 12'h84f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14415; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20559 = 12'h84f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17487; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23631 = 12'h84f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20559; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26703 = 12'h84f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23631; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2127 = io_valid_in ? _GEN_26703 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2127 = 12'h84f == _T_2[11:0] ? image_2127 : _GEN_2126; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5200 = 12'h850 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8272 = 12'h850 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5200; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11344 = 12'h850 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8272; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14416 = 12'h850 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11344; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17488 = 12'h850 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14416; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20560 = 12'h850 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17488; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23632 = 12'h850 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20560; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26704 = 12'h850 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23632; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2128 = io_valid_in ? _GEN_26704 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2128 = 12'h850 == _T_2[11:0] ? image_2128 : _GEN_2127; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5201 = 12'h851 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8273 = 12'h851 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5201; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11345 = 12'h851 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8273; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14417 = 12'h851 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11345; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17489 = 12'h851 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14417; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20561 = 12'h851 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17489; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23633 = 12'h851 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20561; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26705 = 12'h851 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23633; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2129 = io_valid_in ? _GEN_26705 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2129 = 12'h851 == _T_2[11:0] ? image_2129 : _GEN_2128; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5202 = 12'h852 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8274 = 12'h852 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5202; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11346 = 12'h852 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8274; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14418 = 12'h852 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11346; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17490 = 12'h852 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14418; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20562 = 12'h852 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17490; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23634 = 12'h852 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20562; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26706 = 12'h852 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23634; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2130 = io_valid_in ? _GEN_26706 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2130 = 12'h852 == _T_2[11:0] ? image_2130 : _GEN_2129; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5203 = 12'h853 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8275 = 12'h853 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5203; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11347 = 12'h853 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8275; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14419 = 12'h853 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11347; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17491 = 12'h853 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14419; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20563 = 12'h853 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17491; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23635 = 12'h853 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20563; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26707 = 12'h853 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23635; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2131 = io_valid_in ? _GEN_26707 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2131 = 12'h853 == _T_2[11:0] ? image_2131 : _GEN_2130; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5204 = 12'h854 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8276 = 12'h854 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5204; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11348 = 12'h854 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8276; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14420 = 12'h854 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11348; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17492 = 12'h854 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14420; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20564 = 12'h854 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17492; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23636 = 12'h854 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20564; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26708 = 12'h854 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23636; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2132 = io_valid_in ? _GEN_26708 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2132 = 12'h854 == _T_2[11:0] ? image_2132 : _GEN_2131; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5205 = 12'h855 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8277 = 12'h855 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5205; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11349 = 12'h855 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8277; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14421 = 12'h855 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11349; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17493 = 12'h855 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14421; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20565 = 12'h855 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17493; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23637 = 12'h855 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20565; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26709 = 12'h855 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23637; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2133 = io_valid_in ? _GEN_26709 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2133 = 12'h855 == _T_2[11:0] ? image_2133 : _GEN_2132; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5206 = 12'h856 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8278 = 12'h856 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5206; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11350 = 12'h856 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8278; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14422 = 12'h856 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11350; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17494 = 12'h856 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14422; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20566 = 12'h856 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17494; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23638 = 12'h856 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20566; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26710 = 12'h856 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23638; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2134 = io_valid_in ? _GEN_26710 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2134 = 12'h856 == _T_2[11:0] ? image_2134 : _GEN_2133; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5207 = 12'h857 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8279 = 12'h857 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5207; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11351 = 12'h857 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8279; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14423 = 12'h857 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11351; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17495 = 12'h857 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14423; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20567 = 12'h857 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17495; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23639 = 12'h857 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20567; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26711 = 12'h857 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23639; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2135 = io_valid_in ? _GEN_26711 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2135 = 12'h857 == _T_2[11:0] ? image_2135 : _GEN_2134; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5208 = 12'h858 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8280 = 12'h858 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5208; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11352 = 12'h858 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8280; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14424 = 12'h858 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11352; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17496 = 12'h858 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14424; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20568 = 12'h858 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17496; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23640 = 12'h858 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20568; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26712 = 12'h858 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23640; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2136 = io_valid_in ? _GEN_26712 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2136 = 12'h858 == _T_2[11:0] ? image_2136 : _GEN_2135; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5209 = 12'h859 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8281 = 12'h859 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5209; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11353 = 12'h859 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8281; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14425 = 12'h859 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11353; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17497 = 12'h859 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14425; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20569 = 12'h859 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17497; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23641 = 12'h859 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20569; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26713 = 12'h859 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23641; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2137 = io_valid_in ? _GEN_26713 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2137 = 12'h859 == _T_2[11:0] ? image_2137 : _GEN_2136; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5210 = 12'h85a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8282 = 12'h85a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5210; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11354 = 12'h85a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8282; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14426 = 12'h85a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11354; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17498 = 12'h85a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14426; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20570 = 12'h85a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17498; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23642 = 12'h85a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20570; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26714 = 12'h85a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23642; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2138 = io_valid_in ? _GEN_26714 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2138 = 12'h85a == _T_2[11:0] ? image_2138 : _GEN_2137; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5211 = 12'h85b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8283 = 12'h85b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5211; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11355 = 12'h85b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8283; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14427 = 12'h85b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11355; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17499 = 12'h85b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14427; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20571 = 12'h85b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17499; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23643 = 12'h85b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20571; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26715 = 12'h85b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23643; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2139 = io_valid_in ? _GEN_26715 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2139 = 12'h85b == _T_2[11:0] ? image_2139 : _GEN_2138; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5212 = 12'h85c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8284 = 12'h85c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5212; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11356 = 12'h85c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8284; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14428 = 12'h85c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11356; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17500 = 12'h85c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14428; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20572 = 12'h85c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17500; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23644 = 12'h85c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20572; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26716 = 12'h85c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23644; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2140 = io_valid_in ? _GEN_26716 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2140 = 12'h85c == _T_2[11:0] ? image_2140 : _GEN_2139; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5213 = 12'h85d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8285 = 12'h85d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5213; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11357 = 12'h85d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8285; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14429 = 12'h85d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11357; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17501 = 12'h85d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14429; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20573 = 12'h85d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17501; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23645 = 12'h85d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20573; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26717 = 12'h85d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23645; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2141 = io_valid_in ? _GEN_26717 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2141 = 12'h85d == _T_2[11:0] ? image_2141 : _GEN_2140; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5214 = 12'h85e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8286 = 12'h85e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5214; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11358 = 12'h85e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8286; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14430 = 12'h85e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11358; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17502 = 12'h85e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14430; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20574 = 12'h85e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17502; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23646 = 12'h85e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20574; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26718 = 12'h85e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23646; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2142 = io_valid_in ? _GEN_26718 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2142 = 12'h85e == _T_2[11:0] ? image_2142 : _GEN_2141; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5215 = 12'h85f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8287 = 12'h85f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5215; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11359 = 12'h85f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8287; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14431 = 12'h85f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11359; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17503 = 12'h85f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14431; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20575 = 12'h85f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17503; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23647 = 12'h85f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20575; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26719 = 12'h85f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23647; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2143 = io_valid_in ? _GEN_26719 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2143 = 12'h85f == _T_2[11:0] ? image_2143 : _GEN_2142; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5216 = 12'h860 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8288 = 12'h860 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5216; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11360 = 12'h860 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8288; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14432 = 12'h860 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11360; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17504 = 12'h860 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14432; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20576 = 12'h860 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17504; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23648 = 12'h860 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20576; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26720 = 12'h860 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23648; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2144 = io_valid_in ? _GEN_26720 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2144 = 12'h860 == _T_2[11:0] ? image_2144 : _GEN_2143; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5217 = 12'h861 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8289 = 12'h861 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5217; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11361 = 12'h861 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8289; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14433 = 12'h861 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11361; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17505 = 12'h861 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14433; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20577 = 12'h861 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17505; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23649 = 12'h861 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20577; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26721 = 12'h861 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23649; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2145 = io_valid_in ? _GEN_26721 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2145 = 12'h861 == _T_2[11:0] ? image_2145 : _GEN_2144; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5218 = 12'h862 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8290 = 12'h862 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5218; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11362 = 12'h862 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8290; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14434 = 12'h862 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11362; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17506 = 12'h862 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14434; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20578 = 12'h862 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17506; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23650 = 12'h862 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20578; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26722 = 12'h862 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23650; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2146 = io_valid_in ? _GEN_26722 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2146 = 12'h862 == _T_2[11:0] ? image_2146 : _GEN_2145; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5219 = 12'h863 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8291 = 12'h863 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5219; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11363 = 12'h863 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8291; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14435 = 12'h863 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11363; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17507 = 12'h863 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14435; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20579 = 12'h863 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17507; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23651 = 12'h863 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20579; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26723 = 12'h863 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23651; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2147 = io_valid_in ? _GEN_26723 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2147 = 12'h863 == _T_2[11:0] ? image_2147 : _GEN_2146; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5220 = 12'h864 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8292 = 12'h864 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5220; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11364 = 12'h864 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8292; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14436 = 12'h864 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11364; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17508 = 12'h864 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14436; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20580 = 12'h864 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17508; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23652 = 12'h864 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20580; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26724 = 12'h864 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23652; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2148 = io_valid_in ? _GEN_26724 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2148 = 12'h864 == _T_2[11:0] ? image_2148 : _GEN_2147; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5221 = 12'h865 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8293 = 12'h865 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5221; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11365 = 12'h865 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8293; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14437 = 12'h865 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11365; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17509 = 12'h865 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14437; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20581 = 12'h865 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17509; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23653 = 12'h865 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20581; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26725 = 12'h865 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23653; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2149 = io_valid_in ? _GEN_26725 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2149 = 12'h865 == _T_2[11:0] ? image_2149 : _GEN_2148; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5222 = 12'h866 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8294 = 12'h866 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5222; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11366 = 12'h866 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8294; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14438 = 12'h866 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11366; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17510 = 12'h866 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14438; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20582 = 12'h866 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17510; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23654 = 12'h866 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20582; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26726 = 12'h866 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23654; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2150 = io_valid_in ? _GEN_26726 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2150 = 12'h866 == _T_2[11:0] ? image_2150 : _GEN_2149; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5223 = 12'h867 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8295 = 12'h867 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5223; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11367 = 12'h867 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8295; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14439 = 12'h867 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11367; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17511 = 12'h867 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14439; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20583 = 12'h867 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17511; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23655 = 12'h867 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20583; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26727 = 12'h867 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23655; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2151 = io_valid_in ? _GEN_26727 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2151 = 12'h867 == _T_2[11:0] ? image_2151 : _GEN_2150; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5224 = 12'h868 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8296 = 12'h868 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5224; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11368 = 12'h868 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8296; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14440 = 12'h868 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11368; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17512 = 12'h868 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14440; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20584 = 12'h868 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17512; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23656 = 12'h868 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20584; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26728 = 12'h868 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23656; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2152 = io_valid_in ? _GEN_26728 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2152 = 12'h868 == _T_2[11:0] ? image_2152 : _GEN_2151; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5225 = 12'h869 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8297 = 12'h869 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5225; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11369 = 12'h869 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8297; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14441 = 12'h869 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11369; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17513 = 12'h869 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14441; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20585 = 12'h869 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17513; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23657 = 12'h869 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20585; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26729 = 12'h869 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23657; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2153 = io_valid_in ? _GEN_26729 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2153 = 12'h869 == _T_2[11:0] ? image_2153 : _GEN_2152; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5226 = 12'h86a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8298 = 12'h86a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5226; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11370 = 12'h86a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8298; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14442 = 12'h86a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11370; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17514 = 12'h86a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14442; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20586 = 12'h86a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17514; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23658 = 12'h86a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20586; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26730 = 12'h86a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23658; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2154 = io_valid_in ? _GEN_26730 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2154 = 12'h86a == _T_2[11:0] ? image_2154 : _GEN_2153; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5227 = 12'h86b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8299 = 12'h86b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5227; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11371 = 12'h86b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8299; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14443 = 12'h86b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11371; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17515 = 12'h86b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14443; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20587 = 12'h86b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17515; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23659 = 12'h86b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20587; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26731 = 12'h86b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23659; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2155 = io_valid_in ? _GEN_26731 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2155 = 12'h86b == _T_2[11:0] ? image_2155 : _GEN_2154; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5228 = 12'h86c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8300 = 12'h86c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5228; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11372 = 12'h86c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8300; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14444 = 12'h86c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11372; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17516 = 12'h86c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14444; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20588 = 12'h86c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17516; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23660 = 12'h86c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20588; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26732 = 12'h86c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23660; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2156 = io_valid_in ? _GEN_26732 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2156 = 12'h86c == _T_2[11:0] ? image_2156 : _GEN_2155; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5229 = 12'h86d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8301 = 12'h86d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5229; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11373 = 12'h86d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8301; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14445 = 12'h86d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11373; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17517 = 12'h86d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14445; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20589 = 12'h86d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17517; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23661 = 12'h86d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20589; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26733 = 12'h86d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23661; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2157 = io_valid_in ? _GEN_26733 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2157 = 12'h86d == _T_2[11:0] ? image_2157 : _GEN_2156; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5230 = 12'h86e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8302 = 12'h86e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5230; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11374 = 12'h86e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8302; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14446 = 12'h86e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11374; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17518 = 12'h86e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14446; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20590 = 12'h86e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17518; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23662 = 12'h86e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20590; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26734 = 12'h86e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23662; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2158 = io_valid_in ? _GEN_26734 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2158 = 12'h86e == _T_2[11:0] ? image_2158 : _GEN_2157; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5231 = 12'h86f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8303 = 12'h86f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5231; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11375 = 12'h86f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8303; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14447 = 12'h86f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11375; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17519 = 12'h86f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14447; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20591 = 12'h86f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17519; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23663 = 12'h86f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20591; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26735 = 12'h86f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23663; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2159 = io_valid_in ? _GEN_26735 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2159 = 12'h86f == _T_2[11:0] ? image_2159 : _GEN_2158; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5232 = 12'h870 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8304 = 12'h870 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5232; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11376 = 12'h870 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8304; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14448 = 12'h870 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11376; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17520 = 12'h870 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14448; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20592 = 12'h870 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17520; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23664 = 12'h870 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20592; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26736 = 12'h870 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23664; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2160 = io_valid_in ? _GEN_26736 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2160 = 12'h870 == _T_2[11:0] ? image_2160 : _GEN_2159; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5233 = 12'h871 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8305 = 12'h871 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5233; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11377 = 12'h871 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8305; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14449 = 12'h871 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11377; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17521 = 12'h871 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14449; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20593 = 12'h871 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17521; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23665 = 12'h871 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20593; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26737 = 12'h871 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23665; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2161 = io_valid_in ? _GEN_26737 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2161 = 12'h871 == _T_2[11:0] ? image_2161 : _GEN_2160; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5234 = 12'h872 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8306 = 12'h872 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5234; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11378 = 12'h872 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8306; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14450 = 12'h872 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11378; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17522 = 12'h872 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14450; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20594 = 12'h872 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17522; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23666 = 12'h872 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20594; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26738 = 12'h872 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23666; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2162 = io_valid_in ? _GEN_26738 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2162 = 12'h872 == _T_2[11:0] ? image_2162 : _GEN_2161; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5235 = 12'h873 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8307 = 12'h873 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5235; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11379 = 12'h873 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8307; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14451 = 12'h873 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11379; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17523 = 12'h873 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14451; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20595 = 12'h873 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17523; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23667 = 12'h873 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20595; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26739 = 12'h873 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23667; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2163 = io_valid_in ? _GEN_26739 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2163 = 12'h873 == _T_2[11:0] ? image_2163 : _GEN_2162; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5236 = 12'h874 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8308 = 12'h874 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5236; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11380 = 12'h874 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8308; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14452 = 12'h874 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11380; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17524 = 12'h874 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14452; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20596 = 12'h874 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17524; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23668 = 12'h874 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20596; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26740 = 12'h874 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23668; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2164 = io_valid_in ? _GEN_26740 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2164 = 12'h874 == _T_2[11:0] ? image_2164 : _GEN_2163; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5237 = 12'h875 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8309 = 12'h875 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5237; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11381 = 12'h875 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8309; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14453 = 12'h875 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11381; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17525 = 12'h875 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14453; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20597 = 12'h875 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17525; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23669 = 12'h875 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20597; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26741 = 12'h875 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23669; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2165 = io_valid_in ? _GEN_26741 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2165 = 12'h875 == _T_2[11:0] ? image_2165 : _GEN_2164; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5238 = 12'h876 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8310 = 12'h876 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5238; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11382 = 12'h876 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8310; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14454 = 12'h876 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11382; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17526 = 12'h876 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14454; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20598 = 12'h876 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17526; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23670 = 12'h876 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20598; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26742 = 12'h876 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23670; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2166 = io_valid_in ? _GEN_26742 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2166 = 12'h876 == _T_2[11:0] ? image_2166 : _GEN_2165; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5239 = 12'h877 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8311 = 12'h877 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5239; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11383 = 12'h877 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8311; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14455 = 12'h877 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11383; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17527 = 12'h877 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14455; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20599 = 12'h877 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17527; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23671 = 12'h877 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20599; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26743 = 12'h877 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23671; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2167 = io_valid_in ? _GEN_26743 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2167 = 12'h877 == _T_2[11:0] ? image_2167 : _GEN_2166; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5240 = 12'h878 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8312 = 12'h878 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5240; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11384 = 12'h878 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8312; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14456 = 12'h878 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11384; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17528 = 12'h878 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14456; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20600 = 12'h878 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17528; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23672 = 12'h878 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20600; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26744 = 12'h878 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23672; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2168 = io_valid_in ? _GEN_26744 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2168 = 12'h878 == _T_2[11:0] ? image_2168 : _GEN_2167; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5241 = 12'h879 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8313 = 12'h879 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5241; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11385 = 12'h879 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8313; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14457 = 12'h879 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11385; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17529 = 12'h879 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14457; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20601 = 12'h879 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17529; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23673 = 12'h879 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20601; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26745 = 12'h879 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23673; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2169 = io_valid_in ? _GEN_26745 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2169 = 12'h879 == _T_2[11:0] ? image_2169 : _GEN_2168; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5242 = 12'h87a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8314 = 12'h87a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5242; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11386 = 12'h87a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8314; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14458 = 12'h87a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11386; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17530 = 12'h87a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14458; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20602 = 12'h87a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17530; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23674 = 12'h87a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20602; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26746 = 12'h87a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23674; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2170 = io_valid_in ? _GEN_26746 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2170 = 12'h87a == _T_2[11:0] ? image_2170 : _GEN_2169; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5243 = 12'h87b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8315 = 12'h87b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5243; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11387 = 12'h87b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8315; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14459 = 12'h87b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11387; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17531 = 12'h87b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14459; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20603 = 12'h87b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17531; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23675 = 12'h87b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20603; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26747 = 12'h87b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23675; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2171 = io_valid_in ? _GEN_26747 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2171 = 12'h87b == _T_2[11:0] ? image_2171 : _GEN_2170; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5244 = 12'h87c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8316 = 12'h87c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5244; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11388 = 12'h87c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8316; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14460 = 12'h87c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11388; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17532 = 12'h87c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14460; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20604 = 12'h87c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17532; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23676 = 12'h87c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20604; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26748 = 12'h87c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23676; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2172 = io_valid_in ? _GEN_26748 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2172 = 12'h87c == _T_2[11:0] ? image_2172 : _GEN_2171; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5245 = 12'h87d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8317 = 12'h87d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5245; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11389 = 12'h87d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8317; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14461 = 12'h87d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11389; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17533 = 12'h87d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14461; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20605 = 12'h87d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17533; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23677 = 12'h87d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20605; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26749 = 12'h87d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23677; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2173 = io_valid_in ? _GEN_26749 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2173 = 12'h87d == _T_2[11:0] ? image_2173 : _GEN_2172; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5246 = 12'h87e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8318 = 12'h87e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5246; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11390 = 12'h87e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8318; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14462 = 12'h87e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11390; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17534 = 12'h87e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14462; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20606 = 12'h87e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17534; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23678 = 12'h87e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20606; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26750 = 12'h87e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23678; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2174 = io_valid_in ? _GEN_26750 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2174 = 12'h87e == _T_2[11:0] ? image_2174 : _GEN_2173; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5247 = 12'h87f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8319 = 12'h87f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5247; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11391 = 12'h87f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8319; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14463 = 12'h87f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11391; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17535 = 12'h87f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14463; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20607 = 12'h87f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17535; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23679 = 12'h87f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20607; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26751 = 12'h87f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23679; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2175 = io_valid_in ? _GEN_26751 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2175 = 12'h87f == _T_2[11:0] ? image_2175 : _GEN_2174; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5248 = 12'h880 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8320 = 12'h880 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5248; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11392 = 12'h880 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8320; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14464 = 12'h880 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11392; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17536 = 12'h880 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14464; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20608 = 12'h880 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17536; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23680 = 12'h880 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20608; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26752 = 12'h880 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23680; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2176 = io_valid_in ? _GEN_26752 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2176 = 12'h880 == _T_2[11:0] ? image_2176 : _GEN_2175; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5249 = 12'h881 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8321 = 12'h881 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5249; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11393 = 12'h881 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8321; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14465 = 12'h881 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11393; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17537 = 12'h881 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14465; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20609 = 12'h881 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17537; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23681 = 12'h881 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20609; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26753 = 12'h881 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23681; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2177 = io_valid_in ? _GEN_26753 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2177 = 12'h881 == _T_2[11:0] ? image_2177 : _GEN_2176; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5250 = 12'h882 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8322 = 12'h882 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5250; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11394 = 12'h882 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8322; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14466 = 12'h882 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11394; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17538 = 12'h882 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14466; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20610 = 12'h882 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17538; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23682 = 12'h882 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20610; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26754 = 12'h882 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23682; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2178 = io_valid_in ? _GEN_26754 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2178 = 12'h882 == _T_2[11:0] ? image_2178 : _GEN_2177; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5251 = 12'h883 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8323 = 12'h883 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5251; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11395 = 12'h883 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8323; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14467 = 12'h883 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11395; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17539 = 12'h883 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14467; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20611 = 12'h883 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17539; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23683 = 12'h883 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20611; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26755 = 12'h883 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23683; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2179 = io_valid_in ? _GEN_26755 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2179 = 12'h883 == _T_2[11:0] ? image_2179 : _GEN_2178; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5252 = 12'h884 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8324 = 12'h884 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5252; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11396 = 12'h884 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8324; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14468 = 12'h884 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11396; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17540 = 12'h884 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14468; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20612 = 12'h884 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17540; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23684 = 12'h884 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20612; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26756 = 12'h884 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23684; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2180 = io_valid_in ? _GEN_26756 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2180 = 12'h884 == _T_2[11:0] ? image_2180 : _GEN_2179; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5253 = 12'h885 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8325 = 12'h885 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5253; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11397 = 12'h885 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8325; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14469 = 12'h885 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11397; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17541 = 12'h885 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14469; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20613 = 12'h885 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17541; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23685 = 12'h885 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20613; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26757 = 12'h885 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23685; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2181 = io_valid_in ? _GEN_26757 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2181 = 12'h885 == _T_2[11:0] ? image_2181 : _GEN_2180; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5254 = 12'h886 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8326 = 12'h886 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5254; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11398 = 12'h886 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8326; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14470 = 12'h886 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11398; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17542 = 12'h886 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14470; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20614 = 12'h886 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17542; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23686 = 12'h886 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20614; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26758 = 12'h886 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23686; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2182 = io_valid_in ? _GEN_26758 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2182 = 12'h886 == _T_2[11:0] ? image_2182 : _GEN_2181; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5255 = 12'h887 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8327 = 12'h887 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5255; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11399 = 12'h887 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8327; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14471 = 12'h887 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11399; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17543 = 12'h887 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14471; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20615 = 12'h887 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17543; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23687 = 12'h887 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20615; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26759 = 12'h887 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23687; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2183 = io_valid_in ? _GEN_26759 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2183 = 12'h887 == _T_2[11:0] ? image_2183 : _GEN_2182; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5256 = 12'h888 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8328 = 12'h888 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5256; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11400 = 12'h888 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8328; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14472 = 12'h888 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11400; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17544 = 12'h888 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14472; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20616 = 12'h888 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17544; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23688 = 12'h888 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20616; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26760 = 12'h888 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23688; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2184 = io_valid_in ? _GEN_26760 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2184 = 12'h888 == _T_2[11:0] ? image_2184 : _GEN_2183; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5257 = 12'h889 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8329 = 12'h889 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5257; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11401 = 12'h889 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8329; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14473 = 12'h889 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11401; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17545 = 12'h889 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14473; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20617 = 12'h889 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17545; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23689 = 12'h889 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20617; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26761 = 12'h889 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23689; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2185 = io_valid_in ? _GEN_26761 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2185 = 12'h889 == _T_2[11:0] ? image_2185 : _GEN_2184; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5258 = 12'h88a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8330 = 12'h88a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5258; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11402 = 12'h88a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8330; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14474 = 12'h88a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11402; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17546 = 12'h88a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14474; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20618 = 12'h88a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17546; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23690 = 12'h88a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20618; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26762 = 12'h88a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23690; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2186 = io_valid_in ? _GEN_26762 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2186 = 12'h88a == _T_2[11:0] ? image_2186 : _GEN_2185; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5259 = 12'h88b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8331 = 12'h88b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5259; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11403 = 12'h88b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8331; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14475 = 12'h88b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11403; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17547 = 12'h88b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14475; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20619 = 12'h88b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17547; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23691 = 12'h88b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20619; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26763 = 12'h88b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23691; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2187 = io_valid_in ? _GEN_26763 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2187 = 12'h88b == _T_2[11:0] ? image_2187 : _GEN_2186; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5260 = 12'h88c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8332 = 12'h88c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5260; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11404 = 12'h88c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8332; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14476 = 12'h88c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11404; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17548 = 12'h88c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14476; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20620 = 12'h88c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17548; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23692 = 12'h88c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20620; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26764 = 12'h88c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23692; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2188 = io_valid_in ? _GEN_26764 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2188 = 12'h88c == _T_2[11:0] ? image_2188 : _GEN_2187; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5261 = 12'h88d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8333 = 12'h88d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5261; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11405 = 12'h88d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8333; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14477 = 12'h88d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11405; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17549 = 12'h88d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14477; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20621 = 12'h88d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17549; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23693 = 12'h88d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20621; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26765 = 12'h88d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23693; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2189 = io_valid_in ? _GEN_26765 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2189 = 12'h88d == _T_2[11:0] ? image_2189 : _GEN_2188; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5262 = 12'h88e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8334 = 12'h88e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5262; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11406 = 12'h88e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8334; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14478 = 12'h88e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11406; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17550 = 12'h88e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14478; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20622 = 12'h88e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17550; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23694 = 12'h88e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20622; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26766 = 12'h88e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23694; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2190 = io_valid_in ? _GEN_26766 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2190 = 12'h88e == _T_2[11:0] ? image_2190 : _GEN_2189; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5263 = 12'h88f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8335 = 12'h88f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5263; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11407 = 12'h88f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8335; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14479 = 12'h88f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11407; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17551 = 12'h88f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14479; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20623 = 12'h88f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17551; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23695 = 12'h88f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20623; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26767 = 12'h88f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23695; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2191 = io_valid_in ? _GEN_26767 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2191 = 12'h88f == _T_2[11:0] ? image_2191 : _GEN_2190; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5264 = 12'h890 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8336 = 12'h890 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5264; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11408 = 12'h890 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8336; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14480 = 12'h890 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11408; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17552 = 12'h890 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14480; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20624 = 12'h890 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17552; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23696 = 12'h890 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20624; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26768 = 12'h890 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23696; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2192 = io_valid_in ? _GEN_26768 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2192 = 12'h890 == _T_2[11:0] ? image_2192 : _GEN_2191; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5265 = 12'h891 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8337 = 12'h891 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5265; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11409 = 12'h891 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8337; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14481 = 12'h891 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11409; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17553 = 12'h891 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14481; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20625 = 12'h891 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17553; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23697 = 12'h891 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20625; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26769 = 12'h891 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23697; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2193 = io_valid_in ? _GEN_26769 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2193 = 12'h891 == _T_2[11:0] ? image_2193 : _GEN_2192; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5266 = 12'h892 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8338 = 12'h892 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5266; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11410 = 12'h892 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8338; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14482 = 12'h892 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11410; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17554 = 12'h892 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14482; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20626 = 12'h892 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17554; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23698 = 12'h892 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20626; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26770 = 12'h892 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23698; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2194 = io_valid_in ? _GEN_26770 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2194 = 12'h892 == _T_2[11:0] ? image_2194 : _GEN_2193; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5267 = 12'h893 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8339 = 12'h893 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5267; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11411 = 12'h893 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8339; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14483 = 12'h893 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11411; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17555 = 12'h893 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14483; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20627 = 12'h893 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17555; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23699 = 12'h893 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20627; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26771 = 12'h893 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23699; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2195 = io_valid_in ? _GEN_26771 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2195 = 12'h893 == _T_2[11:0] ? image_2195 : _GEN_2194; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5268 = 12'h894 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8340 = 12'h894 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5268; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11412 = 12'h894 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8340; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14484 = 12'h894 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11412; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17556 = 12'h894 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14484; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20628 = 12'h894 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17556; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23700 = 12'h894 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20628; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26772 = 12'h894 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23700; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2196 = io_valid_in ? _GEN_26772 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2196 = 12'h894 == _T_2[11:0] ? image_2196 : _GEN_2195; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5269 = 12'h895 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8341 = 12'h895 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5269; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11413 = 12'h895 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8341; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14485 = 12'h895 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11413; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17557 = 12'h895 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14485; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20629 = 12'h895 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17557; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23701 = 12'h895 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20629; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26773 = 12'h895 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23701; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2197 = io_valid_in ? _GEN_26773 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2197 = 12'h895 == _T_2[11:0] ? image_2197 : _GEN_2196; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5270 = 12'h896 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8342 = 12'h896 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5270; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11414 = 12'h896 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8342; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14486 = 12'h896 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11414; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17558 = 12'h896 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14486; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20630 = 12'h896 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17558; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23702 = 12'h896 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20630; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26774 = 12'h896 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23702; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2198 = io_valid_in ? _GEN_26774 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2198 = 12'h896 == _T_2[11:0] ? image_2198 : _GEN_2197; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5271 = 12'h897 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8343 = 12'h897 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5271; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11415 = 12'h897 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8343; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14487 = 12'h897 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11415; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17559 = 12'h897 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14487; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20631 = 12'h897 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17559; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23703 = 12'h897 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20631; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26775 = 12'h897 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23703; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2199 = io_valid_in ? _GEN_26775 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2199 = 12'h897 == _T_2[11:0] ? image_2199 : _GEN_2198; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5272 = 12'h898 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8344 = 12'h898 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5272; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11416 = 12'h898 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8344; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14488 = 12'h898 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11416; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17560 = 12'h898 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14488; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20632 = 12'h898 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17560; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23704 = 12'h898 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20632; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26776 = 12'h898 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23704; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2200 = io_valid_in ? _GEN_26776 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2200 = 12'h898 == _T_2[11:0] ? image_2200 : _GEN_2199; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5273 = 12'h899 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8345 = 12'h899 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5273; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11417 = 12'h899 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8345; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14489 = 12'h899 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11417; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17561 = 12'h899 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14489; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20633 = 12'h899 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17561; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23705 = 12'h899 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20633; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26777 = 12'h899 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23705; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2201 = io_valid_in ? _GEN_26777 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2201 = 12'h899 == _T_2[11:0] ? image_2201 : _GEN_2200; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5274 = 12'h89a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8346 = 12'h89a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5274; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11418 = 12'h89a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8346; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14490 = 12'h89a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11418; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17562 = 12'h89a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14490; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20634 = 12'h89a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17562; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23706 = 12'h89a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20634; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26778 = 12'h89a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23706; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2202 = io_valid_in ? _GEN_26778 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2202 = 12'h89a == _T_2[11:0] ? image_2202 : _GEN_2201; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5275 = 12'h89b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8347 = 12'h89b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5275; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11419 = 12'h89b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8347; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14491 = 12'h89b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11419; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17563 = 12'h89b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14491; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20635 = 12'h89b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17563; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23707 = 12'h89b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20635; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26779 = 12'h89b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23707; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2203 = io_valid_in ? _GEN_26779 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2203 = 12'h89b == _T_2[11:0] ? image_2203 : _GEN_2202; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5276 = 12'h89c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8348 = 12'h89c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5276; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11420 = 12'h89c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8348; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14492 = 12'h89c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11420; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17564 = 12'h89c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14492; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20636 = 12'h89c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17564; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23708 = 12'h89c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20636; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26780 = 12'h89c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23708; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2204 = io_valid_in ? _GEN_26780 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2204 = 12'h89c == _T_2[11:0] ? image_2204 : _GEN_2203; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5277 = 12'h89d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8349 = 12'h89d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5277; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11421 = 12'h89d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8349; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14493 = 12'h89d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11421; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17565 = 12'h89d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14493; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20637 = 12'h89d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17565; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23709 = 12'h89d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20637; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26781 = 12'h89d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23709; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2205 = io_valid_in ? _GEN_26781 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2205 = 12'h89d == _T_2[11:0] ? image_2205 : _GEN_2204; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5278 = 12'h89e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8350 = 12'h89e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5278; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11422 = 12'h89e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8350; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14494 = 12'h89e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11422; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17566 = 12'h89e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14494; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20638 = 12'h89e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17566; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23710 = 12'h89e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20638; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26782 = 12'h89e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23710; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2206 = io_valid_in ? _GEN_26782 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2206 = 12'h89e == _T_2[11:0] ? image_2206 : _GEN_2205; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5279 = 12'h89f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8351 = 12'h89f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5279; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11423 = 12'h89f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8351; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14495 = 12'h89f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11423; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17567 = 12'h89f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14495; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20639 = 12'h89f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17567; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23711 = 12'h89f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20639; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26783 = 12'h89f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23711; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2207 = io_valid_in ? _GEN_26783 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2207 = 12'h89f == _T_2[11:0] ? image_2207 : _GEN_2206; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5280 = 12'h8a0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8352 = 12'h8a0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5280; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11424 = 12'h8a0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8352; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14496 = 12'h8a0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11424; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17568 = 12'h8a0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14496; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20640 = 12'h8a0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17568; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23712 = 12'h8a0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20640; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26784 = 12'h8a0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23712; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2208 = io_valid_in ? _GEN_26784 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2208 = 12'h8a0 == _T_2[11:0] ? image_2208 : _GEN_2207; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5281 = 12'h8a1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8353 = 12'h8a1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5281; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11425 = 12'h8a1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8353; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14497 = 12'h8a1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11425; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17569 = 12'h8a1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14497; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20641 = 12'h8a1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17569; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23713 = 12'h8a1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20641; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26785 = 12'h8a1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23713; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2209 = io_valid_in ? _GEN_26785 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2209 = 12'h8a1 == _T_2[11:0] ? image_2209 : _GEN_2208; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5282 = 12'h8a2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8354 = 12'h8a2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5282; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11426 = 12'h8a2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8354; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14498 = 12'h8a2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11426; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17570 = 12'h8a2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14498; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20642 = 12'h8a2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17570; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23714 = 12'h8a2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20642; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26786 = 12'h8a2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23714; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2210 = io_valid_in ? _GEN_26786 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2210 = 12'h8a2 == _T_2[11:0] ? image_2210 : _GEN_2209; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5283 = 12'h8a3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8355 = 12'h8a3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5283; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11427 = 12'h8a3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8355; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14499 = 12'h8a3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11427; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17571 = 12'h8a3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14499; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20643 = 12'h8a3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17571; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23715 = 12'h8a3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20643; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26787 = 12'h8a3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23715; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2211 = io_valid_in ? _GEN_26787 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2211 = 12'h8a3 == _T_2[11:0] ? image_2211 : _GEN_2210; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5284 = 12'h8a4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8356 = 12'h8a4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5284; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11428 = 12'h8a4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8356; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14500 = 12'h8a4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11428; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17572 = 12'h8a4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14500; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20644 = 12'h8a4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17572; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23716 = 12'h8a4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20644; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26788 = 12'h8a4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23716; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2212 = io_valid_in ? _GEN_26788 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2212 = 12'h8a4 == _T_2[11:0] ? image_2212 : _GEN_2211; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5285 = 12'h8a5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8357 = 12'h8a5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5285; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11429 = 12'h8a5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8357; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14501 = 12'h8a5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11429; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17573 = 12'h8a5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14501; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20645 = 12'h8a5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17573; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23717 = 12'h8a5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20645; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26789 = 12'h8a5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23717; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2213 = io_valid_in ? _GEN_26789 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2213 = 12'h8a5 == _T_2[11:0] ? image_2213 : _GEN_2212; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5286 = 12'h8a6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8358 = 12'h8a6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5286; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11430 = 12'h8a6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8358; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14502 = 12'h8a6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11430; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17574 = 12'h8a6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14502; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20646 = 12'h8a6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17574; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23718 = 12'h8a6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20646; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26790 = 12'h8a6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23718; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2214 = io_valid_in ? _GEN_26790 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2214 = 12'h8a6 == _T_2[11:0] ? image_2214 : _GEN_2213; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5287 = 12'h8a7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8359 = 12'h8a7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5287; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11431 = 12'h8a7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8359; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14503 = 12'h8a7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11431; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17575 = 12'h8a7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14503; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20647 = 12'h8a7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17575; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23719 = 12'h8a7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20647; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26791 = 12'h8a7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23719; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2215 = io_valid_in ? _GEN_26791 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2215 = 12'h8a7 == _T_2[11:0] ? image_2215 : _GEN_2214; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5288 = 12'h8a8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8360 = 12'h8a8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5288; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11432 = 12'h8a8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8360; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14504 = 12'h8a8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11432; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17576 = 12'h8a8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14504; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20648 = 12'h8a8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17576; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23720 = 12'h8a8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20648; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26792 = 12'h8a8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23720; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2216 = io_valid_in ? _GEN_26792 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2216 = 12'h8a8 == _T_2[11:0] ? image_2216 : _GEN_2215; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5289 = 12'h8a9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8361 = 12'h8a9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5289; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11433 = 12'h8a9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8361; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14505 = 12'h8a9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11433; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17577 = 12'h8a9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14505; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20649 = 12'h8a9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17577; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23721 = 12'h8a9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20649; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26793 = 12'h8a9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23721; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2217 = io_valid_in ? _GEN_26793 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2217 = 12'h8a9 == _T_2[11:0] ? image_2217 : _GEN_2216; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5290 = 12'h8aa == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8362 = 12'h8aa == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5290; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11434 = 12'h8aa == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8362; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14506 = 12'h8aa == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11434; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17578 = 12'h8aa == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14506; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20650 = 12'h8aa == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17578; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23722 = 12'h8aa == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20650; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26794 = 12'h8aa == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23722; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2218 = io_valid_in ? _GEN_26794 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2218 = 12'h8aa == _T_2[11:0] ? image_2218 : _GEN_2217; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5291 = 12'h8ab == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8363 = 12'h8ab == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5291; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11435 = 12'h8ab == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8363; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14507 = 12'h8ab == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11435; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17579 = 12'h8ab == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14507; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20651 = 12'h8ab == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17579; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23723 = 12'h8ab == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20651; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26795 = 12'h8ab == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23723; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2219 = io_valid_in ? _GEN_26795 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2219 = 12'h8ab == _T_2[11:0] ? image_2219 : _GEN_2218; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5292 = 12'h8ac == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8364 = 12'h8ac == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5292; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11436 = 12'h8ac == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8364; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14508 = 12'h8ac == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11436; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17580 = 12'h8ac == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14508; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20652 = 12'h8ac == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17580; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23724 = 12'h8ac == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20652; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26796 = 12'h8ac == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23724; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2220 = io_valid_in ? _GEN_26796 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2220 = 12'h8ac == _T_2[11:0] ? image_2220 : _GEN_2219; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5293 = 12'h8ad == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8365 = 12'h8ad == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5293; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11437 = 12'h8ad == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8365; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14509 = 12'h8ad == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11437; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17581 = 12'h8ad == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14509; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20653 = 12'h8ad == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17581; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23725 = 12'h8ad == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20653; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26797 = 12'h8ad == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23725; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2221 = io_valid_in ? _GEN_26797 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2221 = 12'h8ad == _T_2[11:0] ? image_2221 : _GEN_2220; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5294 = 12'h8ae == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8366 = 12'h8ae == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5294; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11438 = 12'h8ae == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8366; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14510 = 12'h8ae == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11438; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17582 = 12'h8ae == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14510; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20654 = 12'h8ae == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17582; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23726 = 12'h8ae == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20654; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26798 = 12'h8ae == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23726; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2222 = io_valid_in ? _GEN_26798 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2222 = 12'h8ae == _T_2[11:0] ? image_2222 : _GEN_2221; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5295 = 12'h8af == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8367 = 12'h8af == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5295; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11439 = 12'h8af == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8367; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14511 = 12'h8af == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11439; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17583 = 12'h8af == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14511; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20655 = 12'h8af == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17583; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23727 = 12'h8af == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20655; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26799 = 12'h8af == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23727; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2223 = io_valid_in ? _GEN_26799 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2223 = 12'h8af == _T_2[11:0] ? image_2223 : _GEN_2222; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5296 = 12'h8b0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8368 = 12'h8b0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5296; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11440 = 12'h8b0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8368; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14512 = 12'h8b0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11440; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17584 = 12'h8b0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14512; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20656 = 12'h8b0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17584; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23728 = 12'h8b0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20656; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26800 = 12'h8b0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23728; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2224 = io_valid_in ? _GEN_26800 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2224 = 12'h8b0 == _T_2[11:0] ? image_2224 : _GEN_2223; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5297 = 12'h8b1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8369 = 12'h8b1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5297; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11441 = 12'h8b1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8369; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14513 = 12'h8b1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11441; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17585 = 12'h8b1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14513; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20657 = 12'h8b1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17585; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23729 = 12'h8b1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20657; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26801 = 12'h8b1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23729; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2225 = io_valid_in ? _GEN_26801 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2225 = 12'h8b1 == _T_2[11:0] ? image_2225 : _GEN_2224; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5298 = 12'h8b2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8370 = 12'h8b2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5298; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11442 = 12'h8b2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8370; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14514 = 12'h8b2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11442; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17586 = 12'h8b2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14514; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20658 = 12'h8b2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17586; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23730 = 12'h8b2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20658; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26802 = 12'h8b2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23730; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2226 = io_valid_in ? _GEN_26802 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2226 = 12'h8b2 == _T_2[11:0] ? image_2226 : _GEN_2225; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5299 = 12'h8b3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8371 = 12'h8b3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5299; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11443 = 12'h8b3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8371; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14515 = 12'h8b3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11443; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17587 = 12'h8b3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14515; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20659 = 12'h8b3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17587; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23731 = 12'h8b3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20659; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26803 = 12'h8b3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23731; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2227 = io_valid_in ? _GEN_26803 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2227 = 12'h8b3 == _T_2[11:0] ? image_2227 : _GEN_2226; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5300 = 12'h8b4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8372 = 12'h8b4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5300; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11444 = 12'h8b4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8372; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14516 = 12'h8b4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11444; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17588 = 12'h8b4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14516; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20660 = 12'h8b4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17588; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23732 = 12'h8b4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20660; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26804 = 12'h8b4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23732; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2228 = io_valid_in ? _GEN_26804 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2228 = 12'h8b4 == _T_2[11:0] ? image_2228 : _GEN_2227; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5301 = 12'h8b5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8373 = 12'h8b5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5301; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11445 = 12'h8b5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8373; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14517 = 12'h8b5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11445; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17589 = 12'h8b5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14517; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20661 = 12'h8b5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17589; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23733 = 12'h8b5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20661; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26805 = 12'h8b5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23733; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2229 = io_valid_in ? _GEN_26805 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2229 = 12'h8b5 == _T_2[11:0] ? image_2229 : _GEN_2228; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5302 = 12'h8b6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8374 = 12'h8b6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5302; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11446 = 12'h8b6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8374; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14518 = 12'h8b6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11446; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17590 = 12'h8b6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14518; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20662 = 12'h8b6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17590; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23734 = 12'h8b6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20662; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26806 = 12'h8b6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23734; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2230 = io_valid_in ? _GEN_26806 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2230 = 12'h8b6 == _T_2[11:0] ? image_2230 : _GEN_2229; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5303 = 12'h8b7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8375 = 12'h8b7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5303; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11447 = 12'h8b7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8375; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14519 = 12'h8b7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11447; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17591 = 12'h8b7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14519; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20663 = 12'h8b7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17591; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23735 = 12'h8b7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20663; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26807 = 12'h8b7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23735; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2231 = io_valid_in ? _GEN_26807 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2231 = 12'h8b7 == _T_2[11:0] ? image_2231 : _GEN_2230; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5304 = 12'h8b8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8376 = 12'h8b8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5304; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11448 = 12'h8b8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8376; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14520 = 12'h8b8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11448; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17592 = 12'h8b8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14520; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20664 = 12'h8b8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17592; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23736 = 12'h8b8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20664; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26808 = 12'h8b8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23736; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2232 = io_valid_in ? _GEN_26808 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2232 = 12'h8b8 == _T_2[11:0] ? image_2232 : _GEN_2231; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5305 = 12'h8b9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8377 = 12'h8b9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5305; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11449 = 12'h8b9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8377; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14521 = 12'h8b9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11449; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17593 = 12'h8b9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14521; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20665 = 12'h8b9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17593; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23737 = 12'h8b9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20665; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26809 = 12'h8b9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23737; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2233 = io_valid_in ? _GEN_26809 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2233 = 12'h8b9 == _T_2[11:0] ? image_2233 : _GEN_2232; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5306 = 12'h8ba == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8378 = 12'h8ba == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5306; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11450 = 12'h8ba == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8378; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14522 = 12'h8ba == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11450; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17594 = 12'h8ba == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14522; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20666 = 12'h8ba == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17594; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23738 = 12'h8ba == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20666; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26810 = 12'h8ba == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23738; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2234 = io_valid_in ? _GEN_26810 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2234 = 12'h8ba == _T_2[11:0] ? image_2234 : _GEN_2233; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5307 = 12'h8bb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8379 = 12'h8bb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5307; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11451 = 12'h8bb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8379; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14523 = 12'h8bb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11451; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17595 = 12'h8bb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14523; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20667 = 12'h8bb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17595; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23739 = 12'h8bb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20667; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26811 = 12'h8bb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23739; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2235 = io_valid_in ? _GEN_26811 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2235 = 12'h8bb == _T_2[11:0] ? image_2235 : _GEN_2234; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5308 = 12'h8bc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8380 = 12'h8bc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5308; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11452 = 12'h8bc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8380; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14524 = 12'h8bc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11452; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17596 = 12'h8bc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14524; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20668 = 12'h8bc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17596; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23740 = 12'h8bc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20668; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26812 = 12'h8bc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23740; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2236 = io_valid_in ? _GEN_26812 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2236 = 12'h8bc == _T_2[11:0] ? image_2236 : _GEN_2235; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5309 = 12'h8bd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8381 = 12'h8bd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5309; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11453 = 12'h8bd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8381; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14525 = 12'h8bd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11453; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17597 = 12'h8bd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14525; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20669 = 12'h8bd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17597; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23741 = 12'h8bd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20669; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26813 = 12'h8bd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23741; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2237 = io_valid_in ? _GEN_26813 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2237 = 12'h8bd == _T_2[11:0] ? image_2237 : _GEN_2236; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5310 = 12'h8be == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8382 = 12'h8be == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5310; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11454 = 12'h8be == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8382; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14526 = 12'h8be == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11454; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17598 = 12'h8be == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14526; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20670 = 12'h8be == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17598; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23742 = 12'h8be == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20670; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26814 = 12'h8be == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23742; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2238 = io_valid_in ? _GEN_26814 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2238 = 12'h8be == _T_2[11:0] ? image_2238 : _GEN_2237; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5311 = 12'h8bf == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8383 = 12'h8bf == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5311; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11455 = 12'h8bf == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8383; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14527 = 12'h8bf == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11455; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17599 = 12'h8bf == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14527; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20671 = 12'h8bf == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17599; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23743 = 12'h8bf == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20671; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26815 = 12'h8bf == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23743; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2239 = io_valid_in ? _GEN_26815 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2239 = 12'h8bf == _T_2[11:0] ? image_2239 : _GEN_2238; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5312 = 12'h8c0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8384 = 12'h8c0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5312; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11456 = 12'h8c0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8384; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14528 = 12'h8c0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11456; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17600 = 12'h8c0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14528; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20672 = 12'h8c0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17600; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23744 = 12'h8c0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20672; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26816 = 12'h8c0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23744; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2240 = io_valid_in ? _GEN_26816 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2240 = 12'h8c0 == _T_2[11:0] ? image_2240 : _GEN_2239; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5313 = 12'h8c1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8385 = 12'h8c1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5313; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11457 = 12'h8c1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8385; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14529 = 12'h8c1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11457; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17601 = 12'h8c1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14529; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20673 = 12'h8c1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17601; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23745 = 12'h8c1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20673; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26817 = 12'h8c1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23745; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2241 = io_valid_in ? _GEN_26817 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2241 = 12'h8c1 == _T_2[11:0] ? image_2241 : _GEN_2240; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5314 = 12'h8c2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8386 = 12'h8c2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5314; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11458 = 12'h8c2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8386; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14530 = 12'h8c2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11458; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17602 = 12'h8c2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14530; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20674 = 12'h8c2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17602; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23746 = 12'h8c2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20674; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26818 = 12'h8c2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23746; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2242 = io_valid_in ? _GEN_26818 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2242 = 12'h8c2 == _T_2[11:0] ? image_2242 : _GEN_2241; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5315 = 12'h8c3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8387 = 12'h8c3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5315; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11459 = 12'h8c3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8387; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14531 = 12'h8c3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11459; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17603 = 12'h8c3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14531; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20675 = 12'h8c3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17603; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23747 = 12'h8c3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20675; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26819 = 12'h8c3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23747; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2243 = io_valid_in ? _GEN_26819 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2243 = 12'h8c3 == _T_2[11:0] ? image_2243 : _GEN_2242; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5316 = 12'h8c4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8388 = 12'h8c4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5316; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11460 = 12'h8c4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8388; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14532 = 12'h8c4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11460; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17604 = 12'h8c4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14532; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20676 = 12'h8c4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17604; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23748 = 12'h8c4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20676; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26820 = 12'h8c4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23748; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2244 = io_valid_in ? _GEN_26820 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2244 = 12'h8c4 == _T_2[11:0] ? image_2244 : _GEN_2243; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5317 = 12'h8c5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8389 = 12'h8c5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5317; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11461 = 12'h8c5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8389; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14533 = 12'h8c5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11461; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17605 = 12'h8c5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14533; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20677 = 12'h8c5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17605; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23749 = 12'h8c5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20677; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26821 = 12'h8c5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23749; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2245 = io_valid_in ? _GEN_26821 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2245 = 12'h8c5 == _T_2[11:0] ? image_2245 : _GEN_2244; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5318 = 12'h8c6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8390 = 12'h8c6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5318; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11462 = 12'h8c6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8390; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14534 = 12'h8c6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11462; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17606 = 12'h8c6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14534; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20678 = 12'h8c6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17606; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23750 = 12'h8c6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20678; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26822 = 12'h8c6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23750; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2246 = io_valid_in ? _GEN_26822 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2246 = 12'h8c6 == _T_2[11:0] ? image_2246 : _GEN_2245; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5319 = 12'h8c7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8391 = 12'h8c7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5319; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11463 = 12'h8c7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8391; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14535 = 12'h8c7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11463; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17607 = 12'h8c7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14535; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20679 = 12'h8c7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17607; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23751 = 12'h8c7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20679; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26823 = 12'h8c7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23751; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2247 = io_valid_in ? _GEN_26823 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2247 = 12'h8c7 == _T_2[11:0] ? image_2247 : _GEN_2246; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5320 = 12'h8c8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8392 = 12'h8c8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5320; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11464 = 12'h8c8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8392; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14536 = 12'h8c8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11464; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17608 = 12'h8c8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14536; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20680 = 12'h8c8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17608; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23752 = 12'h8c8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20680; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26824 = 12'h8c8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23752; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2248 = io_valid_in ? _GEN_26824 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2248 = 12'h8c8 == _T_2[11:0] ? image_2248 : _GEN_2247; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5321 = 12'h8c9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8393 = 12'h8c9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5321; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11465 = 12'h8c9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8393; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14537 = 12'h8c9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11465; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17609 = 12'h8c9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14537; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20681 = 12'h8c9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17609; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23753 = 12'h8c9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20681; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26825 = 12'h8c9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23753; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2249 = io_valid_in ? _GEN_26825 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2249 = 12'h8c9 == _T_2[11:0] ? image_2249 : _GEN_2248; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5322 = 12'h8ca == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8394 = 12'h8ca == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5322; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11466 = 12'h8ca == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8394; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14538 = 12'h8ca == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11466; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17610 = 12'h8ca == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14538; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20682 = 12'h8ca == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17610; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23754 = 12'h8ca == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20682; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26826 = 12'h8ca == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23754; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2250 = io_valid_in ? _GEN_26826 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2250 = 12'h8ca == _T_2[11:0] ? image_2250 : _GEN_2249; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5323 = 12'h8cb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8395 = 12'h8cb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5323; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11467 = 12'h8cb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8395; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14539 = 12'h8cb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11467; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17611 = 12'h8cb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14539; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20683 = 12'h8cb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17611; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23755 = 12'h8cb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20683; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26827 = 12'h8cb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23755; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2251 = io_valid_in ? _GEN_26827 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2251 = 12'h8cb == _T_2[11:0] ? image_2251 : _GEN_2250; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5324 = 12'h8cc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8396 = 12'h8cc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5324; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11468 = 12'h8cc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8396; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14540 = 12'h8cc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11468; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17612 = 12'h8cc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14540; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20684 = 12'h8cc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17612; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23756 = 12'h8cc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20684; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26828 = 12'h8cc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23756; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2252 = io_valid_in ? _GEN_26828 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2252 = 12'h8cc == _T_2[11:0] ? image_2252 : _GEN_2251; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5325 = 12'h8cd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8397 = 12'h8cd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5325; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11469 = 12'h8cd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8397; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14541 = 12'h8cd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11469; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17613 = 12'h8cd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14541; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20685 = 12'h8cd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17613; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23757 = 12'h8cd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20685; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26829 = 12'h8cd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23757; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2253 = io_valid_in ? _GEN_26829 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2253 = 12'h8cd == _T_2[11:0] ? image_2253 : _GEN_2252; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5326 = 12'h8ce == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8398 = 12'h8ce == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5326; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11470 = 12'h8ce == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8398; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14542 = 12'h8ce == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11470; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17614 = 12'h8ce == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14542; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20686 = 12'h8ce == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17614; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23758 = 12'h8ce == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20686; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26830 = 12'h8ce == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23758; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2254 = io_valid_in ? _GEN_26830 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2254 = 12'h8ce == _T_2[11:0] ? image_2254 : _GEN_2253; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5327 = 12'h8cf == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8399 = 12'h8cf == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5327; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11471 = 12'h8cf == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8399; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14543 = 12'h8cf == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11471; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17615 = 12'h8cf == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14543; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20687 = 12'h8cf == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17615; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23759 = 12'h8cf == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20687; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26831 = 12'h8cf == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23759; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2255 = io_valid_in ? _GEN_26831 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2255 = 12'h8cf == _T_2[11:0] ? image_2255 : _GEN_2254; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5328 = 12'h8d0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8400 = 12'h8d0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5328; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11472 = 12'h8d0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8400; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14544 = 12'h8d0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11472; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17616 = 12'h8d0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14544; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20688 = 12'h8d0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17616; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23760 = 12'h8d0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20688; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26832 = 12'h8d0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23760; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2256 = io_valid_in ? _GEN_26832 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2256 = 12'h8d0 == _T_2[11:0] ? image_2256 : _GEN_2255; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5329 = 12'h8d1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8401 = 12'h8d1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5329; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11473 = 12'h8d1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8401; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14545 = 12'h8d1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11473; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17617 = 12'h8d1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14545; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20689 = 12'h8d1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17617; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23761 = 12'h8d1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20689; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26833 = 12'h8d1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23761; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2257 = io_valid_in ? _GEN_26833 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2257 = 12'h8d1 == _T_2[11:0] ? image_2257 : _GEN_2256; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5330 = 12'h8d2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8402 = 12'h8d2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5330; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11474 = 12'h8d2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8402; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14546 = 12'h8d2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11474; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17618 = 12'h8d2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14546; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20690 = 12'h8d2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17618; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23762 = 12'h8d2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20690; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26834 = 12'h8d2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23762; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2258 = io_valid_in ? _GEN_26834 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2258 = 12'h8d2 == _T_2[11:0] ? image_2258 : _GEN_2257; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5331 = 12'h8d3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8403 = 12'h8d3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5331; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11475 = 12'h8d3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8403; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14547 = 12'h8d3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11475; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17619 = 12'h8d3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14547; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20691 = 12'h8d3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17619; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23763 = 12'h8d3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20691; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26835 = 12'h8d3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23763; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2259 = io_valid_in ? _GEN_26835 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2259 = 12'h8d3 == _T_2[11:0] ? image_2259 : _GEN_2258; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5332 = 12'h8d4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8404 = 12'h8d4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5332; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11476 = 12'h8d4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8404; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14548 = 12'h8d4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11476; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17620 = 12'h8d4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14548; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20692 = 12'h8d4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17620; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23764 = 12'h8d4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20692; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26836 = 12'h8d4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23764; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2260 = io_valid_in ? _GEN_26836 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2260 = 12'h8d4 == _T_2[11:0] ? image_2260 : _GEN_2259; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5333 = 12'h8d5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8405 = 12'h8d5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5333; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11477 = 12'h8d5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8405; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14549 = 12'h8d5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11477; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17621 = 12'h8d5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14549; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20693 = 12'h8d5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17621; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23765 = 12'h8d5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20693; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26837 = 12'h8d5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23765; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2261 = io_valid_in ? _GEN_26837 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2261 = 12'h8d5 == _T_2[11:0] ? image_2261 : _GEN_2260; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5334 = 12'h8d6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8406 = 12'h8d6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5334; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11478 = 12'h8d6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8406; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14550 = 12'h8d6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11478; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17622 = 12'h8d6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14550; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20694 = 12'h8d6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17622; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23766 = 12'h8d6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20694; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26838 = 12'h8d6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23766; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2262 = io_valid_in ? _GEN_26838 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2262 = 12'h8d6 == _T_2[11:0] ? image_2262 : _GEN_2261; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5335 = 12'h8d7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8407 = 12'h8d7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5335; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11479 = 12'h8d7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8407; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14551 = 12'h8d7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11479; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17623 = 12'h8d7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14551; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20695 = 12'h8d7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17623; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23767 = 12'h8d7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20695; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26839 = 12'h8d7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23767; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2263 = io_valid_in ? _GEN_26839 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2263 = 12'h8d7 == _T_2[11:0] ? image_2263 : _GEN_2262; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5336 = 12'h8d8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8408 = 12'h8d8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5336; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11480 = 12'h8d8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8408; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14552 = 12'h8d8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11480; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17624 = 12'h8d8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14552; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20696 = 12'h8d8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17624; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23768 = 12'h8d8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20696; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26840 = 12'h8d8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23768; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2264 = io_valid_in ? _GEN_26840 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2264 = 12'h8d8 == _T_2[11:0] ? image_2264 : _GEN_2263; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5337 = 12'h8d9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8409 = 12'h8d9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5337; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11481 = 12'h8d9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8409; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14553 = 12'h8d9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11481; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17625 = 12'h8d9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14553; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20697 = 12'h8d9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17625; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23769 = 12'h8d9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20697; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26841 = 12'h8d9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23769; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2265 = io_valid_in ? _GEN_26841 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2265 = 12'h8d9 == _T_2[11:0] ? image_2265 : _GEN_2264; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5338 = 12'h8da == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8410 = 12'h8da == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5338; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11482 = 12'h8da == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8410; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14554 = 12'h8da == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11482; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17626 = 12'h8da == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14554; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20698 = 12'h8da == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17626; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23770 = 12'h8da == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20698; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26842 = 12'h8da == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23770; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2266 = io_valid_in ? _GEN_26842 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2266 = 12'h8da == _T_2[11:0] ? image_2266 : _GEN_2265; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5339 = 12'h8db == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8411 = 12'h8db == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5339; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11483 = 12'h8db == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8411; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14555 = 12'h8db == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11483; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17627 = 12'h8db == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14555; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20699 = 12'h8db == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17627; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23771 = 12'h8db == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20699; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26843 = 12'h8db == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23771; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2267 = io_valid_in ? _GEN_26843 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2267 = 12'h8db == _T_2[11:0] ? image_2267 : _GEN_2266; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5340 = 12'h8dc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8412 = 12'h8dc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5340; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11484 = 12'h8dc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8412; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14556 = 12'h8dc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11484; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17628 = 12'h8dc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14556; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20700 = 12'h8dc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17628; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23772 = 12'h8dc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20700; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26844 = 12'h8dc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23772; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2268 = io_valid_in ? _GEN_26844 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2268 = 12'h8dc == _T_2[11:0] ? image_2268 : _GEN_2267; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5341 = 12'h8dd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8413 = 12'h8dd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5341; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11485 = 12'h8dd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8413; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14557 = 12'h8dd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11485; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17629 = 12'h8dd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14557; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20701 = 12'h8dd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17629; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23773 = 12'h8dd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20701; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26845 = 12'h8dd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23773; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2269 = io_valid_in ? _GEN_26845 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2269 = 12'h8dd == _T_2[11:0] ? image_2269 : _GEN_2268; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5342 = 12'h8de == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8414 = 12'h8de == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5342; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11486 = 12'h8de == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8414; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14558 = 12'h8de == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11486; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17630 = 12'h8de == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14558; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20702 = 12'h8de == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17630; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23774 = 12'h8de == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20702; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26846 = 12'h8de == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23774; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2270 = io_valid_in ? _GEN_26846 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2270 = 12'h8de == _T_2[11:0] ? image_2270 : _GEN_2269; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5343 = 12'h8df == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8415 = 12'h8df == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5343; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11487 = 12'h8df == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8415; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14559 = 12'h8df == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11487; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17631 = 12'h8df == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14559; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20703 = 12'h8df == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17631; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23775 = 12'h8df == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20703; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26847 = 12'h8df == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23775; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2271 = io_valid_in ? _GEN_26847 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2271 = 12'h8df == _T_2[11:0] ? image_2271 : _GEN_2270; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5344 = 12'h8e0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8416 = 12'h8e0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5344; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11488 = 12'h8e0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8416; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14560 = 12'h8e0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11488; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17632 = 12'h8e0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14560; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20704 = 12'h8e0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17632; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23776 = 12'h8e0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20704; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26848 = 12'h8e0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23776; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2272 = io_valid_in ? _GEN_26848 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2272 = 12'h8e0 == _T_2[11:0] ? image_2272 : _GEN_2271; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5345 = 12'h8e1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8417 = 12'h8e1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5345; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11489 = 12'h8e1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8417; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14561 = 12'h8e1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11489; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17633 = 12'h8e1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14561; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20705 = 12'h8e1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17633; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23777 = 12'h8e1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20705; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26849 = 12'h8e1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23777; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2273 = io_valid_in ? _GEN_26849 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2273 = 12'h8e1 == _T_2[11:0] ? image_2273 : _GEN_2272; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5346 = 12'h8e2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8418 = 12'h8e2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5346; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11490 = 12'h8e2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8418; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14562 = 12'h8e2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11490; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17634 = 12'h8e2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14562; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20706 = 12'h8e2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17634; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23778 = 12'h8e2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20706; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26850 = 12'h8e2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23778; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2274 = io_valid_in ? _GEN_26850 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2274 = 12'h8e2 == _T_2[11:0] ? image_2274 : _GEN_2273; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5347 = 12'h8e3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8419 = 12'h8e3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5347; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11491 = 12'h8e3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8419; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14563 = 12'h8e3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11491; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17635 = 12'h8e3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14563; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20707 = 12'h8e3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17635; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23779 = 12'h8e3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20707; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26851 = 12'h8e3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23779; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2275 = io_valid_in ? _GEN_26851 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2275 = 12'h8e3 == _T_2[11:0] ? image_2275 : _GEN_2274; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5348 = 12'h8e4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8420 = 12'h8e4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5348; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11492 = 12'h8e4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8420; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14564 = 12'h8e4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11492; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17636 = 12'h8e4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14564; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20708 = 12'h8e4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17636; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23780 = 12'h8e4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20708; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26852 = 12'h8e4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23780; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2276 = io_valid_in ? _GEN_26852 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2276 = 12'h8e4 == _T_2[11:0] ? image_2276 : _GEN_2275; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5349 = 12'h8e5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8421 = 12'h8e5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5349; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11493 = 12'h8e5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8421; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14565 = 12'h8e5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11493; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17637 = 12'h8e5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14565; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20709 = 12'h8e5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17637; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23781 = 12'h8e5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20709; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26853 = 12'h8e5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23781; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2277 = io_valid_in ? _GEN_26853 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2277 = 12'h8e5 == _T_2[11:0] ? image_2277 : _GEN_2276; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5350 = 12'h8e6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8422 = 12'h8e6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5350; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11494 = 12'h8e6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8422; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14566 = 12'h8e6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11494; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17638 = 12'h8e6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14566; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20710 = 12'h8e6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17638; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23782 = 12'h8e6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20710; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26854 = 12'h8e6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23782; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2278 = io_valid_in ? _GEN_26854 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2278 = 12'h8e6 == _T_2[11:0] ? image_2278 : _GEN_2277; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5351 = 12'h8e7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8423 = 12'h8e7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5351; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11495 = 12'h8e7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8423; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14567 = 12'h8e7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11495; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17639 = 12'h8e7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14567; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20711 = 12'h8e7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17639; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23783 = 12'h8e7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20711; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26855 = 12'h8e7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23783; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2279 = io_valid_in ? _GEN_26855 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2279 = 12'h8e7 == _T_2[11:0] ? image_2279 : _GEN_2278; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5352 = 12'h8e8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8424 = 12'h8e8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5352; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11496 = 12'h8e8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8424; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14568 = 12'h8e8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11496; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17640 = 12'h8e8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14568; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20712 = 12'h8e8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17640; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23784 = 12'h8e8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20712; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26856 = 12'h8e8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23784; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2280 = io_valid_in ? _GEN_26856 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2280 = 12'h8e8 == _T_2[11:0] ? image_2280 : _GEN_2279; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5353 = 12'h8e9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8425 = 12'h8e9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5353; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11497 = 12'h8e9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8425; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14569 = 12'h8e9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11497; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17641 = 12'h8e9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14569; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20713 = 12'h8e9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17641; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23785 = 12'h8e9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20713; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26857 = 12'h8e9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23785; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2281 = io_valid_in ? _GEN_26857 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2281 = 12'h8e9 == _T_2[11:0] ? image_2281 : _GEN_2280; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5354 = 12'h8ea == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8426 = 12'h8ea == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5354; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11498 = 12'h8ea == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8426; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14570 = 12'h8ea == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11498; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17642 = 12'h8ea == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14570; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20714 = 12'h8ea == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17642; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23786 = 12'h8ea == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20714; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26858 = 12'h8ea == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23786; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2282 = io_valid_in ? _GEN_26858 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2282 = 12'h8ea == _T_2[11:0] ? image_2282 : _GEN_2281; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5355 = 12'h8eb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8427 = 12'h8eb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5355; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11499 = 12'h8eb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8427; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14571 = 12'h8eb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11499; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17643 = 12'h8eb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14571; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20715 = 12'h8eb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17643; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23787 = 12'h8eb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20715; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26859 = 12'h8eb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23787; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2283 = io_valid_in ? _GEN_26859 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2283 = 12'h8eb == _T_2[11:0] ? image_2283 : _GEN_2282; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5356 = 12'h8ec == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8428 = 12'h8ec == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5356; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11500 = 12'h8ec == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8428; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14572 = 12'h8ec == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11500; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17644 = 12'h8ec == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14572; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20716 = 12'h8ec == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17644; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23788 = 12'h8ec == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20716; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26860 = 12'h8ec == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23788; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2284 = io_valid_in ? _GEN_26860 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2284 = 12'h8ec == _T_2[11:0] ? image_2284 : _GEN_2283; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5357 = 12'h8ed == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8429 = 12'h8ed == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5357; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11501 = 12'h8ed == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8429; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14573 = 12'h8ed == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11501; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17645 = 12'h8ed == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14573; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20717 = 12'h8ed == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17645; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23789 = 12'h8ed == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20717; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26861 = 12'h8ed == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23789; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2285 = io_valid_in ? _GEN_26861 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2285 = 12'h8ed == _T_2[11:0] ? image_2285 : _GEN_2284; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5358 = 12'h8ee == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8430 = 12'h8ee == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5358; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11502 = 12'h8ee == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8430; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14574 = 12'h8ee == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11502; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17646 = 12'h8ee == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14574; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20718 = 12'h8ee == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17646; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23790 = 12'h8ee == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20718; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26862 = 12'h8ee == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23790; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2286 = io_valid_in ? _GEN_26862 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2286 = 12'h8ee == _T_2[11:0] ? image_2286 : _GEN_2285; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5359 = 12'h8ef == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8431 = 12'h8ef == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5359; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11503 = 12'h8ef == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8431; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14575 = 12'h8ef == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11503; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17647 = 12'h8ef == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14575; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20719 = 12'h8ef == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17647; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23791 = 12'h8ef == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20719; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26863 = 12'h8ef == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23791; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2287 = io_valid_in ? _GEN_26863 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2287 = 12'h8ef == _T_2[11:0] ? image_2287 : _GEN_2286; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5360 = 12'h8f0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8432 = 12'h8f0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5360; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11504 = 12'h8f0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8432; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14576 = 12'h8f0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11504; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17648 = 12'h8f0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14576; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20720 = 12'h8f0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17648; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23792 = 12'h8f0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20720; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26864 = 12'h8f0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23792; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2288 = io_valid_in ? _GEN_26864 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2288 = 12'h8f0 == _T_2[11:0] ? image_2288 : _GEN_2287; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5361 = 12'h8f1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8433 = 12'h8f1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5361; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11505 = 12'h8f1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8433; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14577 = 12'h8f1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11505; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17649 = 12'h8f1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14577; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20721 = 12'h8f1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17649; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23793 = 12'h8f1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20721; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26865 = 12'h8f1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23793; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2289 = io_valid_in ? _GEN_26865 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2289 = 12'h8f1 == _T_2[11:0] ? image_2289 : _GEN_2288; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5362 = 12'h8f2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8434 = 12'h8f2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5362; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11506 = 12'h8f2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8434; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14578 = 12'h8f2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11506; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17650 = 12'h8f2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14578; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20722 = 12'h8f2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17650; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23794 = 12'h8f2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20722; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26866 = 12'h8f2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23794; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2290 = io_valid_in ? _GEN_26866 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2290 = 12'h8f2 == _T_2[11:0] ? image_2290 : _GEN_2289; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5363 = 12'h8f3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8435 = 12'h8f3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5363; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11507 = 12'h8f3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8435; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14579 = 12'h8f3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11507; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17651 = 12'h8f3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14579; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20723 = 12'h8f3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17651; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23795 = 12'h8f3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20723; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26867 = 12'h8f3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23795; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2291 = io_valid_in ? _GEN_26867 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2291 = 12'h8f3 == _T_2[11:0] ? image_2291 : _GEN_2290; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5364 = 12'h8f4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8436 = 12'h8f4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5364; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11508 = 12'h8f4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8436; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14580 = 12'h8f4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11508; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17652 = 12'h8f4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14580; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20724 = 12'h8f4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17652; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23796 = 12'h8f4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20724; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26868 = 12'h8f4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23796; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2292 = io_valid_in ? _GEN_26868 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2292 = 12'h8f4 == _T_2[11:0] ? image_2292 : _GEN_2291; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5365 = 12'h8f5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8437 = 12'h8f5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5365; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11509 = 12'h8f5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8437; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14581 = 12'h8f5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11509; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17653 = 12'h8f5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14581; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20725 = 12'h8f5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17653; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23797 = 12'h8f5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20725; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26869 = 12'h8f5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23797; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2293 = io_valid_in ? _GEN_26869 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2293 = 12'h8f5 == _T_2[11:0] ? image_2293 : _GEN_2292; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5366 = 12'h8f6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8438 = 12'h8f6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5366; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11510 = 12'h8f6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8438; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14582 = 12'h8f6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11510; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17654 = 12'h8f6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14582; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20726 = 12'h8f6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17654; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23798 = 12'h8f6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20726; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26870 = 12'h8f6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23798; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2294 = io_valid_in ? _GEN_26870 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2294 = 12'h8f6 == _T_2[11:0] ? image_2294 : _GEN_2293; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5367 = 12'h8f7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8439 = 12'h8f7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5367; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11511 = 12'h8f7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8439; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14583 = 12'h8f7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11511; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17655 = 12'h8f7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14583; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20727 = 12'h8f7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17655; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23799 = 12'h8f7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20727; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26871 = 12'h8f7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23799; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2295 = io_valid_in ? _GEN_26871 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2295 = 12'h8f7 == _T_2[11:0] ? image_2295 : _GEN_2294; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5368 = 12'h8f8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8440 = 12'h8f8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5368; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11512 = 12'h8f8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8440; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14584 = 12'h8f8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11512; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17656 = 12'h8f8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14584; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20728 = 12'h8f8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17656; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23800 = 12'h8f8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20728; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26872 = 12'h8f8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23800; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2296 = io_valid_in ? _GEN_26872 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2296 = 12'h8f8 == _T_2[11:0] ? image_2296 : _GEN_2295; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5369 = 12'h8f9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8441 = 12'h8f9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5369; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11513 = 12'h8f9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8441; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14585 = 12'h8f9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11513; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17657 = 12'h8f9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14585; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20729 = 12'h8f9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17657; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23801 = 12'h8f9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20729; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26873 = 12'h8f9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23801; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2297 = io_valid_in ? _GEN_26873 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2297 = 12'h8f9 == _T_2[11:0] ? image_2297 : _GEN_2296; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5370 = 12'h8fa == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8442 = 12'h8fa == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5370; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11514 = 12'h8fa == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8442; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14586 = 12'h8fa == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11514; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17658 = 12'h8fa == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14586; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20730 = 12'h8fa == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17658; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23802 = 12'h8fa == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20730; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26874 = 12'h8fa == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23802; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2298 = io_valid_in ? _GEN_26874 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2298 = 12'h8fa == _T_2[11:0] ? image_2298 : _GEN_2297; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5371 = 12'h8fb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8443 = 12'h8fb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5371; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11515 = 12'h8fb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8443; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14587 = 12'h8fb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11515; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17659 = 12'h8fb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14587; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20731 = 12'h8fb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17659; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23803 = 12'h8fb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20731; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26875 = 12'h8fb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23803; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2299 = io_valid_in ? _GEN_26875 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2299 = 12'h8fb == _T_2[11:0] ? image_2299 : _GEN_2298; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5372 = 12'h8fc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8444 = 12'h8fc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5372; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11516 = 12'h8fc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8444; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14588 = 12'h8fc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11516; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17660 = 12'h8fc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14588; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20732 = 12'h8fc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17660; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23804 = 12'h8fc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20732; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26876 = 12'h8fc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23804; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2300 = io_valid_in ? _GEN_26876 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2300 = 12'h8fc == _T_2[11:0] ? image_2300 : _GEN_2299; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5373 = 12'h8fd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8445 = 12'h8fd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5373; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11517 = 12'h8fd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8445; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14589 = 12'h8fd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11517; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17661 = 12'h8fd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14589; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20733 = 12'h8fd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17661; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23805 = 12'h8fd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20733; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26877 = 12'h8fd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23805; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2301 = io_valid_in ? _GEN_26877 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2301 = 12'h8fd == _T_2[11:0] ? image_2301 : _GEN_2300; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5374 = 12'h8fe == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8446 = 12'h8fe == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5374; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11518 = 12'h8fe == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8446; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14590 = 12'h8fe == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11518; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17662 = 12'h8fe == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14590; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20734 = 12'h8fe == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17662; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23806 = 12'h8fe == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20734; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26878 = 12'h8fe == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23806; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2302 = io_valid_in ? _GEN_26878 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2302 = 12'h8fe == _T_2[11:0] ? image_2302 : _GEN_2301; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5375 = 12'h8ff == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8447 = 12'h8ff == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5375; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11519 = 12'h8ff == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8447; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14591 = 12'h8ff == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11519; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17663 = 12'h8ff == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14591; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20735 = 12'h8ff == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17663; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23807 = 12'h8ff == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20735; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26879 = 12'h8ff == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23807; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2303 = io_valid_in ? _GEN_26879 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2303 = 12'h8ff == _T_2[11:0] ? image_2303 : _GEN_2302; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5376 = 12'h900 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8448 = 12'h900 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5376; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11520 = 12'h900 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8448; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14592 = 12'h900 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11520; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17664 = 12'h900 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14592; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20736 = 12'h900 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17664; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23808 = 12'h900 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20736; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26880 = 12'h900 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23808; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2304 = io_valid_in ? _GEN_26880 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2304 = 12'h900 == _T_2[11:0] ? image_2304 : _GEN_2303; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5377 = 12'h901 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8449 = 12'h901 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5377; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11521 = 12'h901 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8449; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14593 = 12'h901 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11521; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17665 = 12'h901 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14593; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20737 = 12'h901 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17665; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23809 = 12'h901 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20737; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26881 = 12'h901 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23809; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2305 = io_valid_in ? _GEN_26881 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2305 = 12'h901 == _T_2[11:0] ? image_2305 : _GEN_2304; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5378 = 12'h902 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8450 = 12'h902 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5378; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11522 = 12'h902 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8450; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14594 = 12'h902 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11522; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17666 = 12'h902 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14594; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20738 = 12'h902 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17666; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23810 = 12'h902 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20738; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26882 = 12'h902 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23810; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2306 = io_valid_in ? _GEN_26882 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2306 = 12'h902 == _T_2[11:0] ? image_2306 : _GEN_2305; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5379 = 12'h903 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8451 = 12'h903 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5379; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11523 = 12'h903 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8451; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14595 = 12'h903 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11523; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17667 = 12'h903 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14595; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20739 = 12'h903 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17667; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23811 = 12'h903 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20739; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26883 = 12'h903 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23811; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2307 = io_valid_in ? _GEN_26883 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2307 = 12'h903 == _T_2[11:0] ? image_2307 : _GEN_2306; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5380 = 12'h904 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8452 = 12'h904 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5380; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11524 = 12'h904 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8452; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14596 = 12'h904 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11524; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17668 = 12'h904 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14596; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20740 = 12'h904 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17668; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23812 = 12'h904 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20740; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26884 = 12'h904 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23812; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2308 = io_valid_in ? _GEN_26884 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2308 = 12'h904 == _T_2[11:0] ? image_2308 : _GEN_2307; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5381 = 12'h905 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8453 = 12'h905 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5381; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11525 = 12'h905 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8453; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14597 = 12'h905 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11525; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17669 = 12'h905 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14597; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20741 = 12'h905 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17669; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23813 = 12'h905 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20741; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26885 = 12'h905 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23813; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2309 = io_valid_in ? _GEN_26885 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2309 = 12'h905 == _T_2[11:0] ? image_2309 : _GEN_2308; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5382 = 12'h906 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8454 = 12'h906 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5382; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11526 = 12'h906 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8454; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14598 = 12'h906 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11526; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17670 = 12'h906 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14598; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20742 = 12'h906 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17670; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23814 = 12'h906 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20742; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26886 = 12'h906 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23814; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2310 = io_valid_in ? _GEN_26886 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2310 = 12'h906 == _T_2[11:0] ? image_2310 : _GEN_2309; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5383 = 12'h907 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8455 = 12'h907 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5383; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11527 = 12'h907 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8455; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14599 = 12'h907 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11527; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17671 = 12'h907 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14599; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20743 = 12'h907 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17671; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23815 = 12'h907 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20743; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26887 = 12'h907 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23815; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2311 = io_valid_in ? _GEN_26887 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2311 = 12'h907 == _T_2[11:0] ? image_2311 : _GEN_2310; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5384 = 12'h908 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8456 = 12'h908 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5384; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11528 = 12'h908 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8456; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14600 = 12'h908 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11528; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17672 = 12'h908 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14600; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20744 = 12'h908 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17672; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23816 = 12'h908 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20744; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26888 = 12'h908 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23816; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2312 = io_valid_in ? _GEN_26888 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2312 = 12'h908 == _T_2[11:0] ? image_2312 : _GEN_2311; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5385 = 12'h909 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8457 = 12'h909 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5385; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11529 = 12'h909 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8457; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14601 = 12'h909 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11529; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17673 = 12'h909 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14601; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20745 = 12'h909 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17673; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23817 = 12'h909 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20745; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26889 = 12'h909 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23817; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2313 = io_valid_in ? _GEN_26889 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2313 = 12'h909 == _T_2[11:0] ? image_2313 : _GEN_2312; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5386 = 12'h90a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8458 = 12'h90a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5386; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11530 = 12'h90a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8458; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14602 = 12'h90a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11530; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17674 = 12'h90a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14602; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20746 = 12'h90a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17674; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23818 = 12'h90a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20746; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26890 = 12'h90a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23818; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2314 = io_valid_in ? _GEN_26890 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2314 = 12'h90a == _T_2[11:0] ? image_2314 : _GEN_2313; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5387 = 12'h90b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8459 = 12'h90b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5387; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11531 = 12'h90b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8459; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14603 = 12'h90b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11531; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17675 = 12'h90b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14603; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20747 = 12'h90b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17675; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23819 = 12'h90b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20747; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26891 = 12'h90b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23819; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2315 = io_valid_in ? _GEN_26891 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2315 = 12'h90b == _T_2[11:0] ? image_2315 : _GEN_2314; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5388 = 12'h90c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8460 = 12'h90c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5388; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11532 = 12'h90c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8460; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14604 = 12'h90c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11532; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17676 = 12'h90c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14604; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20748 = 12'h90c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17676; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23820 = 12'h90c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20748; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26892 = 12'h90c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23820; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2316 = io_valid_in ? _GEN_26892 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2316 = 12'h90c == _T_2[11:0] ? image_2316 : _GEN_2315; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5389 = 12'h90d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8461 = 12'h90d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5389; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11533 = 12'h90d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8461; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14605 = 12'h90d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11533; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17677 = 12'h90d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14605; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20749 = 12'h90d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17677; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23821 = 12'h90d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20749; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26893 = 12'h90d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23821; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2317 = io_valid_in ? _GEN_26893 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2317 = 12'h90d == _T_2[11:0] ? image_2317 : _GEN_2316; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5390 = 12'h90e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8462 = 12'h90e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5390; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11534 = 12'h90e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8462; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14606 = 12'h90e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11534; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17678 = 12'h90e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14606; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20750 = 12'h90e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17678; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23822 = 12'h90e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20750; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26894 = 12'h90e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23822; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2318 = io_valid_in ? _GEN_26894 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2318 = 12'h90e == _T_2[11:0] ? image_2318 : _GEN_2317; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5391 = 12'h90f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8463 = 12'h90f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5391; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11535 = 12'h90f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8463; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14607 = 12'h90f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11535; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17679 = 12'h90f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14607; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20751 = 12'h90f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17679; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23823 = 12'h90f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20751; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26895 = 12'h90f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23823; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2319 = io_valid_in ? _GEN_26895 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2319 = 12'h90f == _T_2[11:0] ? image_2319 : _GEN_2318; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5392 = 12'h910 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8464 = 12'h910 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5392; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11536 = 12'h910 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8464; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14608 = 12'h910 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11536; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17680 = 12'h910 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14608; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20752 = 12'h910 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17680; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23824 = 12'h910 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20752; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26896 = 12'h910 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23824; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2320 = io_valid_in ? _GEN_26896 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2320 = 12'h910 == _T_2[11:0] ? image_2320 : _GEN_2319; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5393 = 12'h911 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8465 = 12'h911 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5393; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11537 = 12'h911 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8465; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14609 = 12'h911 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11537; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17681 = 12'h911 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14609; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20753 = 12'h911 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17681; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23825 = 12'h911 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20753; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26897 = 12'h911 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23825; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2321 = io_valid_in ? _GEN_26897 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2321 = 12'h911 == _T_2[11:0] ? image_2321 : _GEN_2320; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5394 = 12'h912 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8466 = 12'h912 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5394; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11538 = 12'h912 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8466; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14610 = 12'h912 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11538; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17682 = 12'h912 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14610; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20754 = 12'h912 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17682; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23826 = 12'h912 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20754; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26898 = 12'h912 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23826; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2322 = io_valid_in ? _GEN_26898 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2322 = 12'h912 == _T_2[11:0] ? image_2322 : _GEN_2321; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5395 = 12'h913 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8467 = 12'h913 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5395; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11539 = 12'h913 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8467; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14611 = 12'h913 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11539; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17683 = 12'h913 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14611; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20755 = 12'h913 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17683; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23827 = 12'h913 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20755; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26899 = 12'h913 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23827; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2323 = io_valid_in ? _GEN_26899 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2323 = 12'h913 == _T_2[11:0] ? image_2323 : _GEN_2322; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5396 = 12'h914 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8468 = 12'h914 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5396; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11540 = 12'h914 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8468; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14612 = 12'h914 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11540; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17684 = 12'h914 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14612; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20756 = 12'h914 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17684; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23828 = 12'h914 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20756; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26900 = 12'h914 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23828; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2324 = io_valid_in ? _GEN_26900 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2324 = 12'h914 == _T_2[11:0] ? image_2324 : _GEN_2323; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5397 = 12'h915 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8469 = 12'h915 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5397; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11541 = 12'h915 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8469; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14613 = 12'h915 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11541; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17685 = 12'h915 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14613; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20757 = 12'h915 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17685; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23829 = 12'h915 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20757; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26901 = 12'h915 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23829; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2325 = io_valid_in ? _GEN_26901 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2325 = 12'h915 == _T_2[11:0] ? image_2325 : _GEN_2324; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5398 = 12'h916 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8470 = 12'h916 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5398; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11542 = 12'h916 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8470; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14614 = 12'h916 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11542; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17686 = 12'h916 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14614; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20758 = 12'h916 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17686; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23830 = 12'h916 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20758; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26902 = 12'h916 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23830; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2326 = io_valid_in ? _GEN_26902 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2326 = 12'h916 == _T_2[11:0] ? image_2326 : _GEN_2325; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5399 = 12'h917 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8471 = 12'h917 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5399; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11543 = 12'h917 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8471; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14615 = 12'h917 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11543; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17687 = 12'h917 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14615; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20759 = 12'h917 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17687; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23831 = 12'h917 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20759; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26903 = 12'h917 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23831; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2327 = io_valid_in ? _GEN_26903 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2327 = 12'h917 == _T_2[11:0] ? image_2327 : _GEN_2326; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5400 = 12'h918 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8472 = 12'h918 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5400; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11544 = 12'h918 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8472; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14616 = 12'h918 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11544; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17688 = 12'h918 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14616; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20760 = 12'h918 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17688; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23832 = 12'h918 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20760; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26904 = 12'h918 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23832; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2328 = io_valid_in ? _GEN_26904 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2328 = 12'h918 == _T_2[11:0] ? image_2328 : _GEN_2327; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5401 = 12'h919 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8473 = 12'h919 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5401; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11545 = 12'h919 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8473; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14617 = 12'h919 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11545; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17689 = 12'h919 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14617; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20761 = 12'h919 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17689; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23833 = 12'h919 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20761; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26905 = 12'h919 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23833; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2329 = io_valid_in ? _GEN_26905 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2329 = 12'h919 == _T_2[11:0] ? image_2329 : _GEN_2328; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5402 = 12'h91a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8474 = 12'h91a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5402; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11546 = 12'h91a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8474; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14618 = 12'h91a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11546; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17690 = 12'h91a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14618; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20762 = 12'h91a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17690; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23834 = 12'h91a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20762; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26906 = 12'h91a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23834; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2330 = io_valid_in ? _GEN_26906 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2330 = 12'h91a == _T_2[11:0] ? image_2330 : _GEN_2329; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5403 = 12'h91b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8475 = 12'h91b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5403; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11547 = 12'h91b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8475; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14619 = 12'h91b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11547; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17691 = 12'h91b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14619; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20763 = 12'h91b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17691; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23835 = 12'h91b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20763; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26907 = 12'h91b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23835; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2331 = io_valid_in ? _GEN_26907 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2331 = 12'h91b == _T_2[11:0] ? image_2331 : _GEN_2330; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5404 = 12'h91c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8476 = 12'h91c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5404; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11548 = 12'h91c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8476; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14620 = 12'h91c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11548; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17692 = 12'h91c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14620; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20764 = 12'h91c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17692; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23836 = 12'h91c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20764; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26908 = 12'h91c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23836; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2332 = io_valid_in ? _GEN_26908 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2332 = 12'h91c == _T_2[11:0] ? image_2332 : _GEN_2331; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5405 = 12'h91d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8477 = 12'h91d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5405; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11549 = 12'h91d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8477; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14621 = 12'h91d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11549; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17693 = 12'h91d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14621; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20765 = 12'h91d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17693; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23837 = 12'h91d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20765; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26909 = 12'h91d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23837; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2333 = io_valid_in ? _GEN_26909 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2333 = 12'h91d == _T_2[11:0] ? image_2333 : _GEN_2332; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5406 = 12'h91e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8478 = 12'h91e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5406; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11550 = 12'h91e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8478; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14622 = 12'h91e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11550; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17694 = 12'h91e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14622; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20766 = 12'h91e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17694; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23838 = 12'h91e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20766; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26910 = 12'h91e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23838; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2334 = io_valid_in ? _GEN_26910 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2334 = 12'h91e == _T_2[11:0] ? image_2334 : _GEN_2333; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5407 = 12'h91f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8479 = 12'h91f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5407; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11551 = 12'h91f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8479; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14623 = 12'h91f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11551; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17695 = 12'h91f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14623; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20767 = 12'h91f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17695; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23839 = 12'h91f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20767; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26911 = 12'h91f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23839; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2335 = io_valid_in ? _GEN_26911 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2335 = 12'h91f == _T_2[11:0] ? image_2335 : _GEN_2334; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5408 = 12'h920 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8480 = 12'h920 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5408; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11552 = 12'h920 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8480; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14624 = 12'h920 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11552; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17696 = 12'h920 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14624; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20768 = 12'h920 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17696; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23840 = 12'h920 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20768; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26912 = 12'h920 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23840; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2336 = io_valid_in ? _GEN_26912 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2336 = 12'h920 == _T_2[11:0] ? image_2336 : _GEN_2335; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5409 = 12'h921 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8481 = 12'h921 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5409; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11553 = 12'h921 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8481; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14625 = 12'h921 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11553; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17697 = 12'h921 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14625; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20769 = 12'h921 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17697; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23841 = 12'h921 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20769; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26913 = 12'h921 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23841; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2337 = io_valid_in ? _GEN_26913 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2337 = 12'h921 == _T_2[11:0] ? image_2337 : _GEN_2336; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5410 = 12'h922 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8482 = 12'h922 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5410; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11554 = 12'h922 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8482; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14626 = 12'h922 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11554; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17698 = 12'h922 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14626; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20770 = 12'h922 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17698; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23842 = 12'h922 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20770; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26914 = 12'h922 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23842; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2338 = io_valid_in ? _GEN_26914 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2338 = 12'h922 == _T_2[11:0] ? image_2338 : _GEN_2337; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5411 = 12'h923 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8483 = 12'h923 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5411; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11555 = 12'h923 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8483; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14627 = 12'h923 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11555; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17699 = 12'h923 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14627; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20771 = 12'h923 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17699; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23843 = 12'h923 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20771; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26915 = 12'h923 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23843; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2339 = io_valid_in ? _GEN_26915 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2339 = 12'h923 == _T_2[11:0] ? image_2339 : _GEN_2338; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5412 = 12'h924 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8484 = 12'h924 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5412; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11556 = 12'h924 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8484; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14628 = 12'h924 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11556; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17700 = 12'h924 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14628; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20772 = 12'h924 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17700; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23844 = 12'h924 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20772; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26916 = 12'h924 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23844; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2340 = io_valid_in ? _GEN_26916 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2340 = 12'h924 == _T_2[11:0] ? image_2340 : _GEN_2339; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5413 = 12'h925 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8485 = 12'h925 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5413; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11557 = 12'h925 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8485; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14629 = 12'h925 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11557; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17701 = 12'h925 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14629; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20773 = 12'h925 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17701; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23845 = 12'h925 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20773; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26917 = 12'h925 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23845; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2341 = io_valid_in ? _GEN_26917 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2341 = 12'h925 == _T_2[11:0] ? image_2341 : _GEN_2340; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5414 = 12'h926 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8486 = 12'h926 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5414; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11558 = 12'h926 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8486; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14630 = 12'h926 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11558; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17702 = 12'h926 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14630; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20774 = 12'h926 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17702; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23846 = 12'h926 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20774; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26918 = 12'h926 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23846; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2342 = io_valid_in ? _GEN_26918 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2342 = 12'h926 == _T_2[11:0] ? image_2342 : _GEN_2341; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5415 = 12'h927 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8487 = 12'h927 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5415; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11559 = 12'h927 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8487; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14631 = 12'h927 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11559; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17703 = 12'h927 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14631; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20775 = 12'h927 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17703; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23847 = 12'h927 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20775; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26919 = 12'h927 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23847; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2343 = io_valid_in ? _GEN_26919 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2343 = 12'h927 == _T_2[11:0] ? image_2343 : _GEN_2342; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5416 = 12'h928 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8488 = 12'h928 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5416; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11560 = 12'h928 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8488; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14632 = 12'h928 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11560; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17704 = 12'h928 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14632; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20776 = 12'h928 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17704; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23848 = 12'h928 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20776; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26920 = 12'h928 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23848; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2344 = io_valid_in ? _GEN_26920 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2344 = 12'h928 == _T_2[11:0] ? image_2344 : _GEN_2343; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5417 = 12'h929 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8489 = 12'h929 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5417; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11561 = 12'h929 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8489; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14633 = 12'h929 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11561; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17705 = 12'h929 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14633; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20777 = 12'h929 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17705; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23849 = 12'h929 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20777; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26921 = 12'h929 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23849; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2345 = io_valid_in ? _GEN_26921 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2345 = 12'h929 == _T_2[11:0] ? image_2345 : _GEN_2344; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5418 = 12'h92a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8490 = 12'h92a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5418; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11562 = 12'h92a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8490; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14634 = 12'h92a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11562; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17706 = 12'h92a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14634; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20778 = 12'h92a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17706; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23850 = 12'h92a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20778; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26922 = 12'h92a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23850; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2346 = io_valid_in ? _GEN_26922 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2346 = 12'h92a == _T_2[11:0] ? image_2346 : _GEN_2345; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5419 = 12'h92b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8491 = 12'h92b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5419; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11563 = 12'h92b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8491; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14635 = 12'h92b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11563; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17707 = 12'h92b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14635; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20779 = 12'h92b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17707; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23851 = 12'h92b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20779; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26923 = 12'h92b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23851; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2347 = io_valid_in ? _GEN_26923 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2347 = 12'h92b == _T_2[11:0] ? image_2347 : _GEN_2346; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5420 = 12'h92c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8492 = 12'h92c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5420; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11564 = 12'h92c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8492; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14636 = 12'h92c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11564; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17708 = 12'h92c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14636; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20780 = 12'h92c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17708; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23852 = 12'h92c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20780; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26924 = 12'h92c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23852; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2348 = io_valid_in ? _GEN_26924 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2348 = 12'h92c == _T_2[11:0] ? image_2348 : _GEN_2347; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5421 = 12'h92d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8493 = 12'h92d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5421; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11565 = 12'h92d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8493; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14637 = 12'h92d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11565; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17709 = 12'h92d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14637; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20781 = 12'h92d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17709; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23853 = 12'h92d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20781; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26925 = 12'h92d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23853; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2349 = io_valid_in ? _GEN_26925 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2349 = 12'h92d == _T_2[11:0] ? image_2349 : _GEN_2348; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5422 = 12'h92e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8494 = 12'h92e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5422; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11566 = 12'h92e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8494; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14638 = 12'h92e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11566; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17710 = 12'h92e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14638; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20782 = 12'h92e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17710; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23854 = 12'h92e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20782; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26926 = 12'h92e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23854; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2350 = io_valid_in ? _GEN_26926 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2350 = 12'h92e == _T_2[11:0] ? image_2350 : _GEN_2349; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5423 = 12'h92f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8495 = 12'h92f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5423; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11567 = 12'h92f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8495; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14639 = 12'h92f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11567; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17711 = 12'h92f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14639; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20783 = 12'h92f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17711; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23855 = 12'h92f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20783; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26927 = 12'h92f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23855; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2351 = io_valid_in ? _GEN_26927 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2351 = 12'h92f == _T_2[11:0] ? image_2351 : _GEN_2350; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5424 = 12'h930 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8496 = 12'h930 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5424; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11568 = 12'h930 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8496; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14640 = 12'h930 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11568; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17712 = 12'h930 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14640; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20784 = 12'h930 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17712; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23856 = 12'h930 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20784; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26928 = 12'h930 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23856; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2352 = io_valid_in ? _GEN_26928 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2352 = 12'h930 == _T_2[11:0] ? image_2352 : _GEN_2351; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5425 = 12'h931 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8497 = 12'h931 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5425; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11569 = 12'h931 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8497; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14641 = 12'h931 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11569; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17713 = 12'h931 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14641; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20785 = 12'h931 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17713; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23857 = 12'h931 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20785; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26929 = 12'h931 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23857; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2353 = io_valid_in ? _GEN_26929 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2353 = 12'h931 == _T_2[11:0] ? image_2353 : _GEN_2352; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5426 = 12'h932 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8498 = 12'h932 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5426; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11570 = 12'h932 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8498; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14642 = 12'h932 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11570; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17714 = 12'h932 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14642; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20786 = 12'h932 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17714; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23858 = 12'h932 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20786; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26930 = 12'h932 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23858; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2354 = io_valid_in ? _GEN_26930 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2354 = 12'h932 == _T_2[11:0] ? image_2354 : _GEN_2353; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5427 = 12'h933 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8499 = 12'h933 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5427; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11571 = 12'h933 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8499; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14643 = 12'h933 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11571; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17715 = 12'h933 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14643; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20787 = 12'h933 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17715; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23859 = 12'h933 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20787; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26931 = 12'h933 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23859; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2355 = io_valid_in ? _GEN_26931 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2355 = 12'h933 == _T_2[11:0] ? image_2355 : _GEN_2354; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5428 = 12'h934 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8500 = 12'h934 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5428; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11572 = 12'h934 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8500; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14644 = 12'h934 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11572; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17716 = 12'h934 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14644; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20788 = 12'h934 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17716; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23860 = 12'h934 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20788; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26932 = 12'h934 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23860; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2356 = io_valid_in ? _GEN_26932 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2356 = 12'h934 == _T_2[11:0] ? image_2356 : _GEN_2355; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5429 = 12'h935 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8501 = 12'h935 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5429; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11573 = 12'h935 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8501; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14645 = 12'h935 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11573; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17717 = 12'h935 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14645; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20789 = 12'h935 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17717; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23861 = 12'h935 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20789; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26933 = 12'h935 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23861; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2357 = io_valid_in ? _GEN_26933 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2357 = 12'h935 == _T_2[11:0] ? image_2357 : _GEN_2356; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5430 = 12'h936 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8502 = 12'h936 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5430; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11574 = 12'h936 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8502; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14646 = 12'h936 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11574; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17718 = 12'h936 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14646; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20790 = 12'h936 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17718; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23862 = 12'h936 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20790; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26934 = 12'h936 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23862; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2358 = io_valid_in ? _GEN_26934 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2358 = 12'h936 == _T_2[11:0] ? image_2358 : _GEN_2357; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5431 = 12'h937 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8503 = 12'h937 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5431; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11575 = 12'h937 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8503; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14647 = 12'h937 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11575; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17719 = 12'h937 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14647; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20791 = 12'h937 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17719; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23863 = 12'h937 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20791; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26935 = 12'h937 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23863; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2359 = io_valid_in ? _GEN_26935 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2359 = 12'h937 == _T_2[11:0] ? image_2359 : _GEN_2358; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5432 = 12'h938 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8504 = 12'h938 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5432; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11576 = 12'h938 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8504; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14648 = 12'h938 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11576; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17720 = 12'h938 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14648; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20792 = 12'h938 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17720; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23864 = 12'h938 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20792; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26936 = 12'h938 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23864; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2360 = io_valid_in ? _GEN_26936 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2360 = 12'h938 == _T_2[11:0] ? image_2360 : _GEN_2359; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5433 = 12'h939 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8505 = 12'h939 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5433; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11577 = 12'h939 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8505; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14649 = 12'h939 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11577; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17721 = 12'h939 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14649; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20793 = 12'h939 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17721; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23865 = 12'h939 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20793; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26937 = 12'h939 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23865; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2361 = io_valid_in ? _GEN_26937 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2361 = 12'h939 == _T_2[11:0] ? image_2361 : _GEN_2360; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5434 = 12'h93a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8506 = 12'h93a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5434; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11578 = 12'h93a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8506; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14650 = 12'h93a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11578; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17722 = 12'h93a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14650; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20794 = 12'h93a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17722; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23866 = 12'h93a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20794; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26938 = 12'h93a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23866; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2362 = io_valid_in ? _GEN_26938 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2362 = 12'h93a == _T_2[11:0] ? image_2362 : _GEN_2361; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5435 = 12'h93b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8507 = 12'h93b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5435; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11579 = 12'h93b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8507; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14651 = 12'h93b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11579; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17723 = 12'h93b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14651; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20795 = 12'h93b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17723; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23867 = 12'h93b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20795; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26939 = 12'h93b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23867; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2363 = io_valid_in ? _GEN_26939 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2363 = 12'h93b == _T_2[11:0] ? image_2363 : _GEN_2362; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5436 = 12'h93c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8508 = 12'h93c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5436; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11580 = 12'h93c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8508; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14652 = 12'h93c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11580; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17724 = 12'h93c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14652; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20796 = 12'h93c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17724; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23868 = 12'h93c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20796; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26940 = 12'h93c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23868; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2364 = io_valid_in ? _GEN_26940 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2364 = 12'h93c == _T_2[11:0] ? image_2364 : _GEN_2363; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5437 = 12'h93d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8509 = 12'h93d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5437; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11581 = 12'h93d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8509; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14653 = 12'h93d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11581; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17725 = 12'h93d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14653; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20797 = 12'h93d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17725; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23869 = 12'h93d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20797; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26941 = 12'h93d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23869; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2365 = io_valid_in ? _GEN_26941 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2365 = 12'h93d == _T_2[11:0] ? image_2365 : _GEN_2364; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5438 = 12'h93e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8510 = 12'h93e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5438; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11582 = 12'h93e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8510; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14654 = 12'h93e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11582; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17726 = 12'h93e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14654; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20798 = 12'h93e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17726; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23870 = 12'h93e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20798; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26942 = 12'h93e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23870; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2366 = io_valid_in ? _GEN_26942 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2366 = 12'h93e == _T_2[11:0] ? image_2366 : _GEN_2365; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5439 = 12'h93f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8511 = 12'h93f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5439; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11583 = 12'h93f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8511; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14655 = 12'h93f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11583; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17727 = 12'h93f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14655; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20799 = 12'h93f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17727; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23871 = 12'h93f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20799; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26943 = 12'h93f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23871; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2367 = io_valid_in ? _GEN_26943 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2367 = 12'h93f == _T_2[11:0] ? image_2367 : _GEN_2366; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5440 = 12'h940 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8512 = 12'h940 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5440; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11584 = 12'h940 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8512; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14656 = 12'h940 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11584; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17728 = 12'h940 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14656; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20800 = 12'h940 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17728; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23872 = 12'h940 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20800; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26944 = 12'h940 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23872; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2368 = io_valid_in ? _GEN_26944 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2368 = 12'h940 == _T_2[11:0] ? image_2368 : _GEN_2367; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5441 = 12'h941 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8513 = 12'h941 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5441; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11585 = 12'h941 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8513; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14657 = 12'h941 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11585; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17729 = 12'h941 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14657; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20801 = 12'h941 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17729; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23873 = 12'h941 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20801; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26945 = 12'h941 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23873; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2369 = io_valid_in ? _GEN_26945 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2369 = 12'h941 == _T_2[11:0] ? image_2369 : _GEN_2368; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5442 = 12'h942 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8514 = 12'h942 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5442; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11586 = 12'h942 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8514; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14658 = 12'h942 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11586; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17730 = 12'h942 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14658; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20802 = 12'h942 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17730; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23874 = 12'h942 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20802; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26946 = 12'h942 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23874; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2370 = io_valid_in ? _GEN_26946 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2370 = 12'h942 == _T_2[11:0] ? image_2370 : _GEN_2369; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5443 = 12'h943 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8515 = 12'h943 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5443; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11587 = 12'h943 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8515; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14659 = 12'h943 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11587; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17731 = 12'h943 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14659; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20803 = 12'h943 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17731; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23875 = 12'h943 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20803; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26947 = 12'h943 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23875; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2371 = io_valid_in ? _GEN_26947 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2371 = 12'h943 == _T_2[11:0] ? image_2371 : _GEN_2370; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5444 = 12'h944 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8516 = 12'h944 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5444; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11588 = 12'h944 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8516; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14660 = 12'h944 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11588; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17732 = 12'h944 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14660; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20804 = 12'h944 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17732; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23876 = 12'h944 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20804; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26948 = 12'h944 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23876; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2372 = io_valid_in ? _GEN_26948 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2372 = 12'h944 == _T_2[11:0] ? image_2372 : _GEN_2371; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5445 = 12'h945 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8517 = 12'h945 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5445; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11589 = 12'h945 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8517; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14661 = 12'h945 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11589; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17733 = 12'h945 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14661; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20805 = 12'h945 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17733; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23877 = 12'h945 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20805; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26949 = 12'h945 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23877; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2373 = io_valid_in ? _GEN_26949 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2373 = 12'h945 == _T_2[11:0] ? image_2373 : _GEN_2372; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5446 = 12'h946 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8518 = 12'h946 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5446; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11590 = 12'h946 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8518; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14662 = 12'h946 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11590; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17734 = 12'h946 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14662; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20806 = 12'h946 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17734; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23878 = 12'h946 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20806; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26950 = 12'h946 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23878; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2374 = io_valid_in ? _GEN_26950 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2374 = 12'h946 == _T_2[11:0] ? image_2374 : _GEN_2373; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5447 = 12'h947 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8519 = 12'h947 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5447; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11591 = 12'h947 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8519; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14663 = 12'h947 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11591; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17735 = 12'h947 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14663; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20807 = 12'h947 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17735; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23879 = 12'h947 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20807; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26951 = 12'h947 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23879; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2375 = io_valid_in ? _GEN_26951 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2375 = 12'h947 == _T_2[11:0] ? image_2375 : _GEN_2374; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5448 = 12'h948 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8520 = 12'h948 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5448; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11592 = 12'h948 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8520; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14664 = 12'h948 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11592; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17736 = 12'h948 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14664; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20808 = 12'h948 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17736; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23880 = 12'h948 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20808; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26952 = 12'h948 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23880; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2376 = io_valid_in ? _GEN_26952 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2376 = 12'h948 == _T_2[11:0] ? image_2376 : _GEN_2375; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5449 = 12'h949 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8521 = 12'h949 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5449; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11593 = 12'h949 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8521; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14665 = 12'h949 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11593; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17737 = 12'h949 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14665; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20809 = 12'h949 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17737; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23881 = 12'h949 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20809; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26953 = 12'h949 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23881; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2377 = io_valid_in ? _GEN_26953 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2377 = 12'h949 == _T_2[11:0] ? image_2377 : _GEN_2376; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5450 = 12'h94a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8522 = 12'h94a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5450; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11594 = 12'h94a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8522; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14666 = 12'h94a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11594; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17738 = 12'h94a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14666; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20810 = 12'h94a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17738; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23882 = 12'h94a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20810; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26954 = 12'h94a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23882; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2378 = io_valid_in ? _GEN_26954 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2378 = 12'h94a == _T_2[11:0] ? image_2378 : _GEN_2377; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5451 = 12'h94b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8523 = 12'h94b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5451; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11595 = 12'h94b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8523; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14667 = 12'h94b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11595; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17739 = 12'h94b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14667; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20811 = 12'h94b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17739; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23883 = 12'h94b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20811; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26955 = 12'h94b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23883; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2379 = io_valid_in ? _GEN_26955 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2379 = 12'h94b == _T_2[11:0] ? image_2379 : _GEN_2378; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5452 = 12'h94c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8524 = 12'h94c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5452; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11596 = 12'h94c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8524; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14668 = 12'h94c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11596; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17740 = 12'h94c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14668; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20812 = 12'h94c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17740; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23884 = 12'h94c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20812; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26956 = 12'h94c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23884; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2380 = io_valid_in ? _GEN_26956 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2380 = 12'h94c == _T_2[11:0] ? image_2380 : _GEN_2379; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5453 = 12'h94d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8525 = 12'h94d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5453; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11597 = 12'h94d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8525; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14669 = 12'h94d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11597; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17741 = 12'h94d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14669; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20813 = 12'h94d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17741; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23885 = 12'h94d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20813; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26957 = 12'h94d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23885; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2381 = io_valid_in ? _GEN_26957 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2381 = 12'h94d == _T_2[11:0] ? image_2381 : _GEN_2380; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5454 = 12'h94e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8526 = 12'h94e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5454; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11598 = 12'h94e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8526; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14670 = 12'h94e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11598; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17742 = 12'h94e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14670; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20814 = 12'h94e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17742; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23886 = 12'h94e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20814; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26958 = 12'h94e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23886; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2382 = io_valid_in ? _GEN_26958 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2382 = 12'h94e == _T_2[11:0] ? image_2382 : _GEN_2381; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5455 = 12'h94f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8527 = 12'h94f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5455; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11599 = 12'h94f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8527; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14671 = 12'h94f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11599; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17743 = 12'h94f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14671; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20815 = 12'h94f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17743; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23887 = 12'h94f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20815; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26959 = 12'h94f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23887; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2383 = io_valid_in ? _GEN_26959 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2383 = 12'h94f == _T_2[11:0] ? image_2383 : _GEN_2382; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5456 = 12'h950 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8528 = 12'h950 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5456; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11600 = 12'h950 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8528; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14672 = 12'h950 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11600; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17744 = 12'h950 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14672; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20816 = 12'h950 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17744; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23888 = 12'h950 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20816; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26960 = 12'h950 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23888; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2384 = io_valid_in ? _GEN_26960 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2384 = 12'h950 == _T_2[11:0] ? image_2384 : _GEN_2383; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5457 = 12'h951 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8529 = 12'h951 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5457; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11601 = 12'h951 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8529; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14673 = 12'h951 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11601; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17745 = 12'h951 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14673; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20817 = 12'h951 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17745; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23889 = 12'h951 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20817; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26961 = 12'h951 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23889; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2385 = io_valid_in ? _GEN_26961 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2385 = 12'h951 == _T_2[11:0] ? image_2385 : _GEN_2384; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5458 = 12'h952 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8530 = 12'h952 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5458; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11602 = 12'h952 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8530; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14674 = 12'h952 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11602; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17746 = 12'h952 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14674; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20818 = 12'h952 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17746; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23890 = 12'h952 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20818; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26962 = 12'h952 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23890; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2386 = io_valid_in ? _GEN_26962 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2386 = 12'h952 == _T_2[11:0] ? image_2386 : _GEN_2385; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5459 = 12'h953 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8531 = 12'h953 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5459; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11603 = 12'h953 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8531; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14675 = 12'h953 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11603; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17747 = 12'h953 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14675; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20819 = 12'h953 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17747; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23891 = 12'h953 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20819; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26963 = 12'h953 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23891; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2387 = io_valid_in ? _GEN_26963 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2387 = 12'h953 == _T_2[11:0] ? image_2387 : _GEN_2386; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5460 = 12'h954 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8532 = 12'h954 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5460; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11604 = 12'h954 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8532; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14676 = 12'h954 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11604; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17748 = 12'h954 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14676; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20820 = 12'h954 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17748; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23892 = 12'h954 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20820; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26964 = 12'h954 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23892; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2388 = io_valid_in ? _GEN_26964 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2388 = 12'h954 == _T_2[11:0] ? image_2388 : _GEN_2387; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5461 = 12'h955 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8533 = 12'h955 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5461; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11605 = 12'h955 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8533; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14677 = 12'h955 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11605; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17749 = 12'h955 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14677; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20821 = 12'h955 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17749; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23893 = 12'h955 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20821; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26965 = 12'h955 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23893; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2389 = io_valid_in ? _GEN_26965 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2389 = 12'h955 == _T_2[11:0] ? image_2389 : _GEN_2388; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5462 = 12'h956 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8534 = 12'h956 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5462; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11606 = 12'h956 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8534; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14678 = 12'h956 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11606; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17750 = 12'h956 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14678; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20822 = 12'h956 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17750; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23894 = 12'h956 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20822; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26966 = 12'h956 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23894; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2390 = io_valid_in ? _GEN_26966 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2390 = 12'h956 == _T_2[11:0] ? image_2390 : _GEN_2389; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5463 = 12'h957 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8535 = 12'h957 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5463; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11607 = 12'h957 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8535; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14679 = 12'h957 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11607; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17751 = 12'h957 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14679; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20823 = 12'h957 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17751; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23895 = 12'h957 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20823; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26967 = 12'h957 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23895; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2391 = io_valid_in ? _GEN_26967 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2391 = 12'h957 == _T_2[11:0] ? image_2391 : _GEN_2390; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5464 = 12'h958 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8536 = 12'h958 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5464; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11608 = 12'h958 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8536; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14680 = 12'h958 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11608; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17752 = 12'h958 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14680; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20824 = 12'h958 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17752; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23896 = 12'h958 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20824; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26968 = 12'h958 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23896; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2392 = io_valid_in ? _GEN_26968 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2392 = 12'h958 == _T_2[11:0] ? image_2392 : _GEN_2391; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5465 = 12'h959 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8537 = 12'h959 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5465; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11609 = 12'h959 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8537; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14681 = 12'h959 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11609; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17753 = 12'h959 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14681; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20825 = 12'h959 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17753; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23897 = 12'h959 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20825; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26969 = 12'h959 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23897; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2393 = io_valid_in ? _GEN_26969 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2393 = 12'h959 == _T_2[11:0] ? image_2393 : _GEN_2392; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5466 = 12'h95a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8538 = 12'h95a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5466; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11610 = 12'h95a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8538; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14682 = 12'h95a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11610; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17754 = 12'h95a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14682; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20826 = 12'h95a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17754; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23898 = 12'h95a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20826; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26970 = 12'h95a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23898; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2394 = io_valid_in ? _GEN_26970 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2394 = 12'h95a == _T_2[11:0] ? image_2394 : _GEN_2393; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5467 = 12'h95b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8539 = 12'h95b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5467; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11611 = 12'h95b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8539; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14683 = 12'h95b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11611; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17755 = 12'h95b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14683; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20827 = 12'h95b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17755; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23899 = 12'h95b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20827; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26971 = 12'h95b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23899; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2395 = io_valid_in ? _GEN_26971 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2395 = 12'h95b == _T_2[11:0] ? image_2395 : _GEN_2394; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5468 = 12'h95c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8540 = 12'h95c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5468; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11612 = 12'h95c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8540; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14684 = 12'h95c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11612; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17756 = 12'h95c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14684; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20828 = 12'h95c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17756; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23900 = 12'h95c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20828; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26972 = 12'h95c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23900; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2396 = io_valid_in ? _GEN_26972 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2396 = 12'h95c == _T_2[11:0] ? image_2396 : _GEN_2395; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5469 = 12'h95d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8541 = 12'h95d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5469; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11613 = 12'h95d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8541; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14685 = 12'h95d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11613; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17757 = 12'h95d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14685; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20829 = 12'h95d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17757; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23901 = 12'h95d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20829; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26973 = 12'h95d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23901; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2397 = io_valid_in ? _GEN_26973 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2397 = 12'h95d == _T_2[11:0] ? image_2397 : _GEN_2396; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5470 = 12'h95e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8542 = 12'h95e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5470; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11614 = 12'h95e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8542; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14686 = 12'h95e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11614; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17758 = 12'h95e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14686; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20830 = 12'h95e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17758; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23902 = 12'h95e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20830; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26974 = 12'h95e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23902; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2398 = io_valid_in ? _GEN_26974 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2398 = 12'h95e == _T_2[11:0] ? image_2398 : _GEN_2397; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5471 = 12'h95f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8543 = 12'h95f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5471; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11615 = 12'h95f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8543; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14687 = 12'h95f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11615; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17759 = 12'h95f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14687; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20831 = 12'h95f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17759; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23903 = 12'h95f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20831; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26975 = 12'h95f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23903; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2399 = io_valid_in ? _GEN_26975 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2399 = 12'h95f == _T_2[11:0] ? image_2399 : _GEN_2398; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5472 = 12'h960 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8544 = 12'h960 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5472; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11616 = 12'h960 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8544; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14688 = 12'h960 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11616; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17760 = 12'h960 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14688; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20832 = 12'h960 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17760; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23904 = 12'h960 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20832; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26976 = 12'h960 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23904; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2400 = io_valid_in ? _GEN_26976 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2400 = 12'h960 == _T_2[11:0] ? image_2400 : _GEN_2399; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5473 = 12'h961 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8545 = 12'h961 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5473; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11617 = 12'h961 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8545; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14689 = 12'h961 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11617; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17761 = 12'h961 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14689; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20833 = 12'h961 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17761; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23905 = 12'h961 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20833; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26977 = 12'h961 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23905; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2401 = io_valid_in ? _GEN_26977 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2401 = 12'h961 == _T_2[11:0] ? image_2401 : _GEN_2400; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5474 = 12'h962 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8546 = 12'h962 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5474; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11618 = 12'h962 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8546; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14690 = 12'h962 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11618; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17762 = 12'h962 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14690; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20834 = 12'h962 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17762; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23906 = 12'h962 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20834; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26978 = 12'h962 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23906; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2402 = io_valid_in ? _GEN_26978 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2402 = 12'h962 == _T_2[11:0] ? image_2402 : _GEN_2401; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5475 = 12'h963 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8547 = 12'h963 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5475; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11619 = 12'h963 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8547; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14691 = 12'h963 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11619; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17763 = 12'h963 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14691; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20835 = 12'h963 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17763; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23907 = 12'h963 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20835; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26979 = 12'h963 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23907; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2403 = io_valid_in ? _GEN_26979 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2403 = 12'h963 == _T_2[11:0] ? image_2403 : _GEN_2402; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5476 = 12'h964 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8548 = 12'h964 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5476; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11620 = 12'h964 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8548; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14692 = 12'h964 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11620; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17764 = 12'h964 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14692; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20836 = 12'h964 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17764; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23908 = 12'h964 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20836; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26980 = 12'h964 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23908; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2404 = io_valid_in ? _GEN_26980 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2404 = 12'h964 == _T_2[11:0] ? image_2404 : _GEN_2403; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5477 = 12'h965 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8549 = 12'h965 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5477; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11621 = 12'h965 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8549; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14693 = 12'h965 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11621; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17765 = 12'h965 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14693; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20837 = 12'h965 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17765; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23909 = 12'h965 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20837; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26981 = 12'h965 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23909; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2405 = io_valid_in ? _GEN_26981 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2405 = 12'h965 == _T_2[11:0] ? image_2405 : _GEN_2404; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5478 = 12'h966 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8550 = 12'h966 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5478; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11622 = 12'h966 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8550; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14694 = 12'h966 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11622; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17766 = 12'h966 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14694; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20838 = 12'h966 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17766; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23910 = 12'h966 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20838; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26982 = 12'h966 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23910; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2406 = io_valid_in ? _GEN_26982 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2406 = 12'h966 == _T_2[11:0] ? image_2406 : _GEN_2405; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5479 = 12'h967 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8551 = 12'h967 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5479; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11623 = 12'h967 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8551; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14695 = 12'h967 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11623; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17767 = 12'h967 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14695; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20839 = 12'h967 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17767; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23911 = 12'h967 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20839; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26983 = 12'h967 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23911; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2407 = io_valid_in ? _GEN_26983 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2407 = 12'h967 == _T_2[11:0] ? image_2407 : _GEN_2406; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5480 = 12'h968 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8552 = 12'h968 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5480; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11624 = 12'h968 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8552; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14696 = 12'h968 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11624; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17768 = 12'h968 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14696; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20840 = 12'h968 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17768; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23912 = 12'h968 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20840; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26984 = 12'h968 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23912; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2408 = io_valid_in ? _GEN_26984 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2408 = 12'h968 == _T_2[11:0] ? image_2408 : _GEN_2407; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5481 = 12'h969 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8553 = 12'h969 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5481; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11625 = 12'h969 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8553; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14697 = 12'h969 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11625; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17769 = 12'h969 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14697; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20841 = 12'h969 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17769; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23913 = 12'h969 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20841; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26985 = 12'h969 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23913; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2409 = io_valid_in ? _GEN_26985 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2409 = 12'h969 == _T_2[11:0] ? image_2409 : _GEN_2408; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5482 = 12'h96a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8554 = 12'h96a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5482; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11626 = 12'h96a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8554; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14698 = 12'h96a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11626; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17770 = 12'h96a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14698; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20842 = 12'h96a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17770; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23914 = 12'h96a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20842; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26986 = 12'h96a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23914; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2410 = io_valid_in ? _GEN_26986 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2410 = 12'h96a == _T_2[11:0] ? image_2410 : _GEN_2409; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5483 = 12'h96b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8555 = 12'h96b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5483; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11627 = 12'h96b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8555; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14699 = 12'h96b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11627; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17771 = 12'h96b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14699; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20843 = 12'h96b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17771; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23915 = 12'h96b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20843; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26987 = 12'h96b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23915; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2411 = io_valid_in ? _GEN_26987 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2411 = 12'h96b == _T_2[11:0] ? image_2411 : _GEN_2410; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5484 = 12'h96c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8556 = 12'h96c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5484; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11628 = 12'h96c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8556; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14700 = 12'h96c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11628; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17772 = 12'h96c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14700; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20844 = 12'h96c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17772; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23916 = 12'h96c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20844; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26988 = 12'h96c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23916; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2412 = io_valid_in ? _GEN_26988 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2412 = 12'h96c == _T_2[11:0] ? image_2412 : _GEN_2411; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5485 = 12'h96d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8557 = 12'h96d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5485; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11629 = 12'h96d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8557; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14701 = 12'h96d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11629; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17773 = 12'h96d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14701; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20845 = 12'h96d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17773; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23917 = 12'h96d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20845; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26989 = 12'h96d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23917; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2413 = io_valid_in ? _GEN_26989 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2413 = 12'h96d == _T_2[11:0] ? image_2413 : _GEN_2412; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5486 = 12'h96e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8558 = 12'h96e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5486; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11630 = 12'h96e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8558; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14702 = 12'h96e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11630; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17774 = 12'h96e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14702; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20846 = 12'h96e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17774; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23918 = 12'h96e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20846; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26990 = 12'h96e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23918; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2414 = io_valid_in ? _GEN_26990 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2414 = 12'h96e == _T_2[11:0] ? image_2414 : _GEN_2413; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5487 = 12'h96f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8559 = 12'h96f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5487; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11631 = 12'h96f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8559; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14703 = 12'h96f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11631; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17775 = 12'h96f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14703; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20847 = 12'h96f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17775; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23919 = 12'h96f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20847; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26991 = 12'h96f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23919; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2415 = io_valid_in ? _GEN_26991 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2415 = 12'h96f == _T_2[11:0] ? image_2415 : _GEN_2414; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5488 = 12'h970 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8560 = 12'h970 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5488; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11632 = 12'h970 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8560; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14704 = 12'h970 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11632; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17776 = 12'h970 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14704; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20848 = 12'h970 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17776; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23920 = 12'h970 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20848; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26992 = 12'h970 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23920; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2416 = io_valid_in ? _GEN_26992 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2416 = 12'h970 == _T_2[11:0] ? image_2416 : _GEN_2415; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5489 = 12'h971 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8561 = 12'h971 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5489; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11633 = 12'h971 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8561; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14705 = 12'h971 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11633; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17777 = 12'h971 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14705; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20849 = 12'h971 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17777; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23921 = 12'h971 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20849; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26993 = 12'h971 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23921; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2417 = io_valid_in ? _GEN_26993 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2417 = 12'h971 == _T_2[11:0] ? image_2417 : _GEN_2416; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5490 = 12'h972 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8562 = 12'h972 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5490; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11634 = 12'h972 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8562; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14706 = 12'h972 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11634; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17778 = 12'h972 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14706; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20850 = 12'h972 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17778; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23922 = 12'h972 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20850; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26994 = 12'h972 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23922; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2418 = io_valid_in ? _GEN_26994 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2418 = 12'h972 == _T_2[11:0] ? image_2418 : _GEN_2417; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5491 = 12'h973 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8563 = 12'h973 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5491; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11635 = 12'h973 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8563; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14707 = 12'h973 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11635; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17779 = 12'h973 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14707; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20851 = 12'h973 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17779; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23923 = 12'h973 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20851; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26995 = 12'h973 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23923; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2419 = io_valid_in ? _GEN_26995 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2419 = 12'h973 == _T_2[11:0] ? image_2419 : _GEN_2418; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5492 = 12'h974 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8564 = 12'h974 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5492; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11636 = 12'h974 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8564; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14708 = 12'h974 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11636; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17780 = 12'h974 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14708; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20852 = 12'h974 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17780; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23924 = 12'h974 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20852; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26996 = 12'h974 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23924; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2420 = io_valid_in ? _GEN_26996 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2420 = 12'h974 == _T_2[11:0] ? image_2420 : _GEN_2419; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5493 = 12'h975 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8565 = 12'h975 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5493; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11637 = 12'h975 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8565; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14709 = 12'h975 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11637; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17781 = 12'h975 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14709; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20853 = 12'h975 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17781; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23925 = 12'h975 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20853; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26997 = 12'h975 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23925; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2421 = io_valid_in ? _GEN_26997 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2421 = 12'h975 == _T_2[11:0] ? image_2421 : _GEN_2420; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5494 = 12'h976 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8566 = 12'h976 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5494; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11638 = 12'h976 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8566; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14710 = 12'h976 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11638; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17782 = 12'h976 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14710; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20854 = 12'h976 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17782; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23926 = 12'h976 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20854; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26998 = 12'h976 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23926; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2422 = io_valid_in ? _GEN_26998 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2422 = 12'h976 == _T_2[11:0] ? image_2422 : _GEN_2421; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5495 = 12'h977 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8567 = 12'h977 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5495; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11639 = 12'h977 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8567; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14711 = 12'h977 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11639; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17783 = 12'h977 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14711; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20855 = 12'h977 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17783; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23927 = 12'h977 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20855; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_26999 = 12'h977 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23927; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2423 = io_valid_in ? _GEN_26999 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2423 = 12'h977 == _T_2[11:0] ? image_2423 : _GEN_2422; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5496 = 12'h978 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8568 = 12'h978 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5496; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11640 = 12'h978 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8568; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14712 = 12'h978 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11640; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17784 = 12'h978 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14712; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20856 = 12'h978 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17784; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23928 = 12'h978 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20856; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27000 = 12'h978 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23928; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2424 = io_valid_in ? _GEN_27000 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2424 = 12'h978 == _T_2[11:0] ? image_2424 : _GEN_2423; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5497 = 12'h979 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8569 = 12'h979 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5497; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11641 = 12'h979 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8569; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14713 = 12'h979 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11641; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17785 = 12'h979 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14713; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20857 = 12'h979 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17785; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23929 = 12'h979 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20857; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27001 = 12'h979 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23929; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2425 = io_valid_in ? _GEN_27001 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2425 = 12'h979 == _T_2[11:0] ? image_2425 : _GEN_2424; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5498 = 12'h97a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8570 = 12'h97a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5498; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11642 = 12'h97a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8570; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14714 = 12'h97a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11642; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17786 = 12'h97a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14714; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20858 = 12'h97a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17786; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23930 = 12'h97a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20858; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27002 = 12'h97a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23930; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2426 = io_valid_in ? _GEN_27002 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2426 = 12'h97a == _T_2[11:0] ? image_2426 : _GEN_2425; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5499 = 12'h97b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8571 = 12'h97b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5499; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11643 = 12'h97b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8571; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14715 = 12'h97b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11643; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17787 = 12'h97b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14715; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20859 = 12'h97b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17787; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23931 = 12'h97b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20859; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27003 = 12'h97b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23931; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2427 = io_valid_in ? _GEN_27003 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2427 = 12'h97b == _T_2[11:0] ? image_2427 : _GEN_2426; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5500 = 12'h97c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8572 = 12'h97c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5500; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11644 = 12'h97c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8572; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14716 = 12'h97c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11644; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17788 = 12'h97c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14716; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20860 = 12'h97c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17788; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23932 = 12'h97c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20860; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27004 = 12'h97c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23932; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2428 = io_valid_in ? _GEN_27004 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2428 = 12'h97c == _T_2[11:0] ? image_2428 : _GEN_2427; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5501 = 12'h97d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8573 = 12'h97d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5501; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11645 = 12'h97d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8573; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14717 = 12'h97d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11645; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17789 = 12'h97d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14717; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20861 = 12'h97d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17789; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23933 = 12'h97d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20861; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27005 = 12'h97d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23933; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2429 = io_valid_in ? _GEN_27005 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2429 = 12'h97d == _T_2[11:0] ? image_2429 : _GEN_2428; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5502 = 12'h97e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8574 = 12'h97e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5502; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11646 = 12'h97e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8574; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14718 = 12'h97e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11646; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17790 = 12'h97e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14718; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20862 = 12'h97e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17790; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23934 = 12'h97e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20862; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27006 = 12'h97e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23934; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2430 = io_valid_in ? _GEN_27006 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2430 = 12'h97e == _T_2[11:0] ? image_2430 : _GEN_2429; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5503 = 12'h97f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8575 = 12'h97f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5503; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11647 = 12'h97f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8575; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14719 = 12'h97f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11647; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17791 = 12'h97f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14719; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20863 = 12'h97f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17791; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23935 = 12'h97f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20863; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27007 = 12'h97f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23935; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2431 = io_valid_in ? _GEN_27007 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2431 = 12'h97f == _T_2[11:0] ? image_2431 : _GEN_2430; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5504 = 12'h980 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8576 = 12'h980 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5504; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11648 = 12'h980 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8576; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14720 = 12'h980 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11648; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17792 = 12'h980 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14720; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20864 = 12'h980 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17792; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23936 = 12'h980 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20864; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27008 = 12'h980 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23936; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2432 = io_valid_in ? _GEN_27008 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2432 = 12'h980 == _T_2[11:0] ? image_2432 : _GEN_2431; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5505 = 12'h981 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8577 = 12'h981 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5505; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11649 = 12'h981 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8577; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14721 = 12'h981 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11649; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17793 = 12'h981 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14721; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20865 = 12'h981 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17793; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23937 = 12'h981 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20865; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27009 = 12'h981 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23937; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2433 = io_valid_in ? _GEN_27009 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2433 = 12'h981 == _T_2[11:0] ? image_2433 : _GEN_2432; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5506 = 12'h982 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8578 = 12'h982 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5506; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11650 = 12'h982 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8578; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14722 = 12'h982 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11650; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17794 = 12'h982 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14722; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20866 = 12'h982 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17794; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23938 = 12'h982 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20866; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27010 = 12'h982 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23938; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2434 = io_valid_in ? _GEN_27010 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2434 = 12'h982 == _T_2[11:0] ? image_2434 : _GEN_2433; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5507 = 12'h983 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8579 = 12'h983 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5507; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11651 = 12'h983 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8579; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14723 = 12'h983 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11651; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17795 = 12'h983 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14723; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20867 = 12'h983 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17795; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23939 = 12'h983 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20867; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27011 = 12'h983 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23939; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2435 = io_valid_in ? _GEN_27011 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2435 = 12'h983 == _T_2[11:0] ? image_2435 : _GEN_2434; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5508 = 12'h984 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8580 = 12'h984 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5508; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11652 = 12'h984 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8580; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14724 = 12'h984 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11652; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17796 = 12'h984 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14724; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20868 = 12'h984 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17796; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23940 = 12'h984 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20868; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27012 = 12'h984 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23940; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2436 = io_valid_in ? _GEN_27012 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2436 = 12'h984 == _T_2[11:0] ? image_2436 : _GEN_2435; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5509 = 12'h985 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8581 = 12'h985 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5509; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11653 = 12'h985 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8581; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14725 = 12'h985 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11653; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17797 = 12'h985 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14725; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20869 = 12'h985 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17797; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23941 = 12'h985 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20869; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27013 = 12'h985 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23941; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2437 = io_valid_in ? _GEN_27013 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2437 = 12'h985 == _T_2[11:0] ? image_2437 : _GEN_2436; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5510 = 12'h986 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8582 = 12'h986 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5510; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11654 = 12'h986 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8582; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14726 = 12'h986 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11654; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17798 = 12'h986 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14726; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20870 = 12'h986 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17798; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23942 = 12'h986 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20870; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27014 = 12'h986 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23942; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2438 = io_valid_in ? _GEN_27014 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2438 = 12'h986 == _T_2[11:0] ? image_2438 : _GEN_2437; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5511 = 12'h987 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8583 = 12'h987 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5511; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11655 = 12'h987 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8583; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14727 = 12'h987 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11655; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17799 = 12'h987 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14727; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20871 = 12'h987 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17799; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23943 = 12'h987 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20871; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27015 = 12'h987 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23943; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2439 = io_valid_in ? _GEN_27015 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2439 = 12'h987 == _T_2[11:0] ? image_2439 : _GEN_2438; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5512 = 12'h988 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8584 = 12'h988 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5512; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11656 = 12'h988 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8584; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14728 = 12'h988 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11656; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17800 = 12'h988 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14728; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20872 = 12'h988 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17800; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23944 = 12'h988 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20872; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27016 = 12'h988 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23944; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2440 = io_valid_in ? _GEN_27016 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2440 = 12'h988 == _T_2[11:0] ? image_2440 : _GEN_2439; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5513 = 12'h989 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8585 = 12'h989 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5513; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11657 = 12'h989 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8585; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14729 = 12'h989 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11657; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17801 = 12'h989 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14729; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20873 = 12'h989 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17801; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23945 = 12'h989 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20873; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27017 = 12'h989 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23945; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2441 = io_valid_in ? _GEN_27017 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2441 = 12'h989 == _T_2[11:0] ? image_2441 : _GEN_2440; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5514 = 12'h98a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8586 = 12'h98a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5514; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11658 = 12'h98a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8586; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14730 = 12'h98a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11658; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17802 = 12'h98a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14730; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20874 = 12'h98a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17802; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23946 = 12'h98a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20874; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27018 = 12'h98a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23946; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2442 = io_valid_in ? _GEN_27018 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2442 = 12'h98a == _T_2[11:0] ? image_2442 : _GEN_2441; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5515 = 12'h98b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8587 = 12'h98b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5515; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11659 = 12'h98b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8587; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14731 = 12'h98b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11659; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17803 = 12'h98b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14731; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20875 = 12'h98b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17803; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23947 = 12'h98b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20875; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27019 = 12'h98b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23947; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2443 = io_valid_in ? _GEN_27019 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2443 = 12'h98b == _T_2[11:0] ? image_2443 : _GEN_2442; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5516 = 12'h98c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8588 = 12'h98c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5516; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11660 = 12'h98c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8588; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14732 = 12'h98c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11660; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17804 = 12'h98c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14732; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20876 = 12'h98c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17804; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23948 = 12'h98c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20876; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27020 = 12'h98c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23948; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2444 = io_valid_in ? _GEN_27020 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2444 = 12'h98c == _T_2[11:0] ? image_2444 : _GEN_2443; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5517 = 12'h98d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8589 = 12'h98d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5517; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11661 = 12'h98d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8589; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14733 = 12'h98d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11661; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17805 = 12'h98d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14733; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20877 = 12'h98d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17805; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23949 = 12'h98d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20877; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27021 = 12'h98d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23949; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2445 = io_valid_in ? _GEN_27021 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2445 = 12'h98d == _T_2[11:0] ? image_2445 : _GEN_2444; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5518 = 12'h98e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8590 = 12'h98e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5518; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11662 = 12'h98e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8590; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14734 = 12'h98e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11662; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17806 = 12'h98e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14734; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20878 = 12'h98e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17806; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23950 = 12'h98e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20878; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27022 = 12'h98e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23950; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2446 = io_valid_in ? _GEN_27022 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2446 = 12'h98e == _T_2[11:0] ? image_2446 : _GEN_2445; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5519 = 12'h98f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8591 = 12'h98f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5519; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11663 = 12'h98f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8591; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14735 = 12'h98f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11663; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17807 = 12'h98f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14735; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20879 = 12'h98f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17807; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23951 = 12'h98f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20879; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27023 = 12'h98f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23951; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2447 = io_valid_in ? _GEN_27023 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2447 = 12'h98f == _T_2[11:0] ? image_2447 : _GEN_2446; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5520 = 12'h990 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8592 = 12'h990 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5520; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11664 = 12'h990 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8592; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14736 = 12'h990 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11664; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17808 = 12'h990 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14736; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20880 = 12'h990 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17808; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23952 = 12'h990 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20880; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27024 = 12'h990 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23952; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2448 = io_valid_in ? _GEN_27024 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2448 = 12'h990 == _T_2[11:0] ? image_2448 : _GEN_2447; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5521 = 12'h991 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8593 = 12'h991 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5521; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11665 = 12'h991 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8593; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14737 = 12'h991 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11665; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17809 = 12'h991 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14737; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20881 = 12'h991 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17809; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23953 = 12'h991 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20881; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27025 = 12'h991 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23953; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2449 = io_valid_in ? _GEN_27025 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2449 = 12'h991 == _T_2[11:0] ? image_2449 : _GEN_2448; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5522 = 12'h992 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8594 = 12'h992 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5522; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11666 = 12'h992 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8594; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14738 = 12'h992 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11666; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17810 = 12'h992 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14738; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20882 = 12'h992 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17810; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23954 = 12'h992 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20882; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27026 = 12'h992 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23954; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2450 = io_valid_in ? _GEN_27026 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2450 = 12'h992 == _T_2[11:0] ? image_2450 : _GEN_2449; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5523 = 12'h993 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8595 = 12'h993 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5523; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11667 = 12'h993 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8595; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14739 = 12'h993 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11667; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17811 = 12'h993 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14739; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20883 = 12'h993 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17811; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23955 = 12'h993 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20883; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27027 = 12'h993 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23955; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2451 = io_valid_in ? _GEN_27027 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2451 = 12'h993 == _T_2[11:0] ? image_2451 : _GEN_2450; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5524 = 12'h994 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8596 = 12'h994 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5524; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11668 = 12'h994 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8596; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14740 = 12'h994 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11668; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17812 = 12'h994 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14740; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20884 = 12'h994 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17812; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23956 = 12'h994 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20884; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27028 = 12'h994 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23956; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2452 = io_valid_in ? _GEN_27028 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2452 = 12'h994 == _T_2[11:0] ? image_2452 : _GEN_2451; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5525 = 12'h995 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8597 = 12'h995 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5525; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11669 = 12'h995 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8597; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14741 = 12'h995 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11669; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17813 = 12'h995 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14741; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20885 = 12'h995 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17813; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23957 = 12'h995 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20885; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27029 = 12'h995 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23957; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2453 = io_valid_in ? _GEN_27029 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2453 = 12'h995 == _T_2[11:0] ? image_2453 : _GEN_2452; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5526 = 12'h996 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8598 = 12'h996 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5526; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11670 = 12'h996 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8598; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14742 = 12'h996 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11670; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17814 = 12'h996 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14742; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20886 = 12'h996 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17814; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23958 = 12'h996 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20886; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27030 = 12'h996 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23958; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2454 = io_valid_in ? _GEN_27030 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2454 = 12'h996 == _T_2[11:0] ? image_2454 : _GEN_2453; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5527 = 12'h997 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8599 = 12'h997 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5527; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11671 = 12'h997 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8599; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14743 = 12'h997 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11671; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17815 = 12'h997 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14743; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20887 = 12'h997 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17815; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23959 = 12'h997 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20887; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27031 = 12'h997 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23959; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2455 = io_valid_in ? _GEN_27031 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2455 = 12'h997 == _T_2[11:0] ? image_2455 : _GEN_2454; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5528 = 12'h998 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8600 = 12'h998 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5528; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11672 = 12'h998 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8600; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14744 = 12'h998 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11672; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17816 = 12'h998 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14744; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20888 = 12'h998 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17816; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23960 = 12'h998 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20888; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27032 = 12'h998 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23960; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2456 = io_valid_in ? _GEN_27032 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2456 = 12'h998 == _T_2[11:0] ? image_2456 : _GEN_2455; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5529 = 12'h999 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8601 = 12'h999 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5529; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11673 = 12'h999 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8601; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14745 = 12'h999 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11673; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17817 = 12'h999 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14745; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20889 = 12'h999 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17817; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23961 = 12'h999 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20889; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27033 = 12'h999 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23961; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2457 = io_valid_in ? _GEN_27033 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2457 = 12'h999 == _T_2[11:0] ? image_2457 : _GEN_2456; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5530 = 12'h99a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8602 = 12'h99a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5530; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11674 = 12'h99a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8602; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14746 = 12'h99a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11674; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17818 = 12'h99a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14746; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20890 = 12'h99a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17818; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23962 = 12'h99a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20890; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27034 = 12'h99a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23962; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2458 = io_valid_in ? _GEN_27034 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2458 = 12'h99a == _T_2[11:0] ? image_2458 : _GEN_2457; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5531 = 12'h99b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8603 = 12'h99b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5531; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11675 = 12'h99b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8603; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14747 = 12'h99b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11675; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17819 = 12'h99b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14747; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20891 = 12'h99b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17819; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23963 = 12'h99b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20891; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27035 = 12'h99b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23963; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2459 = io_valid_in ? _GEN_27035 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2459 = 12'h99b == _T_2[11:0] ? image_2459 : _GEN_2458; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5532 = 12'h99c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8604 = 12'h99c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5532; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11676 = 12'h99c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8604; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14748 = 12'h99c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11676; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17820 = 12'h99c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14748; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20892 = 12'h99c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17820; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23964 = 12'h99c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20892; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27036 = 12'h99c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23964; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2460 = io_valid_in ? _GEN_27036 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2460 = 12'h99c == _T_2[11:0] ? image_2460 : _GEN_2459; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5533 = 12'h99d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8605 = 12'h99d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5533; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11677 = 12'h99d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8605; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14749 = 12'h99d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11677; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17821 = 12'h99d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14749; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20893 = 12'h99d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17821; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23965 = 12'h99d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20893; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27037 = 12'h99d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23965; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2461 = io_valid_in ? _GEN_27037 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2461 = 12'h99d == _T_2[11:0] ? image_2461 : _GEN_2460; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5534 = 12'h99e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8606 = 12'h99e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5534; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11678 = 12'h99e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8606; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14750 = 12'h99e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11678; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17822 = 12'h99e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14750; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20894 = 12'h99e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17822; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23966 = 12'h99e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20894; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27038 = 12'h99e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23966; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2462 = io_valid_in ? _GEN_27038 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2462 = 12'h99e == _T_2[11:0] ? image_2462 : _GEN_2461; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5535 = 12'h99f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8607 = 12'h99f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5535; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11679 = 12'h99f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8607; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14751 = 12'h99f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11679; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17823 = 12'h99f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14751; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20895 = 12'h99f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17823; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23967 = 12'h99f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20895; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27039 = 12'h99f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23967; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2463 = io_valid_in ? _GEN_27039 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2463 = 12'h99f == _T_2[11:0] ? image_2463 : _GEN_2462; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5536 = 12'h9a0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8608 = 12'h9a0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5536; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11680 = 12'h9a0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8608; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14752 = 12'h9a0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11680; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17824 = 12'h9a0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14752; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20896 = 12'h9a0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17824; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23968 = 12'h9a0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20896; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27040 = 12'h9a0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23968; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2464 = io_valid_in ? _GEN_27040 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2464 = 12'h9a0 == _T_2[11:0] ? image_2464 : _GEN_2463; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5537 = 12'h9a1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8609 = 12'h9a1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5537; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11681 = 12'h9a1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8609; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14753 = 12'h9a1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11681; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17825 = 12'h9a1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14753; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20897 = 12'h9a1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17825; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23969 = 12'h9a1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20897; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27041 = 12'h9a1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23969; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2465 = io_valid_in ? _GEN_27041 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2465 = 12'h9a1 == _T_2[11:0] ? image_2465 : _GEN_2464; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5538 = 12'h9a2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8610 = 12'h9a2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5538; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11682 = 12'h9a2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8610; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14754 = 12'h9a2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11682; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17826 = 12'h9a2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14754; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20898 = 12'h9a2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17826; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23970 = 12'h9a2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20898; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27042 = 12'h9a2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23970; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2466 = io_valid_in ? _GEN_27042 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2466 = 12'h9a2 == _T_2[11:0] ? image_2466 : _GEN_2465; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5539 = 12'h9a3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8611 = 12'h9a3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5539; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11683 = 12'h9a3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8611; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14755 = 12'h9a3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11683; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17827 = 12'h9a3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14755; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20899 = 12'h9a3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17827; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23971 = 12'h9a3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20899; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27043 = 12'h9a3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23971; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2467 = io_valid_in ? _GEN_27043 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2467 = 12'h9a3 == _T_2[11:0] ? image_2467 : _GEN_2466; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5540 = 12'h9a4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8612 = 12'h9a4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5540; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11684 = 12'h9a4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8612; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14756 = 12'h9a4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11684; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17828 = 12'h9a4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14756; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20900 = 12'h9a4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17828; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23972 = 12'h9a4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20900; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27044 = 12'h9a4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23972; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2468 = io_valid_in ? _GEN_27044 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2468 = 12'h9a4 == _T_2[11:0] ? image_2468 : _GEN_2467; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5541 = 12'h9a5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8613 = 12'h9a5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5541; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11685 = 12'h9a5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8613; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14757 = 12'h9a5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11685; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17829 = 12'h9a5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14757; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20901 = 12'h9a5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17829; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23973 = 12'h9a5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20901; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27045 = 12'h9a5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23973; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2469 = io_valid_in ? _GEN_27045 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2469 = 12'h9a5 == _T_2[11:0] ? image_2469 : _GEN_2468; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5542 = 12'h9a6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8614 = 12'h9a6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5542; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11686 = 12'h9a6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8614; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14758 = 12'h9a6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11686; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17830 = 12'h9a6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14758; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20902 = 12'h9a6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17830; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23974 = 12'h9a6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20902; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27046 = 12'h9a6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23974; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2470 = io_valid_in ? _GEN_27046 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2470 = 12'h9a6 == _T_2[11:0] ? image_2470 : _GEN_2469; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5543 = 12'h9a7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8615 = 12'h9a7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5543; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11687 = 12'h9a7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8615; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14759 = 12'h9a7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11687; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17831 = 12'h9a7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14759; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20903 = 12'h9a7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17831; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23975 = 12'h9a7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20903; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27047 = 12'h9a7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23975; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2471 = io_valid_in ? _GEN_27047 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2471 = 12'h9a7 == _T_2[11:0] ? image_2471 : _GEN_2470; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5544 = 12'h9a8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8616 = 12'h9a8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5544; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11688 = 12'h9a8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8616; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14760 = 12'h9a8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11688; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17832 = 12'h9a8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14760; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20904 = 12'h9a8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17832; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23976 = 12'h9a8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20904; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27048 = 12'h9a8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23976; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2472 = io_valid_in ? _GEN_27048 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2472 = 12'h9a8 == _T_2[11:0] ? image_2472 : _GEN_2471; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5545 = 12'h9a9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8617 = 12'h9a9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5545; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11689 = 12'h9a9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8617; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14761 = 12'h9a9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11689; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17833 = 12'h9a9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14761; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20905 = 12'h9a9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17833; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23977 = 12'h9a9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20905; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27049 = 12'h9a9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23977; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2473 = io_valid_in ? _GEN_27049 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2473 = 12'h9a9 == _T_2[11:0] ? image_2473 : _GEN_2472; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5546 = 12'h9aa == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8618 = 12'h9aa == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5546; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11690 = 12'h9aa == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8618; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14762 = 12'h9aa == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11690; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17834 = 12'h9aa == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14762; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20906 = 12'h9aa == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17834; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23978 = 12'h9aa == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20906; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27050 = 12'h9aa == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23978; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2474 = io_valid_in ? _GEN_27050 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2474 = 12'h9aa == _T_2[11:0] ? image_2474 : _GEN_2473; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5547 = 12'h9ab == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8619 = 12'h9ab == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5547; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11691 = 12'h9ab == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8619; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14763 = 12'h9ab == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11691; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17835 = 12'h9ab == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14763; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20907 = 12'h9ab == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17835; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23979 = 12'h9ab == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20907; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27051 = 12'h9ab == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23979; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2475 = io_valid_in ? _GEN_27051 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2475 = 12'h9ab == _T_2[11:0] ? image_2475 : _GEN_2474; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5548 = 12'h9ac == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8620 = 12'h9ac == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5548; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11692 = 12'h9ac == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8620; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14764 = 12'h9ac == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11692; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17836 = 12'h9ac == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14764; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20908 = 12'h9ac == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17836; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23980 = 12'h9ac == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20908; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27052 = 12'h9ac == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23980; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2476 = io_valid_in ? _GEN_27052 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2476 = 12'h9ac == _T_2[11:0] ? image_2476 : _GEN_2475; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5549 = 12'h9ad == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8621 = 12'h9ad == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5549; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11693 = 12'h9ad == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8621; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14765 = 12'h9ad == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11693; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17837 = 12'h9ad == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14765; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20909 = 12'h9ad == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17837; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23981 = 12'h9ad == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20909; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27053 = 12'h9ad == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23981; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2477 = io_valid_in ? _GEN_27053 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2477 = 12'h9ad == _T_2[11:0] ? image_2477 : _GEN_2476; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5550 = 12'h9ae == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8622 = 12'h9ae == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5550; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11694 = 12'h9ae == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8622; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14766 = 12'h9ae == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11694; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17838 = 12'h9ae == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14766; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20910 = 12'h9ae == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17838; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23982 = 12'h9ae == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20910; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27054 = 12'h9ae == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23982; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2478 = io_valid_in ? _GEN_27054 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2478 = 12'h9ae == _T_2[11:0] ? image_2478 : _GEN_2477; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5551 = 12'h9af == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8623 = 12'h9af == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5551; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11695 = 12'h9af == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8623; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14767 = 12'h9af == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11695; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17839 = 12'h9af == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14767; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20911 = 12'h9af == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17839; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23983 = 12'h9af == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20911; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27055 = 12'h9af == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23983; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2479 = io_valid_in ? _GEN_27055 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2479 = 12'h9af == _T_2[11:0] ? image_2479 : _GEN_2478; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5552 = 12'h9b0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8624 = 12'h9b0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5552; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11696 = 12'h9b0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8624; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14768 = 12'h9b0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11696; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17840 = 12'h9b0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14768; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20912 = 12'h9b0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17840; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23984 = 12'h9b0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20912; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27056 = 12'h9b0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23984; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2480 = io_valid_in ? _GEN_27056 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2480 = 12'h9b0 == _T_2[11:0] ? image_2480 : _GEN_2479; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5553 = 12'h9b1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8625 = 12'h9b1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5553; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11697 = 12'h9b1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8625; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14769 = 12'h9b1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11697; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17841 = 12'h9b1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14769; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20913 = 12'h9b1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17841; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23985 = 12'h9b1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20913; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27057 = 12'h9b1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23985; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2481 = io_valid_in ? _GEN_27057 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2481 = 12'h9b1 == _T_2[11:0] ? image_2481 : _GEN_2480; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5554 = 12'h9b2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8626 = 12'h9b2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5554; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11698 = 12'h9b2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8626; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14770 = 12'h9b2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11698; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17842 = 12'h9b2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14770; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20914 = 12'h9b2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17842; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23986 = 12'h9b2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20914; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27058 = 12'h9b2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23986; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2482 = io_valid_in ? _GEN_27058 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2482 = 12'h9b2 == _T_2[11:0] ? image_2482 : _GEN_2481; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5555 = 12'h9b3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8627 = 12'h9b3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5555; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11699 = 12'h9b3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8627; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14771 = 12'h9b3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11699; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17843 = 12'h9b3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14771; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20915 = 12'h9b3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17843; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23987 = 12'h9b3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20915; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27059 = 12'h9b3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23987; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2483 = io_valid_in ? _GEN_27059 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2483 = 12'h9b3 == _T_2[11:0] ? image_2483 : _GEN_2482; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5556 = 12'h9b4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8628 = 12'h9b4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5556; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11700 = 12'h9b4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8628; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14772 = 12'h9b4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11700; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17844 = 12'h9b4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14772; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20916 = 12'h9b4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17844; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23988 = 12'h9b4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20916; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27060 = 12'h9b4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23988; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2484 = io_valid_in ? _GEN_27060 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2484 = 12'h9b4 == _T_2[11:0] ? image_2484 : _GEN_2483; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5557 = 12'h9b5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8629 = 12'h9b5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5557; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11701 = 12'h9b5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8629; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14773 = 12'h9b5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11701; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17845 = 12'h9b5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14773; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20917 = 12'h9b5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17845; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23989 = 12'h9b5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20917; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27061 = 12'h9b5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23989; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2485 = io_valid_in ? _GEN_27061 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2485 = 12'h9b5 == _T_2[11:0] ? image_2485 : _GEN_2484; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5558 = 12'h9b6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8630 = 12'h9b6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5558; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11702 = 12'h9b6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8630; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14774 = 12'h9b6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11702; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17846 = 12'h9b6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14774; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20918 = 12'h9b6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17846; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23990 = 12'h9b6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20918; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27062 = 12'h9b6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23990; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2486 = io_valid_in ? _GEN_27062 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2486 = 12'h9b6 == _T_2[11:0] ? image_2486 : _GEN_2485; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5559 = 12'h9b7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8631 = 12'h9b7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5559; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11703 = 12'h9b7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8631; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14775 = 12'h9b7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11703; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17847 = 12'h9b7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14775; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20919 = 12'h9b7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17847; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23991 = 12'h9b7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20919; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27063 = 12'h9b7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23991; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2487 = io_valid_in ? _GEN_27063 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2487 = 12'h9b7 == _T_2[11:0] ? image_2487 : _GEN_2486; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5560 = 12'h9b8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8632 = 12'h9b8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5560; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11704 = 12'h9b8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8632; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14776 = 12'h9b8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11704; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17848 = 12'h9b8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14776; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20920 = 12'h9b8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17848; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23992 = 12'h9b8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20920; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27064 = 12'h9b8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23992; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2488 = io_valid_in ? _GEN_27064 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2488 = 12'h9b8 == _T_2[11:0] ? image_2488 : _GEN_2487; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5561 = 12'h9b9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8633 = 12'h9b9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5561; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11705 = 12'h9b9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8633; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14777 = 12'h9b9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11705; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17849 = 12'h9b9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14777; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20921 = 12'h9b9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17849; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23993 = 12'h9b9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20921; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27065 = 12'h9b9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23993; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2489 = io_valid_in ? _GEN_27065 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2489 = 12'h9b9 == _T_2[11:0] ? image_2489 : _GEN_2488; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5562 = 12'h9ba == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8634 = 12'h9ba == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5562; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11706 = 12'h9ba == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8634; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14778 = 12'h9ba == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11706; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17850 = 12'h9ba == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14778; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20922 = 12'h9ba == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17850; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23994 = 12'h9ba == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20922; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27066 = 12'h9ba == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23994; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2490 = io_valid_in ? _GEN_27066 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2490 = 12'h9ba == _T_2[11:0] ? image_2490 : _GEN_2489; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5563 = 12'h9bb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8635 = 12'h9bb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5563; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11707 = 12'h9bb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8635; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14779 = 12'h9bb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11707; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17851 = 12'h9bb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14779; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20923 = 12'h9bb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17851; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23995 = 12'h9bb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20923; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27067 = 12'h9bb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23995; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2491 = io_valid_in ? _GEN_27067 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2491 = 12'h9bb == _T_2[11:0] ? image_2491 : _GEN_2490; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5564 = 12'h9bc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8636 = 12'h9bc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5564; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11708 = 12'h9bc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8636; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14780 = 12'h9bc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11708; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17852 = 12'h9bc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14780; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20924 = 12'h9bc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17852; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23996 = 12'h9bc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20924; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27068 = 12'h9bc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23996; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2492 = io_valid_in ? _GEN_27068 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2492 = 12'h9bc == _T_2[11:0] ? image_2492 : _GEN_2491; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5565 = 12'h9bd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8637 = 12'h9bd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5565; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11709 = 12'h9bd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8637; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14781 = 12'h9bd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11709; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17853 = 12'h9bd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14781; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20925 = 12'h9bd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17853; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23997 = 12'h9bd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20925; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27069 = 12'h9bd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23997; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2493 = io_valid_in ? _GEN_27069 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2493 = 12'h9bd == _T_2[11:0] ? image_2493 : _GEN_2492; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5566 = 12'h9be == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8638 = 12'h9be == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5566; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11710 = 12'h9be == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8638; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14782 = 12'h9be == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11710; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17854 = 12'h9be == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14782; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20926 = 12'h9be == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17854; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23998 = 12'h9be == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20926; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27070 = 12'h9be == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23998; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2494 = io_valid_in ? _GEN_27070 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2494 = 12'h9be == _T_2[11:0] ? image_2494 : _GEN_2493; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5567 = 12'h9bf == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8639 = 12'h9bf == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5567; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11711 = 12'h9bf == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8639; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14783 = 12'h9bf == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11711; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17855 = 12'h9bf == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14783; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20927 = 12'h9bf == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17855; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_23999 = 12'h9bf == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20927; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27071 = 12'h9bf == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_23999; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2495 = io_valid_in ? _GEN_27071 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2495 = 12'h9bf == _T_2[11:0] ? image_2495 : _GEN_2494; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5568 = 12'h9c0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8640 = 12'h9c0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5568; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11712 = 12'h9c0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8640; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14784 = 12'h9c0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11712; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17856 = 12'h9c0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14784; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20928 = 12'h9c0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17856; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24000 = 12'h9c0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20928; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27072 = 12'h9c0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24000; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2496 = io_valid_in ? _GEN_27072 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2496 = 12'h9c0 == _T_2[11:0] ? image_2496 : _GEN_2495; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5569 = 12'h9c1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8641 = 12'h9c1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5569; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11713 = 12'h9c1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8641; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14785 = 12'h9c1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11713; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17857 = 12'h9c1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14785; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20929 = 12'h9c1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17857; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24001 = 12'h9c1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20929; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27073 = 12'h9c1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24001; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2497 = io_valid_in ? _GEN_27073 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2497 = 12'h9c1 == _T_2[11:0] ? image_2497 : _GEN_2496; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5570 = 12'h9c2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8642 = 12'h9c2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5570; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11714 = 12'h9c2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8642; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14786 = 12'h9c2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11714; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17858 = 12'h9c2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14786; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20930 = 12'h9c2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17858; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24002 = 12'h9c2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20930; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27074 = 12'h9c2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24002; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2498 = io_valid_in ? _GEN_27074 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2498 = 12'h9c2 == _T_2[11:0] ? image_2498 : _GEN_2497; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5571 = 12'h9c3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8643 = 12'h9c3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5571; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11715 = 12'h9c3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8643; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14787 = 12'h9c3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11715; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17859 = 12'h9c3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14787; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20931 = 12'h9c3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17859; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24003 = 12'h9c3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20931; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27075 = 12'h9c3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24003; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2499 = io_valid_in ? _GEN_27075 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2499 = 12'h9c3 == _T_2[11:0] ? image_2499 : _GEN_2498; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5572 = 12'h9c4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8644 = 12'h9c4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5572; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11716 = 12'h9c4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8644; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14788 = 12'h9c4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11716; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17860 = 12'h9c4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14788; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20932 = 12'h9c4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17860; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24004 = 12'h9c4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20932; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27076 = 12'h9c4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24004; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2500 = io_valid_in ? _GEN_27076 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2500 = 12'h9c4 == _T_2[11:0] ? image_2500 : _GEN_2499; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5573 = 12'h9c5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8645 = 12'h9c5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5573; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11717 = 12'h9c5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8645; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14789 = 12'h9c5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11717; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17861 = 12'h9c5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14789; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20933 = 12'h9c5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17861; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24005 = 12'h9c5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20933; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27077 = 12'h9c5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24005; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2501 = io_valid_in ? _GEN_27077 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2501 = 12'h9c5 == _T_2[11:0] ? image_2501 : _GEN_2500; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5574 = 12'h9c6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8646 = 12'h9c6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5574; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11718 = 12'h9c6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8646; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14790 = 12'h9c6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11718; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17862 = 12'h9c6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14790; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20934 = 12'h9c6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17862; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24006 = 12'h9c6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20934; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27078 = 12'h9c6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24006; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2502 = io_valid_in ? _GEN_27078 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2502 = 12'h9c6 == _T_2[11:0] ? image_2502 : _GEN_2501; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5575 = 12'h9c7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8647 = 12'h9c7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5575; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11719 = 12'h9c7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8647; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14791 = 12'h9c7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11719; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17863 = 12'h9c7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14791; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20935 = 12'h9c7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17863; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24007 = 12'h9c7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20935; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27079 = 12'h9c7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24007; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2503 = io_valid_in ? _GEN_27079 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2503 = 12'h9c7 == _T_2[11:0] ? image_2503 : _GEN_2502; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5576 = 12'h9c8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8648 = 12'h9c8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5576; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11720 = 12'h9c8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8648; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14792 = 12'h9c8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11720; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17864 = 12'h9c8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14792; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20936 = 12'h9c8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17864; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24008 = 12'h9c8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20936; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27080 = 12'h9c8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24008; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2504 = io_valid_in ? _GEN_27080 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2504 = 12'h9c8 == _T_2[11:0] ? image_2504 : _GEN_2503; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5577 = 12'h9c9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8649 = 12'h9c9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5577; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11721 = 12'h9c9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8649; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14793 = 12'h9c9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11721; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17865 = 12'h9c9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14793; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20937 = 12'h9c9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17865; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24009 = 12'h9c9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20937; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27081 = 12'h9c9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24009; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2505 = io_valid_in ? _GEN_27081 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2505 = 12'h9c9 == _T_2[11:0] ? image_2505 : _GEN_2504; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5578 = 12'h9ca == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8650 = 12'h9ca == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5578; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11722 = 12'h9ca == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8650; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14794 = 12'h9ca == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11722; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17866 = 12'h9ca == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14794; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20938 = 12'h9ca == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17866; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24010 = 12'h9ca == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20938; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27082 = 12'h9ca == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24010; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2506 = io_valid_in ? _GEN_27082 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2506 = 12'h9ca == _T_2[11:0] ? image_2506 : _GEN_2505; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5579 = 12'h9cb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8651 = 12'h9cb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5579; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11723 = 12'h9cb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8651; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14795 = 12'h9cb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11723; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17867 = 12'h9cb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14795; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20939 = 12'h9cb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17867; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24011 = 12'h9cb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20939; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27083 = 12'h9cb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24011; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2507 = io_valid_in ? _GEN_27083 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2507 = 12'h9cb == _T_2[11:0] ? image_2507 : _GEN_2506; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5580 = 12'h9cc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8652 = 12'h9cc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5580; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11724 = 12'h9cc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8652; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14796 = 12'h9cc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11724; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17868 = 12'h9cc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14796; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20940 = 12'h9cc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17868; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24012 = 12'h9cc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20940; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27084 = 12'h9cc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24012; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2508 = io_valid_in ? _GEN_27084 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2508 = 12'h9cc == _T_2[11:0] ? image_2508 : _GEN_2507; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5581 = 12'h9cd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8653 = 12'h9cd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5581; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11725 = 12'h9cd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8653; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14797 = 12'h9cd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11725; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17869 = 12'h9cd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14797; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20941 = 12'h9cd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17869; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24013 = 12'h9cd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20941; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27085 = 12'h9cd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24013; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2509 = io_valid_in ? _GEN_27085 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2509 = 12'h9cd == _T_2[11:0] ? image_2509 : _GEN_2508; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5582 = 12'h9ce == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8654 = 12'h9ce == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5582; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11726 = 12'h9ce == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8654; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14798 = 12'h9ce == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11726; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17870 = 12'h9ce == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14798; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20942 = 12'h9ce == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17870; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24014 = 12'h9ce == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20942; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27086 = 12'h9ce == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24014; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2510 = io_valid_in ? _GEN_27086 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2510 = 12'h9ce == _T_2[11:0] ? image_2510 : _GEN_2509; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5583 = 12'h9cf == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8655 = 12'h9cf == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5583; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11727 = 12'h9cf == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8655; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14799 = 12'h9cf == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11727; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17871 = 12'h9cf == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14799; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20943 = 12'h9cf == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17871; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24015 = 12'h9cf == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20943; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27087 = 12'h9cf == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24015; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2511 = io_valid_in ? _GEN_27087 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2511 = 12'h9cf == _T_2[11:0] ? image_2511 : _GEN_2510; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5584 = 12'h9d0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8656 = 12'h9d0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5584; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11728 = 12'h9d0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8656; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14800 = 12'h9d0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11728; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17872 = 12'h9d0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14800; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20944 = 12'h9d0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17872; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24016 = 12'h9d0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20944; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27088 = 12'h9d0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24016; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2512 = io_valid_in ? _GEN_27088 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2512 = 12'h9d0 == _T_2[11:0] ? image_2512 : _GEN_2511; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5585 = 12'h9d1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8657 = 12'h9d1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5585; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11729 = 12'h9d1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8657; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14801 = 12'h9d1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11729; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17873 = 12'h9d1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14801; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20945 = 12'h9d1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17873; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24017 = 12'h9d1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20945; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27089 = 12'h9d1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24017; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2513 = io_valid_in ? _GEN_27089 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2513 = 12'h9d1 == _T_2[11:0] ? image_2513 : _GEN_2512; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5586 = 12'h9d2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8658 = 12'h9d2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5586; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11730 = 12'h9d2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8658; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14802 = 12'h9d2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11730; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17874 = 12'h9d2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14802; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20946 = 12'h9d2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17874; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24018 = 12'h9d2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20946; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27090 = 12'h9d2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24018; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2514 = io_valid_in ? _GEN_27090 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2514 = 12'h9d2 == _T_2[11:0] ? image_2514 : _GEN_2513; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5587 = 12'h9d3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8659 = 12'h9d3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5587; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11731 = 12'h9d3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8659; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14803 = 12'h9d3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11731; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17875 = 12'h9d3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14803; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20947 = 12'h9d3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17875; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24019 = 12'h9d3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20947; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27091 = 12'h9d3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24019; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2515 = io_valid_in ? _GEN_27091 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2515 = 12'h9d3 == _T_2[11:0] ? image_2515 : _GEN_2514; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5588 = 12'h9d4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8660 = 12'h9d4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5588; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11732 = 12'h9d4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8660; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14804 = 12'h9d4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11732; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17876 = 12'h9d4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14804; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20948 = 12'h9d4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17876; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24020 = 12'h9d4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20948; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27092 = 12'h9d4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24020; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2516 = io_valid_in ? _GEN_27092 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2516 = 12'h9d4 == _T_2[11:0] ? image_2516 : _GEN_2515; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5589 = 12'h9d5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8661 = 12'h9d5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5589; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11733 = 12'h9d5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8661; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14805 = 12'h9d5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11733; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17877 = 12'h9d5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14805; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20949 = 12'h9d5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17877; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24021 = 12'h9d5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20949; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27093 = 12'h9d5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24021; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2517 = io_valid_in ? _GEN_27093 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2517 = 12'h9d5 == _T_2[11:0] ? image_2517 : _GEN_2516; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5590 = 12'h9d6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8662 = 12'h9d6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5590; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11734 = 12'h9d6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8662; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14806 = 12'h9d6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11734; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17878 = 12'h9d6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14806; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20950 = 12'h9d6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17878; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24022 = 12'h9d6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20950; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27094 = 12'h9d6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24022; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2518 = io_valid_in ? _GEN_27094 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2518 = 12'h9d6 == _T_2[11:0] ? image_2518 : _GEN_2517; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5591 = 12'h9d7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8663 = 12'h9d7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5591; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11735 = 12'h9d7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8663; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14807 = 12'h9d7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11735; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17879 = 12'h9d7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14807; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20951 = 12'h9d7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17879; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24023 = 12'h9d7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20951; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27095 = 12'h9d7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24023; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2519 = io_valid_in ? _GEN_27095 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2519 = 12'h9d7 == _T_2[11:0] ? image_2519 : _GEN_2518; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5592 = 12'h9d8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8664 = 12'h9d8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5592; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11736 = 12'h9d8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8664; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14808 = 12'h9d8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11736; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17880 = 12'h9d8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14808; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20952 = 12'h9d8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17880; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24024 = 12'h9d8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20952; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27096 = 12'h9d8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24024; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2520 = io_valid_in ? _GEN_27096 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2520 = 12'h9d8 == _T_2[11:0] ? image_2520 : _GEN_2519; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5593 = 12'h9d9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8665 = 12'h9d9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5593; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11737 = 12'h9d9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8665; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14809 = 12'h9d9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11737; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17881 = 12'h9d9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14809; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20953 = 12'h9d9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17881; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24025 = 12'h9d9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20953; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27097 = 12'h9d9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24025; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2521 = io_valid_in ? _GEN_27097 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2521 = 12'h9d9 == _T_2[11:0] ? image_2521 : _GEN_2520; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5594 = 12'h9da == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8666 = 12'h9da == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5594; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11738 = 12'h9da == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8666; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14810 = 12'h9da == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11738; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17882 = 12'h9da == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14810; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20954 = 12'h9da == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17882; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24026 = 12'h9da == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20954; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27098 = 12'h9da == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24026; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2522 = io_valid_in ? _GEN_27098 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2522 = 12'h9da == _T_2[11:0] ? image_2522 : _GEN_2521; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5595 = 12'h9db == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8667 = 12'h9db == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5595; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11739 = 12'h9db == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8667; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14811 = 12'h9db == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11739; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17883 = 12'h9db == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14811; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20955 = 12'h9db == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17883; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24027 = 12'h9db == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20955; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27099 = 12'h9db == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24027; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2523 = io_valid_in ? _GEN_27099 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2523 = 12'h9db == _T_2[11:0] ? image_2523 : _GEN_2522; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5596 = 12'h9dc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8668 = 12'h9dc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5596; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11740 = 12'h9dc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8668; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14812 = 12'h9dc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11740; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17884 = 12'h9dc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14812; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20956 = 12'h9dc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17884; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24028 = 12'h9dc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20956; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27100 = 12'h9dc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24028; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2524 = io_valid_in ? _GEN_27100 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2524 = 12'h9dc == _T_2[11:0] ? image_2524 : _GEN_2523; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5597 = 12'h9dd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8669 = 12'h9dd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5597; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11741 = 12'h9dd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8669; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14813 = 12'h9dd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11741; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17885 = 12'h9dd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14813; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20957 = 12'h9dd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17885; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24029 = 12'h9dd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20957; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27101 = 12'h9dd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24029; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2525 = io_valid_in ? _GEN_27101 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2525 = 12'h9dd == _T_2[11:0] ? image_2525 : _GEN_2524; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5598 = 12'h9de == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8670 = 12'h9de == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5598; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11742 = 12'h9de == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8670; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14814 = 12'h9de == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11742; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17886 = 12'h9de == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14814; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20958 = 12'h9de == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17886; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24030 = 12'h9de == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20958; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27102 = 12'h9de == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24030; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2526 = io_valid_in ? _GEN_27102 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2526 = 12'h9de == _T_2[11:0] ? image_2526 : _GEN_2525; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5599 = 12'h9df == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8671 = 12'h9df == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5599; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11743 = 12'h9df == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8671; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14815 = 12'h9df == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11743; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17887 = 12'h9df == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14815; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20959 = 12'h9df == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17887; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24031 = 12'h9df == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20959; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27103 = 12'h9df == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24031; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2527 = io_valid_in ? _GEN_27103 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2527 = 12'h9df == _T_2[11:0] ? image_2527 : _GEN_2526; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5600 = 12'h9e0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8672 = 12'h9e0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5600; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11744 = 12'h9e0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8672; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14816 = 12'h9e0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11744; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17888 = 12'h9e0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14816; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20960 = 12'h9e0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17888; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24032 = 12'h9e0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20960; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27104 = 12'h9e0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24032; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2528 = io_valid_in ? _GEN_27104 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2528 = 12'h9e0 == _T_2[11:0] ? image_2528 : _GEN_2527; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5601 = 12'h9e1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8673 = 12'h9e1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5601; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11745 = 12'h9e1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8673; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14817 = 12'h9e1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11745; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17889 = 12'h9e1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14817; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20961 = 12'h9e1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17889; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24033 = 12'h9e1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20961; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27105 = 12'h9e1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24033; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2529 = io_valid_in ? _GEN_27105 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2529 = 12'h9e1 == _T_2[11:0] ? image_2529 : _GEN_2528; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5602 = 12'h9e2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8674 = 12'h9e2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5602; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11746 = 12'h9e2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8674; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14818 = 12'h9e2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11746; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17890 = 12'h9e2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14818; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20962 = 12'h9e2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17890; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24034 = 12'h9e2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20962; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27106 = 12'h9e2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24034; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2530 = io_valid_in ? _GEN_27106 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2530 = 12'h9e2 == _T_2[11:0] ? image_2530 : _GEN_2529; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5603 = 12'h9e3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8675 = 12'h9e3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5603; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11747 = 12'h9e3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8675; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14819 = 12'h9e3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11747; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17891 = 12'h9e3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14819; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20963 = 12'h9e3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17891; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24035 = 12'h9e3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20963; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27107 = 12'h9e3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24035; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2531 = io_valid_in ? _GEN_27107 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2531 = 12'h9e3 == _T_2[11:0] ? image_2531 : _GEN_2530; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5604 = 12'h9e4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8676 = 12'h9e4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5604; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11748 = 12'h9e4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8676; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14820 = 12'h9e4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11748; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17892 = 12'h9e4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14820; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20964 = 12'h9e4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17892; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24036 = 12'h9e4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20964; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27108 = 12'h9e4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24036; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2532 = io_valid_in ? _GEN_27108 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2532 = 12'h9e4 == _T_2[11:0] ? image_2532 : _GEN_2531; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5605 = 12'h9e5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8677 = 12'h9e5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5605; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11749 = 12'h9e5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8677; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14821 = 12'h9e5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11749; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17893 = 12'h9e5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14821; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20965 = 12'h9e5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17893; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24037 = 12'h9e5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20965; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27109 = 12'h9e5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24037; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2533 = io_valid_in ? _GEN_27109 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2533 = 12'h9e5 == _T_2[11:0] ? image_2533 : _GEN_2532; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5606 = 12'h9e6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8678 = 12'h9e6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5606; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11750 = 12'h9e6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8678; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14822 = 12'h9e6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11750; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17894 = 12'h9e6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14822; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20966 = 12'h9e6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17894; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24038 = 12'h9e6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20966; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27110 = 12'h9e6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24038; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2534 = io_valid_in ? _GEN_27110 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2534 = 12'h9e6 == _T_2[11:0] ? image_2534 : _GEN_2533; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5607 = 12'h9e7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8679 = 12'h9e7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5607; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11751 = 12'h9e7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8679; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14823 = 12'h9e7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11751; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17895 = 12'h9e7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14823; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20967 = 12'h9e7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17895; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24039 = 12'h9e7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20967; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27111 = 12'h9e7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24039; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2535 = io_valid_in ? _GEN_27111 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2535 = 12'h9e7 == _T_2[11:0] ? image_2535 : _GEN_2534; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5608 = 12'h9e8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8680 = 12'h9e8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5608; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11752 = 12'h9e8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8680; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14824 = 12'h9e8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11752; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17896 = 12'h9e8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14824; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20968 = 12'h9e8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17896; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24040 = 12'h9e8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20968; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27112 = 12'h9e8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24040; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2536 = io_valid_in ? _GEN_27112 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2536 = 12'h9e8 == _T_2[11:0] ? image_2536 : _GEN_2535; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5609 = 12'h9e9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8681 = 12'h9e9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5609; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11753 = 12'h9e9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8681; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14825 = 12'h9e9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11753; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17897 = 12'h9e9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14825; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20969 = 12'h9e9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17897; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24041 = 12'h9e9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20969; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27113 = 12'h9e9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24041; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2537 = io_valid_in ? _GEN_27113 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2537 = 12'h9e9 == _T_2[11:0] ? image_2537 : _GEN_2536; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5610 = 12'h9ea == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8682 = 12'h9ea == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5610; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11754 = 12'h9ea == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8682; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14826 = 12'h9ea == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11754; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17898 = 12'h9ea == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14826; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20970 = 12'h9ea == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17898; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24042 = 12'h9ea == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20970; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27114 = 12'h9ea == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24042; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2538 = io_valid_in ? _GEN_27114 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2538 = 12'h9ea == _T_2[11:0] ? image_2538 : _GEN_2537; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5611 = 12'h9eb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8683 = 12'h9eb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5611; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11755 = 12'h9eb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8683; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14827 = 12'h9eb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11755; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17899 = 12'h9eb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14827; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20971 = 12'h9eb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17899; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24043 = 12'h9eb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20971; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27115 = 12'h9eb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24043; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2539 = io_valid_in ? _GEN_27115 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2539 = 12'h9eb == _T_2[11:0] ? image_2539 : _GEN_2538; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5612 = 12'h9ec == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8684 = 12'h9ec == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5612; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11756 = 12'h9ec == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8684; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14828 = 12'h9ec == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11756; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17900 = 12'h9ec == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14828; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20972 = 12'h9ec == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17900; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24044 = 12'h9ec == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20972; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27116 = 12'h9ec == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24044; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2540 = io_valid_in ? _GEN_27116 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2540 = 12'h9ec == _T_2[11:0] ? image_2540 : _GEN_2539; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5613 = 12'h9ed == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8685 = 12'h9ed == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5613; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11757 = 12'h9ed == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8685; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14829 = 12'h9ed == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11757; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17901 = 12'h9ed == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14829; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20973 = 12'h9ed == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17901; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24045 = 12'h9ed == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20973; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27117 = 12'h9ed == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24045; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2541 = io_valid_in ? _GEN_27117 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2541 = 12'h9ed == _T_2[11:0] ? image_2541 : _GEN_2540; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5614 = 12'h9ee == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8686 = 12'h9ee == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5614; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11758 = 12'h9ee == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8686; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14830 = 12'h9ee == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11758; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17902 = 12'h9ee == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14830; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20974 = 12'h9ee == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17902; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24046 = 12'h9ee == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20974; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27118 = 12'h9ee == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24046; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2542 = io_valid_in ? _GEN_27118 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2542 = 12'h9ee == _T_2[11:0] ? image_2542 : _GEN_2541; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5615 = 12'h9ef == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8687 = 12'h9ef == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5615; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11759 = 12'h9ef == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8687; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14831 = 12'h9ef == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11759; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17903 = 12'h9ef == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14831; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20975 = 12'h9ef == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17903; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24047 = 12'h9ef == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20975; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27119 = 12'h9ef == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24047; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2543 = io_valid_in ? _GEN_27119 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2543 = 12'h9ef == _T_2[11:0] ? image_2543 : _GEN_2542; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5616 = 12'h9f0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8688 = 12'h9f0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5616; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11760 = 12'h9f0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8688; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14832 = 12'h9f0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11760; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17904 = 12'h9f0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14832; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20976 = 12'h9f0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17904; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24048 = 12'h9f0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20976; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27120 = 12'h9f0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24048; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2544 = io_valid_in ? _GEN_27120 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2544 = 12'h9f0 == _T_2[11:0] ? image_2544 : _GEN_2543; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5617 = 12'h9f1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8689 = 12'h9f1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5617; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11761 = 12'h9f1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8689; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14833 = 12'h9f1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11761; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17905 = 12'h9f1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14833; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20977 = 12'h9f1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17905; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24049 = 12'h9f1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20977; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27121 = 12'h9f1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24049; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2545 = io_valid_in ? _GEN_27121 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2545 = 12'h9f1 == _T_2[11:0] ? image_2545 : _GEN_2544; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5618 = 12'h9f2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8690 = 12'h9f2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5618; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11762 = 12'h9f2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8690; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14834 = 12'h9f2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11762; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17906 = 12'h9f2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14834; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20978 = 12'h9f2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17906; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24050 = 12'h9f2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20978; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27122 = 12'h9f2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24050; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2546 = io_valid_in ? _GEN_27122 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2546 = 12'h9f2 == _T_2[11:0] ? image_2546 : _GEN_2545; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5619 = 12'h9f3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8691 = 12'h9f3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5619; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11763 = 12'h9f3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8691; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14835 = 12'h9f3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11763; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17907 = 12'h9f3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14835; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20979 = 12'h9f3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17907; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24051 = 12'h9f3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20979; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27123 = 12'h9f3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24051; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2547 = io_valid_in ? _GEN_27123 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2547 = 12'h9f3 == _T_2[11:0] ? image_2547 : _GEN_2546; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5620 = 12'h9f4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8692 = 12'h9f4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5620; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11764 = 12'h9f4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8692; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14836 = 12'h9f4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11764; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17908 = 12'h9f4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14836; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20980 = 12'h9f4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17908; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24052 = 12'h9f4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20980; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27124 = 12'h9f4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24052; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2548 = io_valid_in ? _GEN_27124 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2548 = 12'h9f4 == _T_2[11:0] ? image_2548 : _GEN_2547; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5621 = 12'h9f5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8693 = 12'h9f5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5621; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11765 = 12'h9f5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8693; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14837 = 12'h9f5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11765; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17909 = 12'h9f5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14837; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20981 = 12'h9f5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17909; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24053 = 12'h9f5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20981; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27125 = 12'h9f5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24053; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2549 = io_valid_in ? _GEN_27125 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2549 = 12'h9f5 == _T_2[11:0] ? image_2549 : _GEN_2548; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5622 = 12'h9f6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8694 = 12'h9f6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5622; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11766 = 12'h9f6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8694; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14838 = 12'h9f6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11766; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17910 = 12'h9f6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14838; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20982 = 12'h9f6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17910; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24054 = 12'h9f6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20982; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27126 = 12'h9f6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24054; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2550 = io_valid_in ? _GEN_27126 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2550 = 12'h9f6 == _T_2[11:0] ? image_2550 : _GEN_2549; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5623 = 12'h9f7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8695 = 12'h9f7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5623; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11767 = 12'h9f7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8695; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14839 = 12'h9f7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11767; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17911 = 12'h9f7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14839; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20983 = 12'h9f7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17911; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24055 = 12'h9f7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20983; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27127 = 12'h9f7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24055; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2551 = io_valid_in ? _GEN_27127 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2551 = 12'h9f7 == _T_2[11:0] ? image_2551 : _GEN_2550; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5624 = 12'h9f8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8696 = 12'h9f8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5624; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11768 = 12'h9f8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8696; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14840 = 12'h9f8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11768; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17912 = 12'h9f8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14840; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20984 = 12'h9f8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17912; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24056 = 12'h9f8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20984; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27128 = 12'h9f8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24056; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2552 = io_valid_in ? _GEN_27128 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2552 = 12'h9f8 == _T_2[11:0] ? image_2552 : _GEN_2551; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5625 = 12'h9f9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8697 = 12'h9f9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5625; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11769 = 12'h9f9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8697; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14841 = 12'h9f9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11769; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17913 = 12'h9f9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14841; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20985 = 12'h9f9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17913; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24057 = 12'h9f9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20985; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27129 = 12'h9f9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24057; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2553 = io_valid_in ? _GEN_27129 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2553 = 12'h9f9 == _T_2[11:0] ? image_2553 : _GEN_2552; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5626 = 12'h9fa == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8698 = 12'h9fa == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5626; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11770 = 12'h9fa == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8698; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14842 = 12'h9fa == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11770; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17914 = 12'h9fa == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14842; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20986 = 12'h9fa == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17914; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24058 = 12'h9fa == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20986; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27130 = 12'h9fa == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24058; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2554 = io_valid_in ? _GEN_27130 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2554 = 12'h9fa == _T_2[11:0] ? image_2554 : _GEN_2553; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5627 = 12'h9fb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8699 = 12'h9fb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5627; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11771 = 12'h9fb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8699; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14843 = 12'h9fb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11771; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17915 = 12'h9fb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14843; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20987 = 12'h9fb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17915; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24059 = 12'h9fb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20987; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27131 = 12'h9fb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24059; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2555 = io_valid_in ? _GEN_27131 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2555 = 12'h9fb == _T_2[11:0] ? image_2555 : _GEN_2554; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5628 = 12'h9fc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8700 = 12'h9fc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5628; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11772 = 12'h9fc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8700; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14844 = 12'h9fc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11772; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17916 = 12'h9fc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14844; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20988 = 12'h9fc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17916; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24060 = 12'h9fc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20988; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27132 = 12'h9fc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24060; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2556 = io_valid_in ? _GEN_27132 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2556 = 12'h9fc == _T_2[11:0] ? image_2556 : _GEN_2555; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5629 = 12'h9fd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8701 = 12'h9fd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5629; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11773 = 12'h9fd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8701; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14845 = 12'h9fd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11773; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17917 = 12'h9fd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14845; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20989 = 12'h9fd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17917; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24061 = 12'h9fd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20989; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27133 = 12'h9fd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24061; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2557 = io_valid_in ? _GEN_27133 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2557 = 12'h9fd == _T_2[11:0] ? image_2557 : _GEN_2556; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5630 = 12'h9fe == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8702 = 12'h9fe == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5630; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11774 = 12'h9fe == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8702; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14846 = 12'h9fe == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11774; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17918 = 12'h9fe == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14846; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20990 = 12'h9fe == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17918; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24062 = 12'h9fe == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20990; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27134 = 12'h9fe == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24062; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2558 = io_valid_in ? _GEN_27134 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2558 = 12'h9fe == _T_2[11:0] ? image_2558 : _GEN_2557; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5631 = 12'h9ff == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8703 = 12'h9ff == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5631; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11775 = 12'h9ff == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8703; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14847 = 12'h9ff == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11775; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17919 = 12'h9ff == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14847; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20991 = 12'h9ff == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17919; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24063 = 12'h9ff == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20991; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27135 = 12'h9ff == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24063; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2559 = io_valid_in ? _GEN_27135 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2559 = 12'h9ff == _T_2[11:0] ? image_2559 : _GEN_2558; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5632 = 12'ha00 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8704 = 12'ha00 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5632; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11776 = 12'ha00 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8704; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14848 = 12'ha00 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11776; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17920 = 12'ha00 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14848; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20992 = 12'ha00 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17920; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24064 = 12'ha00 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20992; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27136 = 12'ha00 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24064; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2560 = io_valid_in ? _GEN_27136 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2560 = 12'ha00 == _T_2[11:0] ? image_2560 : _GEN_2559; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5633 = 12'ha01 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8705 = 12'ha01 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5633; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11777 = 12'ha01 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8705; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14849 = 12'ha01 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11777; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17921 = 12'ha01 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14849; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20993 = 12'ha01 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17921; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24065 = 12'ha01 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20993; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27137 = 12'ha01 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24065; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2561 = io_valid_in ? _GEN_27137 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2561 = 12'ha01 == _T_2[11:0] ? image_2561 : _GEN_2560; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5634 = 12'ha02 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8706 = 12'ha02 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5634; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11778 = 12'ha02 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8706; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14850 = 12'ha02 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11778; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17922 = 12'ha02 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14850; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20994 = 12'ha02 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17922; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24066 = 12'ha02 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20994; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27138 = 12'ha02 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24066; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2562 = io_valid_in ? _GEN_27138 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2562 = 12'ha02 == _T_2[11:0] ? image_2562 : _GEN_2561; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5635 = 12'ha03 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8707 = 12'ha03 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5635; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11779 = 12'ha03 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8707; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14851 = 12'ha03 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11779; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17923 = 12'ha03 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14851; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20995 = 12'ha03 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17923; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24067 = 12'ha03 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20995; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27139 = 12'ha03 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24067; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2563 = io_valid_in ? _GEN_27139 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2563 = 12'ha03 == _T_2[11:0] ? image_2563 : _GEN_2562; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5636 = 12'ha04 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8708 = 12'ha04 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5636; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11780 = 12'ha04 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8708; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14852 = 12'ha04 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11780; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17924 = 12'ha04 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14852; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20996 = 12'ha04 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17924; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24068 = 12'ha04 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20996; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27140 = 12'ha04 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24068; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2564 = io_valid_in ? _GEN_27140 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2564 = 12'ha04 == _T_2[11:0] ? image_2564 : _GEN_2563; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5637 = 12'ha05 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8709 = 12'ha05 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5637; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11781 = 12'ha05 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8709; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14853 = 12'ha05 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11781; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17925 = 12'ha05 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14853; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20997 = 12'ha05 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17925; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24069 = 12'ha05 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20997; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27141 = 12'ha05 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24069; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2565 = io_valid_in ? _GEN_27141 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2565 = 12'ha05 == _T_2[11:0] ? image_2565 : _GEN_2564; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5638 = 12'ha06 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8710 = 12'ha06 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5638; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11782 = 12'ha06 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8710; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14854 = 12'ha06 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11782; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17926 = 12'ha06 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14854; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20998 = 12'ha06 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17926; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24070 = 12'ha06 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20998; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27142 = 12'ha06 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24070; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2566 = io_valid_in ? _GEN_27142 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2566 = 12'ha06 == _T_2[11:0] ? image_2566 : _GEN_2565; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5639 = 12'ha07 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8711 = 12'ha07 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5639; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11783 = 12'ha07 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8711; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14855 = 12'ha07 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11783; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17927 = 12'ha07 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14855; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_20999 = 12'ha07 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17927; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24071 = 12'ha07 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_20999; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27143 = 12'ha07 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24071; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2567 = io_valid_in ? _GEN_27143 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2567 = 12'ha07 == _T_2[11:0] ? image_2567 : _GEN_2566; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5640 = 12'ha08 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8712 = 12'ha08 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5640; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11784 = 12'ha08 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8712; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14856 = 12'ha08 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11784; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17928 = 12'ha08 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14856; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21000 = 12'ha08 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17928; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24072 = 12'ha08 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21000; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27144 = 12'ha08 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24072; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2568 = io_valid_in ? _GEN_27144 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2568 = 12'ha08 == _T_2[11:0] ? image_2568 : _GEN_2567; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5641 = 12'ha09 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8713 = 12'ha09 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5641; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11785 = 12'ha09 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8713; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14857 = 12'ha09 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11785; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17929 = 12'ha09 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14857; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21001 = 12'ha09 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17929; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24073 = 12'ha09 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21001; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27145 = 12'ha09 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24073; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2569 = io_valid_in ? _GEN_27145 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2569 = 12'ha09 == _T_2[11:0] ? image_2569 : _GEN_2568; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5642 = 12'ha0a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8714 = 12'ha0a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5642; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11786 = 12'ha0a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8714; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14858 = 12'ha0a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11786; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17930 = 12'ha0a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14858; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21002 = 12'ha0a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17930; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24074 = 12'ha0a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21002; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27146 = 12'ha0a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24074; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2570 = io_valid_in ? _GEN_27146 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2570 = 12'ha0a == _T_2[11:0] ? image_2570 : _GEN_2569; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5643 = 12'ha0b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8715 = 12'ha0b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5643; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11787 = 12'ha0b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8715; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14859 = 12'ha0b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11787; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17931 = 12'ha0b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14859; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21003 = 12'ha0b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17931; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24075 = 12'ha0b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21003; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27147 = 12'ha0b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24075; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2571 = io_valid_in ? _GEN_27147 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2571 = 12'ha0b == _T_2[11:0] ? image_2571 : _GEN_2570; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5644 = 12'ha0c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8716 = 12'ha0c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5644; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11788 = 12'ha0c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8716; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14860 = 12'ha0c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11788; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17932 = 12'ha0c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14860; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21004 = 12'ha0c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17932; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24076 = 12'ha0c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21004; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27148 = 12'ha0c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24076; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2572 = io_valid_in ? _GEN_27148 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2572 = 12'ha0c == _T_2[11:0] ? image_2572 : _GEN_2571; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5645 = 12'ha0d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8717 = 12'ha0d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5645; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11789 = 12'ha0d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8717; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14861 = 12'ha0d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11789; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17933 = 12'ha0d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14861; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21005 = 12'ha0d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17933; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24077 = 12'ha0d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21005; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27149 = 12'ha0d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24077; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2573 = io_valid_in ? _GEN_27149 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2573 = 12'ha0d == _T_2[11:0] ? image_2573 : _GEN_2572; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5646 = 12'ha0e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8718 = 12'ha0e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5646; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11790 = 12'ha0e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8718; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14862 = 12'ha0e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11790; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17934 = 12'ha0e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14862; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21006 = 12'ha0e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17934; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24078 = 12'ha0e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21006; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27150 = 12'ha0e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24078; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2574 = io_valid_in ? _GEN_27150 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2574 = 12'ha0e == _T_2[11:0] ? image_2574 : _GEN_2573; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5647 = 12'ha0f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8719 = 12'ha0f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5647; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11791 = 12'ha0f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8719; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14863 = 12'ha0f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11791; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17935 = 12'ha0f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14863; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21007 = 12'ha0f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17935; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24079 = 12'ha0f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21007; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27151 = 12'ha0f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24079; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2575 = io_valid_in ? _GEN_27151 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2575 = 12'ha0f == _T_2[11:0] ? image_2575 : _GEN_2574; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5648 = 12'ha10 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8720 = 12'ha10 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5648; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11792 = 12'ha10 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8720; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14864 = 12'ha10 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11792; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17936 = 12'ha10 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14864; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21008 = 12'ha10 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17936; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24080 = 12'ha10 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21008; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27152 = 12'ha10 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24080; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2576 = io_valid_in ? _GEN_27152 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2576 = 12'ha10 == _T_2[11:0] ? image_2576 : _GEN_2575; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5649 = 12'ha11 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8721 = 12'ha11 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5649; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11793 = 12'ha11 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8721; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14865 = 12'ha11 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11793; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17937 = 12'ha11 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14865; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21009 = 12'ha11 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17937; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24081 = 12'ha11 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21009; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27153 = 12'ha11 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24081; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2577 = io_valid_in ? _GEN_27153 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2577 = 12'ha11 == _T_2[11:0] ? image_2577 : _GEN_2576; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5650 = 12'ha12 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8722 = 12'ha12 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5650; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11794 = 12'ha12 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8722; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14866 = 12'ha12 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11794; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17938 = 12'ha12 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14866; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21010 = 12'ha12 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17938; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24082 = 12'ha12 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21010; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27154 = 12'ha12 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24082; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2578 = io_valid_in ? _GEN_27154 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2578 = 12'ha12 == _T_2[11:0] ? image_2578 : _GEN_2577; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5651 = 12'ha13 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8723 = 12'ha13 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5651; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11795 = 12'ha13 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8723; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14867 = 12'ha13 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11795; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17939 = 12'ha13 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14867; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21011 = 12'ha13 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17939; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24083 = 12'ha13 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21011; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27155 = 12'ha13 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24083; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2579 = io_valid_in ? _GEN_27155 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2579 = 12'ha13 == _T_2[11:0] ? image_2579 : _GEN_2578; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5652 = 12'ha14 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8724 = 12'ha14 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5652; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11796 = 12'ha14 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8724; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14868 = 12'ha14 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11796; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17940 = 12'ha14 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14868; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21012 = 12'ha14 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17940; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24084 = 12'ha14 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21012; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27156 = 12'ha14 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24084; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2580 = io_valid_in ? _GEN_27156 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2580 = 12'ha14 == _T_2[11:0] ? image_2580 : _GEN_2579; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5653 = 12'ha15 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8725 = 12'ha15 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5653; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11797 = 12'ha15 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8725; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14869 = 12'ha15 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11797; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17941 = 12'ha15 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14869; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21013 = 12'ha15 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17941; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24085 = 12'ha15 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21013; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27157 = 12'ha15 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24085; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2581 = io_valid_in ? _GEN_27157 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2581 = 12'ha15 == _T_2[11:0] ? image_2581 : _GEN_2580; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5654 = 12'ha16 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8726 = 12'ha16 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5654; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11798 = 12'ha16 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8726; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14870 = 12'ha16 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11798; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17942 = 12'ha16 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14870; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21014 = 12'ha16 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17942; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24086 = 12'ha16 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21014; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27158 = 12'ha16 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24086; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2582 = io_valid_in ? _GEN_27158 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2582 = 12'ha16 == _T_2[11:0] ? image_2582 : _GEN_2581; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5655 = 12'ha17 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8727 = 12'ha17 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5655; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11799 = 12'ha17 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8727; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14871 = 12'ha17 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11799; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17943 = 12'ha17 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14871; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21015 = 12'ha17 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17943; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24087 = 12'ha17 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21015; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27159 = 12'ha17 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24087; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2583 = io_valid_in ? _GEN_27159 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2583 = 12'ha17 == _T_2[11:0] ? image_2583 : _GEN_2582; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5656 = 12'ha18 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8728 = 12'ha18 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5656; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11800 = 12'ha18 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8728; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14872 = 12'ha18 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11800; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17944 = 12'ha18 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14872; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21016 = 12'ha18 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17944; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24088 = 12'ha18 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21016; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27160 = 12'ha18 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24088; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2584 = io_valid_in ? _GEN_27160 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2584 = 12'ha18 == _T_2[11:0] ? image_2584 : _GEN_2583; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5657 = 12'ha19 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8729 = 12'ha19 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5657; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11801 = 12'ha19 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8729; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14873 = 12'ha19 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11801; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17945 = 12'ha19 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14873; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21017 = 12'ha19 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17945; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24089 = 12'ha19 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21017; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27161 = 12'ha19 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24089; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2585 = io_valid_in ? _GEN_27161 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2585 = 12'ha19 == _T_2[11:0] ? image_2585 : _GEN_2584; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5658 = 12'ha1a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8730 = 12'ha1a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5658; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11802 = 12'ha1a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8730; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14874 = 12'ha1a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11802; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17946 = 12'ha1a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14874; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21018 = 12'ha1a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17946; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24090 = 12'ha1a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21018; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27162 = 12'ha1a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24090; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2586 = io_valid_in ? _GEN_27162 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2586 = 12'ha1a == _T_2[11:0] ? image_2586 : _GEN_2585; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5659 = 12'ha1b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8731 = 12'ha1b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5659; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11803 = 12'ha1b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8731; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14875 = 12'ha1b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11803; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17947 = 12'ha1b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14875; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21019 = 12'ha1b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17947; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24091 = 12'ha1b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21019; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27163 = 12'ha1b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24091; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2587 = io_valid_in ? _GEN_27163 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2587 = 12'ha1b == _T_2[11:0] ? image_2587 : _GEN_2586; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5660 = 12'ha1c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8732 = 12'ha1c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5660; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11804 = 12'ha1c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8732; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14876 = 12'ha1c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11804; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17948 = 12'ha1c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14876; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21020 = 12'ha1c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17948; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24092 = 12'ha1c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21020; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27164 = 12'ha1c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24092; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2588 = io_valid_in ? _GEN_27164 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2588 = 12'ha1c == _T_2[11:0] ? image_2588 : _GEN_2587; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5661 = 12'ha1d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8733 = 12'ha1d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5661; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11805 = 12'ha1d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8733; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14877 = 12'ha1d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11805; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17949 = 12'ha1d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14877; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21021 = 12'ha1d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17949; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24093 = 12'ha1d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21021; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27165 = 12'ha1d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24093; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2589 = io_valid_in ? _GEN_27165 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2589 = 12'ha1d == _T_2[11:0] ? image_2589 : _GEN_2588; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5662 = 12'ha1e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8734 = 12'ha1e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5662; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11806 = 12'ha1e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8734; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14878 = 12'ha1e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11806; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17950 = 12'ha1e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14878; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21022 = 12'ha1e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17950; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24094 = 12'ha1e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21022; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27166 = 12'ha1e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24094; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2590 = io_valid_in ? _GEN_27166 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2590 = 12'ha1e == _T_2[11:0] ? image_2590 : _GEN_2589; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5663 = 12'ha1f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8735 = 12'ha1f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5663; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11807 = 12'ha1f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8735; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14879 = 12'ha1f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11807; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17951 = 12'ha1f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14879; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21023 = 12'ha1f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17951; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24095 = 12'ha1f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21023; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27167 = 12'ha1f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24095; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2591 = io_valid_in ? _GEN_27167 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2591 = 12'ha1f == _T_2[11:0] ? image_2591 : _GEN_2590; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5664 = 12'ha20 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8736 = 12'ha20 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5664; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11808 = 12'ha20 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8736; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14880 = 12'ha20 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11808; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17952 = 12'ha20 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14880; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21024 = 12'ha20 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17952; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24096 = 12'ha20 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21024; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27168 = 12'ha20 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24096; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2592 = io_valid_in ? _GEN_27168 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2592 = 12'ha20 == _T_2[11:0] ? image_2592 : _GEN_2591; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5665 = 12'ha21 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8737 = 12'ha21 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5665; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11809 = 12'ha21 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8737; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14881 = 12'ha21 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11809; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17953 = 12'ha21 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14881; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21025 = 12'ha21 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17953; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24097 = 12'ha21 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21025; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27169 = 12'ha21 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24097; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2593 = io_valid_in ? _GEN_27169 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2593 = 12'ha21 == _T_2[11:0] ? image_2593 : _GEN_2592; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5666 = 12'ha22 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8738 = 12'ha22 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5666; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11810 = 12'ha22 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8738; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14882 = 12'ha22 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11810; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17954 = 12'ha22 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14882; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21026 = 12'ha22 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17954; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24098 = 12'ha22 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21026; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27170 = 12'ha22 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24098; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2594 = io_valid_in ? _GEN_27170 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2594 = 12'ha22 == _T_2[11:0] ? image_2594 : _GEN_2593; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5667 = 12'ha23 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8739 = 12'ha23 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5667; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11811 = 12'ha23 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8739; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14883 = 12'ha23 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11811; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17955 = 12'ha23 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14883; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21027 = 12'ha23 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17955; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24099 = 12'ha23 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21027; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27171 = 12'ha23 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24099; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2595 = io_valid_in ? _GEN_27171 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2595 = 12'ha23 == _T_2[11:0] ? image_2595 : _GEN_2594; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5668 = 12'ha24 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8740 = 12'ha24 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5668; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11812 = 12'ha24 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8740; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14884 = 12'ha24 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11812; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17956 = 12'ha24 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14884; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21028 = 12'ha24 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17956; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24100 = 12'ha24 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21028; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27172 = 12'ha24 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24100; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2596 = io_valid_in ? _GEN_27172 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2596 = 12'ha24 == _T_2[11:0] ? image_2596 : _GEN_2595; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5669 = 12'ha25 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8741 = 12'ha25 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5669; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11813 = 12'ha25 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8741; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14885 = 12'ha25 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11813; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17957 = 12'ha25 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14885; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21029 = 12'ha25 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17957; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24101 = 12'ha25 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21029; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27173 = 12'ha25 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24101; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2597 = io_valid_in ? _GEN_27173 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2597 = 12'ha25 == _T_2[11:0] ? image_2597 : _GEN_2596; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5670 = 12'ha26 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8742 = 12'ha26 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5670; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11814 = 12'ha26 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8742; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14886 = 12'ha26 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11814; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17958 = 12'ha26 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14886; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21030 = 12'ha26 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17958; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24102 = 12'ha26 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21030; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27174 = 12'ha26 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24102; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2598 = io_valid_in ? _GEN_27174 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2598 = 12'ha26 == _T_2[11:0] ? image_2598 : _GEN_2597; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5671 = 12'ha27 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8743 = 12'ha27 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5671; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11815 = 12'ha27 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8743; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14887 = 12'ha27 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11815; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17959 = 12'ha27 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14887; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21031 = 12'ha27 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17959; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24103 = 12'ha27 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21031; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27175 = 12'ha27 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24103; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2599 = io_valid_in ? _GEN_27175 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2599 = 12'ha27 == _T_2[11:0] ? image_2599 : _GEN_2598; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5672 = 12'ha28 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8744 = 12'ha28 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5672; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11816 = 12'ha28 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8744; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14888 = 12'ha28 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11816; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17960 = 12'ha28 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14888; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21032 = 12'ha28 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17960; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24104 = 12'ha28 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21032; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27176 = 12'ha28 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24104; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2600 = io_valid_in ? _GEN_27176 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2600 = 12'ha28 == _T_2[11:0] ? image_2600 : _GEN_2599; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5673 = 12'ha29 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8745 = 12'ha29 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5673; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11817 = 12'ha29 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8745; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14889 = 12'ha29 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11817; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17961 = 12'ha29 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14889; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21033 = 12'ha29 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17961; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24105 = 12'ha29 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21033; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27177 = 12'ha29 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24105; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2601 = io_valid_in ? _GEN_27177 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2601 = 12'ha29 == _T_2[11:0] ? image_2601 : _GEN_2600; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5674 = 12'ha2a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8746 = 12'ha2a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5674; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11818 = 12'ha2a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8746; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14890 = 12'ha2a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11818; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17962 = 12'ha2a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14890; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21034 = 12'ha2a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17962; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24106 = 12'ha2a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21034; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27178 = 12'ha2a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24106; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2602 = io_valid_in ? _GEN_27178 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2602 = 12'ha2a == _T_2[11:0] ? image_2602 : _GEN_2601; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5675 = 12'ha2b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8747 = 12'ha2b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5675; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11819 = 12'ha2b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8747; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14891 = 12'ha2b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11819; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17963 = 12'ha2b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14891; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21035 = 12'ha2b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17963; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24107 = 12'ha2b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21035; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27179 = 12'ha2b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24107; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2603 = io_valid_in ? _GEN_27179 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2603 = 12'ha2b == _T_2[11:0] ? image_2603 : _GEN_2602; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5676 = 12'ha2c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8748 = 12'ha2c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5676; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11820 = 12'ha2c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8748; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14892 = 12'ha2c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11820; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17964 = 12'ha2c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14892; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21036 = 12'ha2c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17964; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24108 = 12'ha2c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21036; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27180 = 12'ha2c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24108; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2604 = io_valid_in ? _GEN_27180 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2604 = 12'ha2c == _T_2[11:0] ? image_2604 : _GEN_2603; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5677 = 12'ha2d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8749 = 12'ha2d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5677; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11821 = 12'ha2d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8749; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14893 = 12'ha2d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11821; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17965 = 12'ha2d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14893; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21037 = 12'ha2d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17965; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24109 = 12'ha2d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21037; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27181 = 12'ha2d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24109; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2605 = io_valid_in ? _GEN_27181 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2605 = 12'ha2d == _T_2[11:0] ? image_2605 : _GEN_2604; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5678 = 12'ha2e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8750 = 12'ha2e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5678; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11822 = 12'ha2e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8750; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14894 = 12'ha2e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11822; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17966 = 12'ha2e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14894; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21038 = 12'ha2e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17966; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24110 = 12'ha2e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21038; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27182 = 12'ha2e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24110; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2606 = io_valid_in ? _GEN_27182 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2606 = 12'ha2e == _T_2[11:0] ? image_2606 : _GEN_2605; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5679 = 12'ha2f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8751 = 12'ha2f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5679; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11823 = 12'ha2f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8751; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14895 = 12'ha2f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11823; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17967 = 12'ha2f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14895; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21039 = 12'ha2f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17967; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24111 = 12'ha2f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21039; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27183 = 12'ha2f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24111; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2607 = io_valid_in ? _GEN_27183 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2607 = 12'ha2f == _T_2[11:0] ? image_2607 : _GEN_2606; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5680 = 12'ha30 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8752 = 12'ha30 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5680; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11824 = 12'ha30 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8752; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14896 = 12'ha30 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11824; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17968 = 12'ha30 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14896; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21040 = 12'ha30 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17968; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24112 = 12'ha30 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21040; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27184 = 12'ha30 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24112; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2608 = io_valid_in ? _GEN_27184 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2608 = 12'ha30 == _T_2[11:0] ? image_2608 : _GEN_2607; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5681 = 12'ha31 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8753 = 12'ha31 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5681; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11825 = 12'ha31 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8753; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14897 = 12'ha31 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11825; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17969 = 12'ha31 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14897; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21041 = 12'ha31 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17969; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24113 = 12'ha31 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21041; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27185 = 12'ha31 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24113; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2609 = io_valid_in ? _GEN_27185 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2609 = 12'ha31 == _T_2[11:0] ? image_2609 : _GEN_2608; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5682 = 12'ha32 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8754 = 12'ha32 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5682; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11826 = 12'ha32 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8754; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14898 = 12'ha32 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11826; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17970 = 12'ha32 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14898; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21042 = 12'ha32 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17970; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24114 = 12'ha32 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21042; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27186 = 12'ha32 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24114; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2610 = io_valid_in ? _GEN_27186 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2610 = 12'ha32 == _T_2[11:0] ? image_2610 : _GEN_2609; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5683 = 12'ha33 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8755 = 12'ha33 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5683; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11827 = 12'ha33 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8755; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14899 = 12'ha33 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11827; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17971 = 12'ha33 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14899; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21043 = 12'ha33 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17971; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24115 = 12'ha33 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21043; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27187 = 12'ha33 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24115; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2611 = io_valid_in ? _GEN_27187 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2611 = 12'ha33 == _T_2[11:0] ? image_2611 : _GEN_2610; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5684 = 12'ha34 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8756 = 12'ha34 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5684; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11828 = 12'ha34 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8756; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14900 = 12'ha34 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11828; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17972 = 12'ha34 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14900; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21044 = 12'ha34 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17972; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24116 = 12'ha34 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21044; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27188 = 12'ha34 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24116; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2612 = io_valid_in ? _GEN_27188 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2612 = 12'ha34 == _T_2[11:0] ? image_2612 : _GEN_2611; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5685 = 12'ha35 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8757 = 12'ha35 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5685; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11829 = 12'ha35 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8757; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14901 = 12'ha35 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11829; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17973 = 12'ha35 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14901; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21045 = 12'ha35 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17973; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24117 = 12'ha35 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21045; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27189 = 12'ha35 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24117; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2613 = io_valid_in ? _GEN_27189 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2613 = 12'ha35 == _T_2[11:0] ? image_2613 : _GEN_2612; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5686 = 12'ha36 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8758 = 12'ha36 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5686; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11830 = 12'ha36 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8758; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14902 = 12'ha36 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11830; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17974 = 12'ha36 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14902; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21046 = 12'ha36 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17974; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24118 = 12'ha36 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21046; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27190 = 12'ha36 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24118; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2614 = io_valid_in ? _GEN_27190 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2614 = 12'ha36 == _T_2[11:0] ? image_2614 : _GEN_2613; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5687 = 12'ha37 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8759 = 12'ha37 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5687; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11831 = 12'ha37 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8759; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14903 = 12'ha37 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11831; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17975 = 12'ha37 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14903; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21047 = 12'ha37 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17975; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24119 = 12'ha37 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21047; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27191 = 12'ha37 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24119; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2615 = io_valid_in ? _GEN_27191 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2615 = 12'ha37 == _T_2[11:0] ? image_2615 : _GEN_2614; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5688 = 12'ha38 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8760 = 12'ha38 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5688; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11832 = 12'ha38 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8760; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14904 = 12'ha38 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11832; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17976 = 12'ha38 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14904; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21048 = 12'ha38 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17976; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24120 = 12'ha38 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21048; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27192 = 12'ha38 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24120; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2616 = io_valid_in ? _GEN_27192 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2616 = 12'ha38 == _T_2[11:0] ? image_2616 : _GEN_2615; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5689 = 12'ha39 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8761 = 12'ha39 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5689; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11833 = 12'ha39 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8761; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14905 = 12'ha39 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11833; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17977 = 12'ha39 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14905; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21049 = 12'ha39 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17977; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24121 = 12'ha39 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21049; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27193 = 12'ha39 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24121; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2617 = io_valid_in ? _GEN_27193 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2617 = 12'ha39 == _T_2[11:0] ? image_2617 : _GEN_2616; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5690 = 12'ha3a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8762 = 12'ha3a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5690; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11834 = 12'ha3a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8762; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14906 = 12'ha3a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11834; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17978 = 12'ha3a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14906; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21050 = 12'ha3a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17978; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24122 = 12'ha3a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21050; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27194 = 12'ha3a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24122; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2618 = io_valid_in ? _GEN_27194 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2618 = 12'ha3a == _T_2[11:0] ? image_2618 : _GEN_2617; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5691 = 12'ha3b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8763 = 12'ha3b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5691; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11835 = 12'ha3b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8763; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14907 = 12'ha3b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11835; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17979 = 12'ha3b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14907; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21051 = 12'ha3b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17979; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24123 = 12'ha3b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21051; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27195 = 12'ha3b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24123; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2619 = io_valid_in ? _GEN_27195 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2619 = 12'ha3b == _T_2[11:0] ? image_2619 : _GEN_2618; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5692 = 12'ha3c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8764 = 12'ha3c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5692; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11836 = 12'ha3c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8764; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14908 = 12'ha3c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11836; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17980 = 12'ha3c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14908; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21052 = 12'ha3c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17980; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24124 = 12'ha3c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21052; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27196 = 12'ha3c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24124; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2620 = io_valid_in ? _GEN_27196 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2620 = 12'ha3c == _T_2[11:0] ? image_2620 : _GEN_2619; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5693 = 12'ha3d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8765 = 12'ha3d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5693; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11837 = 12'ha3d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8765; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14909 = 12'ha3d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11837; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17981 = 12'ha3d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14909; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21053 = 12'ha3d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17981; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24125 = 12'ha3d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21053; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27197 = 12'ha3d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24125; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2621 = io_valid_in ? _GEN_27197 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2621 = 12'ha3d == _T_2[11:0] ? image_2621 : _GEN_2620; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5694 = 12'ha3e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8766 = 12'ha3e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5694; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11838 = 12'ha3e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8766; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14910 = 12'ha3e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11838; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17982 = 12'ha3e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14910; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21054 = 12'ha3e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17982; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24126 = 12'ha3e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21054; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27198 = 12'ha3e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24126; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2622 = io_valid_in ? _GEN_27198 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2622 = 12'ha3e == _T_2[11:0] ? image_2622 : _GEN_2621; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5695 = 12'ha3f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8767 = 12'ha3f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5695; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11839 = 12'ha3f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8767; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14911 = 12'ha3f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11839; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17983 = 12'ha3f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14911; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21055 = 12'ha3f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17983; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24127 = 12'ha3f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21055; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27199 = 12'ha3f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24127; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2623 = io_valid_in ? _GEN_27199 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2623 = 12'ha3f == _T_2[11:0] ? image_2623 : _GEN_2622; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5696 = 12'ha40 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8768 = 12'ha40 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5696; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11840 = 12'ha40 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8768; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14912 = 12'ha40 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11840; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17984 = 12'ha40 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14912; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21056 = 12'ha40 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17984; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24128 = 12'ha40 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21056; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27200 = 12'ha40 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24128; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2624 = io_valid_in ? _GEN_27200 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2624 = 12'ha40 == _T_2[11:0] ? image_2624 : _GEN_2623; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5697 = 12'ha41 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8769 = 12'ha41 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5697; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11841 = 12'ha41 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8769; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14913 = 12'ha41 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11841; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17985 = 12'ha41 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14913; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21057 = 12'ha41 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17985; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24129 = 12'ha41 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21057; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27201 = 12'ha41 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24129; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2625 = io_valid_in ? _GEN_27201 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2625 = 12'ha41 == _T_2[11:0] ? image_2625 : _GEN_2624; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5698 = 12'ha42 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8770 = 12'ha42 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5698; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11842 = 12'ha42 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8770; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14914 = 12'ha42 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11842; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17986 = 12'ha42 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14914; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21058 = 12'ha42 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17986; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24130 = 12'ha42 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21058; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27202 = 12'ha42 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24130; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2626 = io_valid_in ? _GEN_27202 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2626 = 12'ha42 == _T_2[11:0] ? image_2626 : _GEN_2625; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5699 = 12'ha43 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8771 = 12'ha43 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5699; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11843 = 12'ha43 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8771; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14915 = 12'ha43 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11843; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17987 = 12'ha43 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14915; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21059 = 12'ha43 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17987; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24131 = 12'ha43 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21059; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27203 = 12'ha43 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24131; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2627 = io_valid_in ? _GEN_27203 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2627 = 12'ha43 == _T_2[11:0] ? image_2627 : _GEN_2626; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5700 = 12'ha44 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8772 = 12'ha44 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5700; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11844 = 12'ha44 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8772; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14916 = 12'ha44 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11844; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17988 = 12'ha44 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14916; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21060 = 12'ha44 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17988; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24132 = 12'ha44 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21060; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27204 = 12'ha44 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24132; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2628 = io_valid_in ? _GEN_27204 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2628 = 12'ha44 == _T_2[11:0] ? image_2628 : _GEN_2627; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5701 = 12'ha45 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8773 = 12'ha45 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5701; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11845 = 12'ha45 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8773; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14917 = 12'ha45 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11845; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17989 = 12'ha45 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14917; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21061 = 12'ha45 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17989; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24133 = 12'ha45 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21061; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27205 = 12'ha45 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24133; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2629 = io_valid_in ? _GEN_27205 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2629 = 12'ha45 == _T_2[11:0] ? image_2629 : _GEN_2628; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5702 = 12'ha46 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8774 = 12'ha46 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5702; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11846 = 12'ha46 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8774; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14918 = 12'ha46 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11846; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17990 = 12'ha46 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14918; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21062 = 12'ha46 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17990; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24134 = 12'ha46 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21062; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27206 = 12'ha46 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24134; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2630 = io_valid_in ? _GEN_27206 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2630 = 12'ha46 == _T_2[11:0] ? image_2630 : _GEN_2629; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5703 = 12'ha47 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8775 = 12'ha47 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5703; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11847 = 12'ha47 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8775; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14919 = 12'ha47 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11847; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17991 = 12'ha47 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14919; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21063 = 12'ha47 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17991; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24135 = 12'ha47 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21063; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27207 = 12'ha47 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24135; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2631 = io_valid_in ? _GEN_27207 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2631 = 12'ha47 == _T_2[11:0] ? image_2631 : _GEN_2630; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5704 = 12'ha48 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8776 = 12'ha48 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5704; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11848 = 12'ha48 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8776; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14920 = 12'ha48 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11848; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17992 = 12'ha48 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14920; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21064 = 12'ha48 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17992; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24136 = 12'ha48 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21064; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27208 = 12'ha48 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24136; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2632 = io_valid_in ? _GEN_27208 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2632 = 12'ha48 == _T_2[11:0] ? image_2632 : _GEN_2631; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5705 = 12'ha49 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8777 = 12'ha49 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5705; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11849 = 12'ha49 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8777; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14921 = 12'ha49 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11849; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17993 = 12'ha49 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14921; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21065 = 12'ha49 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17993; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24137 = 12'ha49 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21065; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27209 = 12'ha49 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24137; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2633 = io_valid_in ? _GEN_27209 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2633 = 12'ha49 == _T_2[11:0] ? image_2633 : _GEN_2632; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5706 = 12'ha4a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8778 = 12'ha4a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5706; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11850 = 12'ha4a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8778; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14922 = 12'ha4a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11850; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17994 = 12'ha4a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14922; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21066 = 12'ha4a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17994; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24138 = 12'ha4a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21066; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27210 = 12'ha4a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24138; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2634 = io_valid_in ? _GEN_27210 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2634 = 12'ha4a == _T_2[11:0] ? image_2634 : _GEN_2633; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5707 = 12'ha4b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8779 = 12'ha4b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5707; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11851 = 12'ha4b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8779; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14923 = 12'ha4b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11851; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17995 = 12'ha4b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14923; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21067 = 12'ha4b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17995; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24139 = 12'ha4b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21067; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27211 = 12'ha4b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24139; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2635 = io_valid_in ? _GEN_27211 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2635 = 12'ha4b == _T_2[11:0] ? image_2635 : _GEN_2634; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5708 = 12'ha4c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8780 = 12'ha4c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5708; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11852 = 12'ha4c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8780; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14924 = 12'ha4c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11852; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17996 = 12'ha4c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14924; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21068 = 12'ha4c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17996; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24140 = 12'ha4c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21068; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27212 = 12'ha4c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24140; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2636 = io_valid_in ? _GEN_27212 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2636 = 12'ha4c == _T_2[11:0] ? image_2636 : _GEN_2635; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5709 = 12'ha4d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8781 = 12'ha4d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5709; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11853 = 12'ha4d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8781; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14925 = 12'ha4d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11853; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17997 = 12'ha4d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14925; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21069 = 12'ha4d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17997; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24141 = 12'ha4d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21069; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27213 = 12'ha4d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24141; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2637 = io_valid_in ? _GEN_27213 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2637 = 12'ha4d == _T_2[11:0] ? image_2637 : _GEN_2636; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5710 = 12'ha4e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8782 = 12'ha4e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5710; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11854 = 12'ha4e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8782; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14926 = 12'ha4e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11854; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17998 = 12'ha4e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14926; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21070 = 12'ha4e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17998; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24142 = 12'ha4e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21070; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27214 = 12'ha4e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24142; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2638 = io_valid_in ? _GEN_27214 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2638 = 12'ha4e == _T_2[11:0] ? image_2638 : _GEN_2637; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5711 = 12'ha4f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8783 = 12'ha4f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5711; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11855 = 12'ha4f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8783; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14927 = 12'ha4f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11855; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_17999 = 12'ha4f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14927; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21071 = 12'ha4f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_17999; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24143 = 12'ha4f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21071; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27215 = 12'ha4f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24143; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2639 = io_valid_in ? _GEN_27215 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2639 = 12'ha4f == _T_2[11:0] ? image_2639 : _GEN_2638; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5712 = 12'ha50 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8784 = 12'ha50 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5712; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11856 = 12'ha50 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8784; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14928 = 12'ha50 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11856; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18000 = 12'ha50 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14928; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21072 = 12'ha50 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18000; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24144 = 12'ha50 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21072; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27216 = 12'ha50 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24144; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2640 = io_valid_in ? _GEN_27216 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2640 = 12'ha50 == _T_2[11:0] ? image_2640 : _GEN_2639; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5713 = 12'ha51 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8785 = 12'ha51 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5713; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11857 = 12'ha51 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8785; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14929 = 12'ha51 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11857; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18001 = 12'ha51 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14929; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21073 = 12'ha51 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18001; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24145 = 12'ha51 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21073; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27217 = 12'ha51 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24145; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2641 = io_valid_in ? _GEN_27217 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2641 = 12'ha51 == _T_2[11:0] ? image_2641 : _GEN_2640; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5714 = 12'ha52 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8786 = 12'ha52 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5714; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11858 = 12'ha52 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8786; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14930 = 12'ha52 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11858; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18002 = 12'ha52 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14930; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21074 = 12'ha52 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18002; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24146 = 12'ha52 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21074; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27218 = 12'ha52 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24146; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2642 = io_valid_in ? _GEN_27218 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2642 = 12'ha52 == _T_2[11:0] ? image_2642 : _GEN_2641; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5715 = 12'ha53 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8787 = 12'ha53 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5715; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11859 = 12'ha53 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8787; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14931 = 12'ha53 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11859; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18003 = 12'ha53 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14931; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21075 = 12'ha53 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18003; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24147 = 12'ha53 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21075; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27219 = 12'ha53 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24147; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2643 = io_valid_in ? _GEN_27219 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2643 = 12'ha53 == _T_2[11:0] ? image_2643 : _GEN_2642; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5716 = 12'ha54 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8788 = 12'ha54 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5716; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11860 = 12'ha54 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8788; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14932 = 12'ha54 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11860; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18004 = 12'ha54 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14932; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21076 = 12'ha54 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18004; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24148 = 12'ha54 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21076; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27220 = 12'ha54 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24148; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2644 = io_valid_in ? _GEN_27220 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2644 = 12'ha54 == _T_2[11:0] ? image_2644 : _GEN_2643; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5717 = 12'ha55 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8789 = 12'ha55 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5717; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11861 = 12'ha55 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8789; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14933 = 12'ha55 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11861; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18005 = 12'ha55 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14933; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21077 = 12'ha55 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18005; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24149 = 12'ha55 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21077; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27221 = 12'ha55 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24149; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2645 = io_valid_in ? _GEN_27221 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2645 = 12'ha55 == _T_2[11:0] ? image_2645 : _GEN_2644; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5718 = 12'ha56 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8790 = 12'ha56 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5718; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11862 = 12'ha56 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8790; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14934 = 12'ha56 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11862; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18006 = 12'ha56 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14934; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21078 = 12'ha56 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18006; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24150 = 12'ha56 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21078; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27222 = 12'ha56 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24150; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2646 = io_valid_in ? _GEN_27222 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2646 = 12'ha56 == _T_2[11:0] ? image_2646 : _GEN_2645; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5719 = 12'ha57 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8791 = 12'ha57 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5719; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11863 = 12'ha57 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8791; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14935 = 12'ha57 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11863; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18007 = 12'ha57 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14935; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21079 = 12'ha57 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18007; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24151 = 12'ha57 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21079; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27223 = 12'ha57 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24151; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2647 = io_valid_in ? _GEN_27223 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2647 = 12'ha57 == _T_2[11:0] ? image_2647 : _GEN_2646; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5720 = 12'ha58 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8792 = 12'ha58 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5720; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11864 = 12'ha58 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8792; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14936 = 12'ha58 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11864; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18008 = 12'ha58 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14936; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21080 = 12'ha58 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18008; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24152 = 12'ha58 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21080; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27224 = 12'ha58 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24152; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2648 = io_valid_in ? _GEN_27224 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2648 = 12'ha58 == _T_2[11:0] ? image_2648 : _GEN_2647; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5721 = 12'ha59 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8793 = 12'ha59 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5721; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11865 = 12'ha59 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8793; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14937 = 12'ha59 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11865; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18009 = 12'ha59 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14937; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21081 = 12'ha59 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18009; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24153 = 12'ha59 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21081; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27225 = 12'ha59 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24153; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2649 = io_valid_in ? _GEN_27225 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2649 = 12'ha59 == _T_2[11:0] ? image_2649 : _GEN_2648; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5722 = 12'ha5a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8794 = 12'ha5a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5722; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11866 = 12'ha5a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8794; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14938 = 12'ha5a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11866; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18010 = 12'ha5a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14938; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21082 = 12'ha5a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18010; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24154 = 12'ha5a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21082; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27226 = 12'ha5a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24154; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2650 = io_valid_in ? _GEN_27226 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2650 = 12'ha5a == _T_2[11:0] ? image_2650 : _GEN_2649; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5723 = 12'ha5b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8795 = 12'ha5b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5723; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11867 = 12'ha5b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8795; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14939 = 12'ha5b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11867; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18011 = 12'ha5b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14939; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21083 = 12'ha5b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18011; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24155 = 12'ha5b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21083; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27227 = 12'ha5b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24155; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2651 = io_valid_in ? _GEN_27227 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2651 = 12'ha5b == _T_2[11:0] ? image_2651 : _GEN_2650; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5724 = 12'ha5c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8796 = 12'ha5c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5724; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11868 = 12'ha5c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8796; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14940 = 12'ha5c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11868; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18012 = 12'ha5c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14940; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21084 = 12'ha5c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18012; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24156 = 12'ha5c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21084; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27228 = 12'ha5c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24156; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2652 = io_valid_in ? _GEN_27228 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2652 = 12'ha5c == _T_2[11:0] ? image_2652 : _GEN_2651; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5725 = 12'ha5d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8797 = 12'ha5d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5725; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11869 = 12'ha5d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8797; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14941 = 12'ha5d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11869; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18013 = 12'ha5d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14941; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21085 = 12'ha5d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18013; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24157 = 12'ha5d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21085; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27229 = 12'ha5d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24157; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2653 = io_valid_in ? _GEN_27229 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2653 = 12'ha5d == _T_2[11:0] ? image_2653 : _GEN_2652; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5726 = 12'ha5e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8798 = 12'ha5e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5726; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11870 = 12'ha5e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8798; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14942 = 12'ha5e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11870; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18014 = 12'ha5e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14942; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21086 = 12'ha5e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18014; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24158 = 12'ha5e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21086; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27230 = 12'ha5e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24158; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2654 = io_valid_in ? _GEN_27230 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2654 = 12'ha5e == _T_2[11:0] ? image_2654 : _GEN_2653; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5727 = 12'ha5f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8799 = 12'ha5f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5727; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11871 = 12'ha5f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8799; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14943 = 12'ha5f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11871; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18015 = 12'ha5f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14943; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21087 = 12'ha5f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18015; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24159 = 12'ha5f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21087; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27231 = 12'ha5f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24159; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2655 = io_valid_in ? _GEN_27231 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2655 = 12'ha5f == _T_2[11:0] ? image_2655 : _GEN_2654; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5728 = 12'ha60 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8800 = 12'ha60 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5728; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11872 = 12'ha60 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8800; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14944 = 12'ha60 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11872; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18016 = 12'ha60 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14944; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21088 = 12'ha60 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18016; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24160 = 12'ha60 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21088; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27232 = 12'ha60 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24160; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2656 = io_valid_in ? _GEN_27232 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2656 = 12'ha60 == _T_2[11:0] ? image_2656 : _GEN_2655; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5729 = 12'ha61 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8801 = 12'ha61 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5729; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11873 = 12'ha61 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8801; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14945 = 12'ha61 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11873; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18017 = 12'ha61 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14945; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21089 = 12'ha61 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18017; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24161 = 12'ha61 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21089; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27233 = 12'ha61 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24161; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2657 = io_valid_in ? _GEN_27233 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2657 = 12'ha61 == _T_2[11:0] ? image_2657 : _GEN_2656; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5730 = 12'ha62 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8802 = 12'ha62 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5730; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11874 = 12'ha62 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8802; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14946 = 12'ha62 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11874; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18018 = 12'ha62 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14946; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21090 = 12'ha62 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18018; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24162 = 12'ha62 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21090; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27234 = 12'ha62 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24162; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2658 = io_valid_in ? _GEN_27234 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2658 = 12'ha62 == _T_2[11:0] ? image_2658 : _GEN_2657; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5731 = 12'ha63 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8803 = 12'ha63 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5731; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11875 = 12'ha63 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8803; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14947 = 12'ha63 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11875; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18019 = 12'ha63 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14947; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21091 = 12'ha63 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18019; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24163 = 12'ha63 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21091; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27235 = 12'ha63 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24163; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2659 = io_valid_in ? _GEN_27235 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2659 = 12'ha63 == _T_2[11:0] ? image_2659 : _GEN_2658; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5732 = 12'ha64 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8804 = 12'ha64 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5732; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11876 = 12'ha64 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8804; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14948 = 12'ha64 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11876; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18020 = 12'ha64 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14948; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21092 = 12'ha64 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18020; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24164 = 12'ha64 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21092; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27236 = 12'ha64 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24164; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2660 = io_valid_in ? _GEN_27236 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2660 = 12'ha64 == _T_2[11:0] ? image_2660 : _GEN_2659; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5733 = 12'ha65 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8805 = 12'ha65 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5733; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11877 = 12'ha65 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8805; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14949 = 12'ha65 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11877; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18021 = 12'ha65 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14949; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21093 = 12'ha65 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18021; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24165 = 12'ha65 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21093; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27237 = 12'ha65 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24165; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2661 = io_valid_in ? _GEN_27237 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2661 = 12'ha65 == _T_2[11:0] ? image_2661 : _GEN_2660; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5734 = 12'ha66 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8806 = 12'ha66 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5734; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11878 = 12'ha66 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8806; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14950 = 12'ha66 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11878; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18022 = 12'ha66 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14950; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21094 = 12'ha66 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18022; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24166 = 12'ha66 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21094; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27238 = 12'ha66 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24166; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2662 = io_valid_in ? _GEN_27238 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2662 = 12'ha66 == _T_2[11:0] ? image_2662 : _GEN_2661; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5735 = 12'ha67 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8807 = 12'ha67 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5735; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11879 = 12'ha67 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8807; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14951 = 12'ha67 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11879; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18023 = 12'ha67 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14951; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21095 = 12'ha67 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18023; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24167 = 12'ha67 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21095; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27239 = 12'ha67 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24167; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2663 = io_valid_in ? _GEN_27239 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2663 = 12'ha67 == _T_2[11:0] ? image_2663 : _GEN_2662; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5736 = 12'ha68 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8808 = 12'ha68 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5736; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11880 = 12'ha68 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8808; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14952 = 12'ha68 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11880; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18024 = 12'ha68 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14952; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21096 = 12'ha68 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18024; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24168 = 12'ha68 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21096; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27240 = 12'ha68 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24168; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2664 = io_valid_in ? _GEN_27240 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2664 = 12'ha68 == _T_2[11:0] ? image_2664 : _GEN_2663; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5737 = 12'ha69 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8809 = 12'ha69 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5737; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11881 = 12'ha69 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8809; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14953 = 12'ha69 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11881; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18025 = 12'ha69 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14953; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21097 = 12'ha69 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18025; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24169 = 12'ha69 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21097; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27241 = 12'ha69 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24169; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2665 = io_valid_in ? _GEN_27241 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2665 = 12'ha69 == _T_2[11:0] ? image_2665 : _GEN_2664; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5738 = 12'ha6a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8810 = 12'ha6a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5738; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11882 = 12'ha6a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8810; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14954 = 12'ha6a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11882; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18026 = 12'ha6a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14954; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21098 = 12'ha6a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18026; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24170 = 12'ha6a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21098; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27242 = 12'ha6a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24170; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2666 = io_valid_in ? _GEN_27242 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2666 = 12'ha6a == _T_2[11:0] ? image_2666 : _GEN_2665; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5739 = 12'ha6b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8811 = 12'ha6b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5739; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11883 = 12'ha6b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8811; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14955 = 12'ha6b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11883; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18027 = 12'ha6b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14955; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21099 = 12'ha6b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18027; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24171 = 12'ha6b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21099; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27243 = 12'ha6b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24171; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2667 = io_valid_in ? _GEN_27243 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2667 = 12'ha6b == _T_2[11:0] ? image_2667 : _GEN_2666; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5740 = 12'ha6c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8812 = 12'ha6c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5740; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11884 = 12'ha6c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8812; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14956 = 12'ha6c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11884; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18028 = 12'ha6c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14956; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21100 = 12'ha6c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18028; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24172 = 12'ha6c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21100; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27244 = 12'ha6c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24172; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2668 = io_valid_in ? _GEN_27244 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2668 = 12'ha6c == _T_2[11:0] ? image_2668 : _GEN_2667; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5741 = 12'ha6d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8813 = 12'ha6d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5741; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11885 = 12'ha6d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8813; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14957 = 12'ha6d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11885; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18029 = 12'ha6d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14957; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21101 = 12'ha6d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18029; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24173 = 12'ha6d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21101; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27245 = 12'ha6d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24173; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2669 = io_valid_in ? _GEN_27245 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2669 = 12'ha6d == _T_2[11:0] ? image_2669 : _GEN_2668; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5742 = 12'ha6e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8814 = 12'ha6e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5742; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11886 = 12'ha6e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8814; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14958 = 12'ha6e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11886; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18030 = 12'ha6e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14958; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21102 = 12'ha6e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18030; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24174 = 12'ha6e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21102; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27246 = 12'ha6e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24174; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2670 = io_valid_in ? _GEN_27246 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2670 = 12'ha6e == _T_2[11:0] ? image_2670 : _GEN_2669; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5743 = 12'ha6f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8815 = 12'ha6f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5743; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11887 = 12'ha6f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8815; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14959 = 12'ha6f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11887; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18031 = 12'ha6f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14959; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21103 = 12'ha6f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18031; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24175 = 12'ha6f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21103; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27247 = 12'ha6f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24175; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2671 = io_valid_in ? _GEN_27247 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2671 = 12'ha6f == _T_2[11:0] ? image_2671 : _GEN_2670; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5744 = 12'ha70 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8816 = 12'ha70 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5744; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11888 = 12'ha70 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8816; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14960 = 12'ha70 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11888; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18032 = 12'ha70 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14960; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21104 = 12'ha70 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18032; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24176 = 12'ha70 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21104; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27248 = 12'ha70 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24176; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2672 = io_valid_in ? _GEN_27248 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2672 = 12'ha70 == _T_2[11:0] ? image_2672 : _GEN_2671; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5745 = 12'ha71 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8817 = 12'ha71 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5745; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11889 = 12'ha71 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8817; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14961 = 12'ha71 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11889; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18033 = 12'ha71 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14961; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21105 = 12'ha71 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18033; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24177 = 12'ha71 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21105; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27249 = 12'ha71 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24177; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2673 = io_valid_in ? _GEN_27249 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2673 = 12'ha71 == _T_2[11:0] ? image_2673 : _GEN_2672; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5746 = 12'ha72 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8818 = 12'ha72 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5746; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11890 = 12'ha72 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8818; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14962 = 12'ha72 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11890; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18034 = 12'ha72 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14962; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21106 = 12'ha72 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18034; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24178 = 12'ha72 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21106; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27250 = 12'ha72 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24178; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2674 = io_valid_in ? _GEN_27250 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2674 = 12'ha72 == _T_2[11:0] ? image_2674 : _GEN_2673; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5747 = 12'ha73 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8819 = 12'ha73 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5747; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11891 = 12'ha73 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8819; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14963 = 12'ha73 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11891; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18035 = 12'ha73 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14963; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21107 = 12'ha73 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18035; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24179 = 12'ha73 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21107; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27251 = 12'ha73 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24179; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2675 = io_valid_in ? _GEN_27251 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2675 = 12'ha73 == _T_2[11:0] ? image_2675 : _GEN_2674; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5748 = 12'ha74 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8820 = 12'ha74 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5748; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11892 = 12'ha74 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8820; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14964 = 12'ha74 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11892; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18036 = 12'ha74 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14964; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21108 = 12'ha74 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18036; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24180 = 12'ha74 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21108; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27252 = 12'ha74 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24180; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2676 = io_valid_in ? _GEN_27252 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2676 = 12'ha74 == _T_2[11:0] ? image_2676 : _GEN_2675; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5749 = 12'ha75 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8821 = 12'ha75 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5749; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11893 = 12'ha75 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8821; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14965 = 12'ha75 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11893; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18037 = 12'ha75 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14965; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21109 = 12'ha75 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18037; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24181 = 12'ha75 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21109; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27253 = 12'ha75 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24181; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2677 = io_valid_in ? _GEN_27253 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2677 = 12'ha75 == _T_2[11:0] ? image_2677 : _GEN_2676; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5750 = 12'ha76 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8822 = 12'ha76 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5750; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11894 = 12'ha76 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8822; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14966 = 12'ha76 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11894; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18038 = 12'ha76 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14966; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21110 = 12'ha76 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18038; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24182 = 12'ha76 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21110; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27254 = 12'ha76 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24182; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2678 = io_valid_in ? _GEN_27254 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2678 = 12'ha76 == _T_2[11:0] ? image_2678 : _GEN_2677; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5751 = 12'ha77 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8823 = 12'ha77 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5751; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11895 = 12'ha77 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8823; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14967 = 12'ha77 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11895; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18039 = 12'ha77 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14967; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21111 = 12'ha77 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18039; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24183 = 12'ha77 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21111; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27255 = 12'ha77 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24183; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2679 = io_valid_in ? _GEN_27255 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2679 = 12'ha77 == _T_2[11:0] ? image_2679 : _GEN_2678; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5752 = 12'ha78 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8824 = 12'ha78 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5752; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11896 = 12'ha78 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8824; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14968 = 12'ha78 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11896; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18040 = 12'ha78 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14968; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21112 = 12'ha78 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18040; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24184 = 12'ha78 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21112; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27256 = 12'ha78 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24184; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2680 = io_valid_in ? _GEN_27256 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2680 = 12'ha78 == _T_2[11:0] ? image_2680 : _GEN_2679; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5753 = 12'ha79 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8825 = 12'ha79 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5753; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11897 = 12'ha79 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8825; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14969 = 12'ha79 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11897; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18041 = 12'ha79 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14969; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21113 = 12'ha79 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18041; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24185 = 12'ha79 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21113; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27257 = 12'ha79 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24185; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2681 = io_valid_in ? _GEN_27257 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2681 = 12'ha79 == _T_2[11:0] ? image_2681 : _GEN_2680; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5754 = 12'ha7a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8826 = 12'ha7a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5754; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11898 = 12'ha7a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8826; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14970 = 12'ha7a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11898; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18042 = 12'ha7a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14970; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21114 = 12'ha7a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18042; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24186 = 12'ha7a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21114; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27258 = 12'ha7a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24186; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2682 = io_valid_in ? _GEN_27258 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2682 = 12'ha7a == _T_2[11:0] ? image_2682 : _GEN_2681; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5755 = 12'ha7b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8827 = 12'ha7b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5755; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11899 = 12'ha7b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8827; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14971 = 12'ha7b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11899; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18043 = 12'ha7b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14971; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21115 = 12'ha7b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18043; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24187 = 12'ha7b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21115; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27259 = 12'ha7b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24187; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2683 = io_valid_in ? _GEN_27259 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2683 = 12'ha7b == _T_2[11:0] ? image_2683 : _GEN_2682; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5756 = 12'ha7c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8828 = 12'ha7c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5756; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11900 = 12'ha7c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8828; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14972 = 12'ha7c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11900; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18044 = 12'ha7c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14972; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21116 = 12'ha7c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18044; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24188 = 12'ha7c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21116; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27260 = 12'ha7c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24188; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2684 = io_valid_in ? _GEN_27260 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2684 = 12'ha7c == _T_2[11:0] ? image_2684 : _GEN_2683; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5757 = 12'ha7d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8829 = 12'ha7d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5757; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11901 = 12'ha7d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8829; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14973 = 12'ha7d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11901; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18045 = 12'ha7d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14973; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21117 = 12'ha7d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18045; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24189 = 12'ha7d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21117; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27261 = 12'ha7d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24189; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2685 = io_valid_in ? _GEN_27261 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2685 = 12'ha7d == _T_2[11:0] ? image_2685 : _GEN_2684; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5758 = 12'ha7e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8830 = 12'ha7e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5758; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11902 = 12'ha7e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8830; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14974 = 12'ha7e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11902; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18046 = 12'ha7e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14974; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21118 = 12'ha7e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18046; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24190 = 12'ha7e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21118; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27262 = 12'ha7e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24190; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2686 = io_valid_in ? _GEN_27262 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2686 = 12'ha7e == _T_2[11:0] ? image_2686 : _GEN_2685; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5759 = 12'ha7f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8831 = 12'ha7f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5759; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11903 = 12'ha7f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8831; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14975 = 12'ha7f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11903; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18047 = 12'ha7f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14975; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21119 = 12'ha7f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18047; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24191 = 12'ha7f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21119; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27263 = 12'ha7f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24191; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2687 = io_valid_in ? _GEN_27263 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2687 = 12'ha7f == _T_2[11:0] ? image_2687 : _GEN_2686; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5760 = 12'ha80 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8832 = 12'ha80 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5760; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11904 = 12'ha80 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8832; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14976 = 12'ha80 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11904; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18048 = 12'ha80 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14976; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21120 = 12'ha80 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18048; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24192 = 12'ha80 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21120; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27264 = 12'ha80 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24192; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2688 = io_valid_in ? _GEN_27264 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2688 = 12'ha80 == _T_2[11:0] ? image_2688 : _GEN_2687; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5761 = 12'ha81 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8833 = 12'ha81 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5761; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11905 = 12'ha81 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8833; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14977 = 12'ha81 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11905; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18049 = 12'ha81 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14977; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21121 = 12'ha81 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18049; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24193 = 12'ha81 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21121; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27265 = 12'ha81 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24193; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2689 = io_valid_in ? _GEN_27265 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2689 = 12'ha81 == _T_2[11:0] ? image_2689 : _GEN_2688; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5762 = 12'ha82 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8834 = 12'ha82 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5762; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11906 = 12'ha82 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8834; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14978 = 12'ha82 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11906; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18050 = 12'ha82 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14978; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21122 = 12'ha82 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18050; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24194 = 12'ha82 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21122; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27266 = 12'ha82 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24194; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2690 = io_valid_in ? _GEN_27266 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2690 = 12'ha82 == _T_2[11:0] ? image_2690 : _GEN_2689; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5763 = 12'ha83 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8835 = 12'ha83 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5763; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11907 = 12'ha83 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8835; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14979 = 12'ha83 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11907; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18051 = 12'ha83 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14979; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21123 = 12'ha83 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18051; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24195 = 12'ha83 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21123; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27267 = 12'ha83 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24195; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2691 = io_valid_in ? _GEN_27267 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2691 = 12'ha83 == _T_2[11:0] ? image_2691 : _GEN_2690; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5764 = 12'ha84 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8836 = 12'ha84 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5764; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11908 = 12'ha84 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8836; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14980 = 12'ha84 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11908; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18052 = 12'ha84 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14980; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21124 = 12'ha84 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18052; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24196 = 12'ha84 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21124; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27268 = 12'ha84 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24196; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2692 = io_valid_in ? _GEN_27268 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2692 = 12'ha84 == _T_2[11:0] ? image_2692 : _GEN_2691; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5765 = 12'ha85 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8837 = 12'ha85 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5765; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11909 = 12'ha85 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8837; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14981 = 12'ha85 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11909; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18053 = 12'ha85 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14981; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21125 = 12'ha85 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18053; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24197 = 12'ha85 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21125; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27269 = 12'ha85 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24197; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2693 = io_valid_in ? _GEN_27269 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2693 = 12'ha85 == _T_2[11:0] ? image_2693 : _GEN_2692; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5766 = 12'ha86 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8838 = 12'ha86 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5766; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11910 = 12'ha86 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8838; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14982 = 12'ha86 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11910; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18054 = 12'ha86 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14982; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21126 = 12'ha86 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18054; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24198 = 12'ha86 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21126; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27270 = 12'ha86 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24198; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2694 = io_valid_in ? _GEN_27270 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2694 = 12'ha86 == _T_2[11:0] ? image_2694 : _GEN_2693; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5767 = 12'ha87 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8839 = 12'ha87 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5767; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11911 = 12'ha87 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8839; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14983 = 12'ha87 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11911; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18055 = 12'ha87 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14983; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21127 = 12'ha87 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18055; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24199 = 12'ha87 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21127; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27271 = 12'ha87 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24199; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2695 = io_valid_in ? _GEN_27271 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2695 = 12'ha87 == _T_2[11:0] ? image_2695 : _GEN_2694; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5768 = 12'ha88 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8840 = 12'ha88 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5768; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11912 = 12'ha88 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8840; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14984 = 12'ha88 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11912; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18056 = 12'ha88 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14984; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21128 = 12'ha88 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18056; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24200 = 12'ha88 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21128; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27272 = 12'ha88 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24200; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2696 = io_valid_in ? _GEN_27272 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2696 = 12'ha88 == _T_2[11:0] ? image_2696 : _GEN_2695; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5769 = 12'ha89 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8841 = 12'ha89 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5769; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11913 = 12'ha89 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8841; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14985 = 12'ha89 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11913; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18057 = 12'ha89 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14985; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21129 = 12'ha89 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18057; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24201 = 12'ha89 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21129; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27273 = 12'ha89 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24201; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2697 = io_valid_in ? _GEN_27273 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2697 = 12'ha89 == _T_2[11:0] ? image_2697 : _GEN_2696; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5770 = 12'ha8a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8842 = 12'ha8a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5770; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11914 = 12'ha8a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8842; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14986 = 12'ha8a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11914; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18058 = 12'ha8a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14986; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21130 = 12'ha8a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18058; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24202 = 12'ha8a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21130; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27274 = 12'ha8a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24202; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2698 = io_valid_in ? _GEN_27274 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2698 = 12'ha8a == _T_2[11:0] ? image_2698 : _GEN_2697; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5771 = 12'ha8b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8843 = 12'ha8b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5771; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11915 = 12'ha8b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8843; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14987 = 12'ha8b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11915; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18059 = 12'ha8b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14987; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21131 = 12'ha8b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18059; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24203 = 12'ha8b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21131; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27275 = 12'ha8b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24203; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2699 = io_valid_in ? _GEN_27275 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2699 = 12'ha8b == _T_2[11:0] ? image_2699 : _GEN_2698; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5772 = 12'ha8c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8844 = 12'ha8c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5772; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11916 = 12'ha8c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8844; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14988 = 12'ha8c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11916; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18060 = 12'ha8c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14988; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21132 = 12'ha8c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18060; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24204 = 12'ha8c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21132; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27276 = 12'ha8c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24204; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2700 = io_valid_in ? _GEN_27276 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2700 = 12'ha8c == _T_2[11:0] ? image_2700 : _GEN_2699; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5773 = 12'ha8d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8845 = 12'ha8d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5773; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11917 = 12'ha8d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8845; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14989 = 12'ha8d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11917; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18061 = 12'ha8d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14989; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21133 = 12'ha8d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18061; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24205 = 12'ha8d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21133; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27277 = 12'ha8d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24205; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2701 = io_valid_in ? _GEN_27277 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2701 = 12'ha8d == _T_2[11:0] ? image_2701 : _GEN_2700; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5774 = 12'ha8e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8846 = 12'ha8e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5774; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11918 = 12'ha8e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8846; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14990 = 12'ha8e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11918; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18062 = 12'ha8e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14990; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21134 = 12'ha8e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18062; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24206 = 12'ha8e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21134; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27278 = 12'ha8e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24206; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2702 = io_valid_in ? _GEN_27278 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2702 = 12'ha8e == _T_2[11:0] ? image_2702 : _GEN_2701; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5775 = 12'ha8f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8847 = 12'ha8f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5775; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11919 = 12'ha8f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8847; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14991 = 12'ha8f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11919; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18063 = 12'ha8f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14991; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21135 = 12'ha8f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18063; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24207 = 12'ha8f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21135; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27279 = 12'ha8f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24207; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2703 = io_valid_in ? _GEN_27279 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2703 = 12'ha8f == _T_2[11:0] ? image_2703 : _GEN_2702; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5776 = 12'ha90 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8848 = 12'ha90 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5776; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11920 = 12'ha90 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8848; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14992 = 12'ha90 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11920; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18064 = 12'ha90 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14992; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21136 = 12'ha90 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18064; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24208 = 12'ha90 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21136; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27280 = 12'ha90 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24208; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2704 = io_valid_in ? _GEN_27280 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2704 = 12'ha90 == _T_2[11:0] ? image_2704 : _GEN_2703; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5777 = 12'ha91 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8849 = 12'ha91 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5777; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11921 = 12'ha91 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8849; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14993 = 12'ha91 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11921; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18065 = 12'ha91 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14993; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21137 = 12'ha91 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18065; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24209 = 12'ha91 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21137; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27281 = 12'ha91 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24209; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2705 = io_valid_in ? _GEN_27281 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2705 = 12'ha91 == _T_2[11:0] ? image_2705 : _GEN_2704; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5778 = 12'ha92 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8850 = 12'ha92 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5778; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11922 = 12'ha92 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8850; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14994 = 12'ha92 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11922; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18066 = 12'ha92 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14994; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21138 = 12'ha92 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18066; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24210 = 12'ha92 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21138; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27282 = 12'ha92 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24210; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2706 = io_valid_in ? _GEN_27282 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2706 = 12'ha92 == _T_2[11:0] ? image_2706 : _GEN_2705; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5779 = 12'ha93 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8851 = 12'ha93 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5779; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11923 = 12'ha93 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8851; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14995 = 12'ha93 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11923; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18067 = 12'ha93 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14995; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21139 = 12'ha93 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18067; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24211 = 12'ha93 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21139; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27283 = 12'ha93 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24211; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2707 = io_valid_in ? _GEN_27283 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2707 = 12'ha93 == _T_2[11:0] ? image_2707 : _GEN_2706; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5780 = 12'ha94 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8852 = 12'ha94 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5780; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11924 = 12'ha94 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8852; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14996 = 12'ha94 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11924; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18068 = 12'ha94 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14996; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21140 = 12'ha94 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18068; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24212 = 12'ha94 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21140; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27284 = 12'ha94 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24212; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2708 = io_valid_in ? _GEN_27284 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2708 = 12'ha94 == _T_2[11:0] ? image_2708 : _GEN_2707; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5781 = 12'ha95 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8853 = 12'ha95 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5781; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11925 = 12'ha95 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8853; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14997 = 12'ha95 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11925; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18069 = 12'ha95 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14997; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21141 = 12'ha95 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18069; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24213 = 12'ha95 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21141; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27285 = 12'ha95 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24213; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2709 = io_valid_in ? _GEN_27285 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2709 = 12'ha95 == _T_2[11:0] ? image_2709 : _GEN_2708; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5782 = 12'ha96 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8854 = 12'ha96 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5782; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11926 = 12'ha96 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8854; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14998 = 12'ha96 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11926; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18070 = 12'ha96 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14998; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21142 = 12'ha96 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18070; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24214 = 12'ha96 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21142; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27286 = 12'ha96 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24214; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2710 = io_valid_in ? _GEN_27286 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2710 = 12'ha96 == _T_2[11:0] ? image_2710 : _GEN_2709; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5783 = 12'ha97 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8855 = 12'ha97 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5783; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11927 = 12'ha97 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8855; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_14999 = 12'ha97 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11927; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18071 = 12'ha97 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_14999; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21143 = 12'ha97 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18071; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24215 = 12'ha97 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21143; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27287 = 12'ha97 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24215; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2711 = io_valid_in ? _GEN_27287 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2711 = 12'ha97 == _T_2[11:0] ? image_2711 : _GEN_2710; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5784 = 12'ha98 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8856 = 12'ha98 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5784; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11928 = 12'ha98 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8856; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15000 = 12'ha98 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11928; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18072 = 12'ha98 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15000; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21144 = 12'ha98 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18072; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24216 = 12'ha98 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21144; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27288 = 12'ha98 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24216; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2712 = io_valid_in ? _GEN_27288 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2712 = 12'ha98 == _T_2[11:0] ? image_2712 : _GEN_2711; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5785 = 12'ha99 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8857 = 12'ha99 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5785; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11929 = 12'ha99 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8857; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15001 = 12'ha99 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11929; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18073 = 12'ha99 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15001; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21145 = 12'ha99 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18073; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24217 = 12'ha99 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21145; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27289 = 12'ha99 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24217; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2713 = io_valid_in ? _GEN_27289 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2713 = 12'ha99 == _T_2[11:0] ? image_2713 : _GEN_2712; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5786 = 12'ha9a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8858 = 12'ha9a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5786; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11930 = 12'ha9a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8858; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15002 = 12'ha9a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11930; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18074 = 12'ha9a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15002; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21146 = 12'ha9a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18074; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24218 = 12'ha9a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21146; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27290 = 12'ha9a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24218; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2714 = io_valid_in ? _GEN_27290 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2714 = 12'ha9a == _T_2[11:0] ? image_2714 : _GEN_2713; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5787 = 12'ha9b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8859 = 12'ha9b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5787; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11931 = 12'ha9b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8859; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15003 = 12'ha9b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11931; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18075 = 12'ha9b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15003; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21147 = 12'ha9b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18075; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24219 = 12'ha9b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21147; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27291 = 12'ha9b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24219; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2715 = io_valid_in ? _GEN_27291 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2715 = 12'ha9b == _T_2[11:0] ? image_2715 : _GEN_2714; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5788 = 12'ha9c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8860 = 12'ha9c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5788; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11932 = 12'ha9c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8860; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15004 = 12'ha9c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11932; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18076 = 12'ha9c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15004; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21148 = 12'ha9c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18076; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24220 = 12'ha9c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21148; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27292 = 12'ha9c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24220; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2716 = io_valid_in ? _GEN_27292 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2716 = 12'ha9c == _T_2[11:0] ? image_2716 : _GEN_2715; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5789 = 12'ha9d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8861 = 12'ha9d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5789; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11933 = 12'ha9d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8861; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15005 = 12'ha9d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11933; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18077 = 12'ha9d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15005; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21149 = 12'ha9d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18077; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24221 = 12'ha9d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21149; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27293 = 12'ha9d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24221; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2717 = io_valid_in ? _GEN_27293 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2717 = 12'ha9d == _T_2[11:0] ? image_2717 : _GEN_2716; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5790 = 12'ha9e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8862 = 12'ha9e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5790; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11934 = 12'ha9e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8862; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15006 = 12'ha9e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11934; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18078 = 12'ha9e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15006; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21150 = 12'ha9e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18078; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24222 = 12'ha9e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21150; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27294 = 12'ha9e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24222; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2718 = io_valid_in ? _GEN_27294 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2718 = 12'ha9e == _T_2[11:0] ? image_2718 : _GEN_2717; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5791 = 12'ha9f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8863 = 12'ha9f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5791; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11935 = 12'ha9f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8863; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15007 = 12'ha9f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11935; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18079 = 12'ha9f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15007; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21151 = 12'ha9f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18079; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24223 = 12'ha9f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21151; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27295 = 12'ha9f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24223; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2719 = io_valid_in ? _GEN_27295 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2719 = 12'ha9f == _T_2[11:0] ? image_2719 : _GEN_2718; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5792 = 12'haa0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8864 = 12'haa0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5792; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11936 = 12'haa0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8864; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15008 = 12'haa0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11936; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18080 = 12'haa0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15008; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21152 = 12'haa0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18080; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24224 = 12'haa0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21152; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27296 = 12'haa0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24224; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2720 = io_valid_in ? _GEN_27296 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2720 = 12'haa0 == _T_2[11:0] ? image_2720 : _GEN_2719; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5793 = 12'haa1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8865 = 12'haa1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5793; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11937 = 12'haa1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8865; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15009 = 12'haa1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11937; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18081 = 12'haa1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15009; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21153 = 12'haa1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18081; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24225 = 12'haa1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21153; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27297 = 12'haa1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24225; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2721 = io_valid_in ? _GEN_27297 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2721 = 12'haa1 == _T_2[11:0] ? image_2721 : _GEN_2720; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5794 = 12'haa2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8866 = 12'haa2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5794; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11938 = 12'haa2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8866; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15010 = 12'haa2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11938; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18082 = 12'haa2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15010; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21154 = 12'haa2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18082; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24226 = 12'haa2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21154; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27298 = 12'haa2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24226; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2722 = io_valid_in ? _GEN_27298 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2722 = 12'haa2 == _T_2[11:0] ? image_2722 : _GEN_2721; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5795 = 12'haa3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8867 = 12'haa3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5795; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11939 = 12'haa3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8867; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15011 = 12'haa3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11939; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18083 = 12'haa3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15011; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21155 = 12'haa3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18083; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24227 = 12'haa3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21155; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27299 = 12'haa3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24227; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2723 = io_valid_in ? _GEN_27299 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2723 = 12'haa3 == _T_2[11:0] ? image_2723 : _GEN_2722; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5796 = 12'haa4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8868 = 12'haa4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5796; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11940 = 12'haa4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8868; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15012 = 12'haa4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11940; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18084 = 12'haa4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15012; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21156 = 12'haa4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18084; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24228 = 12'haa4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21156; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27300 = 12'haa4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24228; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2724 = io_valid_in ? _GEN_27300 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2724 = 12'haa4 == _T_2[11:0] ? image_2724 : _GEN_2723; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5797 = 12'haa5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8869 = 12'haa5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5797; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11941 = 12'haa5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8869; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15013 = 12'haa5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11941; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18085 = 12'haa5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15013; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21157 = 12'haa5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18085; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24229 = 12'haa5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21157; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27301 = 12'haa5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24229; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2725 = io_valid_in ? _GEN_27301 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2725 = 12'haa5 == _T_2[11:0] ? image_2725 : _GEN_2724; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5798 = 12'haa6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8870 = 12'haa6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5798; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11942 = 12'haa6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8870; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15014 = 12'haa6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11942; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18086 = 12'haa6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15014; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21158 = 12'haa6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18086; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24230 = 12'haa6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21158; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27302 = 12'haa6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24230; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2726 = io_valid_in ? _GEN_27302 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2726 = 12'haa6 == _T_2[11:0] ? image_2726 : _GEN_2725; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5799 = 12'haa7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8871 = 12'haa7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5799; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11943 = 12'haa7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8871; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15015 = 12'haa7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11943; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18087 = 12'haa7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15015; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21159 = 12'haa7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18087; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24231 = 12'haa7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21159; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27303 = 12'haa7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24231; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2727 = io_valid_in ? _GEN_27303 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2727 = 12'haa7 == _T_2[11:0] ? image_2727 : _GEN_2726; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5800 = 12'haa8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8872 = 12'haa8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5800; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11944 = 12'haa8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8872; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15016 = 12'haa8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11944; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18088 = 12'haa8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15016; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21160 = 12'haa8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18088; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24232 = 12'haa8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21160; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27304 = 12'haa8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24232; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2728 = io_valid_in ? _GEN_27304 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2728 = 12'haa8 == _T_2[11:0] ? image_2728 : _GEN_2727; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5801 = 12'haa9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8873 = 12'haa9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5801; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11945 = 12'haa9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8873; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15017 = 12'haa9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11945; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18089 = 12'haa9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15017; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21161 = 12'haa9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18089; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24233 = 12'haa9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21161; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27305 = 12'haa9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24233; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2729 = io_valid_in ? _GEN_27305 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2729 = 12'haa9 == _T_2[11:0] ? image_2729 : _GEN_2728; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5802 = 12'haaa == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8874 = 12'haaa == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5802; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11946 = 12'haaa == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8874; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15018 = 12'haaa == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11946; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18090 = 12'haaa == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15018; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21162 = 12'haaa == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18090; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24234 = 12'haaa == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21162; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27306 = 12'haaa == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24234; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2730 = io_valid_in ? _GEN_27306 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2730 = 12'haaa == _T_2[11:0] ? image_2730 : _GEN_2729; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5803 = 12'haab == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8875 = 12'haab == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5803; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11947 = 12'haab == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8875; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15019 = 12'haab == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11947; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18091 = 12'haab == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15019; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21163 = 12'haab == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18091; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24235 = 12'haab == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21163; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27307 = 12'haab == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24235; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2731 = io_valid_in ? _GEN_27307 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2731 = 12'haab == _T_2[11:0] ? image_2731 : _GEN_2730; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5804 = 12'haac == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8876 = 12'haac == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5804; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11948 = 12'haac == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8876; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15020 = 12'haac == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11948; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18092 = 12'haac == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15020; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21164 = 12'haac == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18092; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24236 = 12'haac == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21164; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27308 = 12'haac == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24236; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2732 = io_valid_in ? _GEN_27308 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2732 = 12'haac == _T_2[11:0] ? image_2732 : _GEN_2731; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5805 = 12'haad == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8877 = 12'haad == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5805; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11949 = 12'haad == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8877; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15021 = 12'haad == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11949; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18093 = 12'haad == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15021; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21165 = 12'haad == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18093; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24237 = 12'haad == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21165; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27309 = 12'haad == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24237; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2733 = io_valid_in ? _GEN_27309 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2733 = 12'haad == _T_2[11:0] ? image_2733 : _GEN_2732; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5806 = 12'haae == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8878 = 12'haae == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5806; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11950 = 12'haae == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8878; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15022 = 12'haae == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11950; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18094 = 12'haae == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15022; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21166 = 12'haae == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18094; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24238 = 12'haae == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21166; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27310 = 12'haae == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24238; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2734 = io_valid_in ? _GEN_27310 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2734 = 12'haae == _T_2[11:0] ? image_2734 : _GEN_2733; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5807 = 12'haaf == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8879 = 12'haaf == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5807; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11951 = 12'haaf == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8879; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15023 = 12'haaf == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11951; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18095 = 12'haaf == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15023; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21167 = 12'haaf == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18095; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24239 = 12'haaf == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21167; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27311 = 12'haaf == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24239; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2735 = io_valid_in ? _GEN_27311 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2735 = 12'haaf == _T_2[11:0] ? image_2735 : _GEN_2734; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5808 = 12'hab0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8880 = 12'hab0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5808; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11952 = 12'hab0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8880; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15024 = 12'hab0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11952; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18096 = 12'hab0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15024; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21168 = 12'hab0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18096; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24240 = 12'hab0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21168; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27312 = 12'hab0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24240; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2736 = io_valid_in ? _GEN_27312 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2736 = 12'hab0 == _T_2[11:0] ? image_2736 : _GEN_2735; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5809 = 12'hab1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8881 = 12'hab1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5809; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11953 = 12'hab1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8881; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15025 = 12'hab1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11953; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18097 = 12'hab1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15025; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21169 = 12'hab1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18097; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24241 = 12'hab1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21169; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27313 = 12'hab1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24241; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2737 = io_valid_in ? _GEN_27313 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2737 = 12'hab1 == _T_2[11:0] ? image_2737 : _GEN_2736; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5810 = 12'hab2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8882 = 12'hab2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5810; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11954 = 12'hab2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8882; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15026 = 12'hab2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11954; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18098 = 12'hab2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15026; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21170 = 12'hab2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18098; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24242 = 12'hab2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21170; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27314 = 12'hab2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24242; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2738 = io_valid_in ? _GEN_27314 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2738 = 12'hab2 == _T_2[11:0] ? image_2738 : _GEN_2737; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5811 = 12'hab3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8883 = 12'hab3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5811; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11955 = 12'hab3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8883; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15027 = 12'hab3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11955; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18099 = 12'hab3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15027; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21171 = 12'hab3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18099; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24243 = 12'hab3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21171; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27315 = 12'hab3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24243; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2739 = io_valid_in ? _GEN_27315 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2739 = 12'hab3 == _T_2[11:0] ? image_2739 : _GEN_2738; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5812 = 12'hab4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8884 = 12'hab4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5812; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11956 = 12'hab4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8884; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15028 = 12'hab4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11956; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18100 = 12'hab4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15028; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21172 = 12'hab4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18100; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24244 = 12'hab4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21172; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27316 = 12'hab4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24244; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2740 = io_valid_in ? _GEN_27316 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2740 = 12'hab4 == _T_2[11:0] ? image_2740 : _GEN_2739; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5813 = 12'hab5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8885 = 12'hab5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5813; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11957 = 12'hab5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8885; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15029 = 12'hab5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11957; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18101 = 12'hab5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15029; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21173 = 12'hab5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18101; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24245 = 12'hab5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21173; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27317 = 12'hab5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24245; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2741 = io_valid_in ? _GEN_27317 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2741 = 12'hab5 == _T_2[11:0] ? image_2741 : _GEN_2740; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5814 = 12'hab6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8886 = 12'hab6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5814; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11958 = 12'hab6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8886; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15030 = 12'hab6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11958; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18102 = 12'hab6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15030; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21174 = 12'hab6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18102; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24246 = 12'hab6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21174; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27318 = 12'hab6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24246; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2742 = io_valid_in ? _GEN_27318 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2742 = 12'hab6 == _T_2[11:0] ? image_2742 : _GEN_2741; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5815 = 12'hab7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8887 = 12'hab7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5815; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11959 = 12'hab7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8887; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15031 = 12'hab7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11959; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18103 = 12'hab7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15031; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21175 = 12'hab7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18103; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24247 = 12'hab7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21175; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27319 = 12'hab7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24247; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2743 = io_valid_in ? _GEN_27319 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2743 = 12'hab7 == _T_2[11:0] ? image_2743 : _GEN_2742; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5816 = 12'hab8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8888 = 12'hab8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5816; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11960 = 12'hab8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8888; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15032 = 12'hab8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11960; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18104 = 12'hab8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15032; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21176 = 12'hab8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18104; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24248 = 12'hab8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21176; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27320 = 12'hab8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24248; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2744 = io_valid_in ? _GEN_27320 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2744 = 12'hab8 == _T_2[11:0] ? image_2744 : _GEN_2743; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5817 = 12'hab9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8889 = 12'hab9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5817; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11961 = 12'hab9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8889; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15033 = 12'hab9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11961; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18105 = 12'hab9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15033; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21177 = 12'hab9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18105; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24249 = 12'hab9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21177; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27321 = 12'hab9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24249; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2745 = io_valid_in ? _GEN_27321 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2745 = 12'hab9 == _T_2[11:0] ? image_2745 : _GEN_2744; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5818 = 12'haba == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8890 = 12'haba == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5818; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11962 = 12'haba == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8890; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15034 = 12'haba == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11962; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18106 = 12'haba == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15034; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21178 = 12'haba == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18106; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24250 = 12'haba == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21178; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27322 = 12'haba == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24250; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2746 = io_valid_in ? _GEN_27322 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2746 = 12'haba == _T_2[11:0] ? image_2746 : _GEN_2745; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5819 = 12'habb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8891 = 12'habb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5819; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11963 = 12'habb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8891; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15035 = 12'habb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11963; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18107 = 12'habb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15035; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21179 = 12'habb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18107; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24251 = 12'habb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21179; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27323 = 12'habb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24251; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2747 = io_valid_in ? _GEN_27323 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2747 = 12'habb == _T_2[11:0] ? image_2747 : _GEN_2746; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5820 = 12'habc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8892 = 12'habc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5820; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11964 = 12'habc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8892; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15036 = 12'habc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11964; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18108 = 12'habc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15036; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21180 = 12'habc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18108; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24252 = 12'habc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21180; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27324 = 12'habc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24252; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2748 = io_valid_in ? _GEN_27324 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2748 = 12'habc == _T_2[11:0] ? image_2748 : _GEN_2747; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5821 = 12'habd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8893 = 12'habd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5821; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11965 = 12'habd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8893; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15037 = 12'habd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11965; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18109 = 12'habd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15037; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21181 = 12'habd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18109; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24253 = 12'habd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21181; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27325 = 12'habd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24253; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2749 = io_valid_in ? _GEN_27325 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2749 = 12'habd == _T_2[11:0] ? image_2749 : _GEN_2748; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5822 = 12'habe == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8894 = 12'habe == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5822; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11966 = 12'habe == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8894; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15038 = 12'habe == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11966; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18110 = 12'habe == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15038; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21182 = 12'habe == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18110; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24254 = 12'habe == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21182; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27326 = 12'habe == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24254; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2750 = io_valid_in ? _GEN_27326 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2750 = 12'habe == _T_2[11:0] ? image_2750 : _GEN_2749; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5823 = 12'habf == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8895 = 12'habf == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5823; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11967 = 12'habf == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8895; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15039 = 12'habf == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11967; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18111 = 12'habf == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15039; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21183 = 12'habf == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18111; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24255 = 12'habf == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21183; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27327 = 12'habf == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24255; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2751 = io_valid_in ? _GEN_27327 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2751 = 12'habf == _T_2[11:0] ? image_2751 : _GEN_2750; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5824 = 12'hac0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8896 = 12'hac0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5824; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11968 = 12'hac0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8896; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15040 = 12'hac0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11968; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18112 = 12'hac0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15040; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21184 = 12'hac0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18112; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24256 = 12'hac0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21184; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27328 = 12'hac0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24256; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2752 = io_valid_in ? _GEN_27328 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2752 = 12'hac0 == _T_2[11:0] ? image_2752 : _GEN_2751; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5825 = 12'hac1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8897 = 12'hac1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5825; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11969 = 12'hac1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8897; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15041 = 12'hac1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11969; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18113 = 12'hac1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15041; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21185 = 12'hac1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18113; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24257 = 12'hac1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21185; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27329 = 12'hac1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24257; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2753 = io_valid_in ? _GEN_27329 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2753 = 12'hac1 == _T_2[11:0] ? image_2753 : _GEN_2752; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5826 = 12'hac2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8898 = 12'hac2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5826; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11970 = 12'hac2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8898; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15042 = 12'hac2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11970; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18114 = 12'hac2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15042; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21186 = 12'hac2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18114; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24258 = 12'hac2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21186; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27330 = 12'hac2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24258; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2754 = io_valid_in ? _GEN_27330 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2754 = 12'hac2 == _T_2[11:0] ? image_2754 : _GEN_2753; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5827 = 12'hac3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8899 = 12'hac3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5827; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11971 = 12'hac3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8899; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15043 = 12'hac3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11971; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18115 = 12'hac3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15043; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21187 = 12'hac3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18115; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24259 = 12'hac3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21187; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27331 = 12'hac3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24259; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2755 = io_valid_in ? _GEN_27331 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2755 = 12'hac3 == _T_2[11:0] ? image_2755 : _GEN_2754; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5828 = 12'hac4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8900 = 12'hac4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5828; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11972 = 12'hac4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8900; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15044 = 12'hac4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11972; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18116 = 12'hac4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15044; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21188 = 12'hac4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18116; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24260 = 12'hac4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21188; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27332 = 12'hac4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24260; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2756 = io_valid_in ? _GEN_27332 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2756 = 12'hac4 == _T_2[11:0] ? image_2756 : _GEN_2755; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5829 = 12'hac5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8901 = 12'hac5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5829; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11973 = 12'hac5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8901; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15045 = 12'hac5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11973; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18117 = 12'hac5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15045; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21189 = 12'hac5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18117; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24261 = 12'hac5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21189; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27333 = 12'hac5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24261; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2757 = io_valid_in ? _GEN_27333 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2757 = 12'hac5 == _T_2[11:0] ? image_2757 : _GEN_2756; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5830 = 12'hac6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8902 = 12'hac6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5830; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11974 = 12'hac6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8902; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15046 = 12'hac6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11974; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18118 = 12'hac6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15046; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21190 = 12'hac6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18118; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24262 = 12'hac6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21190; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27334 = 12'hac6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24262; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2758 = io_valid_in ? _GEN_27334 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2758 = 12'hac6 == _T_2[11:0] ? image_2758 : _GEN_2757; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5831 = 12'hac7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8903 = 12'hac7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5831; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11975 = 12'hac7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8903; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15047 = 12'hac7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11975; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18119 = 12'hac7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15047; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21191 = 12'hac7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18119; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24263 = 12'hac7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21191; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27335 = 12'hac7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24263; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2759 = io_valid_in ? _GEN_27335 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2759 = 12'hac7 == _T_2[11:0] ? image_2759 : _GEN_2758; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5832 = 12'hac8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8904 = 12'hac8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5832; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11976 = 12'hac8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8904; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15048 = 12'hac8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11976; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18120 = 12'hac8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15048; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21192 = 12'hac8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18120; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24264 = 12'hac8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21192; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27336 = 12'hac8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24264; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2760 = io_valid_in ? _GEN_27336 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2760 = 12'hac8 == _T_2[11:0] ? image_2760 : _GEN_2759; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5833 = 12'hac9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8905 = 12'hac9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5833; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11977 = 12'hac9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8905; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15049 = 12'hac9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11977; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18121 = 12'hac9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15049; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21193 = 12'hac9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18121; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24265 = 12'hac9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21193; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27337 = 12'hac9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24265; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2761 = io_valid_in ? _GEN_27337 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2761 = 12'hac9 == _T_2[11:0] ? image_2761 : _GEN_2760; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5834 = 12'haca == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8906 = 12'haca == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5834; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11978 = 12'haca == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8906; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15050 = 12'haca == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11978; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18122 = 12'haca == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15050; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21194 = 12'haca == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18122; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24266 = 12'haca == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21194; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27338 = 12'haca == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24266; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2762 = io_valid_in ? _GEN_27338 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2762 = 12'haca == _T_2[11:0] ? image_2762 : _GEN_2761; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5835 = 12'hacb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8907 = 12'hacb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5835; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11979 = 12'hacb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8907; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15051 = 12'hacb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11979; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18123 = 12'hacb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15051; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21195 = 12'hacb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18123; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24267 = 12'hacb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21195; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27339 = 12'hacb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24267; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2763 = io_valid_in ? _GEN_27339 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2763 = 12'hacb == _T_2[11:0] ? image_2763 : _GEN_2762; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5836 = 12'hacc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8908 = 12'hacc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5836; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11980 = 12'hacc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8908; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15052 = 12'hacc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11980; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18124 = 12'hacc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15052; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21196 = 12'hacc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18124; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24268 = 12'hacc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21196; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27340 = 12'hacc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24268; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2764 = io_valid_in ? _GEN_27340 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2764 = 12'hacc == _T_2[11:0] ? image_2764 : _GEN_2763; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5837 = 12'hacd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8909 = 12'hacd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5837; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11981 = 12'hacd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8909; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15053 = 12'hacd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11981; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18125 = 12'hacd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15053; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21197 = 12'hacd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18125; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24269 = 12'hacd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21197; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27341 = 12'hacd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24269; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2765 = io_valid_in ? _GEN_27341 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2765 = 12'hacd == _T_2[11:0] ? image_2765 : _GEN_2764; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5838 = 12'hace == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8910 = 12'hace == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5838; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11982 = 12'hace == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8910; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15054 = 12'hace == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11982; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18126 = 12'hace == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15054; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21198 = 12'hace == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18126; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24270 = 12'hace == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21198; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27342 = 12'hace == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24270; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2766 = io_valid_in ? _GEN_27342 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2766 = 12'hace == _T_2[11:0] ? image_2766 : _GEN_2765; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5839 = 12'hacf == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8911 = 12'hacf == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5839; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11983 = 12'hacf == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8911; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15055 = 12'hacf == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11983; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18127 = 12'hacf == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15055; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21199 = 12'hacf == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18127; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24271 = 12'hacf == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21199; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27343 = 12'hacf == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24271; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2767 = io_valid_in ? _GEN_27343 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2767 = 12'hacf == _T_2[11:0] ? image_2767 : _GEN_2766; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5840 = 12'had0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8912 = 12'had0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5840; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11984 = 12'had0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8912; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15056 = 12'had0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11984; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18128 = 12'had0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15056; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21200 = 12'had0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18128; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24272 = 12'had0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21200; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27344 = 12'had0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24272; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2768 = io_valid_in ? _GEN_27344 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2768 = 12'had0 == _T_2[11:0] ? image_2768 : _GEN_2767; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5841 = 12'had1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8913 = 12'had1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5841; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11985 = 12'had1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8913; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15057 = 12'had1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11985; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18129 = 12'had1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15057; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21201 = 12'had1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18129; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24273 = 12'had1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21201; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27345 = 12'had1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24273; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2769 = io_valid_in ? _GEN_27345 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2769 = 12'had1 == _T_2[11:0] ? image_2769 : _GEN_2768; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5842 = 12'had2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8914 = 12'had2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5842; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11986 = 12'had2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8914; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15058 = 12'had2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11986; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18130 = 12'had2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15058; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21202 = 12'had2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18130; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24274 = 12'had2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21202; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27346 = 12'had2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24274; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2770 = io_valid_in ? _GEN_27346 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2770 = 12'had2 == _T_2[11:0] ? image_2770 : _GEN_2769; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5843 = 12'had3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8915 = 12'had3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5843; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11987 = 12'had3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8915; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15059 = 12'had3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11987; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18131 = 12'had3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15059; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21203 = 12'had3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18131; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24275 = 12'had3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21203; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27347 = 12'had3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24275; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2771 = io_valid_in ? _GEN_27347 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2771 = 12'had3 == _T_2[11:0] ? image_2771 : _GEN_2770; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5844 = 12'had4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8916 = 12'had4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5844; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11988 = 12'had4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8916; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15060 = 12'had4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11988; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18132 = 12'had4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15060; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21204 = 12'had4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18132; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24276 = 12'had4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21204; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27348 = 12'had4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24276; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2772 = io_valid_in ? _GEN_27348 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2772 = 12'had4 == _T_2[11:0] ? image_2772 : _GEN_2771; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5845 = 12'had5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8917 = 12'had5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5845; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11989 = 12'had5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8917; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15061 = 12'had5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11989; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18133 = 12'had5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15061; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21205 = 12'had5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18133; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24277 = 12'had5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21205; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27349 = 12'had5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24277; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2773 = io_valid_in ? _GEN_27349 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2773 = 12'had5 == _T_2[11:0] ? image_2773 : _GEN_2772; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5846 = 12'had6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8918 = 12'had6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5846; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11990 = 12'had6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8918; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15062 = 12'had6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11990; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18134 = 12'had6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15062; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21206 = 12'had6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18134; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24278 = 12'had6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21206; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27350 = 12'had6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24278; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2774 = io_valid_in ? _GEN_27350 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2774 = 12'had6 == _T_2[11:0] ? image_2774 : _GEN_2773; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5847 = 12'had7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8919 = 12'had7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5847; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11991 = 12'had7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8919; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15063 = 12'had7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11991; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18135 = 12'had7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15063; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21207 = 12'had7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18135; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24279 = 12'had7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21207; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27351 = 12'had7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24279; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2775 = io_valid_in ? _GEN_27351 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2775 = 12'had7 == _T_2[11:0] ? image_2775 : _GEN_2774; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5848 = 12'had8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8920 = 12'had8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5848; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11992 = 12'had8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8920; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15064 = 12'had8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11992; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18136 = 12'had8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15064; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21208 = 12'had8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18136; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24280 = 12'had8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21208; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27352 = 12'had8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24280; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2776 = io_valid_in ? _GEN_27352 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2776 = 12'had8 == _T_2[11:0] ? image_2776 : _GEN_2775; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5849 = 12'had9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8921 = 12'had9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5849; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11993 = 12'had9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8921; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15065 = 12'had9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11993; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18137 = 12'had9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15065; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21209 = 12'had9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18137; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24281 = 12'had9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21209; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27353 = 12'had9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24281; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2777 = io_valid_in ? _GEN_27353 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2777 = 12'had9 == _T_2[11:0] ? image_2777 : _GEN_2776; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5850 = 12'hada == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8922 = 12'hada == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5850; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11994 = 12'hada == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8922; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15066 = 12'hada == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11994; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18138 = 12'hada == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15066; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21210 = 12'hada == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18138; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24282 = 12'hada == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21210; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27354 = 12'hada == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24282; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2778 = io_valid_in ? _GEN_27354 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2778 = 12'hada == _T_2[11:0] ? image_2778 : _GEN_2777; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5851 = 12'hadb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8923 = 12'hadb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5851; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11995 = 12'hadb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8923; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15067 = 12'hadb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11995; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18139 = 12'hadb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15067; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21211 = 12'hadb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18139; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24283 = 12'hadb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21211; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27355 = 12'hadb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24283; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2779 = io_valid_in ? _GEN_27355 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2779 = 12'hadb == _T_2[11:0] ? image_2779 : _GEN_2778; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5852 = 12'hadc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8924 = 12'hadc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5852; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11996 = 12'hadc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8924; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15068 = 12'hadc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11996; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18140 = 12'hadc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15068; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21212 = 12'hadc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18140; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24284 = 12'hadc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21212; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27356 = 12'hadc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24284; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2780 = io_valid_in ? _GEN_27356 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2780 = 12'hadc == _T_2[11:0] ? image_2780 : _GEN_2779; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5853 = 12'hadd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8925 = 12'hadd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5853; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11997 = 12'hadd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8925; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15069 = 12'hadd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11997; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18141 = 12'hadd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15069; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21213 = 12'hadd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18141; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24285 = 12'hadd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21213; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27357 = 12'hadd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24285; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2781 = io_valid_in ? _GEN_27357 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2781 = 12'hadd == _T_2[11:0] ? image_2781 : _GEN_2780; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5854 = 12'hade == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8926 = 12'hade == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5854; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11998 = 12'hade == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8926; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15070 = 12'hade == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11998; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18142 = 12'hade == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15070; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21214 = 12'hade == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18142; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24286 = 12'hade == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21214; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27358 = 12'hade == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24286; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2782 = io_valid_in ? _GEN_27358 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2782 = 12'hade == _T_2[11:0] ? image_2782 : _GEN_2781; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5855 = 12'hadf == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8927 = 12'hadf == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5855; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_11999 = 12'hadf == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8927; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15071 = 12'hadf == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_11999; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18143 = 12'hadf == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15071; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21215 = 12'hadf == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18143; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24287 = 12'hadf == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21215; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27359 = 12'hadf == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24287; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2783 = io_valid_in ? _GEN_27359 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2783 = 12'hadf == _T_2[11:0] ? image_2783 : _GEN_2782; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5856 = 12'hae0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8928 = 12'hae0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5856; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12000 = 12'hae0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8928; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15072 = 12'hae0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12000; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18144 = 12'hae0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15072; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21216 = 12'hae0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18144; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24288 = 12'hae0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21216; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27360 = 12'hae0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24288; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2784 = io_valid_in ? _GEN_27360 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2784 = 12'hae0 == _T_2[11:0] ? image_2784 : _GEN_2783; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5857 = 12'hae1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8929 = 12'hae1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5857; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12001 = 12'hae1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8929; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15073 = 12'hae1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12001; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18145 = 12'hae1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15073; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21217 = 12'hae1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18145; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24289 = 12'hae1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21217; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27361 = 12'hae1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24289; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2785 = io_valid_in ? _GEN_27361 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2785 = 12'hae1 == _T_2[11:0] ? image_2785 : _GEN_2784; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5858 = 12'hae2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8930 = 12'hae2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5858; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12002 = 12'hae2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8930; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15074 = 12'hae2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12002; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18146 = 12'hae2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15074; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21218 = 12'hae2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18146; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24290 = 12'hae2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21218; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27362 = 12'hae2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24290; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2786 = io_valid_in ? _GEN_27362 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2786 = 12'hae2 == _T_2[11:0] ? image_2786 : _GEN_2785; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5859 = 12'hae3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8931 = 12'hae3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5859; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12003 = 12'hae3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8931; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15075 = 12'hae3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12003; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18147 = 12'hae3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15075; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21219 = 12'hae3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18147; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24291 = 12'hae3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21219; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27363 = 12'hae3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24291; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2787 = io_valid_in ? _GEN_27363 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2787 = 12'hae3 == _T_2[11:0] ? image_2787 : _GEN_2786; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5860 = 12'hae4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8932 = 12'hae4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5860; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12004 = 12'hae4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8932; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15076 = 12'hae4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12004; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18148 = 12'hae4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15076; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21220 = 12'hae4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18148; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24292 = 12'hae4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21220; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27364 = 12'hae4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24292; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2788 = io_valid_in ? _GEN_27364 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2788 = 12'hae4 == _T_2[11:0] ? image_2788 : _GEN_2787; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5861 = 12'hae5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8933 = 12'hae5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5861; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12005 = 12'hae5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8933; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15077 = 12'hae5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12005; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18149 = 12'hae5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15077; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21221 = 12'hae5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18149; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24293 = 12'hae5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21221; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27365 = 12'hae5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24293; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2789 = io_valid_in ? _GEN_27365 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2789 = 12'hae5 == _T_2[11:0] ? image_2789 : _GEN_2788; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5862 = 12'hae6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8934 = 12'hae6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5862; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12006 = 12'hae6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8934; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15078 = 12'hae6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12006; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18150 = 12'hae6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15078; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21222 = 12'hae6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18150; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24294 = 12'hae6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21222; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27366 = 12'hae6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24294; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2790 = io_valid_in ? _GEN_27366 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2790 = 12'hae6 == _T_2[11:0] ? image_2790 : _GEN_2789; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5863 = 12'hae7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8935 = 12'hae7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5863; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12007 = 12'hae7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8935; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15079 = 12'hae7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12007; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18151 = 12'hae7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15079; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21223 = 12'hae7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18151; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24295 = 12'hae7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21223; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27367 = 12'hae7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24295; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2791 = io_valid_in ? _GEN_27367 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2791 = 12'hae7 == _T_2[11:0] ? image_2791 : _GEN_2790; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5864 = 12'hae8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8936 = 12'hae8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5864; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12008 = 12'hae8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8936; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15080 = 12'hae8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12008; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18152 = 12'hae8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15080; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21224 = 12'hae8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18152; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24296 = 12'hae8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21224; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27368 = 12'hae8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24296; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2792 = io_valid_in ? _GEN_27368 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2792 = 12'hae8 == _T_2[11:0] ? image_2792 : _GEN_2791; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5865 = 12'hae9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8937 = 12'hae9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5865; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12009 = 12'hae9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8937; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15081 = 12'hae9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12009; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18153 = 12'hae9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15081; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21225 = 12'hae9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18153; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24297 = 12'hae9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21225; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27369 = 12'hae9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24297; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2793 = io_valid_in ? _GEN_27369 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2793 = 12'hae9 == _T_2[11:0] ? image_2793 : _GEN_2792; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5866 = 12'haea == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8938 = 12'haea == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5866; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12010 = 12'haea == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8938; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15082 = 12'haea == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12010; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18154 = 12'haea == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15082; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21226 = 12'haea == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18154; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24298 = 12'haea == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21226; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27370 = 12'haea == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24298; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2794 = io_valid_in ? _GEN_27370 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2794 = 12'haea == _T_2[11:0] ? image_2794 : _GEN_2793; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5867 = 12'haeb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8939 = 12'haeb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5867; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12011 = 12'haeb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8939; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15083 = 12'haeb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12011; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18155 = 12'haeb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15083; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21227 = 12'haeb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18155; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24299 = 12'haeb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21227; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27371 = 12'haeb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24299; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2795 = io_valid_in ? _GEN_27371 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2795 = 12'haeb == _T_2[11:0] ? image_2795 : _GEN_2794; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5868 = 12'haec == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8940 = 12'haec == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5868; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12012 = 12'haec == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8940; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15084 = 12'haec == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12012; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18156 = 12'haec == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15084; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21228 = 12'haec == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18156; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24300 = 12'haec == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21228; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27372 = 12'haec == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24300; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2796 = io_valid_in ? _GEN_27372 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2796 = 12'haec == _T_2[11:0] ? image_2796 : _GEN_2795; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5869 = 12'haed == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8941 = 12'haed == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5869; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12013 = 12'haed == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8941; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15085 = 12'haed == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12013; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18157 = 12'haed == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15085; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21229 = 12'haed == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18157; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24301 = 12'haed == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21229; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27373 = 12'haed == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24301; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2797 = io_valid_in ? _GEN_27373 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2797 = 12'haed == _T_2[11:0] ? image_2797 : _GEN_2796; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5870 = 12'haee == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8942 = 12'haee == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5870; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12014 = 12'haee == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8942; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15086 = 12'haee == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12014; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18158 = 12'haee == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15086; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21230 = 12'haee == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18158; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24302 = 12'haee == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21230; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27374 = 12'haee == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24302; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2798 = io_valid_in ? _GEN_27374 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2798 = 12'haee == _T_2[11:0] ? image_2798 : _GEN_2797; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5871 = 12'haef == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8943 = 12'haef == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5871; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12015 = 12'haef == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8943; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15087 = 12'haef == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12015; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18159 = 12'haef == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15087; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21231 = 12'haef == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18159; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24303 = 12'haef == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21231; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27375 = 12'haef == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24303; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2799 = io_valid_in ? _GEN_27375 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2799 = 12'haef == _T_2[11:0] ? image_2799 : _GEN_2798; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5872 = 12'haf0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8944 = 12'haf0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5872; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12016 = 12'haf0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8944; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15088 = 12'haf0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12016; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18160 = 12'haf0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15088; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21232 = 12'haf0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18160; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24304 = 12'haf0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21232; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27376 = 12'haf0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24304; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2800 = io_valid_in ? _GEN_27376 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2800 = 12'haf0 == _T_2[11:0] ? image_2800 : _GEN_2799; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5873 = 12'haf1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8945 = 12'haf1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5873; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12017 = 12'haf1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8945; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15089 = 12'haf1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12017; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18161 = 12'haf1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15089; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21233 = 12'haf1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18161; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24305 = 12'haf1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21233; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27377 = 12'haf1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24305; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2801 = io_valid_in ? _GEN_27377 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2801 = 12'haf1 == _T_2[11:0] ? image_2801 : _GEN_2800; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5874 = 12'haf2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8946 = 12'haf2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5874; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12018 = 12'haf2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8946; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15090 = 12'haf2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12018; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18162 = 12'haf2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15090; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21234 = 12'haf2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18162; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24306 = 12'haf2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21234; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27378 = 12'haf2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24306; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2802 = io_valid_in ? _GEN_27378 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2802 = 12'haf2 == _T_2[11:0] ? image_2802 : _GEN_2801; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5875 = 12'haf3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8947 = 12'haf3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5875; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12019 = 12'haf3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8947; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15091 = 12'haf3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12019; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18163 = 12'haf3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15091; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21235 = 12'haf3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18163; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24307 = 12'haf3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21235; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27379 = 12'haf3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24307; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2803 = io_valid_in ? _GEN_27379 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2803 = 12'haf3 == _T_2[11:0] ? image_2803 : _GEN_2802; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5876 = 12'haf4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8948 = 12'haf4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5876; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12020 = 12'haf4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8948; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15092 = 12'haf4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12020; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18164 = 12'haf4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15092; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21236 = 12'haf4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18164; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24308 = 12'haf4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21236; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27380 = 12'haf4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24308; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2804 = io_valid_in ? _GEN_27380 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2804 = 12'haf4 == _T_2[11:0] ? image_2804 : _GEN_2803; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5877 = 12'haf5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8949 = 12'haf5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5877; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12021 = 12'haf5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8949; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15093 = 12'haf5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12021; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18165 = 12'haf5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15093; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21237 = 12'haf5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18165; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24309 = 12'haf5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21237; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27381 = 12'haf5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24309; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2805 = io_valid_in ? _GEN_27381 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2805 = 12'haf5 == _T_2[11:0] ? image_2805 : _GEN_2804; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5878 = 12'haf6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8950 = 12'haf6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5878; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12022 = 12'haf6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8950; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15094 = 12'haf6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12022; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18166 = 12'haf6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15094; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21238 = 12'haf6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18166; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24310 = 12'haf6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21238; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27382 = 12'haf6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24310; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2806 = io_valid_in ? _GEN_27382 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2806 = 12'haf6 == _T_2[11:0] ? image_2806 : _GEN_2805; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5879 = 12'haf7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8951 = 12'haf7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5879; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12023 = 12'haf7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8951; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15095 = 12'haf7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12023; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18167 = 12'haf7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15095; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21239 = 12'haf7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18167; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24311 = 12'haf7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21239; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27383 = 12'haf7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24311; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2807 = io_valid_in ? _GEN_27383 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2807 = 12'haf7 == _T_2[11:0] ? image_2807 : _GEN_2806; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5880 = 12'haf8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8952 = 12'haf8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5880; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12024 = 12'haf8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8952; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15096 = 12'haf8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12024; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18168 = 12'haf8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15096; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21240 = 12'haf8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18168; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24312 = 12'haf8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21240; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27384 = 12'haf8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24312; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2808 = io_valid_in ? _GEN_27384 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2808 = 12'haf8 == _T_2[11:0] ? image_2808 : _GEN_2807; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5881 = 12'haf9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8953 = 12'haf9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5881; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12025 = 12'haf9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8953; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15097 = 12'haf9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12025; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18169 = 12'haf9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15097; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21241 = 12'haf9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18169; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24313 = 12'haf9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21241; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27385 = 12'haf9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24313; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2809 = io_valid_in ? _GEN_27385 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2809 = 12'haf9 == _T_2[11:0] ? image_2809 : _GEN_2808; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5882 = 12'hafa == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8954 = 12'hafa == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5882; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12026 = 12'hafa == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8954; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15098 = 12'hafa == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12026; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18170 = 12'hafa == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15098; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21242 = 12'hafa == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18170; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24314 = 12'hafa == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21242; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27386 = 12'hafa == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24314; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2810 = io_valid_in ? _GEN_27386 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2810 = 12'hafa == _T_2[11:0] ? image_2810 : _GEN_2809; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5883 = 12'hafb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8955 = 12'hafb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5883; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12027 = 12'hafb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8955; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15099 = 12'hafb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12027; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18171 = 12'hafb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15099; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21243 = 12'hafb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18171; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24315 = 12'hafb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21243; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27387 = 12'hafb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24315; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2811 = io_valid_in ? _GEN_27387 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2811 = 12'hafb == _T_2[11:0] ? image_2811 : _GEN_2810; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5884 = 12'hafc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8956 = 12'hafc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5884; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12028 = 12'hafc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8956; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15100 = 12'hafc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12028; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18172 = 12'hafc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15100; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21244 = 12'hafc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18172; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24316 = 12'hafc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21244; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27388 = 12'hafc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24316; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2812 = io_valid_in ? _GEN_27388 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2812 = 12'hafc == _T_2[11:0] ? image_2812 : _GEN_2811; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5885 = 12'hafd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8957 = 12'hafd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5885; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12029 = 12'hafd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8957; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15101 = 12'hafd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12029; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18173 = 12'hafd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15101; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21245 = 12'hafd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18173; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24317 = 12'hafd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21245; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27389 = 12'hafd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24317; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2813 = io_valid_in ? _GEN_27389 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2813 = 12'hafd == _T_2[11:0] ? image_2813 : _GEN_2812; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5886 = 12'hafe == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8958 = 12'hafe == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5886; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12030 = 12'hafe == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8958; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15102 = 12'hafe == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12030; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18174 = 12'hafe == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15102; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21246 = 12'hafe == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18174; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24318 = 12'hafe == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21246; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27390 = 12'hafe == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24318; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2814 = io_valid_in ? _GEN_27390 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2814 = 12'hafe == _T_2[11:0] ? image_2814 : _GEN_2813; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5887 = 12'haff == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8959 = 12'haff == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5887; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12031 = 12'haff == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8959; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15103 = 12'haff == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12031; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18175 = 12'haff == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15103; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21247 = 12'haff == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18175; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24319 = 12'haff == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21247; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27391 = 12'haff == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24319; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2815 = io_valid_in ? _GEN_27391 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2815 = 12'haff == _T_2[11:0] ? image_2815 : _GEN_2814; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5888 = 12'hb00 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8960 = 12'hb00 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5888; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12032 = 12'hb00 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8960; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15104 = 12'hb00 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12032; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18176 = 12'hb00 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15104; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21248 = 12'hb00 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18176; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24320 = 12'hb00 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21248; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27392 = 12'hb00 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24320; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2816 = io_valid_in ? _GEN_27392 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2816 = 12'hb00 == _T_2[11:0] ? image_2816 : _GEN_2815; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5889 = 12'hb01 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8961 = 12'hb01 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5889; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12033 = 12'hb01 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8961; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15105 = 12'hb01 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12033; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18177 = 12'hb01 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15105; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21249 = 12'hb01 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18177; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24321 = 12'hb01 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21249; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27393 = 12'hb01 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24321; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2817 = io_valid_in ? _GEN_27393 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2817 = 12'hb01 == _T_2[11:0] ? image_2817 : _GEN_2816; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5890 = 12'hb02 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8962 = 12'hb02 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5890; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12034 = 12'hb02 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8962; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15106 = 12'hb02 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12034; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18178 = 12'hb02 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15106; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21250 = 12'hb02 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18178; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24322 = 12'hb02 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21250; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27394 = 12'hb02 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24322; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2818 = io_valid_in ? _GEN_27394 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2818 = 12'hb02 == _T_2[11:0] ? image_2818 : _GEN_2817; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5891 = 12'hb03 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8963 = 12'hb03 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5891; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12035 = 12'hb03 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8963; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15107 = 12'hb03 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12035; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18179 = 12'hb03 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15107; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21251 = 12'hb03 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18179; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24323 = 12'hb03 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21251; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27395 = 12'hb03 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24323; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2819 = io_valid_in ? _GEN_27395 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2819 = 12'hb03 == _T_2[11:0] ? image_2819 : _GEN_2818; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5892 = 12'hb04 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8964 = 12'hb04 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5892; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12036 = 12'hb04 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8964; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15108 = 12'hb04 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12036; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18180 = 12'hb04 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15108; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21252 = 12'hb04 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18180; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24324 = 12'hb04 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21252; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27396 = 12'hb04 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24324; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2820 = io_valid_in ? _GEN_27396 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2820 = 12'hb04 == _T_2[11:0] ? image_2820 : _GEN_2819; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5893 = 12'hb05 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8965 = 12'hb05 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5893; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12037 = 12'hb05 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8965; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15109 = 12'hb05 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12037; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18181 = 12'hb05 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15109; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21253 = 12'hb05 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18181; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24325 = 12'hb05 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21253; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27397 = 12'hb05 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24325; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2821 = io_valid_in ? _GEN_27397 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2821 = 12'hb05 == _T_2[11:0] ? image_2821 : _GEN_2820; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5894 = 12'hb06 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8966 = 12'hb06 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5894; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12038 = 12'hb06 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8966; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15110 = 12'hb06 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12038; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18182 = 12'hb06 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15110; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21254 = 12'hb06 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18182; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24326 = 12'hb06 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21254; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27398 = 12'hb06 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24326; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2822 = io_valid_in ? _GEN_27398 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2822 = 12'hb06 == _T_2[11:0] ? image_2822 : _GEN_2821; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5895 = 12'hb07 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8967 = 12'hb07 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5895; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12039 = 12'hb07 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8967; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15111 = 12'hb07 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12039; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18183 = 12'hb07 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15111; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21255 = 12'hb07 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18183; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24327 = 12'hb07 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21255; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27399 = 12'hb07 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24327; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2823 = io_valid_in ? _GEN_27399 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2823 = 12'hb07 == _T_2[11:0] ? image_2823 : _GEN_2822; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5896 = 12'hb08 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8968 = 12'hb08 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5896; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12040 = 12'hb08 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8968; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15112 = 12'hb08 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12040; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18184 = 12'hb08 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15112; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21256 = 12'hb08 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18184; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24328 = 12'hb08 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21256; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27400 = 12'hb08 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24328; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2824 = io_valid_in ? _GEN_27400 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2824 = 12'hb08 == _T_2[11:0] ? image_2824 : _GEN_2823; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5897 = 12'hb09 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8969 = 12'hb09 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5897; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12041 = 12'hb09 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8969; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15113 = 12'hb09 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12041; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18185 = 12'hb09 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15113; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21257 = 12'hb09 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18185; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24329 = 12'hb09 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21257; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27401 = 12'hb09 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24329; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2825 = io_valid_in ? _GEN_27401 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2825 = 12'hb09 == _T_2[11:0] ? image_2825 : _GEN_2824; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5898 = 12'hb0a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8970 = 12'hb0a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5898; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12042 = 12'hb0a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8970; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15114 = 12'hb0a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12042; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18186 = 12'hb0a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15114; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21258 = 12'hb0a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18186; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24330 = 12'hb0a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21258; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27402 = 12'hb0a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24330; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2826 = io_valid_in ? _GEN_27402 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2826 = 12'hb0a == _T_2[11:0] ? image_2826 : _GEN_2825; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5899 = 12'hb0b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8971 = 12'hb0b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5899; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12043 = 12'hb0b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8971; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15115 = 12'hb0b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12043; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18187 = 12'hb0b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15115; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21259 = 12'hb0b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18187; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24331 = 12'hb0b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21259; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27403 = 12'hb0b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24331; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2827 = io_valid_in ? _GEN_27403 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2827 = 12'hb0b == _T_2[11:0] ? image_2827 : _GEN_2826; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5900 = 12'hb0c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8972 = 12'hb0c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5900; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12044 = 12'hb0c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8972; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15116 = 12'hb0c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12044; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18188 = 12'hb0c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15116; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21260 = 12'hb0c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18188; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24332 = 12'hb0c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21260; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27404 = 12'hb0c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24332; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2828 = io_valid_in ? _GEN_27404 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2828 = 12'hb0c == _T_2[11:0] ? image_2828 : _GEN_2827; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5901 = 12'hb0d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8973 = 12'hb0d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5901; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12045 = 12'hb0d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8973; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15117 = 12'hb0d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12045; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18189 = 12'hb0d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15117; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21261 = 12'hb0d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18189; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24333 = 12'hb0d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21261; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27405 = 12'hb0d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24333; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2829 = io_valid_in ? _GEN_27405 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2829 = 12'hb0d == _T_2[11:0] ? image_2829 : _GEN_2828; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5902 = 12'hb0e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8974 = 12'hb0e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5902; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12046 = 12'hb0e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8974; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15118 = 12'hb0e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12046; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18190 = 12'hb0e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15118; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21262 = 12'hb0e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18190; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24334 = 12'hb0e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21262; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27406 = 12'hb0e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24334; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2830 = io_valid_in ? _GEN_27406 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2830 = 12'hb0e == _T_2[11:0] ? image_2830 : _GEN_2829; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5903 = 12'hb0f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8975 = 12'hb0f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5903; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12047 = 12'hb0f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8975; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15119 = 12'hb0f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12047; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18191 = 12'hb0f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15119; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21263 = 12'hb0f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18191; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24335 = 12'hb0f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21263; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27407 = 12'hb0f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24335; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2831 = io_valid_in ? _GEN_27407 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2831 = 12'hb0f == _T_2[11:0] ? image_2831 : _GEN_2830; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5904 = 12'hb10 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8976 = 12'hb10 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5904; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12048 = 12'hb10 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8976; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15120 = 12'hb10 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12048; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18192 = 12'hb10 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15120; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21264 = 12'hb10 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18192; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24336 = 12'hb10 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21264; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27408 = 12'hb10 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24336; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2832 = io_valid_in ? _GEN_27408 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2832 = 12'hb10 == _T_2[11:0] ? image_2832 : _GEN_2831; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5905 = 12'hb11 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8977 = 12'hb11 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5905; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12049 = 12'hb11 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8977; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15121 = 12'hb11 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12049; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18193 = 12'hb11 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15121; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21265 = 12'hb11 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18193; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24337 = 12'hb11 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21265; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27409 = 12'hb11 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24337; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2833 = io_valid_in ? _GEN_27409 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2833 = 12'hb11 == _T_2[11:0] ? image_2833 : _GEN_2832; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5906 = 12'hb12 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8978 = 12'hb12 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5906; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12050 = 12'hb12 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8978; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15122 = 12'hb12 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12050; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18194 = 12'hb12 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15122; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21266 = 12'hb12 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18194; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24338 = 12'hb12 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21266; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27410 = 12'hb12 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24338; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2834 = io_valid_in ? _GEN_27410 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2834 = 12'hb12 == _T_2[11:0] ? image_2834 : _GEN_2833; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5907 = 12'hb13 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8979 = 12'hb13 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5907; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12051 = 12'hb13 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8979; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15123 = 12'hb13 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12051; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18195 = 12'hb13 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15123; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21267 = 12'hb13 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18195; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24339 = 12'hb13 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21267; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27411 = 12'hb13 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24339; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2835 = io_valid_in ? _GEN_27411 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2835 = 12'hb13 == _T_2[11:0] ? image_2835 : _GEN_2834; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5908 = 12'hb14 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8980 = 12'hb14 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5908; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12052 = 12'hb14 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8980; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15124 = 12'hb14 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12052; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18196 = 12'hb14 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15124; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21268 = 12'hb14 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18196; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24340 = 12'hb14 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21268; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27412 = 12'hb14 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24340; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2836 = io_valid_in ? _GEN_27412 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2836 = 12'hb14 == _T_2[11:0] ? image_2836 : _GEN_2835; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5909 = 12'hb15 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8981 = 12'hb15 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5909; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12053 = 12'hb15 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8981; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15125 = 12'hb15 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12053; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18197 = 12'hb15 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15125; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21269 = 12'hb15 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18197; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24341 = 12'hb15 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21269; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27413 = 12'hb15 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24341; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2837 = io_valid_in ? _GEN_27413 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2837 = 12'hb15 == _T_2[11:0] ? image_2837 : _GEN_2836; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5910 = 12'hb16 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8982 = 12'hb16 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5910; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12054 = 12'hb16 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8982; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15126 = 12'hb16 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12054; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18198 = 12'hb16 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15126; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21270 = 12'hb16 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18198; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24342 = 12'hb16 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21270; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27414 = 12'hb16 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24342; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2838 = io_valid_in ? _GEN_27414 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2838 = 12'hb16 == _T_2[11:0] ? image_2838 : _GEN_2837; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5911 = 12'hb17 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8983 = 12'hb17 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5911; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12055 = 12'hb17 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8983; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15127 = 12'hb17 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12055; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18199 = 12'hb17 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15127; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21271 = 12'hb17 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18199; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24343 = 12'hb17 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21271; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27415 = 12'hb17 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24343; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2839 = io_valid_in ? _GEN_27415 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2839 = 12'hb17 == _T_2[11:0] ? image_2839 : _GEN_2838; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5912 = 12'hb18 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8984 = 12'hb18 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5912; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12056 = 12'hb18 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8984; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15128 = 12'hb18 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12056; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18200 = 12'hb18 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15128; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21272 = 12'hb18 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18200; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24344 = 12'hb18 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21272; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27416 = 12'hb18 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24344; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2840 = io_valid_in ? _GEN_27416 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2840 = 12'hb18 == _T_2[11:0] ? image_2840 : _GEN_2839; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5913 = 12'hb19 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8985 = 12'hb19 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5913; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12057 = 12'hb19 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8985; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15129 = 12'hb19 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12057; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18201 = 12'hb19 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15129; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21273 = 12'hb19 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18201; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24345 = 12'hb19 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21273; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27417 = 12'hb19 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24345; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2841 = io_valid_in ? _GEN_27417 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2841 = 12'hb19 == _T_2[11:0] ? image_2841 : _GEN_2840; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5914 = 12'hb1a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8986 = 12'hb1a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5914; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12058 = 12'hb1a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8986; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15130 = 12'hb1a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12058; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18202 = 12'hb1a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15130; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21274 = 12'hb1a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18202; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24346 = 12'hb1a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21274; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27418 = 12'hb1a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24346; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2842 = io_valid_in ? _GEN_27418 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2842 = 12'hb1a == _T_2[11:0] ? image_2842 : _GEN_2841; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5915 = 12'hb1b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8987 = 12'hb1b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5915; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12059 = 12'hb1b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8987; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15131 = 12'hb1b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12059; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18203 = 12'hb1b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15131; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21275 = 12'hb1b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18203; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24347 = 12'hb1b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21275; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27419 = 12'hb1b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24347; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2843 = io_valid_in ? _GEN_27419 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2843 = 12'hb1b == _T_2[11:0] ? image_2843 : _GEN_2842; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5916 = 12'hb1c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8988 = 12'hb1c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5916; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12060 = 12'hb1c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8988; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15132 = 12'hb1c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12060; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18204 = 12'hb1c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15132; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21276 = 12'hb1c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18204; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24348 = 12'hb1c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21276; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27420 = 12'hb1c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24348; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2844 = io_valid_in ? _GEN_27420 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2844 = 12'hb1c == _T_2[11:0] ? image_2844 : _GEN_2843; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5917 = 12'hb1d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8989 = 12'hb1d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5917; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12061 = 12'hb1d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8989; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15133 = 12'hb1d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12061; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18205 = 12'hb1d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15133; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21277 = 12'hb1d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18205; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24349 = 12'hb1d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21277; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27421 = 12'hb1d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24349; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2845 = io_valid_in ? _GEN_27421 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2845 = 12'hb1d == _T_2[11:0] ? image_2845 : _GEN_2844; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5918 = 12'hb1e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8990 = 12'hb1e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5918; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12062 = 12'hb1e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8990; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15134 = 12'hb1e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12062; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18206 = 12'hb1e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15134; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21278 = 12'hb1e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18206; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24350 = 12'hb1e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21278; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27422 = 12'hb1e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24350; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2846 = io_valid_in ? _GEN_27422 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2846 = 12'hb1e == _T_2[11:0] ? image_2846 : _GEN_2845; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5919 = 12'hb1f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8991 = 12'hb1f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5919; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12063 = 12'hb1f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8991; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15135 = 12'hb1f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12063; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18207 = 12'hb1f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15135; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21279 = 12'hb1f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18207; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24351 = 12'hb1f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21279; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27423 = 12'hb1f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24351; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2847 = io_valid_in ? _GEN_27423 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2847 = 12'hb1f == _T_2[11:0] ? image_2847 : _GEN_2846; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5920 = 12'hb20 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8992 = 12'hb20 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5920; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12064 = 12'hb20 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8992; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15136 = 12'hb20 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12064; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18208 = 12'hb20 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15136; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21280 = 12'hb20 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18208; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24352 = 12'hb20 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21280; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27424 = 12'hb20 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24352; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2848 = io_valid_in ? _GEN_27424 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2848 = 12'hb20 == _T_2[11:0] ? image_2848 : _GEN_2847; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5921 = 12'hb21 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8993 = 12'hb21 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5921; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12065 = 12'hb21 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8993; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15137 = 12'hb21 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12065; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18209 = 12'hb21 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15137; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21281 = 12'hb21 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18209; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24353 = 12'hb21 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21281; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27425 = 12'hb21 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24353; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2849 = io_valid_in ? _GEN_27425 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2849 = 12'hb21 == _T_2[11:0] ? image_2849 : _GEN_2848; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5922 = 12'hb22 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8994 = 12'hb22 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5922; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12066 = 12'hb22 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8994; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15138 = 12'hb22 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12066; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18210 = 12'hb22 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15138; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21282 = 12'hb22 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18210; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24354 = 12'hb22 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21282; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27426 = 12'hb22 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24354; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2850 = io_valid_in ? _GEN_27426 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2850 = 12'hb22 == _T_2[11:0] ? image_2850 : _GEN_2849; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5923 = 12'hb23 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8995 = 12'hb23 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5923; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12067 = 12'hb23 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8995; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15139 = 12'hb23 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12067; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18211 = 12'hb23 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15139; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21283 = 12'hb23 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18211; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24355 = 12'hb23 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21283; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27427 = 12'hb23 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24355; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2851 = io_valid_in ? _GEN_27427 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2851 = 12'hb23 == _T_2[11:0] ? image_2851 : _GEN_2850; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5924 = 12'hb24 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8996 = 12'hb24 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5924; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12068 = 12'hb24 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8996; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15140 = 12'hb24 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12068; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18212 = 12'hb24 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15140; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21284 = 12'hb24 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18212; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24356 = 12'hb24 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21284; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27428 = 12'hb24 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24356; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2852 = io_valid_in ? _GEN_27428 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2852 = 12'hb24 == _T_2[11:0] ? image_2852 : _GEN_2851; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5925 = 12'hb25 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8997 = 12'hb25 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5925; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12069 = 12'hb25 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8997; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15141 = 12'hb25 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12069; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18213 = 12'hb25 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15141; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21285 = 12'hb25 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18213; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24357 = 12'hb25 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21285; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27429 = 12'hb25 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24357; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2853 = io_valid_in ? _GEN_27429 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2853 = 12'hb25 == _T_2[11:0] ? image_2853 : _GEN_2852; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5926 = 12'hb26 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8998 = 12'hb26 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5926; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12070 = 12'hb26 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8998; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15142 = 12'hb26 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12070; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18214 = 12'hb26 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15142; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21286 = 12'hb26 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18214; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24358 = 12'hb26 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21286; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27430 = 12'hb26 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24358; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2854 = io_valid_in ? _GEN_27430 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2854 = 12'hb26 == _T_2[11:0] ? image_2854 : _GEN_2853; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5927 = 12'hb27 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_8999 = 12'hb27 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5927; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12071 = 12'hb27 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_8999; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15143 = 12'hb27 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12071; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18215 = 12'hb27 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15143; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21287 = 12'hb27 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18215; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24359 = 12'hb27 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21287; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27431 = 12'hb27 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24359; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2855 = io_valid_in ? _GEN_27431 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2855 = 12'hb27 == _T_2[11:0] ? image_2855 : _GEN_2854; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5928 = 12'hb28 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9000 = 12'hb28 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5928; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12072 = 12'hb28 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9000; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15144 = 12'hb28 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12072; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18216 = 12'hb28 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15144; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21288 = 12'hb28 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18216; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24360 = 12'hb28 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21288; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27432 = 12'hb28 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24360; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2856 = io_valid_in ? _GEN_27432 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2856 = 12'hb28 == _T_2[11:0] ? image_2856 : _GEN_2855; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5929 = 12'hb29 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9001 = 12'hb29 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5929; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12073 = 12'hb29 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9001; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15145 = 12'hb29 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12073; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18217 = 12'hb29 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15145; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21289 = 12'hb29 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18217; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24361 = 12'hb29 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21289; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27433 = 12'hb29 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24361; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2857 = io_valid_in ? _GEN_27433 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2857 = 12'hb29 == _T_2[11:0] ? image_2857 : _GEN_2856; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5930 = 12'hb2a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9002 = 12'hb2a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5930; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12074 = 12'hb2a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9002; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15146 = 12'hb2a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12074; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18218 = 12'hb2a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15146; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21290 = 12'hb2a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18218; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24362 = 12'hb2a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21290; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27434 = 12'hb2a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24362; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2858 = io_valid_in ? _GEN_27434 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2858 = 12'hb2a == _T_2[11:0] ? image_2858 : _GEN_2857; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5931 = 12'hb2b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9003 = 12'hb2b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5931; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12075 = 12'hb2b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9003; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15147 = 12'hb2b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12075; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18219 = 12'hb2b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15147; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21291 = 12'hb2b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18219; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24363 = 12'hb2b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21291; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27435 = 12'hb2b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24363; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2859 = io_valid_in ? _GEN_27435 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2859 = 12'hb2b == _T_2[11:0] ? image_2859 : _GEN_2858; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5932 = 12'hb2c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9004 = 12'hb2c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5932; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12076 = 12'hb2c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9004; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15148 = 12'hb2c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12076; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18220 = 12'hb2c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15148; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21292 = 12'hb2c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18220; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24364 = 12'hb2c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21292; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27436 = 12'hb2c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24364; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2860 = io_valid_in ? _GEN_27436 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2860 = 12'hb2c == _T_2[11:0] ? image_2860 : _GEN_2859; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5933 = 12'hb2d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9005 = 12'hb2d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5933; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12077 = 12'hb2d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9005; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15149 = 12'hb2d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12077; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18221 = 12'hb2d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15149; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21293 = 12'hb2d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18221; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24365 = 12'hb2d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21293; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27437 = 12'hb2d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24365; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2861 = io_valid_in ? _GEN_27437 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2861 = 12'hb2d == _T_2[11:0] ? image_2861 : _GEN_2860; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5934 = 12'hb2e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9006 = 12'hb2e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5934; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12078 = 12'hb2e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9006; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15150 = 12'hb2e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12078; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18222 = 12'hb2e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15150; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21294 = 12'hb2e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18222; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24366 = 12'hb2e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21294; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27438 = 12'hb2e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24366; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2862 = io_valid_in ? _GEN_27438 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2862 = 12'hb2e == _T_2[11:0] ? image_2862 : _GEN_2861; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5935 = 12'hb2f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9007 = 12'hb2f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5935; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12079 = 12'hb2f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9007; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15151 = 12'hb2f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12079; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18223 = 12'hb2f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15151; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21295 = 12'hb2f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18223; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24367 = 12'hb2f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21295; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27439 = 12'hb2f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24367; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2863 = io_valid_in ? _GEN_27439 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2863 = 12'hb2f == _T_2[11:0] ? image_2863 : _GEN_2862; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5936 = 12'hb30 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9008 = 12'hb30 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5936; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12080 = 12'hb30 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9008; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15152 = 12'hb30 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12080; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18224 = 12'hb30 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15152; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21296 = 12'hb30 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18224; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24368 = 12'hb30 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21296; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27440 = 12'hb30 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24368; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2864 = io_valid_in ? _GEN_27440 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2864 = 12'hb30 == _T_2[11:0] ? image_2864 : _GEN_2863; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5937 = 12'hb31 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9009 = 12'hb31 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5937; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12081 = 12'hb31 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9009; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15153 = 12'hb31 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12081; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18225 = 12'hb31 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15153; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21297 = 12'hb31 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18225; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24369 = 12'hb31 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21297; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27441 = 12'hb31 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24369; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2865 = io_valid_in ? _GEN_27441 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2865 = 12'hb31 == _T_2[11:0] ? image_2865 : _GEN_2864; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5938 = 12'hb32 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9010 = 12'hb32 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5938; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12082 = 12'hb32 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9010; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15154 = 12'hb32 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12082; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18226 = 12'hb32 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15154; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21298 = 12'hb32 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18226; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24370 = 12'hb32 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21298; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27442 = 12'hb32 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24370; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2866 = io_valid_in ? _GEN_27442 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2866 = 12'hb32 == _T_2[11:0] ? image_2866 : _GEN_2865; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5939 = 12'hb33 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9011 = 12'hb33 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5939; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12083 = 12'hb33 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9011; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15155 = 12'hb33 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12083; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18227 = 12'hb33 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15155; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21299 = 12'hb33 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18227; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24371 = 12'hb33 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21299; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27443 = 12'hb33 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24371; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2867 = io_valid_in ? _GEN_27443 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2867 = 12'hb33 == _T_2[11:0] ? image_2867 : _GEN_2866; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5940 = 12'hb34 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9012 = 12'hb34 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5940; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12084 = 12'hb34 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9012; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15156 = 12'hb34 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12084; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18228 = 12'hb34 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15156; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21300 = 12'hb34 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18228; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24372 = 12'hb34 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21300; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27444 = 12'hb34 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24372; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2868 = io_valid_in ? _GEN_27444 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2868 = 12'hb34 == _T_2[11:0] ? image_2868 : _GEN_2867; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5941 = 12'hb35 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9013 = 12'hb35 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5941; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12085 = 12'hb35 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9013; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15157 = 12'hb35 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12085; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18229 = 12'hb35 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15157; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21301 = 12'hb35 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18229; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24373 = 12'hb35 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21301; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27445 = 12'hb35 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24373; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2869 = io_valid_in ? _GEN_27445 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2869 = 12'hb35 == _T_2[11:0] ? image_2869 : _GEN_2868; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5942 = 12'hb36 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9014 = 12'hb36 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5942; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12086 = 12'hb36 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9014; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15158 = 12'hb36 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12086; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18230 = 12'hb36 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15158; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21302 = 12'hb36 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18230; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24374 = 12'hb36 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21302; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27446 = 12'hb36 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24374; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2870 = io_valid_in ? _GEN_27446 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2870 = 12'hb36 == _T_2[11:0] ? image_2870 : _GEN_2869; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5943 = 12'hb37 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9015 = 12'hb37 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5943; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12087 = 12'hb37 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9015; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15159 = 12'hb37 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12087; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18231 = 12'hb37 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15159; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21303 = 12'hb37 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18231; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24375 = 12'hb37 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21303; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27447 = 12'hb37 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24375; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2871 = io_valid_in ? _GEN_27447 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2871 = 12'hb37 == _T_2[11:0] ? image_2871 : _GEN_2870; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5944 = 12'hb38 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9016 = 12'hb38 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5944; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12088 = 12'hb38 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9016; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15160 = 12'hb38 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12088; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18232 = 12'hb38 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15160; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21304 = 12'hb38 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18232; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24376 = 12'hb38 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21304; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27448 = 12'hb38 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24376; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2872 = io_valid_in ? _GEN_27448 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2872 = 12'hb38 == _T_2[11:0] ? image_2872 : _GEN_2871; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5945 = 12'hb39 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9017 = 12'hb39 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5945; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12089 = 12'hb39 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9017; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15161 = 12'hb39 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12089; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18233 = 12'hb39 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15161; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21305 = 12'hb39 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18233; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24377 = 12'hb39 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21305; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27449 = 12'hb39 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24377; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2873 = io_valid_in ? _GEN_27449 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2873 = 12'hb39 == _T_2[11:0] ? image_2873 : _GEN_2872; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5946 = 12'hb3a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9018 = 12'hb3a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5946; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12090 = 12'hb3a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9018; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15162 = 12'hb3a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12090; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18234 = 12'hb3a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15162; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21306 = 12'hb3a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18234; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24378 = 12'hb3a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21306; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27450 = 12'hb3a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24378; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2874 = io_valid_in ? _GEN_27450 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2874 = 12'hb3a == _T_2[11:0] ? image_2874 : _GEN_2873; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5947 = 12'hb3b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9019 = 12'hb3b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5947; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12091 = 12'hb3b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9019; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15163 = 12'hb3b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12091; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18235 = 12'hb3b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15163; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21307 = 12'hb3b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18235; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24379 = 12'hb3b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21307; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27451 = 12'hb3b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24379; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2875 = io_valid_in ? _GEN_27451 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2875 = 12'hb3b == _T_2[11:0] ? image_2875 : _GEN_2874; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5948 = 12'hb3c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9020 = 12'hb3c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5948; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12092 = 12'hb3c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9020; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15164 = 12'hb3c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12092; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18236 = 12'hb3c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15164; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21308 = 12'hb3c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18236; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24380 = 12'hb3c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21308; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27452 = 12'hb3c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24380; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2876 = io_valid_in ? _GEN_27452 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2876 = 12'hb3c == _T_2[11:0] ? image_2876 : _GEN_2875; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5949 = 12'hb3d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9021 = 12'hb3d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5949; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12093 = 12'hb3d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9021; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15165 = 12'hb3d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12093; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18237 = 12'hb3d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15165; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21309 = 12'hb3d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18237; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24381 = 12'hb3d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21309; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27453 = 12'hb3d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24381; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2877 = io_valid_in ? _GEN_27453 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2877 = 12'hb3d == _T_2[11:0] ? image_2877 : _GEN_2876; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5950 = 12'hb3e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9022 = 12'hb3e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5950; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12094 = 12'hb3e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9022; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15166 = 12'hb3e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12094; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18238 = 12'hb3e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15166; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21310 = 12'hb3e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18238; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24382 = 12'hb3e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21310; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27454 = 12'hb3e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24382; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2878 = io_valid_in ? _GEN_27454 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2878 = 12'hb3e == _T_2[11:0] ? image_2878 : _GEN_2877; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5951 = 12'hb3f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9023 = 12'hb3f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5951; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12095 = 12'hb3f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9023; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15167 = 12'hb3f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12095; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18239 = 12'hb3f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15167; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21311 = 12'hb3f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18239; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24383 = 12'hb3f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21311; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27455 = 12'hb3f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24383; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2879 = io_valid_in ? _GEN_27455 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2879 = 12'hb3f == _T_2[11:0] ? image_2879 : _GEN_2878; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5952 = 12'hb40 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9024 = 12'hb40 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5952; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12096 = 12'hb40 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9024; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15168 = 12'hb40 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12096; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18240 = 12'hb40 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15168; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21312 = 12'hb40 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18240; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24384 = 12'hb40 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21312; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27456 = 12'hb40 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24384; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2880 = io_valid_in ? _GEN_27456 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2880 = 12'hb40 == _T_2[11:0] ? image_2880 : _GEN_2879; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5953 = 12'hb41 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9025 = 12'hb41 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5953; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12097 = 12'hb41 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9025; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15169 = 12'hb41 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12097; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18241 = 12'hb41 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15169; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21313 = 12'hb41 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18241; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24385 = 12'hb41 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21313; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27457 = 12'hb41 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24385; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2881 = io_valid_in ? _GEN_27457 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2881 = 12'hb41 == _T_2[11:0] ? image_2881 : _GEN_2880; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5954 = 12'hb42 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9026 = 12'hb42 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5954; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12098 = 12'hb42 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9026; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15170 = 12'hb42 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12098; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18242 = 12'hb42 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15170; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21314 = 12'hb42 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18242; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24386 = 12'hb42 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21314; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27458 = 12'hb42 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24386; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2882 = io_valid_in ? _GEN_27458 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2882 = 12'hb42 == _T_2[11:0] ? image_2882 : _GEN_2881; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5955 = 12'hb43 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9027 = 12'hb43 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5955; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12099 = 12'hb43 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9027; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15171 = 12'hb43 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12099; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18243 = 12'hb43 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15171; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21315 = 12'hb43 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18243; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24387 = 12'hb43 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21315; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27459 = 12'hb43 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24387; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2883 = io_valid_in ? _GEN_27459 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2883 = 12'hb43 == _T_2[11:0] ? image_2883 : _GEN_2882; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5956 = 12'hb44 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9028 = 12'hb44 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5956; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12100 = 12'hb44 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9028; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15172 = 12'hb44 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12100; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18244 = 12'hb44 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15172; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21316 = 12'hb44 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18244; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24388 = 12'hb44 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21316; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27460 = 12'hb44 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24388; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2884 = io_valid_in ? _GEN_27460 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2884 = 12'hb44 == _T_2[11:0] ? image_2884 : _GEN_2883; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5957 = 12'hb45 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9029 = 12'hb45 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5957; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12101 = 12'hb45 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9029; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15173 = 12'hb45 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12101; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18245 = 12'hb45 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15173; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21317 = 12'hb45 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18245; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24389 = 12'hb45 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21317; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27461 = 12'hb45 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24389; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2885 = io_valid_in ? _GEN_27461 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2885 = 12'hb45 == _T_2[11:0] ? image_2885 : _GEN_2884; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5958 = 12'hb46 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9030 = 12'hb46 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5958; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12102 = 12'hb46 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9030; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15174 = 12'hb46 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12102; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18246 = 12'hb46 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15174; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21318 = 12'hb46 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18246; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24390 = 12'hb46 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21318; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27462 = 12'hb46 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24390; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2886 = io_valid_in ? _GEN_27462 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2886 = 12'hb46 == _T_2[11:0] ? image_2886 : _GEN_2885; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5959 = 12'hb47 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9031 = 12'hb47 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5959; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12103 = 12'hb47 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9031; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15175 = 12'hb47 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12103; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18247 = 12'hb47 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15175; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21319 = 12'hb47 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18247; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24391 = 12'hb47 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21319; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27463 = 12'hb47 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24391; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2887 = io_valid_in ? _GEN_27463 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2887 = 12'hb47 == _T_2[11:0] ? image_2887 : _GEN_2886; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5960 = 12'hb48 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9032 = 12'hb48 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5960; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12104 = 12'hb48 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9032; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15176 = 12'hb48 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12104; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18248 = 12'hb48 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15176; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21320 = 12'hb48 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18248; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24392 = 12'hb48 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21320; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27464 = 12'hb48 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24392; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2888 = io_valid_in ? _GEN_27464 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2888 = 12'hb48 == _T_2[11:0] ? image_2888 : _GEN_2887; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5961 = 12'hb49 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9033 = 12'hb49 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5961; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12105 = 12'hb49 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9033; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15177 = 12'hb49 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12105; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18249 = 12'hb49 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15177; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21321 = 12'hb49 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18249; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24393 = 12'hb49 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21321; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27465 = 12'hb49 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24393; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2889 = io_valid_in ? _GEN_27465 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2889 = 12'hb49 == _T_2[11:0] ? image_2889 : _GEN_2888; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5962 = 12'hb4a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9034 = 12'hb4a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5962; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12106 = 12'hb4a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9034; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15178 = 12'hb4a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12106; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18250 = 12'hb4a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15178; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21322 = 12'hb4a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18250; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24394 = 12'hb4a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21322; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27466 = 12'hb4a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24394; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2890 = io_valid_in ? _GEN_27466 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2890 = 12'hb4a == _T_2[11:0] ? image_2890 : _GEN_2889; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5963 = 12'hb4b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9035 = 12'hb4b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5963; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12107 = 12'hb4b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9035; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15179 = 12'hb4b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12107; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18251 = 12'hb4b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15179; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21323 = 12'hb4b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18251; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24395 = 12'hb4b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21323; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27467 = 12'hb4b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24395; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2891 = io_valid_in ? _GEN_27467 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2891 = 12'hb4b == _T_2[11:0] ? image_2891 : _GEN_2890; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5964 = 12'hb4c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9036 = 12'hb4c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5964; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12108 = 12'hb4c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9036; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15180 = 12'hb4c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12108; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18252 = 12'hb4c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15180; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21324 = 12'hb4c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18252; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24396 = 12'hb4c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21324; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27468 = 12'hb4c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24396; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2892 = io_valid_in ? _GEN_27468 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2892 = 12'hb4c == _T_2[11:0] ? image_2892 : _GEN_2891; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5965 = 12'hb4d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9037 = 12'hb4d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5965; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12109 = 12'hb4d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9037; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15181 = 12'hb4d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12109; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18253 = 12'hb4d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15181; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21325 = 12'hb4d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18253; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24397 = 12'hb4d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21325; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27469 = 12'hb4d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24397; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2893 = io_valid_in ? _GEN_27469 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2893 = 12'hb4d == _T_2[11:0] ? image_2893 : _GEN_2892; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5966 = 12'hb4e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9038 = 12'hb4e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5966; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12110 = 12'hb4e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9038; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15182 = 12'hb4e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12110; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18254 = 12'hb4e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15182; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21326 = 12'hb4e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18254; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24398 = 12'hb4e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21326; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27470 = 12'hb4e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24398; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2894 = io_valid_in ? _GEN_27470 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2894 = 12'hb4e == _T_2[11:0] ? image_2894 : _GEN_2893; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5967 = 12'hb4f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9039 = 12'hb4f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5967; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12111 = 12'hb4f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9039; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15183 = 12'hb4f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12111; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18255 = 12'hb4f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15183; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21327 = 12'hb4f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18255; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24399 = 12'hb4f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21327; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27471 = 12'hb4f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24399; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2895 = io_valid_in ? _GEN_27471 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2895 = 12'hb4f == _T_2[11:0] ? image_2895 : _GEN_2894; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5968 = 12'hb50 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9040 = 12'hb50 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5968; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12112 = 12'hb50 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9040; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15184 = 12'hb50 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12112; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18256 = 12'hb50 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15184; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21328 = 12'hb50 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18256; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24400 = 12'hb50 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21328; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27472 = 12'hb50 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24400; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2896 = io_valid_in ? _GEN_27472 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2896 = 12'hb50 == _T_2[11:0] ? image_2896 : _GEN_2895; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5969 = 12'hb51 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9041 = 12'hb51 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5969; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12113 = 12'hb51 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9041; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15185 = 12'hb51 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12113; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18257 = 12'hb51 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15185; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21329 = 12'hb51 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18257; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24401 = 12'hb51 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21329; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27473 = 12'hb51 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24401; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2897 = io_valid_in ? _GEN_27473 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2897 = 12'hb51 == _T_2[11:0] ? image_2897 : _GEN_2896; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5970 = 12'hb52 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9042 = 12'hb52 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5970; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12114 = 12'hb52 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9042; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15186 = 12'hb52 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12114; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18258 = 12'hb52 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15186; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21330 = 12'hb52 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18258; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24402 = 12'hb52 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21330; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27474 = 12'hb52 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24402; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2898 = io_valid_in ? _GEN_27474 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2898 = 12'hb52 == _T_2[11:0] ? image_2898 : _GEN_2897; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5971 = 12'hb53 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9043 = 12'hb53 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5971; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12115 = 12'hb53 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9043; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15187 = 12'hb53 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12115; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18259 = 12'hb53 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15187; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21331 = 12'hb53 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18259; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24403 = 12'hb53 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21331; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27475 = 12'hb53 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24403; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2899 = io_valid_in ? _GEN_27475 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2899 = 12'hb53 == _T_2[11:0] ? image_2899 : _GEN_2898; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5972 = 12'hb54 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9044 = 12'hb54 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5972; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12116 = 12'hb54 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9044; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15188 = 12'hb54 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12116; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18260 = 12'hb54 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15188; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21332 = 12'hb54 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18260; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24404 = 12'hb54 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21332; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27476 = 12'hb54 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24404; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2900 = io_valid_in ? _GEN_27476 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2900 = 12'hb54 == _T_2[11:0] ? image_2900 : _GEN_2899; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5973 = 12'hb55 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9045 = 12'hb55 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5973; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12117 = 12'hb55 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9045; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15189 = 12'hb55 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12117; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18261 = 12'hb55 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15189; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21333 = 12'hb55 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18261; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24405 = 12'hb55 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21333; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27477 = 12'hb55 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24405; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2901 = io_valid_in ? _GEN_27477 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2901 = 12'hb55 == _T_2[11:0] ? image_2901 : _GEN_2900; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5974 = 12'hb56 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9046 = 12'hb56 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5974; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12118 = 12'hb56 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9046; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15190 = 12'hb56 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12118; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18262 = 12'hb56 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15190; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21334 = 12'hb56 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18262; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24406 = 12'hb56 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21334; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27478 = 12'hb56 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24406; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2902 = io_valid_in ? _GEN_27478 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2902 = 12'hb56 == _T_2[11:0] ? image_2902 : _GEN_2901; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5975 = 12'hb57 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9047 = 12'hb57 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5975; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12119 = 12'hb57 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9047; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15191 = 12'hb57 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12119; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18263 = 12'hb57 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15191; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21335 = 12'hb57 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18263; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24407 = 12'hb57 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21335; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27479 = 12'hb57 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24407; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2903 = io_valid_in ? _GEN_27479 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2903 = 12'hb57 == _T_2[11:0] ? image_2903 : _GEN_2902; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5976 = 12'hb58 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9048 = 12'hb58 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5976; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12120 = 12'hb58 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9048; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15192 = 12'hb58 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12120; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18264 = 12'hb58 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15192; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21336 = 12'hb58 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18264; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24408 = 12'hb58 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21336; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27480 = 12'hb58 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24408; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2904 = io_valid_in ? _GEN_27480 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2904 = 12'hb58 == _T_2[11:0] ? image_2904 : _GEN_2903; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5977 = 12'hb59 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9049 = 12'hb59 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5977; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12121 = 12'hb59 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9049; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15193 = 12'hb59 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12121; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18265 = 12'hb59 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15193; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21337 = 12'hb59 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18265; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24409 = 12'hb59 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21337; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27481 = 12'hb59 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24409; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2905 = io_valid_in ? _GEN_27481 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2905 = 12'hb59 == _T_2[11:0] ? image_2905 : _GEN_2904; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5978 = 12'hb5a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9050 = 12'hb5a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5978; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12122 = 12'hb5a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9050; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15194 = 12'hb5a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12122; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18266 = 12'hb5a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15194; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21338 = 12'hb5a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18266; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24410 = 12'hb5a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21338; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27482 = 12'hb5a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24410; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2906 = io_valid_in ? _GEN_27482 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2906 = 12'hb5a == _T_2[11:0] ? image_2906 : _GEN_2905; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5979 = 12'hb5b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9051 = 12'hb5b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5979; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12123 = 12'hb5b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9051; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15195 = 12'hb5b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12123; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18267 = 12'hb5b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15195; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21339 = 12'hb5b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18267; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24411 = 12'hb5b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21339; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27483 = 12'hb5b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24411; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2907 = io_valid_in ? _GEN_27483 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2907 = 12'hb5b == _T_2[11:0] ? image_2907 : _GEN_2906; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5980 = 12'hb5c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9052 = 12'hb5c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5980; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12124 = 12'hb5c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9052; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15196 = 12'hb5c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12124; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18268 = 12'hb5c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15196; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21340 = 12'hb5c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18268; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24412 = 12'hb5c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21340; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27484 = 12'hb5c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24412; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2908 = io_valid_in ? _GEN_27484 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2908 = 12'hb5c == _T_2[11:0] ? image_2908 : _GEN_2907; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5981 = 12'hb5d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9053 = 12'hb5d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5981; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12125 = 12'hb5d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9053; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15197 = 12'hb5d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12125; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18269 = 12'hb5d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15197; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21341 = 12'hb5d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18269; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24413 = 12'hb5d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21341; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27485 = 12'hb5d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24413; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2909 = io_valid_in ? _GEN_27485 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2909 = 12'hb5d == _T_2[11:0] ? image_2909 : _GEN_2908; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5982 = 12'hb5e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9054 = 12'hb5e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5982; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12126 = 12'hb5e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9054; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15198 = 12'hb5e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12126; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18270 = 12'hb5e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15198; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21342 = 12'hb5e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18270; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24414 = 12'hb5e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21342; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27486 = 12'hb5e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24414; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2910 = io_valid_in ? _GEN_27486 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2910 = 12'hb5e == _T_2[11:0] ? image_2910 : _GEN_2909; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5983 = 12'hb5f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9055 = 12'hb5f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5983; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12127 = 12'hb5f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9055; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15199 = 12'hb5f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12127; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18271 = 12'hb5f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15199; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21343 = 12'hb5f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18271; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24415 = 12'hb5f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21343; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27487 = 12'hb5f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24415; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2911 = io_valid_in ? _GEN_27487 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2911 = 12'hb5f == _T_2[11:0] ? image_2911 : _GEN_2910; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5984 = 12'hb60 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9056 = 12'hb60 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5984; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12128 = 12'hb60 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9056; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15200 = 12'hb60 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12128; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18272 = 12'hb60 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15200; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21344 = 12'hb60 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18272; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24416 = 12'hb60 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21344; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27488 = 12'hb60 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24416; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2912 = io_valid_in ? _GEN_27488 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2912 = 12'hb60 == _T_2[11:0] ? image_2912 : _GEN_2911; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5985 = 12'hb61 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9057 = 12'hb61 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5985; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12129 = 12'hb61 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9057; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15201 = 12'hb61 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12129; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18273 = 12'hb61 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15201; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21345 = 12'hb61 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18273; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24417 = 12'hb61 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21345; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27489 = 12'hb61 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24417; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2913 = io_valid_in ? _GEN_27489 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2913 = 12'hb61 == _T_2[11:0] ? image_2913 : _GEN_2912; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5986 = 12'hb62 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9058 = 12'hb62 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5986; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12130 = 12'hb62 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9058; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15202 = 12'hb62 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12130; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18274 = 12'hb62 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15202; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21346 = 12'hb62 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18274; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24418 = 12'hb62 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21346; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27490 = 12'hb62 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24418; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2914 = io_valid_in ? _GEN_27490 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2914 = 12'hb62 == _T_2[11:0] ? image_2914 : _GEN_2913; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5987 = 12'hb63 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9059 = 12'hb63 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5987; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12131 = 12'hb63 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9059; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15203 = 12'hb63 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12131; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18275 = 12'hb63 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15203; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21347 = 12'hb63 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18275; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24419 = 12'hb63 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21347; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27491 = 12'hb63 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24419; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2915 = io_valid_in ? _GEN_27491 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2915 = 12'hb63 == _T_2[11:0] ? image_2915 : _GEN_2914; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5988 = 12'hb64 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9060 = 12'hb64 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5988; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12132 = 12'hb64 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9060; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15204 = 12'hb64 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12132; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18276 = 12'hb64 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15204; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21348 = 12'hb64 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18276; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24420 = 12'hb64 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21348; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27492 = 12'hb64 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24420; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2916 = io_valid_in ? _GEN_27492 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2916 = 12'hb64 == _T_2[11:0] ? image_2916 : _GEN_2915; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5989 = 12'hb65 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9061 = 12'hb65 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5989; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12133 = 12'hb65 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9061; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15205 = 12'hb65 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12133; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18277 = 12'hb65 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15205; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21349 = 12'hb65 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18277; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24421 = 12'hb65 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21349; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27493 = 12'hb65 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24421; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2917 = io_valid_in ? _GEN_27493 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2917 = 12'hb65 == _T_2[11:0] ? image_2917 : _GEN_2916; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5990 = 12'hb66 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9062 = 12'hb66 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5990; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12134 = 12'hb66 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9062; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15206 = 12'hb66 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12134; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18278 = 12'hb66 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15206; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21350 = 12'hb66 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18278; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24422 = 12'hb66 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21350; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27494 = 12'hb66 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24422; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2918 = io_valid_in ? _GEN_27494 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2918 = 12'hb66 == _T_2[11:0] ? image_2918 : _GEN_2917; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5991 = 12'hb67 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9063 = 12'hb67 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5991; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12135 = 12'hb67 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9063; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15207 = 12'hb67 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12135; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18279 = 12'hb67 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15207; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21351 = 12'hb67 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18279; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24423 = 12'hb67 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21351; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27495 = 12'hb67 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24423; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2919 = io_valid_in ? _GEN_27495 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2919 = 12'hb67 == _T_2[11:0] ? image_2919 : _GEN_2918; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5992 = 12'hb68 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9064 = 12'hb68 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5992; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12136 = 12'hb68 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9064; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15208 = 12'hb68 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12136; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18280 = 12'hb68 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15208; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21352 = 12'hb68 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18280; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24424 = 12'hb68 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21352; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27496 = 12'hb68 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24424; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2920 = io_valid_in ? _GEN_27496 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2920 = 12'hb68 == _T_2[11:0] ? image_2920 : _GEN_2919; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5993 = 12'hb69 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9065 = 12'hb69 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5993; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12137 = 12'hb69 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9065; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15209 = 12'hb69 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12137; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18281 = 12'hb69 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15209; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21353 = 12'hb69 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18281; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24425 = 12'hb69 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21353; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27497 = 12'hb69 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24425; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2921 = io_valid_in ? _GEN_27497 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2921 = 12'hb69 == _T_2[11:0] ? image_2921 : _GEN_2920; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5994 = 12'hb6a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9066 = 12'hb6a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5994; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12138 = 12'hb6a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9066; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15210 = 12'hb6a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12138; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18282 = 12'hb6a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15210; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21354 = 12'hb6a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18282; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24426 = 12'hb6a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21354; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27498 = 12'hb6a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24426; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2922 = io_valid_in ? _GEN_27498 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2922 = 12'hb6a == _T_2[11:0] ? image_2922 : _GEN_2921; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5995 = 12'hb6b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9067 = 12'hb6b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5995; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12139 = 12'hb6b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9067; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15211 = 12'hb6b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12139; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18283 = 12'hb6b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15211; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21355 = 12'hb6b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18283; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24427 = 12'hb6b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21355; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27499 = 12'hb6b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24427; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2923 = io_valid_in ? _GEN_27499 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2923 = 12'hb6b == _T_2[11:0] ? image_2923 : _GEN_2922; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5996 = 12'hb6c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9068 = 12'hb6c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5996; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12140 = 12'hb6c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9068; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15212 = 12'hb6c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12140; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18284 = 12'hb6c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15212; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21356 = 12'hb6c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18284; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24428 = 12'hb6c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21356; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27500 = 12'hb6c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24428; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2924 = io_valid_in ? _GEN_27500 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2924 = 12'hb6c == _T_2[11:0] ? image_2924 : _GEN_2923; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5997 = 12'hb6d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9069 = 12'hb6d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5997; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12141 = 12'hb6d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9069; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15213 = 12'hb6d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12141; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18285 = 12'hb6d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15213; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21357 = 12'hb6d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18285; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24429 = 12'hb6d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21357; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27501 = 12'hb6d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24429; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2925 = io_valid_in ? _GEN_27501 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2925 = 12'hb6d == _T_2[11:0] ? image_2925 : _GEN_2924; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5998 = 12'hb6e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9070 = 12'hb6e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5998; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12142 = 12'hb6e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9070; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15214 = 12'hb6e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12142; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18286 = 12'hb6e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15214; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21358 = 12'hb6e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18286; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24430 = 12'hb6e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21358; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27502 = 12'hb6e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24430; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2926 = io_valid_in ? _GEN_27502 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2926 = 12'hb6e == _T_2[11:0] ? image_2926 : _GEN_2925; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_5999 = 12'hb6f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9071 = 12'hb6f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_5999; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12143 = 12'hb6f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9071; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15215 = 12'hb6f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12143; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18287 = 12'hb6f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15215; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21359 = 12'hb6f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18287; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24431 = 12'hb6f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21359; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27503 = 12'hb6f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24431; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2927 = io_valid_in ? _GEN_27503 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2927 = 12'hb6f == _T_2[11:0] ? image_2927 : _GEN_2926; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6000 = 12'hb70 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9072 = 12'hb70 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6000; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12144 = 12'hb70 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9072; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15216 = 12'hb70 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12144; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18288 = 12'hb70 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15216; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21360 = 12'hb70 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18288; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24432 = 12'hb70 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21360; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27504 = 12'hb70 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24432; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2928 = io_valid_in ? _GEN_27504 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2928 = 12'hb70 == _T_2[11:0] ? image_2928 : _GEN_2927; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6001 = 12'hb71 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9073 = 12'hb71 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6001; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12145 = 12'hb71 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9073; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15217 = 12'hb71 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12145; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18289 = 12'hb71 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15217; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21361 = 12'hb71 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18289; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24433 = 12'hb71 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21361; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27505 = 12'hb71 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24433; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2929 = io_valid_in ? _GEN_27505 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2929 = 12'hb71 == _T_2[11:0] ? image_2929 : _GEN_2928; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6002 = 12'hb72 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9074 = 12'hb72 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6002; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12146 = 12'hb72 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9074; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15218 = 12'hb72 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12146; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18290 = 12'hb72 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15218; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21362 = 12'hb72 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18290; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24434 = 12'hb72 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21362; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27506 = 12'hb72 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24434; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2930 = io_valid_in ? _GEN_27506 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2930 = 12'hb72 == _T_2[11:0] ? image_2930 : _GEN_2929; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6003 = 12'hb73 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9075 = 12'hb73 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6003; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12147 = 12'hb73 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9075; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15219 = 12'hb73 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12147; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18291 = 12'hb73 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15219; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21363 = 12'hb73 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18291; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24435 = 12'hb73 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21363; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27507 = 12'hb73 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24435; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2931 = io_valid_in ? _GEN_27507 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2931 = 12'hb73 == _T_2[11:0] ? image_2931 : _GEN_2930; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6004 = 12'hb74 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9076 = 12'hb74 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6004; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12148 = 12'hb74 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9076; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15220 = 12'hb74 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12148; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18292 = 12'hb74 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15220; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21364 = 12'hb74 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18292; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24436 = 12'hb74 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21364; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27508 = 12'hb74 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24436; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2932 = io_valid_in ? _GEN_27508 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2932 = 12'hb74 == _T_2[11:0] ? image_2932 : _GEN_2931; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6005 = 12'hb75 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9077 = 12'hb75 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6005; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12149 = 12'hb75 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9077; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15221 = 12'hb75 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12149; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18293 = 12'hb75 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15221; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21365 = 12'hb75 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18293; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24437 = 12'hb75 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21365; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27509 = 12'hb75 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24437; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2933 = io_valid_in ? _GEN_27509 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2933 = 12'hb75 == _T_2[11:0] ? image_2933 : _GEN_2932; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6006 = 12'hb76 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9078 = 12'hb76 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6006; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12150 = 12'hb76 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9078; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15222 = 12'hb76 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12150; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18294 = 12'hb76 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15222; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21366 = 12'hb76 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18294; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24438 = 12'hb76 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21366; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27510 = 12'hb76 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24438; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2934 = io_valid_in ? _GEN_27510 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2934 = 12'hb76 == _T_2[11:0] ? image_2934 : _GEN_2933; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6007 = 12'hb77 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9079 = 12'hb77 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6007; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12151 = 12'hb77 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9079; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15223 = 12'hb77 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12151; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18295 = 12'hb77 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15223; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21367 = 12'hb77 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18295; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24439 = 12'hb77 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21367; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27511 = 12'hb77 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24439; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2935 = io_valid_in ? _GEN_27511 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2935 = 12'hb77 == _T_2[11:0] ? image_2935 : _GEN_2934; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6008 = 12'hb78 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9080 = 12'hb78 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6008; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12152 = 12'hb78 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9080; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15224 = 12'hb78 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12152; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18296 = 12'hb78 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15224; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21368 = 12'hb78 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18296; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24440 = 12'hb78 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21368; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27512 = 12'hb78 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24440; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2936 = io_valid_in ? _GEN_27512 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2936 = 12'hb78 == _T_2[11:0] ? image_2936 : _GEN_2935; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6009 = 12'hb79 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9081 = 12'hb79 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6009; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12153 = 12'hb79 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9081; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15225 = 12'hb79 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12153; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18297 = 12'hb79 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15225; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21369 = 12'hb79 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18297; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24441 = 12'hb79 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21369; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27513 = 12'hb79 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24441; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2937 = io_valid_in ? _GEN_27513 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2937 = 12'hb79 == _T_2[11:0] ? image_2937 : _GEN_2936; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6010 = 12'hb7a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9082 = 12'hb7a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6010; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12154 = 12'hb7a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9082; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15226 = 12'hb7a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12154; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18298 = 12'hb7a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15226; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21370 = 12'hb7a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18298; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24442 = 12'hb7a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21370; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27514 = 12'hb7a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24442; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2938 = io_valid_in ? _GEN_27514 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2938 = 12'hb7a == _T_2[11:0] ? image_2938 : _GEN_2937; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6011 = 12'hb7b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9083 = 12'hb7b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6011; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12155 = 12'hb7b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9083; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15227 = 12'hb7b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12155; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18299 = 12'hb7b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15227; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21371 = 12'hb7b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18299; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24443 = 12'hb7b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21371; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27515 = 12'hb7b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24443; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2939 = io_valid_in ? _GEN_27515 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2939 = 12'hb7b == _T_2[11:0] ? image_2939 : _GEN_2938; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6012 = 12'hb7c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9084 = 12'hb7c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6012; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12156 = 12'hb7c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9084; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15228 = 12'hb7c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12156; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18300 = 12'hb7c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15228; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21372 = 12'hb7c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18300; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24444 = 12'hb7c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21372; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27516 = 12'hb7c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24444; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2940 = io_valid_in ? _GEN_27516 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2940 = 12'hb7c == _T_2[11:0] ? image_2940 : _GEN_2939; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6013 = 12'hb7d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9085 = 12'hb7d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6013; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12157 = 12'hb7d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9085; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15229 = 12'hb7d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12157; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18301 = 12'hb7d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15229; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21373 = 12'hb7d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18301; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24445 = 12'hb7d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21373; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27517 = 12'hb7d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24445; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2941 = io_valid_in ? _GEN_27517 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2941 = 12'hb7d == _T_2[11:0] ? image_2941 : _GEN_2940; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6014 = 12'hb7e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9086 = 12'hb7e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6014; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12158 = 12'hb7e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9086; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15230 = 12'hb7e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12158; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18302 = 12'hb7e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15230; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21374 = 12'hb7e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18302; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24446 = 12'hb7e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21374; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27518 = 12'hb7e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24446; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2942 = io_valid_in ? _GEN_27518 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2942 = 12'hb7e == _T_2[11:0] ? image_2942 : _GEN_2941; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6015 = 12'hb7f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9087 = 12'hb7f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6015; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12159 = 12'hb7f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9087; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15231 = 12'hb7f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12159; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18303 = 12'hb7f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15231; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21375 = 12'hb7f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18303; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24447 = 12'hb7f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21375; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27519 = 12'hb7f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24447; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2943 = io_valid_in ? _GEN_27519 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2943 = 12'hb7f == _T_2[11:0] ? image_2943 : _GEN_2942; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6016 = 12'hb80 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9088 = 12'hb80 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6016; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12160 = 12'hb80 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9088; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15232 = 12'hb80 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12160; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18304 = 12'hb80 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15232; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21376 = 12'hb80 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18304; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24448 = 12'hb80 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21376; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27520 = 12'hb80 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24448; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2944 = io_valid_in ? _GEN_27520 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2944 = 12'hb80 == _T_2[11:0] ? image_2944 : _GEN_2943; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6017 = 12'hb81 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9089 = 12'hb81 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6017; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12161 = 12'hb81 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9089; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15233 = 12'hb81 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12161; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18305 = 12'hb81 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15233; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21377 = 12'hb81 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18305; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24449 = 12'hb81 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21377; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27521 = 12'hb81 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24449; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2945 = io_valid_in ? _GEN_27521 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2945 = 12'hb81 == _T_2[11:0] ? image_2945 : _GEN_2944; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6018 = 12'hb82 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9090 = 12'hb82 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6018; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12162 = 12'hb82 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9090; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15234 = 12'hb82 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12162; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18306 = 12'hb82 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15234; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21378 = 12'hb82 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18306; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24450 = 12'hb82 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21378; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27522 = 12'hb82 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24450; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2946 = io_valid_in ? _GEN_27522 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2946 = 12'hb82 == _T_2[11:0] ? image_2946 : _GEN_2945; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6019 = 12'hb83 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9091 = 12'hb83 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6019; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12163 = 12'hb83 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9091; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15235 = 12'hb83 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12163; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18307 = 12'hb83 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15235; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21379 = 12'hb83 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18307; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24451 = 12'hb83 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21379; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27523 = 12'hb83 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24451; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2947 = io_valid_in ? _GEN_27523 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2947 = 12'hb83 == _T_2[11:0] ? image_2947 : _GEN_2946; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6020 = 12'hb84 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9092 = 12'hb84 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6020; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12164 = 12'hb84 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9092; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15236 = 12'hb84 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12164; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18308 = 12'hb84 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15236; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21380 = 12'hb84 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18308; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24452 = 12'hb84 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21380; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27524 = 12'hb84 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24452; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2948 = io_valid_in ? _GEN_27524 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2948 = 12'hb84 == _T_2[11:0] ? image_2948 : _GEN_2947; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6021 = 12'hb85 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9093 = 12'hb85 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6021; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12165 = 12'hb85 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9093; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15237 = 12'hb85 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12165; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18309 = 12'hb85 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15237; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21381 = 12'hb85 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18309; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24453 = 12'hb85 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21381; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27525 = 12'hb85 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24453; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2949 = io_valid_in ? _GEN_27525 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2949 = 12'hb85 == _T_2[11:0] ? image_2949 : _GEN_2948; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6022 = 12'hb86 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9094 = 12'hb86 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6022; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12166 = 12'hb86 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9094; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15238 = 12'hb86 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12166; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18310 = 12'hb86 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15238; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21382 = 12'hb86 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18310; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24454 = 12'hb86 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21382; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27526 = 12'hb86 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24454; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2950 = io_valid_in ? _GEN_27526 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2950 = 12'hb86 == _T_2[11:0] ? image_2950 : _GEN_2949; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6023 = 12'hb87 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9095 = 12'hb87 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6023; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12167 = 12'hb87 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9095; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15239 = 12'hb87 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12167; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18311 = 12'hb87 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15239; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21383 = 12'hb87 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18311; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24455 = 12'hb87 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21383; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27527 = 12'hb87 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24455; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2951 = io_valid_in ? _GEN_27527 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2951 = 12'hb87 == _T_2[11:0] ? image_2951 : _GEN_2950; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6024 = 12'hb88 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9096 = 12'hb88 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6024; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12168 = 12'hb88 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9096; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15240 = 12'hb88 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12168; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18312 = 12'hb88 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15240; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21384 = 12'hb88 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18312; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24456 = 12'hb88 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21384; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27528 = 12'hb88 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24456; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2952 = io_valid_in ? _GEN_27528 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2952 = 12'hb88 == _T_2[11:0] ? image_2952 : _GEN_2951; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6025 = 12'hb89 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9097 = 12'hb89 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6025; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12169 = 12'hb89 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9097; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15241 = 12'hb89 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12169; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18313 = 12'hb89 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15241; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21385 = 12'hb89 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18313; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24457 = 12'hb89 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21385; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27529 = 12'hb89 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24457; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2953 = io_valid_in ? _GEN_27529 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2953 = 12'hb89 == _T_2[11:0] ? image_2953 : _GEN_2952; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6026 = 12'hb8a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9098 = 12'hb8a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6026; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12170 = 12'hb8a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9098; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15242 = 12'hb8a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12170; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18314 = 12'hb8a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15242; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21386 = 12'hb8a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18314; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24458 = 12'hb8a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21386; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27530 = 12'hb8a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24458; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2954 = io_valid_in ? _GEN_27530 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2954 = 12'hb8a == _T_2[11:0] ? image_2954 : _GEN_2953; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6027 = 12'hb8b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9099 = 12'hb8b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6027; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12171 = 12'hb8b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9099; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15243 = 12'hb8b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12171; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18315 = 12'hb8b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15243; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21387 = 12'hb8b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18315; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24459 = 12'hb8b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21387; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27531 = 12'hb8b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24459; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2955 = io_valid_in ? _GEN_27531 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2955 = 12'hb8b == _T_2[11:0] ? image_2955 : _GEN_2954; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6028 = 12'hb8c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9100 = 12'hb8c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6028; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12172 = 12'hb8c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9100; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15244 = 12'hb8c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12172; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18316 = 12'hb8c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15244; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21388 = 12'hb8c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18316; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24460 = 12'hb8c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21388; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27532 = 12'hb8c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24460; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2956 = io_valid_in ? _GEN_27532 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2956 = 12'hb8c == _T_2[11:0] ? image_2956 : _GEN_2955; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6029 = 12'hb8d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9101 = 12'hb8d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6029; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12173 = 12'hb8d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9101; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15245 = 12'hb8d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12173; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18317 = 12'hb8d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15245; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21389 = 12'hb8d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18317; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24461 = 12'hb8d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21389; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27533 = 12'hb8d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24461; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2957 = io_valid_in ? _GEN_27533 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2957 = 12'hb8d == _T_2[11:0] ? image_2957 : _GEN_2956; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6030 = 12'hb8e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9102 = 12'hb8e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6030; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12174 = 12'hb8e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9102; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15246 = 12'hb8e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12174; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18318 = 12'hb8e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15246; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21390 = 12'hb8e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18318; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24462 = 12'hb8e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21390; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27534 = 12'hb8e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24462; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2958 = io_valid_in ? _GEN_27534 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2958 = 12'hb8e == _T_2[11:0] ? image_2958 : _GEN_2957; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6031 = 12'hb8f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9103 = 12'hb8f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6031; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12175 = 12'hb8f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9103; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15247 = 12'hb8f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12175; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18319 = 12'hb8f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15247; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21391 = 12'hb8f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18319; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24463 = 12'hb8f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21391; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27535 = 12'hb8f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24463; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2959 = io_valid_in ? _GEN_27535 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2959 = 12'hb8f == _T_2[11:0] ? image_2959 : _GEN_2958; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6032 = 12'hb90 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9104 = 12'hb90 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6032; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12176 = 12'hb90 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9104; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15248 = 12'hb90 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12176; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18320 = 12'hb90 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15248; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21392 = 12'hb90 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18320; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24464 = 12'hb90 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21392; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27536 = 12'hb90 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24464; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2960 = io_valid_in ? _GEN_27536 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2960 = 12'hb90 == _T_2[11:0] ? image_2960 : _GEN_2959; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6033 = 12'hb91 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9105 = 12'hb91 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6033; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12177 = 12'hb91 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9105; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15249 = 12'hb91 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12177; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18321 = 12'hb91 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15249; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21393 = 12'hb91 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18321; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24465 = 12'hb91 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21393; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27537 = 12'hb91 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24465; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2961 = io_valid_in ? _GEN_27537 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2961 = 12'hb91 == _T_2[11:0] ? image_2961 : _GEN_2960; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6034 = 12'hb92 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9106 = 12'hb92 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6034; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12178 = 12'hb92 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9106; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15250 = 12'hb92 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12178; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18322 = 12'hb92 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15250; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21394 = 12'hb92 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18322; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24466 = 12'hb92 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21394; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27538 = 12'hb92 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24466; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2962 = io_valid_in ? _GEN_27538 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2962 = 12'hb92 == _T_2[11:0] ? image_2962 : _GEN_2961; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6035 = 12'hb93 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9107 = 12'hb93 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6035; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12179 = 12'hb93 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9107; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15251 = 12'hb93 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12179; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18323 = 12'hb93 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15251; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21395 = 12'hb93 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18323; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24467 = 12'hb93 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21395; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27539 = 12'hb93 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24467; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2963 = io_valid_in ? _GEN_27539 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2963 = 12'hb93 == _T_2[11:0] ? image_2963 : _GEN_2962; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6036 = 12'hb94 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9108 = 12'hb94 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6036; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12180 = 12'hb94 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9108; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15252 = 12'hb94 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12180; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18324 = 12'hb94 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15252; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21396 = 12'hb94 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18324; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24468 = 12'hb94 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21396; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27540 = 12'hb94 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24468; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2964 = io_valid_in ? _GEN_27540 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2964 = 12'hb94 == _T_2[11:0] ? image_2964 : _GEN_2963; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6037 = 12'hb95 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9109 = 12'hb95 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6037; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12181 = 12'hb95 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9109; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15253 = 12'hb95 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12181; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18325 = 12'hb95 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15253; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21397 = 12'hb95 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18325; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24469 = 12'hb95 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21397; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27541 = 12'hb95 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24469; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2965 = io_valid_in ? _GEN_27541 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2965 = 12'hb95 == _T_2[11:0] ? image_2965 : _GEN_2964; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6038 = 12'hb96 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9110 = 12'hb96 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6038; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12182 = 12'hb96 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9110; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15254 = 12'hb96 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12182; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18326 = 12'hb96 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15254; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21398 = 12'hb96 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18326; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24470 = 12'hb96 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21398; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27542 = 12'hb96 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24470; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2966 = io_valid_in ? _GEN_27542 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2966 = 12'hb96 == _T_2[11:0] ? image_2966 : _GEN_2965; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6039 = 12'hb97 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9111 = 12'hb97 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6039; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12183 = 12'hb97 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9111; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15255 = 12'hb97 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12183; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18327 = 12'hb97 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15255; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21399 = 12'hb97 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18327; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24471 = 12'hb97 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21399; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27543 = 12'hb97 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24471; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2967 = io_valid_in ? _GEN_27543 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2967 = 12'hb97 == _T_2[11:0] ? image_2967 : _GEN_2966; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6040 = 12'hb98 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9112 = 12'hb98 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6040; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12184 = 12'hb98 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9112; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15256 = 12'hb98 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12184; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18328 = 12'hb98 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15256; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21400 = 12'hb98 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18328; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24472 = 12'hb98 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21400; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27544 = 12'hb98 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24472; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2968 = io_valid_in ? _GEN_27544 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2968 = 12'hb98 == _T_2[11:0] ? image_2968 : _GEN_2967; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6041 = 12'hb99 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9113 = 12'hb99 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6041; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12185 = 12'hb99 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9113; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15257 = 12'hb99 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12185; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18329 = 12'hb99 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15257; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21401 = 12'hb99 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18329; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24473 = 12'hb99 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21401; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27545 = 12'hb99 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24473; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2969 = io_valid_in ? _GEN_27545 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2969 = 12'hb99 == _T_2[11:0] ? image_2969 : _GEN_2968; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6042 = 12'hb9a == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9114 = 12'hb9a == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6042; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12186 = 12'hb9a == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9114; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15258 = 12'hb9a == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12186; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18330 = 12'hb9a == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15258; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21402 = 12'hb9a == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18330; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24474 = 12'hb9a == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21402; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27546 = 12'hb9a == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24474; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2970 = io_valid_in ? _GEN_27546 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2970 = 12'hb9a == _T_2[11:0] ? image_2970 : _GEN_2969; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6043 = 12'hb9b == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9115 = 12'hb9b == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6043; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12187 = 12'hb9b == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9115; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15259 = 12'hb9b == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12187; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18331 = 12'hb9b == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15259; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21403 = 12'hb9b == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18331; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24475 = 12'hb9b == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21403; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27547 = 12'hb9b == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24475; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2971 = io_valid_in ? _GEN_27547 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2971 = 12'hb9b == _T_2[11:0] ? image_2971 : _GEN_2970; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6044 = 12'hb9c == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9116 = 12'hb9c == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6044; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12188 = 12'hb9c == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9116; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15260 = 12'hb9c == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12188; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18332 = 12'hb9c == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15260; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21404 = 12'hb9c == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18332; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24476 = 12'hb9c == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21404; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27548 = 12'hb9c == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24476; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2972 = io_valid_in ? _GEN_27548 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2972 = 12'hb9c == _T_2[11:0] ? image_2972 : _GEN_2971; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6045 = 12'hb9d == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9117 = 12'hb9d == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6045; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12189 = 12'hb9d == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9117; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15261 = 12'hb9d == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12189; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18333 = 12'hb9d == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15261; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21405 = 12'hb9d == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18333; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24477 = 12'hb9d == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21405; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27549 = 12'hb9d == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24477; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2973 = io_valid_in ? _GEN_27549 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2973 = 12'hb9d == _T_2[11:0] ? image_2973 : _GEN_2972; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6046 = 12'hb9e == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9118 = 12'hb9e == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6046; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12190 = 12'hb9e == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9118; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15262 = 12'hb9e == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12190; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18334 = 12'hb9e == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15262; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21406 = 12'hb9e == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18334; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24478 = 12'hb9e == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21406; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27550 = 12'hb9e == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24478; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2974 = io_valid_in ? _GEN_27550 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2974 = 12'hb9e == _T_2[11:0] ? image_2974 : _GEN_2973; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6047 = 12'hb9f == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9119 = 12'hb9f == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6047; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12191 = 12'hb9f == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9119; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15263 = 12'hb9f == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12191; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18335 = 12'hb9f == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15263; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21407 = 12'hb9f == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18335; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24479 = 12'hb9f == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21407; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27551 = 12'hb9f == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24479; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2975 = io_valid_in ? _GEN_27551 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2975 = 12'hb9f == _T_2[11:0] ? image_2975 : _GEN_2974; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6048 = 12'hba0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9120 = 12'hba0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6048; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12192 = 12'hba0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9120; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15264 = 12'hba0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12192; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18336 = 12'hba0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15264; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21408 = 12'hba0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18336; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24480 = 12'hba0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21408; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27552 = 12'hba0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24480; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2976 = io_valid_in ? _GEN_27552 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2976 = 12'hba0 == _T_2[11:0] ? image_2976 : _GEN_2975; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6049 = 12'hba1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9121 = 12'hba1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6049; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12193 = 12'hba1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9121; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15265 = 12'hba1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12193; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18337 = 12'hba1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15265; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21409 = 12'hba1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18337; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24481 = 12'hba1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21409; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27553 = 12'hba1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24481; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2977 = io_valid_in ? _GEN_27553 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2977 = 12'hba1 == _T_2[11:0] ? image_2977 : _GEN_2976; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6050 = 12'hba2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9122 = 12'hba2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6050; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12194 = 12'hba2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9122; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15266 = 12'hba2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12194; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18338 = 12'hba2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15266; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21410 = 12'hba2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18338; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24482 = 12'hba2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21410; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27554 = 12'hba2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24482; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2978 = io_valid_in ? _GEN_27554 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2978 = 12'hba2 == _T_2[11:0] ? image_2978 : _GEN_2977; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6051 = 12'hba3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9123 = 12'hba3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6051; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12195 = 12'hba3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9123; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15267 = 12'hba3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12195; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18339 = 12'hba3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15267; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21411 = 12'hba3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18339; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24483 = 12'hba3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21411; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27555 = 12'hba3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24483; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2979 = io_valid_in ? _GEN_27555 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2979 = 12'hba3 == _T_2[11:0] ? image_2979 : _GEN_2978; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6052 = 12'hba4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9124 = 12'hba4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6052; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12196 = 12'hba4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9124; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15268 = 12'hba4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12196; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18340 = 12'hba4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15268; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21412 = 12'hba4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18340; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24484 = 12'hba4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21412; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27556 = 12'hba4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24484; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2980 = io_valid_in ? _GEN_27556 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2980 = 12'hba4 == _T_2[11:0] ? image_2980 : _GEN_2979; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6053 = 12'hba5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9125 = 12'hba5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6053; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12197 = 12'hba5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9125; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15269 = 12'hba5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12197; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18341 = 12'hba5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15269; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21413 = 12'hba5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18341; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24485 = 12'hba5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21413; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27557 = 12'hba5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24485; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2981 = io_valid_in ? _GEN_27557 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2981 = 12'hba5 == _T_2[11:0] ? image_2981 : _GEN_2980; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6054 = 12'hba6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9126 = 12'hba6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6054; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12198 = 12'hba6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9126; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15270 = 12'hba6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12198; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18342 = 12'hba6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15270; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21414 = 12'hba6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18342; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24486 = 12'hba6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21414; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27558 = 12'hba6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24486; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2982 = io_valid_in ? _GEN_27558 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2982 = 12'hba6 == _T_2[11:0] ? image_2982 : _GEN_2981; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6055 = 12'hba7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9127 = 12'hba7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6055; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12199 = 12'hba7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9127; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15271 = 12'hba7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12199; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18343 = 12'hba7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15271; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21415 = 12'hba7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18343; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24487 = 12'hba7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21415; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27559 = 12'hba7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24487; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2983 = io_valid_in ? _GEN_27559 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2983 = 12'hba7 == _T_2[11:0] ? image_2983 : _GEN_2982; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6056 = 12'hba8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9128 = 12'hba8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6056; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12200 = 12'hba8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9128; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15272 = 12'hba8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12200; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18344 = 12'hba8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15272; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21416 = 12'hba8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18344; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24488 = 12'hba8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21416; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27560 = 12'hba8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24488; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2984 = io_valid_in ? _GEN_27560 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2984 = 12'hba8 == _T_2[11:0] ? image_2984 : _GEN_2983; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6057 = 12'hba9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9129 = 12'hba9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6057; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12201 = 12'hba9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9129; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15273 = 12'hba9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12201; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18345 = 12'hba9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15273; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21417 = 12'hba9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18345; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24489 = 12'hba9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21417; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27561 = 12'hba9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24489; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2985 = io_valid_in ? _GEN_27561 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2985 = 12'hba9 == _T_2[11:0] ? image_2985 : _GEN_2984; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6058 = 12'hbaa == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9130 = 12'hbaa == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6058; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12202 = 12'hbaa == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9130; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15274 = 12'hbaa == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12202; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18346 = 12'hbaa == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15274; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21418 = 12'hbaa == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18346; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24490 = 12'hbaa == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21418; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27562 = 12'hbaa == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24490; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2986 = io_valid_in ? _GEN_27562 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2986 = 12'hbaa == _T_2[11:0] ? image_2986 : _GEN_2985; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6059 = 12'hbab == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9131 = 12'hbab == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6059; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12203 = 12'hbab == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9131; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15275 = 12'hbab == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12203; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18347 = 12'hbab == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15275; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21419 = 12'hbab == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18347; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24491 = 12'hbab == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21419; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27563 = 12'hbab == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24491; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2987 = io_valid_in ? _GEN_27563 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2987 = 12'hbab == _T_2[11:0] ? image_2987 : _GEN_2986; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6060 = 12'hbac == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9132 = 12'hbac == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6060; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12204 = 12'hbac == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9132; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15276 = 12'hbac == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12204; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18348 = 12'hbac == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15276; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21420 = 12'hbac == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18348; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24492 = 12'hbac == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21420; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27564 = 12'hbac == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24492; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2988 = io_valid_in ? _GEN_27564 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2988 = 12'hbac == _T_2[11:0] ? image_2988 : _GEN_2987; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6061 = 12'hbad == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9133 = 12'hbad == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6061; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12205 = 12'hbad == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9133; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15277 = 12'hbad == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12205; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18349 = 12'hbad == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15277; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21421 = 12'hbad == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18349; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24493 = 12'hbad == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21421; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27565 = 12'hbad == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24493; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2989 = io_valid_in ? _GEN_27565 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2989 = 12'hbad == _T_2[11:0] ? image_2989 : _GEN_2988; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6062 = 12'hbae == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9134 = 12'hbae == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6062; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12206 = 12'hbae == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9134; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15278 = 12'hbae == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12206; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18350 = 12'hbae == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15278; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21422 = 12'hbae == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18350; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24494 = 12'hbae == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21422; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27566 = 12'hbae == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24494; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2990 = io_valid_in ? _GEN_27566 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2990 = 12'hbae == _T_2[11:0] ? image_2990 : _GEN_2989; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6063 = 12'hbaf == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9135 = 12'hbaf == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6063; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12207 = 12'hbaf == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9135; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15279 = 12'hbaf == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12207; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18351 = 12'hbaf == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15279; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21423 = 12'hbaf == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18351; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24495 = 12'hbaf == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21423; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27567 = 12'hbaf == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24495; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2991 = io_valid_in ? _GEN_27567 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2991 = 12'hbaf == _T_2[11:0] ? image_2991 : _GEN_2990; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6064 = 12'hbb0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9136 = 12'hbb0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6064; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12208 = 12'hbb0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9136; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15280 = 12'hbb0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12208; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18352 = 12'hbb0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15280; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21424 = 12'hbb0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18352; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24496 = 12'hbb0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21424; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27568 = 12'hbb0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24496; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2992 = io_valid_in ? _GEN_27568 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2992 = 12'hbb0 == _T_2[11:0] ? image_2992 : _GEN_2991; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6065 = 12'hbb1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9137 = 12'hbb1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6065; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12209 = 12'hbb1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9137; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15281 = 12'hbb1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12209; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18353 = 12'hbb1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15281; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21425 = 12'hbb1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18353; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24497 = 12'hbb1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21425; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27569 = 12'hbb1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24497; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2993 = io_valid_in ? _GEN_27569 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2993 = 12'hbb1 == _T_2[11:0] ? image_2993 : _GEN_2992; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6066 = 12'hbb2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9138 = 12'hbb2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6066; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12210 = 12'hbb2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9138; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15282 = 12'hbb2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12210; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18354 = 12'hbb2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15282; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21426 = 12'hbb2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18354; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24498 = 12'hbb2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21426; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27570 = 12'hbb2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24498; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2994 = io_valid_in ? _GEN_27570 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2994 = 12'hbb2 == _T_2[11:0] ? image_2994 : _GEN_2993; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6067 = 12'hbb3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9139 = 12'hbb3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6067; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12211 = 12'hbb3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9139; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15283 = 12'hbb3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12211; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18355 = 12'hbb3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15283; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21427 = 12'hbb3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18355; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24499 = 12'hbb3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21427; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27571 = 12'hbb3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24499; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2995 = io_valid_in ? _GEN_27571 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2995 = 12'hbb3 == _T_2[11:0] ? image_2995 : _GEN_2994; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6068 = 12'hbb4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9140 = 12'hbb4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6068; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12212 = 12'hbb4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9140; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15284 = 12'hbb4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12212; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18356 = 12'hbb4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15284; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21428 = 12'hbb4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18356; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24500 = 12'hbb4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21428; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27572 = 12'hbb4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24500; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2996 = io_valid_in ? _GEN_27572 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2996 = 12'hbb4 == _T_2[11:0] ? image_2996 : _GEN_2995; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6069 = 12'hbb5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9141 = 12'hbb5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6069; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12213 = 12'hbb5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9141; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15285 = 12'hbb5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12213; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18357 = 12'hbb5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15285; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21429 = 12'hbb5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18357; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24501 = 12'hbb5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21429; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27573 = 12'hbb5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24501; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2997 = io_valid_in ? _GEN_27573 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2997 = 12'hbb5 == _T_2[11:0] ? image_2997 : _GEN_2996; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6070 = 12'hbb6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9142 = 12'hbb6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6070; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12214 = 12'hbb6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9142; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15286 = 12'hbb6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12214; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18358 = 12'hbb6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15286; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21430 = 12'hbb6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18358; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24502 = 12'hbb6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21430; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27574 = 12'hbb6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24502; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2998 = io_valid_in ? _GEN_27574 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2998 = 12'hbb6 == _T_2[11:0] ? image_2998 : _GEN_2997; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6071 = 12'hbb7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9143 = 12'hbb7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6071; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12215 = 12'hbb7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9143; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15287 = 12'hbb7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12215; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18359 = 12'hbb7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15287; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21431 = 12'hbb7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18359; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24503 = 12'hbb7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21431; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27575 = 12'hbb7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24503; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2999 = io_valid_in ? _GEN_27575 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2999 = 12'hbb7 == _T_2[11:0] ? image_2999 : _GEN_2998; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6072 = 12'hbb8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9144 = 12'hbb8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6072; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12216 = 12'hbb8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9144; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15288 = 12'hbb8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12216; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18360 = 12'hbb8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15288; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21432 = 12'hbb8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18360; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24504 = 12'hbb8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21432; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27576 = 12'hbb8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24504; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3000 = io_valid_in ? _GEN_27576 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3000 = 12'hbb8 == _T_2[11:0] ? image_3000 : _GEN_2999; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6073 = 12'hbb9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9145 = 12'hbb9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6073; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12217 = 12'hbb9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9145; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15289 = 12'hbb9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12217; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18361 = 12'hbb9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15289; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21433 = 12'hbb9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18361; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24505 = 12'hbb9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21433; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27577 = 12'hbb9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24505; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3001 = io_valid_in ? _GEN_27577 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3001 = 12'hbb9 == _T_2[11:0] ? image_3001 : _GEN_3000; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6074 = 12'hbba == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9146 = 12'hbba == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6074; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12218 = 12'hbba == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9146; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15290 = 12'hbba == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12218; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18362 = 12'hbba == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15290; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21434 = 12'hbba == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18362; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24506 = 12'hbba == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21434; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27578 = 12'hbba == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24506; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3002 = io_valid_in ? _GEN_27578 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3002 = 12'hbba == _T_2[11:0] ? image_3002 : _GEN_3001; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6075 = 12'hbbb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9147 = 12'hbbb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6075; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12219 = 12'hbbb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9147; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15291 = 12'hbbb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12219; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18363 = 12'hbbb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15291; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21435 = 12'hbbb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18363; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24507 = 12'hbbb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21435; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27579 = 12'hbbb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24507; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3003 = io_valid_in ? _GEN_27579 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3003 = 12'hbbb == _T_2[11:0] ? image_3003 : _GEN_3002; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6076 = 12'hbbc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9148 = 12'hbbc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6076; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12220 = 12'hbbc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9148; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15292 = 12'hbbc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12220; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18364 = 12'hbbc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15292; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21436 = 12'hbbc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18364; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24508 = 12'hbbc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21436; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27580 = 12'hbbc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24508; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3004 = io_valid_in ? _GEN_27580 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3004 = 12'hbbc == _T_2[11:0] ? image_3004 : _GEN_3003; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6077 = 12'hbbd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9149 = 12'hbbd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6077; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12221 = 12'hbbd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9149; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15293 = 12'hbbd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12221; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18365 = 12'hbbd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15293; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21437 = 12'hbbd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18365; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24509 = 12'hbbd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21437; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27581 = 12'hbbd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24509; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3005 = io_valid_in ? _GEN_27581 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3005 = 12'hbbd == _T_2[11:0] ? image_3005 : _GEN_3004; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6078 = 12'hbbe == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9150 = 12'hbbe == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6078; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12222 = 12'hbbe == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9150; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15294 = 12'hbbe == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12222; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18366 = 12'hbbe == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15294; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21438 = 12'hbbe == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18366; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24510 = 12'hbbe == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21438; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27582 = 12'hbbe == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24510; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3006 = io_valid_in ? _GEN_27582 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3006 = 12'hbbe == _T_2[11:0] ? image_3006 : _GEN_3005; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6079 = 12'hbbf == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9151 = 12'hbbf == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6079; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12223 = 12'hbbf == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9151; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15295 = 12'hbbf == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12223; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18367 = 12'hbbf == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15295; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21439 = 12'hbbf == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18367; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24511 = 12'hbbf == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21439; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27583 = 12'hbbf == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24511; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3007 = io_valid_in ? _GEN_27583 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3007 = 12'hbbf == _T_2[11:0] ? image_3007 : _GEN_3006; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6080 = 12'hbc0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9152 = 12'hbc0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6080; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12224 = 12'hbc0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9152; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15296 = 12'hbc0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12224; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18368 = 12'hbc0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15296; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21440 = 12'hbc0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18368; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24512 = 12'hbc0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21440; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27584 = 12'hbc0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24512; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3008 = io_valid_in ? _GEN_27584 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3008 = 12'hbc0 == _T_2[11:0] ? image_3008 : _GEN_3007; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6081 = 12'hbc1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9153 = 12'hbc1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6081; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12225 = 12'hbc1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9153; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15297 = 12'hbc1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12225; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18369 = 12'hbc1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15297; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21441 = 12'hbc1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18369; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24513 = 12'hbc1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21441; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27585 = 12'hbc1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24513; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3009 = io_valid_in ? _GEN_27585 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3009 = 12'hbc1 == _T_2[11:0] ? image_3009 : _GEN_3008; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6082 = 12'hbc2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9154 = 12'hbc2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6082; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12226 = 12'hbc2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9154; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15298 = 12'hbc2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12226; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18370 = 12'hbc2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15298; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21442 = 12'hbc2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18370; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24514 = 12'hbc2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21442; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27586 = 12'hbc2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24514; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3010 = io_valid_in ? _GEN_27586 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3010 = 12'hbc2 == _T_2[11:0] ? image_3010 : _GEN_3009; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6083 = 12'hbc3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9155 = 12'hbc3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6083; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12227 = 12'hbc3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9155; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15299 = 12'hbc3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12227; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18371 = 12'hbc3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15299; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21443 = 12'hbc3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18371; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24515 = 12'hbc3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21443; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27587 = 12'hbc3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24515; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3011 = io_valid_in ? _GEN_27587 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3011 = 12'hbc3 == _T_2[11:0] ? image_3011 : _GEN_3010; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6084 = 12'hbc4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9156 = 12'hbc4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6084; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12228 = 12'hbc4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9156; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15300 = 12'hbc4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12228; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18372 = 12'hbc4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15300; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21444 = 12'hbc4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18372; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24516 = 12'hbc4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21444; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27588 = 12'hbc4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24516; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3012 = io_valid_in ? _GEN_27588 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3012 = 12'hbc4 == _T_2[11:0] ? image_3012 : _GEN_3011; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6085 = 12'hbc5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9157 = 12'hbc5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6085; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12229 = 12'hbc5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9157; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15301 = 12'hbc5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12229; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18373 = 12'hbc5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15301; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21445 = 12'hbc5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18373; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24517 = 12'hbc5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21445; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27589 = 12'hbc5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24517; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3013 = io_valid_in ? _GEN_27589 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3013 = 12'hbc5 == _T_2[11:0] ? image_3013 : _GEN_3012; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6086 = 12'hbc6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9158 = 12'hbc6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6086; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12230 = 12'hbc6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9158; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15302 = 12'hbc6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12230; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18374 = 12'hbc6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15302; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21446 = 12'hbc6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18374; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24518 = 12'hbc6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21446; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27590 = 12'hbc6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24518; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3014 = io_valid_in ? _GEN_27590 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3014 = 12'hbc6 == _T_2[11:0] ? image_3014 : _GEN_3013; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6087 = 12'hbc7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9159 = 12'hbc7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6087; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12231 = 12'hbc7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9159; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15303 = 12'hbc7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12231; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18375 = 12'hbc7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15303; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21447 = 12'hbc7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18375; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24519 = 12'hbc7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21447; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27591 = 12'hbc7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24519; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3015 = io_valid_in ? _GEN_27591 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3015 = 12'hbc7 == _T_2[11:0] ? image_3015 : _GEN_3014; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6088 = 12'hbc8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9160 = 12'hbc8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6088; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12232 = 12'hbc8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9160; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15304 = 12'hbc8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12232; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18376 = 12'hbc8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15304; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21448 = 12'hbc8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18376; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24520 = 12'hbc8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21448; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27592 = 12'hbc8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24520; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3016 = io_valid_in ? _GEN_27592 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3016 = 12'hbc8 == _T_2[11:0] ? image_3016 : _GEN_3015; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6089 = 12'hbc9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9161 = 12'hbc9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6089; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12233 = 12'hbc9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9161; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15305 = 12'hbc9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12233; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18377 = 12'hbc9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15305; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21449 = 12'hbc9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18377; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24521 = 12'hbc9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21449; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27593 = 12'hbc9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24521; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3017 = io_valid_in ? _GEN_27593 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3017 = 12'hbc9 == _T_2[11:0] ? image_3017 : _GEN_3016; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6090 = 12'hbca == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9162 = 12'hbca == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6090; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12234 = 12'hbca == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9162; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15306 = 12'hbca == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12234; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18378 = 12'hbca == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15306; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21450 = 12'hbca == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18378; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24522 = 12'hbca == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21450; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27594 = 12'hbca == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24522; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3018 = io_valid_in ? _GEN_27594 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3018 = 12'hbca == _T_2[11:0] ? image_3018 : _GEN_3017; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6091 = 12'hbcb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9163 = 12'hbcb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6091; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12235 = 12'hbcb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9163; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15307 = 12'hbcb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12235; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18379 = 12'hbcb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15307; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21451 = 12'hbcb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18379; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24523 = 12'hbcb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21451; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27595 = 12'hbcb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24523; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3019 = io_valid_in ? _GEN_27595 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3019 = 12'hbcb == _T_2[11:0] ? image_3019 : _GEN_3018; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6092 = 12'hbcc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9164 = 12'hbcc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6092; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12236 = 12'hbcc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9164; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15308 = 12'hbcc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12236; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18380 = 12'hbcc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15308; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21452 = 12'hbcc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18380; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24524 = 12'hbcc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21452; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27596 = 12'hbcc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24524; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3020 = io_valid_in ? _GEN_27596 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3020 = 12'hbcc == _T_2[11:0] ? image_3020 : _GEN_3019; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6093 = 12'hbcd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9165 = 12'hbcd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6093; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12237 = 12'hbcd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9165; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15309 = 12'hbcd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12237; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18381 = 12'hbcd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15309; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21453 = 12'hbcd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18381; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24525 = 12'hbcd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21453; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27597 = 12'hbcd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24525; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3021 = io_valid_in ? _GEN_27597 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3021 = 12'hbcd == _T_2[11:0] ? image_3021 : _GEN_3020; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6094 = 12'hbce == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9166 = 12'hbce == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6094; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12238 = 12'hbce == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9166; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15310 = 12'hbce == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12238; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18382 = 12'hbce == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15310; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21454 = 12'hbce == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18382; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24526 = 12'hbce == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21454; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27598 = 12'hbce == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24526; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3022 = io_valid_in ? _GEN_27598 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3022 = 12'hbce == _T_2[11:0] ? image_3022 : _GEN_3021; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6095 = 12'hbcf == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9167 = 12'hbcf == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6095; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12239 = 12'hbcf == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9167; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15311 = 12'hbcf == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12239; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18383 = 12'hbcf == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15311; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21455 = 12'hbcf == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18383; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24527 = 12'hbcf == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21455; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27599 = 12'hbcf == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24527; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3023 = io_valid_in ? _GEN_27599 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3023 = 12'hbcf == _T_2[11:0] ? image_3023 : _GEN_3022; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6096 = 12'hbd0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9168 = 12'hbd0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6096; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12240 = 12'hbd0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9168; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15312 = 12'hbd0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12240; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18384 = 12'hbd0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15312; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21456 = 12'hbd0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18384; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24528 = 12'hbd0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21456; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27600 = 12'hbd0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24528; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3024 = io_valid_in ? _GEN_27600 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3024 = 12'hbd0 == _T_2[11:0] ? image_3024 : _GEN_3023; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6097 = 12'hbd1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9169 = 12'hbd1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6097; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12241 = 12'hbd1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9169; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15313 = 12'hbd1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12241; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18385 = 12'hbd1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15313; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21457 = 12'hbd1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18385; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24529 = 12'hbd1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21457; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27601 = 12'hbd1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24529; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3025 = io_valid_in ? _GEN_27601 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3025 = 12'hbd1 == _T_2[11:0] ? image_3025 : _GEN_3024; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6098 = 12'hbd2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9170 = 12'hbd2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6098; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12242 = 12'hbd2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9170; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15314 = 12'hbd2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12242; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18386 = 12'hbd2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15314; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21458 = 12'hbd2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18386; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24530 = 12'hbd2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21458; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27602 = 12'hbd2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24530; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3026 = io_valid_in ? _GEN_27602 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3026 = 12'hbd2 == _T_2[11:0] ? image_3026 : _GEN_3025; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6099 = 12'hbd3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9171 = 12'hbd3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6099; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12243 = 12'hbd3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9171; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15315 = 12'hbd3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12243; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18387 = 12'hbd3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15315; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21459 = 12'hbd3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18387; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24531 = 12'hbd3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21459; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27603 = 12'hbd3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24531; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3027 = io_valid_in ? _GEN_27603 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3027 = 12'hbd3 == _T_2[11:0] ? image_3027 : _GEN_3026; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6100 = 12'hbd4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9172 = 12'hbd4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6100; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12244 = 12'hbd4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9172; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15316 = 12'hbd4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12244; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18388 = 12'hbd4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15316; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21460 = 12'hbd4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18388; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24532 = 12'hbd4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21460; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27604 = 12'hbd4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24532; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3028 = io_valid_in ? _GEN_27604 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3028 = 12'hbd4 == _T_2[11:0] ? image_3028 : _GEN_3027; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6101 = 12'hbd5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9173 = 12'hbd5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6101; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12245 = 12'hbd5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9173; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15317 = 12'hbd5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12245; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18389 = 12'hbd5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15317; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21461 = 12'hbd5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18389; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24533 = 12'hbd5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21461; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27605 = 12'hbd5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24533; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3029 = io_valid_in ? _GEN_27605 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3029 = 12'hbd5 == _T_2[11:0] ? image_3029 : _GEN_3028; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6102 = 12'hbd6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9174 = 12'hbd6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6102; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12246 = 12'hbd6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9174; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15318 = 12'hbd6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12246; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18390 = 12'hbd6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15318; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21462 = 12'hbd6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18390; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24534 = 12'hbd6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21462; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27606 = 12'hbd6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24534; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3030 = io_valid_in ? _GEN_27606 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3030 = 12'hbd6 == _T_2[11:0] ? image_3030 : _GEN_3029; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6103 = 12'hbd7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9175 = 12'hbd7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6103; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12247 = 12'hbd7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9175; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15319 = 12'hbd7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12247; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18391 = 12'hbd7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15319; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21463 = 12'hbd7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18391; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24535 = 12'hbd7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21463; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27607 = 12'hbd7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24535; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3031 = io_valid_in ? _GEN_27607 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3031 = 12'hbd7 == _T_2[11:0] ? image_3031 : _GEN_3030; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6104 = 12'hbd8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9176 = 12'hbd8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6104; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12248 = 12'hbd8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9176; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15320 = 12'hbd8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12248; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18392 = 12'hbd8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15320; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21464 = 12'hbd8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18392; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24536 = 12'hbd8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21464; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27608 = 12'hbd8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24536; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3032 = io_valid_in ? _GEN_27608 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3032 = 12'hbd8 == _T_2[11:0] ? image_3032 : _GEN_3031; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6105 = 12'hbd9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9177 = 12'hbd9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6105; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12249 = 12'hbd9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9177; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15321 = 12'hbd9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12249; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18393 = 12'hbd9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15321; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21465 = 12'hbd9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18393; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24537 = 12'hbd9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21465; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27609 = 12'hbd9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24537; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3033 = io_valid_in ? _GEN_27609 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3033 = 12'hbd9 == _T_2[11:0] ? image_3033 : _GEN_3032; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6106 = 12'hbda == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9178 = 12'hbda == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6106; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12250 = 12'hbda == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9178; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15322 = 12'hbda == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12250; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18394 = 12'hbda == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15322; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21466 = 12'hbda == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18394; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24538 = 12'hbda == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21466; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27610 = 12'hbda == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24538; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3034 = io_valid_in ? _GEN_27610 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3034 = 12'hbda == _T_2[11:0] ? image_3034 : _GEN_3033; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6107 = 12'hbdb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9179 = 12'hbdb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6107; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12251 = 12'hbdb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9179; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15323 = 12'hbdb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12251; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18395 = 12'hbdb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15323; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21467 = 12'hbdb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18395; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24539 = 12'hbdb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21467; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27611 = 12'hbdb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24539; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3035 = io_valid_in ? _GEN_27611 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3035 = 12'hbdb == _T_2[11:0] ? image_3035 : _GEN_3034; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6108 = 12'hbdc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9180 = 12'hbdc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6108; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12252 = 12'hbdc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9180; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15324 = 12'hbdc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12252; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18396 = 12'hbdc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15324; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21468 = 12'hbdc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18396; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24540 = 12'hbdc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21468; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27612 = 12'hbdc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24540; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3036 = io_valid_in ? _GEN_27612 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3036 = 12'hbdc == _T_2[11:0] ? image_3036 : _GEN_3035; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6109 = 12'hbdd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9181 = 12'hbdd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6109; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12253 = 12'hbdd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9181; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15325 = 12'hbdd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12253; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18397 = 12'hbdd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15325; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21469 = 12'hbdd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18397; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24541 = 12'hbdd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21469; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27613 = 12'hbdd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24541; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3037 = io_valid_in ? _GEN_27613 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3037 = 12'hbdd == _T_2[11:0] ? image_3037 : _GEN_3036; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6110 = 12'hbde == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9182 = 12'hbde == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6110; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12254 = 12'hbde == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9182; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15326 = 12'hbde == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12254; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18398 = 12'hbde == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15326; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21470 = 12'hbde == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18398; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24542 = 12'hbde == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21470; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27614 = 12'hbde == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24542; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3038 = io_valid_in ? _GEN_27614 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3038 = 12'hbde == _T_2[11:0] ? image_3038 : _GEN_3037; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6111 = 12'hbdf == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9183 = 12'hbdf == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6111; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12255 = 12'hbdf == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9183; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15327 = 12'hbdf == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12255; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18399 = 12'hbdf == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15327; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21471 = 12'hbdf == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18399; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24543 = 12'hbdf == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21471; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27615 = 12'hbdf == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24543; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3039 = io_valid_in ? _GEN_27615 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3039 = 12'hbdf == _T_2[11:0] ? image_3039 : _GEN_3038; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6112 = 12'hbe0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9184 = 12'hbe0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6112; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12256 = 12'hbe0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9184; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15328 = 12'hbe0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12256; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18400 = 12'hbe0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15328; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21472 = 12'hbe0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18400; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24544 = 12'hbe0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21472; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27616 = 12'hbe0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24544; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3040 = io_valid_in ? _GEN_27616 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3040 = 12'hbe0 == _T_2[11:0] ? image_3040 : _GEN_3039; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6113 = 12'hbe1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9185 = 12'hbe1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6113; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12257 = 12'hbe1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9185; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15329 = 12'hbe1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12257; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18401 = 12'hbe1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15329; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21473 = 12'hbe1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18401; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24545 = 12'hbe1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21473; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27617 = 12'hbe1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24545; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3041 = io_valid_in ? _GEN_27617 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3041 = 12'hbe1 == _T_2[11:0] ? image_3041 : _GEN_3040; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6114 = 12'hbe2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9186 = 12'hbe2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6114; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12258 = 12'hbe2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9186; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15330 = 12'hbe2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12258; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18402 = 12'hbe2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15330; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21474 = 12'hbe2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18402; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24546 = 12'hbe2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21474; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27618 = 12'hbe2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24546; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3042 = io_valid_in ? _GEN_27618 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3042 = 12'hbe2 == _T_2[11:0] ? image_3042 : _GEN_3041; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6115 = 12'hbe3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9187 = 12'hbe3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6115; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12259 = 12'hbe3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9187; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15331 = 12'hbe3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12259; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18403 = 12'hbe3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15331; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21475 = 12'hbe3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18403; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24547 = 12'hbe3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21475; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27619 = 12'hbe3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24547; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3043 = io_valid_in ? _GEN_27619 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3043 = 12'hbe3 == _T_2[11:0] ? image_3043 : _GEN_3042; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6116 = 12'hbe4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9188 = 12'hbe4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6116; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12260 = 12'hbe4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9188; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15332 = 12'hbe4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12260; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18404 = 12'hbe4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15332; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21476 = 12'hbe4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18404; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24548 = 12'hbe4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21476; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27620 = 12'hbe4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24548; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3044 = io_valid_in ? _GEN_27620 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3044 = 12'hbe4 == _T_2[11:0] ? image_3044 : _GEN_3043; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6117 = 12'hbe5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9189 = 12'hbe5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6117; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12261 = 12'hbe5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9189; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15333 = 12'hbe5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12261; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18405 = 12'hbe5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15333; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21477 = 12'hbe5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18405; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24549 = 12'hbe5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21477; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27621 = 12'hbe5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24549; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3045 = io_valid_in ? _GEN_27621 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3045 = 12'hbe5 == _T_2[11:0] ? image_3045 : _GEN_3044; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6118 = 12'hbe6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9190 = 12'hbe6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6118; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12262 = 12'hbe6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9190; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15334 = 12'hbe6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12262; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18406 = 12'hbe6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15334; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21478 = 12'hbe6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18406; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24550 = 12'hbe6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21478; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27622 = 12'hbe6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24550; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3046 = io_valid_in ? _GEN_27622 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3046 = 12'hbe6 == _T_2[11:0] ? image_3046 : _GEN_3045; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6119 = 12'hbe7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9191 = 12'hbe7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6119; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12263 = 12'hbe7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9191; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15335 = 12'hbe7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12263; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18407 = 12'hbe7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15335; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21479 = 12'hbe7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18407; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24551 = 12'hbe7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21479; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27623 = 12'hbe7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24551; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3047 = io_valid_in ? _GEN_27623 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3047 = 12'hbe7 == _T_2[11:0] ? image_3047 : _GEN_3046; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6120 = 12'hbe8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9192 = 12'hbe8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6120; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12264 = 12'hbe8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9192; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15336 = 12'hbe8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12264; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18408 = 12'hbe8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15336; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21480 = 12'hbe8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18408; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24552 = 12'hbe8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21480; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27624 = 12'hbe8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24552; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3048 = io_valid_in ? _GEN_27624 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3048 = 12'hbe8 == _T_2[11:0] ? image_3048 : _GEN_3047; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6121 = 12'hbe9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9193 = 12'hbe9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6121; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12265 = 12'hbe9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9193; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15337 = 12'hbe9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12265; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18409 = 12'hbe9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15337; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21481 = 12'hbe9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18409; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24553 = 12'hbe9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21481; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27625 = 12'hbe9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24553; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3049 = io_valid_in ? _GEN_27625 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3049 = 12'hbe9 == _T_2[11:0] ? image_3049 : _GEN_3048; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6122 = 12'hbea == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9194 = 12'hbea == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6122; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12266 = 12'hbea == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9194; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15338 = 12'hbea == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12266; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18410 = 12'hbea == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15338; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21482 = 12'hbea == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18410; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24554 = 12'hbea == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21482; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27626 = 12'hbea == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24554; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3050 = io_valid_in ? _GEN_27626 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3050 = 12'hbea == _T_2[11:0] ? image_3050 : _GEN_3049; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6123 = 12'hbeb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9195 = 12'hbeb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6123; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12267 = 12'hbeb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9195; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15339 = 12'hbeb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12267; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18411 = 12'hbeb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15339; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21483 = 12'hbeb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18411; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24555 = 12'hbeb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21483; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27627 = 12'hbeb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24555; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3051 = io_valid_in ? _GEN_27627 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3051 = 12'hbeb == _T_2[11:0] ? image_3051 : _GEN_3050; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6124 = 12'hbec == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9196 = 12'hbec == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6124; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12268 = 12'hbec == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9196; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15340 = 12'hbec == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12268; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18412 = 12'hbec == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15340; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21484 = 12'hbec == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18412; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24556 = 12'hbec == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21484; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27628 = 12'hbec == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24556; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3052 = io_valid_in ? _GEN_27628 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3052 = 12'hbec == _T_2[11:0] ? image_3052 : _GEN_3051; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6125 = 12'hbed == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9197 = 12'hbed == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6125; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12269 = 12'hbed == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9197; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15341 = 12'hbed == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12269; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18413 = 12'hbed == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15341; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21485 = 12'hbed == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18413; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24557 = 12'hbed == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21485; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27629 = 12'hbed == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24557; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3053 = io_valid_in ? _GEN_27629 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3053 = 12'hbed == _T_2[11:0] ? image_3053 : _GEN_3052; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6126 = 12'hbee == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9198 = 12'hbee == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6126; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12270 = 12'hbee == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9198; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15342 = 12'hbee == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12270; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18414 = 12'hbee == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15342; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21486 = 12'hbee == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18414; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24558 = 12'hbee == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21486; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27630 = 12'hbee == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24558; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3054 = io_valid_in ? _GEN_27630 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3054 = 12'hbee == _T_2[11:0] ? image_3054 : _GEN_3053; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6127 = 12'hbef == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9199 = 12'hbef == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6127; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12271 = 12'hbef == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9199; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15343 = 12'hbef == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12271; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18415 = 12'hbef == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15343; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21487 = 12'hbef == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18415; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24559 = 12'hbef == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21487; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27631 = 12'hbef == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24559; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3055 = io_valid_in ? _GEN_27631 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3055 = 12'hbef == _T_2[11:0] ? image_3055 : _GEN_3054; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6128 = 12'hbf0 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9200 = 12'hbf0 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6128; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12272 = 12'hbf0 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9200; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15344 = 12'hbf0 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12272; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18416 = 12'hbf0 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15344; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21488 = 12'hbf0 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18416; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24560 = 12'hbf0 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21488; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27632 = 12'hbf0 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24560; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3056 = io_valid_in ? _GEN_27632 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3056 = 12'hbf0 == _T_2[11:0] ? image_3056 : _GEN_3055; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6129 = 12'hbf1 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9201 = 12'hbf1 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6129; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12273 = 12'hbf1 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9201; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15345 = 12'hbf1 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12273; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18417 = 12'hbf1 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15345; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21489 = 12'hbf1 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18417; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24561 = 12'hbf1 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21489; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27633 = 12'hbf1 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24561; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3057 = io_valid_in ? _GEN_27633 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3057 = 12'hbf1 == _T_2[11:0] ? image_3057 : _GEN_3056; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6130 = 12'hbf2 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9202 = 12'hbf2 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6130; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12274 = 12'hbf2 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9202; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15346 = 12'hbf2 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12274; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18418 = 12'hbf2 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15346; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21490 = 12'hbf2 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18418; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24562 = 12'hbf2 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21490; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27634 = 12'hbf2 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24562; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3058 = io_valid_in ? _GEN_27634 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3058 = 12'hbf2 == _T_2[11:0] ? image_3058 : _GEN_3057; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6131 = 12'hbf3 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9203 = 12'hbf3 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6131; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12275 = 12'hbf3 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9203; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15347 = 12'hbf3 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12275; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18419 = 12'hbf3 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15347; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21491 = 12'hbf3 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18419; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24563 = 12'hbf3 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21491; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27635 = 12'hbf3 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24563; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3059 = io_valid_in ? _GEN_27635 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3059 = 12'hbf3 == _T_2[11:0] ? image_3059 : _GEN_3058; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6132 = 12'hbf4 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9204 = 12'hbf4 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6132; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12276 = 12'hbf4 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9204; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15348 = 12'hbf4 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12276; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18420 = 12'hbf4 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15348; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21492 = 12'hbf4 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18420; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24564 = 12'hbf4 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21492; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27636 = 12'hbf4 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24564; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3060 = io_valid_in ? _GEN_27636 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3060 = 12'hbf4 == _T_2[11:0] ? image_3060 : _GEN_3059; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6133 = 12'hbf5 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9205 = 12'hbf5 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6133; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12277 = 12'hbf5 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9205; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15349 = 12'hbf5 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12277; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18421 = 12'hbf5 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15349; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21493 = 12'hbf5 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18421; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24565 = 12'hbf5 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21493; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27637 = 12'hbf5 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24565; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3061 = io_valid_in ? _GEN_27637 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3061 = 12'hbf5 == _T_2[11:0] ? image_3061 : _GEN_3060; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6134 = 12'hbf6 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9206 = 12'hbf6 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6134; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12278 = 12'hbf6 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9206; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15350 = 12'hbf6 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12278; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18422 = 12'hbf6 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15350; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21494 = 12'hbf6 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18422; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24566 = 12'hbf6 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21494; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27638 = 12'hbf6 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24566; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3062 = io_valid_in ? _GEN_27638 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3062 = 12'hbf6 == _T_2[11:0] ? image_3062 : _GEN_3061; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6135 = 12'hbf7 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9207 = 12'hbf7 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6135; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12279 = 12'hbf7 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9207; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15351 = 12'hbf7 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12279; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18423 = 12'hbf7 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15351; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21495 = 12'hbf7 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18423; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24567 = 12'hbf7 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21495; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27639 = 12'hbf7 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24567; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3063 = io_valid_in ? _GEN_27639 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3063 = 12'hbf7 == _T_2[11:0] ? image_3063 : _GEN_3062; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6136 = 12'hbf8 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9208 = 12'hbf8 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6136; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12280 = 12'hbf8 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9208; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15352 = 12'hbf8 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12280; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18424 = 12'hbf8 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15352; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21496 = 12'hbf8 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18424; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24568 = 12'hbf8 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21496; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27640 = 12'hbf8 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24568; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3064 = io_valid_in ? _GEN_27640 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3064 = 12'hbf8 == _T_2[11:0] ? image_3064 : _GEN_3063; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6137 = 12'hbf9 == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9209 = 12'hbf9 == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6137; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12281 = 12'hbf9 == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9209; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15353 = 12'hbf9 == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12281; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18425 = 12'hbf9 == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15353; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21497 = 12'hbf9 == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18425; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24569 = 12'hbf9 == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21497; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27641 = 12'hbf9 == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24569; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3065 = io_valid_in ? _GEN_27641 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3065 = 12'hbf9 == _T_2[11:0] ? image_3065 : _GEN_3064; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6138 = 12'hbfa == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9210 = 12'hbfa == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6138; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12282 = 12'hbfa == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9210; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15354 = 12'hbfa == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12282; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18426 = 12'hbfa == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15354; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21498 = 12'hbfa == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18426; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24570 = 12'hbfa == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21498; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27642 = 12'hbfa == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24570; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3066 = io_valid_in ? _GEN_27642 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3066 = 12'hbfa == _T_2[11:0] ? image_3066 : _GEN_3065; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6139 = 12'hbfb == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9211 = 12'hbfb == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6139; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12283 = 12'hbfb == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9211; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15355 = 12'hbfb == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12283; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18427 = 12'hbfb == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15355; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21499 = 12'hbfb == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18427; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24571 = 12'hbfb == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21499; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27643 = 12'hbfb == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24571; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3067 = io_valid_in ? _GEN_27643 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3067 = 12'hbfb == _T_2[11:0] ? image_3067 : _GEN_3066; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6140 = 12'hbfc == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9212 = 12'hbfc == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6140; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12284 = 12'hbfc == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9212; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15356 = 12'hbfc == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12284; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18428 = 12'hbfc == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15356; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21500 = 12'hbfc == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18428; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24572 = 12'hbfc == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21500; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27644 = 12'hbfc == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24572; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3068 = io_valid_in ? _GEN_27644 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3068 = 12'hbfc == _T_2[11:0] ? image_3068 : _GEN_3067; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6141 = 12'hbfd == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9213 = 12'hbfd == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6141; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12285 = 12'hbfd == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9213; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15357 = 12'hbfd == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12285; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18429 = 12'hbfd == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15357; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21501 = 12'hbfd == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18429; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24573 = 12'hbfd == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21501; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27645 = 12'hbfd == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24573; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3069 = io_valid_in ? _GEN_27645 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3069 = 12'hbfd == _T_2[11:0] ? image_3069 : _GEN_3068; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6142 = 12'hbfe == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9214 = 12'hbfe == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6142; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12286 = 12'hbfe == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9214; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15358 = 12'hbfe == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12286; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18430 = 12'hbfe == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15358; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21502 = 12'hbfe == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18430; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24574 = 12'hbfe == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21502; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27646 = 12'hbfe == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24574; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3070 = io_valid_in ? _GEN_27646 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3070 = 12'hbfe == _T_2[11:0] ? image_3070 : _GEN_3069; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_6143 = 12'hbff == _T_4[11:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_9215 = 12'hbff == _T_8[11:0] ? io_pixelVal_in_1 : _GEN_6143; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_12287 = 12'hbff == _T_11[11:0] ? io_pixelVal_in_2 : _GEN_9215; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_15359 = 12'hbff == _T_14[11:0] ? io_pixelVal_in_3 : _GEN_12287; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_18431 = 12'hbff == _T_17[11:0] ? io_pixelVal_in_4 : _GEN_15359; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_21503 = 12'hbff == _T_20[11:0] ? io_pixelVal_in_5 : _GEN_18431; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_24575 = 12'hbff == _T_23[11:0] ? io_pixelVal_in_6 : _GEN_21503; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_27647 = 12'hbff == _T_26[11:0] ? io_pixelVal_in_7 : _GEN_24575; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3071 = io_valid_in ? _GEN_27647 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [31:0] _T_29 = pixelIndex + 32'h8; // @[VideoBuffer.scala 37:42]
  wire [12:0] _T_30 = 7'h40 * 7'h30; // @[VideoBuffer.scala 38:42]
  wire [31:0] _GEN_30723 = {{19'd0}, _T_30}; // @[VideoBuffer.scala 38:25]
  wire  _T_31 = pixelIndex == _GEN_30723; // @[VideoBuffer.scala 38:25]
  assign io_pixelVal_out = 12'hbff == _T_2[11:0] ? image_3071 : _GEN_3070; // @[VideoBuffer.scala 29:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pixelIndex = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      pixelIndex <= 32'h0;
    end else if (io_valid_in) begin
      if (_T_31) begin
        pixelIndex <= 32'h0;
      end else begin
        pixelIndex <= _T_29;
      end
    end
  end
endmodule
