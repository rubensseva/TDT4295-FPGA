module DotProd(
  input        clock,
  input        reset,
  input  [7:0] io_dataInA,
  input  [7:0] io_dataInB,
  output [8:0] io_dataOut,
  output       io_outputValid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] countVal; // @[Counter.scala 29:33]
  wire  countReset = countVal == 4'h8; // @[Counter.scala 38:24]
  wire [3:0] _T_2 = countVal + 4'h1; // @[Counter.scala 39:22]
  reg [8:0] accumulator; // @[DotProd.scala 19:28]
  wire [15:0] product = $signed(io_dataInA) * $signed(io_dataInB); // @[DotProd.scala 20:35]
  wire [15:0] _GEN_5 = {{7{accumulator[8]}},accumulator}; // @[DotProd.scala 21:30]
  wire [15:0] _T_6 = $signed(_GEN_5) + $signed(product); // @[DotProd.scala 21:30]
  wire  _T_11 = ~reset; // @[DotProd.scala 29:11]
  wire [15:0] _GEN_4 = countReset ? $signed(16'sh0) : $signed(_T_6); // @[DotProd.scala 25:20]
  assign io_dataOut = _T_6[8:0]; // @[DotProd.scala 23:14]
  assign io_outputValid = countVal == 4'h8; // @[DotProd.scala 26:20 DotProd.scala 31:20]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  countVal = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  accumulator = _RAND_1[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      countVal <= 4'h0;
    end else if (countReset) begin
      countVal <= 4'h0;
    end else begin
      countVal <= _T_2;
    end
    if (reset) begin
      accumulator <= 9'sh0;
    end else begin
      accumulator <= _GEN_4[8:0];
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (countReset & _T_11) begin
          $fwrite(32'h80000002,"VALOUTidghspdolgnfgkln\n"); // @[DotProd.scala 29:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module KernelConvolution(
  input        clock,
  input        reset,
  input  [4:0] io_kernelVal_in,
  input  [3:0] io_pixelVal_in_0,
  input  [3:0] io_pixelVal_in_1,
  input  [3:0] io_pixelVal_in_2,
  input  [3:0] io_pixelVal_in_3,
  input  [3:0] io_pixelVal_in_4,
  input  [3:0] io_pixelVal_in_5,
  input  [3:0] io_pixelVal_in_6,
  input  [3:0] io_pixelVal_in_7,
  output [8:0] io_pixelVal_out_0,
  output [8:0] io_pixelVal_out_1,
  output [8:0] io_pixelVal_out_2,
  output [8:0] io_pixelVal_out_3,
  output [8:0] io_pixelVal_out_4,
  output [8:0] io_pixelVal_out_5,
  output [8:0] io_pixelVal_out_6,
  output [8:0] io_pixelVal_out_7,
  output       io_valid_out
);
  wire  DotProd_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_1_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_1_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_1_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_1_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_1_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_1_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_2_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_2_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_2_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_2_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_2_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_2_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_3_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_3_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_3_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_3_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_3_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_3_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_4_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_4_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_4_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_4_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_4_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_4_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_5_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_5_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_5_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_5_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_5_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_5_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_6_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_6_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_6_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_6_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_6_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_6_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_7_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_7_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_7_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_7_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_7_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_7_io_outputValid; // @[KernelConvolution.scala 21:58]
  DotProd DotProd ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_clock),
    .reset(DotProd_reset),
    .io_dataInA(DotProd_io_dataInA),
    .io_dataInB(DotProd_io_dataInB),
    .io_dataOut(DotProd_io_dataOut),
    .io_outputValid(DotProd_io_outputValid)
  );
  DotProd DotProd_1 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_1_clock),
    .reset(DotProd_1_reset),
    .io_dataInA(DotProd_1_io_dataInA),
    .io_dataInB(DotProd_1_io_dataInB),
    .io_dataOut(DotProd_1_io_dataOut),
    .io_outputValid(DotProd_1_io_outputValid)
  );
  DotProd DotProd_2 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_2_clock),
    .reset(DotProd_2_reset),
    .io_dataInA(DotProd_2_io_dataInA),
    .io_dataInB(DotProd_2_io_dataInB),
    .io_dataOut(DotProd_2_io_dataOut),
    .io_outputValid(DotProd_2_io_outputValid)
  );
  DotProd DotProd_3 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_3_clock),
    .reset(DotProd_3_reset),
    .io_dataInA(DotProd_3_io_dataInA),
    .io_dataInB(DotProd_3_io_dataInB),
    .io_dataOut(DotProd_3_io_dataOut),
    .io_outputValid(DotProd_3_io_outputValid)
  );
  DotProd DotProd_4 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_4_clock),
    .reset(DotProd_4_reset),
    .io_dataInA(DotProd_4_io_dataInA),
    .io_dataInB(DotProd_4_io_dataInB),
    .io_dataOut(DotProd_4_io_dataOut),
    .io_outputValid(DotProd_4_io_outputValid)
  );
  DotProd DotProd_5 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_5_clock),
    .reset(DotProd_5_reset),
    .io_dataInA(DotProd_5_io_dataInA),
    .io_dataInB(DotProd_5_io_dataInB),
    .io_dataOut(DotProd_5_io_dataOut),
    .io_outputValid(DotProd_5_io_outputValid)
  );
  DotProd DotProd_6 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_6_clock),
    .reset(DotProd_6_reset),
    .io_dataInA(DotProd_6_io_dataInA),
    .io_dataInB(DotProd_6_io_dataInB),
    .io_dataOut(DotProd_6_io_dataOut),
    .io_outputValid(DotProd_6_io_outputValid)
  );
  DotProd DotProd_7 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_7_clock),
    .reset(DotProd_7_reset),
    .io_dataInA(DotProd_7_io_dataInA),
    .io_dataInB(DotProd_7_io_dataInB),
    .io_dataOut(DotProd_7_io_dataOut),
    .io_outputValid(DotProd_7_io_outputValid)
  );
  assign io_pixelVal_out_0 = DotProd_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_1 = DotProd_1_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_2 = DotProd_2_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_3 = DotProd_3_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_4 = DotProd_4_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_5 = DotProd_5_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_6 = DotProd_6_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_7 = DotProd_7_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_valid_out = DotProd_io_outputValid; // @[KernelConvolution.scala 35:30]
  assign DotProd_clock = clock;
  assign DotProd_reset = reset;
  assign DotProd_io_dataInA = {{4'd0}, io_pixelVal_in_0}; // @[KernelConvolution.scala 21:32]
  assign DotProd_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_1_clock = clock;
  assign DotProd_1_reset = reset;
  assign DotProd_1_io_dataInA = {{4'd0}, io_pixelVal_in_1}; // @[KernelConvolution.scala 21:32]
  assign DotProd_1_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_2_clock = clock;
  assign DotProd_2_reset = reset;
  assign DotProd_2_io_dataInA = {{4'd0}, io_pixelVal_in_2}; // @[KernelConvolution.scala 21:32]
  assign DotProd_2_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_3_clock = clock;
  assign DotProd_3_reset = reset;
  assign DotProd_3_io_dataInA = {{4'd0}, io_pixelVal_in_3}; // @[KernelConvolution.scala 21:32]
  assign DotProd_3_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_4_clock = clock;
  assign DotProd_4_reset = reset;
  assign DotProd_4_io_dataInA = {{4'd0}, io_pixelVal_in_4}; // @[KernelConvolution.scala 21:32]
  assign DotProd_4_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_5_clock = clock;
  assign DotProd_5_reset = reset;
  assign DotProd_5_io_dataInA = {{4'd0}, io_pixelVal_in_5}; // @[KernelConvolution.scala 21:32]
  assign DotProd_5_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_6_clock = clock;
  assign DotProd_6_reset = reset;
  assign DotProd_6_io_dataInA = {{4'd0}, io_pixelVal_in_6}; // @[KernelConvolution.scala 21:32]
  assign DotProd_6_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_7_clock = clock;
  assign DotProd_7_reset = reset;
  assign DotProd_7_io_dataInA = {{4'd0}, io_pixelVal_in_7}; // @[KernelConvolution.scala 21:32]
  assign DotProd_7_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
endmodule
module Filter(
  input        clock,
  input        reset,
  input  [5:0] io_SPI_filterIndex,
  input        io_SPI_invert,
  input        io_SPI_distort,
  output [3:0] io_pixelVal_out_0,
  output [3:0] io_pixelVal_out_1,
  output [3:0] io_pixelVal_out_2,
  output [3:0] io_pixelVal_out_3,
  output [3:0] io_pixelVal_out_4,
  output [3:0] io_pixelVal_out_5,
  output [3:0] io_pixelVal_out_6,
  output [3:0] io_pixelVal_out_7,
  output       io_valid_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1041;
  reg [31:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1045;
  reg [31:0] _RAND_1046;
  reg [31:0] _RAND_1047;
  reg [31:0] _RAND_1048;
  reg [31:0] _RAND_1049;
  reg [31:0] _RAND_1050;
  reg [31:0] _RAND_1051;
  reg [31:0] _RAND_1052;
  reg [31:0] _RAND_1053;
  reg [31:0] _RAND_1054;
  reg [31:0] _RAND_1055;
  reg [31:0] _RAND_1056;
  reg [31:0] _RAND_1057;
  reg [31:0] _RAND_1058;
  reg [31:0] _RAND_1059;
  reg [31:0] _RAND_1060;
  reg [31:0] _RAND_1061;
  reg [31:0] _RAND_1062;
  reg [31:0] _RAND_1063;
  reg [31:0] _RAND_1064;
  reg [31:0] _RAND_1065;
  reg [31:0] _RAND_1066;
  reg [31:0] _RAND_1067;
  reg [31:0] _RAND_1068;
  reg [31:0] _RAND_1069;
  reg [31:0] _RAND_1070;
  reg [31:0] _RAND_1071;
  reg [31:0] _RAND_1072;
  reg [31:0] _RAND_1073;
  reg [31:0] _RAND_1074;
  reg [31:0] _RAND_1075;
  reg [31:0] _RAND_1076;
  reg [31:0] _RAND_1077;
  reg [31:0] _RAND_1078;
  reg [31:0] _RAND_1079;
  reg [31:0] _RAND_1080;
  reg [31:0] _RAND_1081;
  reg [31:0] _RAND_1082;
  reg [31:0] _RAND_1083;
  reg [31:0] _RAND_1084;
  reg [31:0] _RAND_1085;
  reg [31:0] _RAND_1086;
  reg [31:0] _RAND_1087;
  reg [31:0] _RAND_1088;
  reg [31:0] _RAND_1089;
  reg [31:0] _RAND_1090;
  reg [31:0] _RAND_1091;
  reg [31:0] _RAND_1092;
  reg [31:0] _RAND_1093;
  reg [31:0] _RAND_1094;
  reg [31:0] _RAND_1095;
  reg [31:0] _RAND_1096;
  reg [31:0] _RAND_1097;
  reg [31:0] _RAND_1098;
  reg [31:0] _RAND_1099;
  reg [31:0] _RAND_1100;
  reg [31:0] _RAND_1101;
  reg [31:0] _RAND_1102;
  reg [31:0] _RAND_1103;
  reg [31:0] _RAND_1104;
  reg [31:0] _RAND_1105;
  reg [31:0] _RAND_1106;
  reg [31:0] _RAND_1107;
  reg [31:0] _RAND_1108;
  reg [31:0] _RAND_1109;
  reg [31:0] _RAND_1110;
  reg [31:0] _RAND_1111;
  reg [31:0] _RAND_1112;
  reg [31:0] _RAND_1113;
  reg [31:0] _RAND_1114;
  reg [31:0] _RAND_1115;
  reg [31:0] _RAND_1116;
  reg [31:0] _RAND_1117;
  reg [31:0] _RAND_1118;
  reg [31:0] _RAND_1119;
  reg [31:0] _RAND_1120;
  reg [31:0] _RAND_1121;
  reg [31:0] _RAND_1122;
  reg [31:0] _RAND_1123;
  reg [31:0] _RAND_1124;
  reg [31:0] _RAND_1125;
  reg [31:0] _RAND_1126;
  reg [31:0] _RAND_1127;
  reg [31:0] _RAND_1128;
  reg [31:0] _RAND_1129;
  reg [31:0] _RAND_1130;
  reg [31:0] _RAND_1131;
  reg [31:0] _RAND_1132;
  reg [31:0] _RAND_1133;
  reg [31:0] _RAND_1134;
  reg [31:0] _RAND_1135;
  reg [31:0] _RAND_1136;
  reg [31:0] _RAND_1137;
  reg [31:0] _RAND_1138;
  reg [31:0] _RAND_1139;
  reg [31:0] _RAND_1140;
  reg [31:0] _RAND_1141;
  reg [31:0] _RAND_1142;
  reg [31:0] _RAND_1143;
  reg [31:0] _RAND_1144;
  reg [31:0] _RAND_1145;
  reg [31:0] _RAND_1146;
  reg [31:0] _RAND_1147;
  reg [31:0] _RAND_1148;
  reg [31:0] _RAND_1149;
  reg [31:0] _RAND_1150;
  reg [31:0] _RAND_1151;
  reg [31:0] _RAND_1152;
  reg [31:0] _RAND_1153;
  reg [31:0] _RAND_1154;
  reg [31:0] _RAND_1155;
  reg [31:0] _RAND_1156;
  reg [31:0] _RAND_1157;
  reg [31:0] _RAND_1158;
  reg [31:0] _RAND_1159;
  reg [31:0] _RAND_1160;
  reg [31:0] _RAND_1161;
  reg [31:0] _RAND_1162;
  reg [31:0] _RAND_1163;
  reg [31:0] _RAND_1164;
  reg [31:0] _RAND_1165;
  reg [31:0] _RAND_1166;
  reg [31:0] _RAND_1167;
  reg [31:0] _RAND_1168;
  reg [31:0] _RAND_1169;
  reg [31:0] _RAND_1170;
  reg [31:0] _RAND_1171;
  reg [31:0] _RAND_1172;
  reg [31:0] _RAND_1173;
  reg [31:0] _RAND_1174;
  reg [31:0] _RAND_1175;
  reg [31:0] _RAND_1176;
  reg [31:0] _RAND_1177;
  reg [31:0] _RAND_1178;
  reg [31:0] _RAND_1179;
  reg [31:0] _RAND_1180;
  reg [31:0] _RAND_1181;
  reg [31:0] _RAND_1182;
  reg [31:0] _RAND_1183;
  reg [31:0] _RAND_1184;
  reg [31:0] _RAND_1185;
  reg [31:0] _RAND_1186;
  reg [31:0] _RAND_1187;
  reg [31:0] _RAND_1188;
  reg [31:0] _RAND_1189;
  reg [31:0] _RAND_1190;
  reg [31:0] _RAND_1191;
  reg [31:0] _RAND_1192;
  reg [31:0] _RAND_1193;
  reg [31:0] _RAND_1194;
  reg [31:0] _RAND_1195;
  reg [31:0] _RAND_1196;
  reg [31:0] _RAND_1197;
  reg [31:0] _RAND_1198;
  reg [31:0] _RAND_1199;
  reg [31:0] _RAND_1200;
  reg [31:0] _RAND_1201;
  reg [31:0] _RAND_1202;
  reg [31:0] _RAND_1203;
  reg [31:0] _RAND_1204;
  reg [31:0] _RAND_1205;
  reg [31:0] _RAND_1206;
  reg [31:0] _RAND_1207;
  reg [31:0] _RAND_1208;
  reg [31:0] _RAND_1209;
  reg [31:0] _RAND_1210;
  reg [31:0] _RAND_1211;
  reg [31:0] _RAND_1212;
  reg [31:0] _RAND_1213;
  reg [31:0] _RAND_1214;
  reg [31:0] _RAND_1215;
  reg [31:0] _RAND_1216;
  reg [31:0] _RAND_1217;
  reg [31:0] _RAND_1218;
  reg [31:0] _RAND_1219;
  reg [31:0] _RAND_1220;
  reg [31:0] _RAND_1221;
  reg [31:0] _RAND_1222;
  reg [31:0] _RAND_1223;
  reg [31:0] _RAND_1224;
  reg [31:0] _RAND_1225;
  reg [31:0] _RAND_1226;
  reg [31:0] _RAND_1227;
  reg [31:0] _RAND_1228;
  reg [31:0] _RAND_1229;
  reg [31:0] _RAND_1230;
  reg [31:0] _RAND_1231;
  reg [31:0] _RAND_1232;
  reg [31:0] _RAND_1233;
  reg [31:0] _RAND_1234;
  reg [31:0] _RAND_1235;
  reg [31:0] _RAND_1236;
  reg [31:0] _RAND_1237;
  reg [31:0] _RAND_1238;
  reg [31:0] _RAND_1239;
  reg [31:0] _RAND_1240;
  reg [31:0] _RAND_1241;
  reg [31:0] _RAND_1242;
  reg [31:0] _RAND_1243;
  reg [31:0] _RAND_1244;
  reg [31:0] _RAND_1245;
  reg [31:0] _RAND_1246;
  reg [31:0] _RAND_1247;
  reg [31:0] _RAND_1248;
  reg [31:0] _RAND_1249;
  reg [31:0] _RAND_1250;
  reg [31:0] _RAND_1251;
  reg [31:0] _RAND_1252;
  reg [31:0] _RAND_1253;
  reg [31:0] _RAND_1254;
  reg [31:0] _RAND_1255;
  reg [31:0] _RAND_1256;
  reg [31:0] _RAND_1257;
  reg [31:0] _RAND_1258;
  reg [31:0] _RAND_1259;
  reg [31:0] _RAND_1260;
  reg [31:0] _RAND_1261;
  reg [31:0] _RAND_1262;
  reg [31:0] _RAND_1263;
  reg [31:0] _RAND_1264;
  reg [31:0] _RAND_1265;
  reg [31:0] _RAND_1266;
  reg [31:0] _RAND_1267;
  reg [31:0] _RAND_1268;
  reg [31:0] _RAND_1269;
  reg [31:0] _RAND_1270;
  reg [31:0] _RAND_1271;
  reg [31:0] _RAND_1272;
  reg [31:0] _RAND_1273;
  reg [31:0] _RAND_1274;
  reg [31:0] _RAND_1275;
  reg [31:0] _RAND_1276;
  reg [31:0] _RAND_1277;
  reg [31:0] _RAND_1278;
  reg [31:0] _RAND_1279;
  reg [31:0] _RAND_1280;
  reg [31:0] _RAND_1281;
  reg [31:0] _RAND_1282;
  reg [31:0] _RAND_1283;
  reg [31:0] _RAND_1284;
  reg [31:0] _RAND_1285;
  reg [31:0] _RAND_1286;
  reg [31:0] _RAND_1287;
  reg [31:0] _RAND_1288;
  reg [31:0] _RAND_1289;
  reg [31:0] _RAND_1290;
  reg [31:0] _RAND_1291;
  reg [31:0] _RAND_1292;
  reg [31:0] _RAND_1293;
  reg [31:0] _RAND_1294;
  reg [31:0] _RAND_1295;
  reg [31:0] _RAND_1296;
  reg [31:0] _RAND_1297;
  reg [31:0] _RAND_1298;
  reg [31:0] _RAND_1299;
  reg [31:0] _RAND_1300;
  reg [31:0] _RAND_1301;
  reg [31:0] _RAND_1302;
  reg [31:0] _RAND_1303;
  reg [31:0] _RAND_1304;
  reg [31:0] _RAND_1305;
  reg [31:0] _RAND_1306;
  reg [31:0] _RAND_1307;
  reg [31:0] _RAND_1308;
  reg [31:0] _RAND_1309;
  reg [31:0] _RAND_1310;
  reg [31:0] _RAND_1311;
  reg [31:0] _RAND_1312;
  reg [31:0] _RAND_1313;
  reg [31:0] _RAND_1314;
  reg [31:0] _RAND_1315;
  reg [31:0] _RAND_1316;
  reg [31:0] _RAND_1317;
  reg [31:0] _RAND_1318;
  reg [31:0] _RAND_1319;
  reg [31:0] _RAND_1320;
  reg [31:0] _RAND_1321;
  reg [31:0] _RAND_1322;
  reg [31:0] _RAND_1323;
  reg [31:0] _RAND_1324;
  reg [31:0] _RAND_1325;
  reg [31:0] _RAND_1326;
  reg [31:0] _RAND_1327;
  reg [31:0] _RAND_1328;
  reg [31:0] _RAND_1329;
  reg [31:0] _RAND_1330;
  reg [31:0] _RAND_1331;
  reg [31:0] _RAND_1332;
  reg [31:0] _RAND_1333;
  reg [31:0] _RAND_1334;
  reg [31:0] _RAND_1335;
  reg [31:0] _RAND_1336;
  reg [31:0] _RAND_1337;
  reg [31:0] _RAND_1338;
  reg [31:0] _RAND_1339;
  reg [31:0] _RAND_1340;
  reg [31:0] _RAND_1341;
  reg [31:0] _RAND_1342;
  reg [31:0] _RAND_1343;
  reg [31:0] _RAND_1344;
  reg [31:0] _RAND_1345;
  reg [31:0] _RAND_1346;
  reg [31:0] _RAND_1347;
  reg [31:0] _RAND_1348;
  reg [31:0] _RAND_1349;
  reg [31:0] _RAND_1350;
  reg [31:0] _RAND_1351;
  reg [31:0] _RAND_1352;
  reg [31:0] _RAND_1353;
  reg [31:0] _RAND_1354;
  reg [31:0] _RAND_1355;
  reg [31:0] _RAND_1356;
  reg [31:0] _RAND_1357;
  reg [31:0] _RAND_1358;
  reg [31:0] _RAND_1359;
  reg [31:0] _RAND_1360;
  reg [31:0] _RAND_1361;
  reg [31:0] _RAND_1362;
  reg [31:0] _RAND_1363;
  reg [31:0] _RAND_1364;
  reg [31:0] _RAND_1365;
  reg [31:0] _RAND_1366;
  reg [31:0] _RAND_1367;
  reg [31:0] _RAND_1368;
  reg [31:0] _RAND_1369;
  reg [31:0] _RAND_1370;
  reg [31:0] _RAND_1371;
  reg [31:0] _RAND_1372;
  reg [31:0] _RAND_1373;
  reg [31:0] _RAND_1374;
  reg [31:0] _RAND_1375;
  reg [31:0] _RAND_1376;
  reg [31:0] _RAND_1377;
  reg [31:0] _RAND_1378;
  reg [31:0] _RAND_1379;
  reg [31:0] _RAND_1380;
  reg [31:0] _RAND_1381;
  reg [31:0] _RAND_1382;
  reg [31:0] _RAND_1383;
  reg [31:0] _RAND_1384;
  reg [31:0] _RAND_1385;
  reg [31:0] _RAND_1386;
  reg [31:0] _RAND_1387;
  reg [31:0] _RAND_1388;
  reg [31:0] _RAND_1389;
  reg [31:0] _RAND_1390;
  reg [31:0] _RAND_1391;
  reg [31:0] _RAND_1392;
  reg [31:0] _RAND_1393;
  reg [31:0] _RAND_1394;
  reg [31:0] _RAND_1395;
  reg [31:0] _RAND_1396;
  reg [31:0] _RAND_1397;
  reg [31:0] _RAND_1398;
  reg [31:0] _RAND_1399;
  reg [31:0] _RAND_1400;
  reg [31:0] _RAND_1401;
  reg [31:0] _RAND_1402;
  reg [31:0] _RAND_1403;
  reg [31:0] _RAND_1404;
  reg [31:0] _RAND_1405;
  reg [31:0] _RAND_1406;
  reg [31:0] _RAND_1407;
  reg [31:0] _RAND_1408;
  reg [31:0] _RAND_1409;
  reg [31:0] _RAND_1410;
  reg [31:0] _RAND_1411;
  reg [31:0] _RAND_1412;
  reg [31:0] _RAND_1413;
  reg [31:0] _RAND_1414;
  reg [31:0] _RAND_1415;
  reg [31:0] _RAND_1416;
  reg [31:0] _RAND_1417;
  reg [31:0] _RAND_1418;
  reg [31:0] _RAND_1419;
  reg [31:0] _RAND_1420;
  reg [31:0] _RAND_1421;
  reg [31:0] _RAND_1422;
  reg [31:0] _RAND_1423;
  reg [31:0] _RAND_1424;
  reg [31:0] _RAND_1425;
  reg [31:0] _RAND_1426;
  reg [31:0] _RAND_1427;
  reg [31:0] _RAND_1428;
  reg [31:0] _RAND_1429;
  reg [31:0] _RAND_1430;
  reg [31:0] _RAND_1431;
  reg [31:0] _RAND_1432;
  reg [31:0] _RAND_1433;
  reg [31:0] _RAND_1434;
  reg [31:0] _RAND_1435;
  reg [31:0] _RAND_1436;
  reg [31:0] _RAND_1437;
  reg [31:0] _RAND_1438;
  reg [31:0] _RAND_1439;
  reg [31:0] _RAND_1440;
  reg [31:0] _RAND_1441;
  reg [31:0] _RAND_1442;
  reg [31:0] _RAND_1443;
  reg [31:0] _RAND_1444;
  reg [31:0] _RAND_1445;
  reg [31:0] _RAND_1446;
  reg [31:0] _RAND_1447;
  reg [31:0] _RAND_1448;
  reg [31:0] _RAND_1449;
  reg [31:0] _RAND_1450;
  reg [31:0] _RAND_1451;
  reg [31:0] _RAND_1452;
  reg [31:0] _RAND_1453;
  reg [31:0] _RAND_1454;
  reg [31:0] _RAND_1455;
  reg [31:0] _RAND_1456;
  reg [31:0] _RAND_1457;
  reg [31:0] _RAND_1458;
  reg [31:0] _RAND_1459;
  reg [31:0] _RAND_1460;
  reg [31:0] _RAND_1461;
  reg [31:0] _RAND_1462;
  reg [31:0] _RAND_1463;
  reg [31:0] _RAND_1464;
  reg [31:0] _RAND_1465;
  reg [31:0] _RAND_1466;
  reg [31:0] _RAND_1467;
  reg [31:0] _RAND_1468;
  reg [31:0] _RAND_1469;
  reg [31:0] _RAND_1470;
  reg [31:0] _RAND_1471;
  reg [31:0] _RAND_1472;
  reg [31:0] _RAND_1473;
  reg [31:0] _RAND_1474;
  reg [31:0] _RAND_1475;
  reg [31:0] _RAND_1476;
  reg [31:0] _RAND_1477;
  reg [31:0] _RAND_1478;
  reg [31:0] _RAND_1479;
  reg [31:0] _RAND_1480;
  reg [31:0] _RAND_1481;
  reg [31:0] _RAND_1482;
  reg [31:0] _RAND_1483;
  reg [31:0] _RAND_1484;
  reg [31:0] _RAND_1485;
  reg [31:0] _RAND_1486;
  reg [31:0] _RAND_1487;
  reg [31:0] _RAND_1488;
  reg [31:0] _RAND_1489;
  reg [31:0] _RAND_1490;
  reg [31:0] _RAND_1491;
  reg [31:0] _RAND_1492;
  reg [31:0] _RAND_1493;
  reg [31:0] _RAND_1494;
  reg [31:0] _RAND_1495;
  reg [31:0] _RAND_1496;
  reg [31:0] _RAND_1497;
  reg [31:0] _RAND_1498;
  reg [31:0] _RAND_1499;
  reg [31:0] _RAND_1500;
  reg [31:0] _RAND_1501;
  reg [31:0] _RAND_1502;
  reg [31:0] _RAND_1503;
  reg [31:0] _RAND_1504;
  reg [31:0] _RAND_1505;
  reg [31:0] _RAND_1506;
  reg [31:0] _RAND_1507;
  reg [31:0] _RAND_1508;
  reg [31:0] _RAND_1509;
  reg [31:0] _RAND_1510;
  reg [31:0] _RAND_1511;
  reg [31:0] _RAND_1512;
  reg [31:0] _RAND_1513;
  reg [31:0] _RAND_1514;
  reg [31:0] _RAND_1515;
  reg [31:0] _RAND_1516;
  reg [31:0] _RAND_1517;
  reg [31:0] _RAND_1518;
  reg [31:0] _RAND_1519;
  reg [31:0] _RAND_1520;
  reg [31:0] _RAND_1521;
  reg [31:0] _RAND_1522;
  reg [31:0] _RAND_1523;
  reg [31:0] _RAND_1524;
  reg [31:0] _RAND_1525;
  reg [31:0] _RAND_1526;
  reg [31:0] _RAND_1527;
  reg [31:0] _RAND_1528;
  reg [31:0] _RAND_1529;
  reg [31:0] _RAND_1530;
  reg [31:0] _RAND_1531;
  reg [31:0] _RAND_1532;
  reg [31:0] _RAND_1533;
  reg [31:0] _RAND_1534;
  reg [31:0] _RAND_1535;
  reg [31:0] _RAND_1536;
  reg [31:0] _RAND_1537;
  reg [31:0] _RAND_1538;
  reg [31:0] _RAND_1539;
  reg [31:0] _RAND_1540;
  reg [31:0] _RAND_1541;
  reg [31:0] _RAND_1542;
  reg [31:0] _RAND_1543;
  reg [31:0] _RAND_1544;
  reg [31:0] _RAND_1545;
  reg [31:0] _RAND_1546;
  reg [31:0] _RAND_1547;
  reg [31:0] _RAND_1548;
  reg [31:0] _RAND_1549;
  reg [31:0] _RAND_1550;
  reg [31:0] _RAND_1551;
  reg [31:0] _RAND_1552;
  reg [31:0] _RAND_1553;
  reg [31:0] _RAND_1554;
  reg [31:0] _RAND_1555;
  reg [31:0] _RAND_1556;
  reg [31:0] _RAND_1557;
  reg [31:0] _RAND_1558;
  reg [31:0] _RAND_1559;
  reg [31:0] _RAND_1560;
  reg [31:0] _RAND_1561;
  reg [31:0] _RAND_1562;
  reg [31:0] _RAND_1563;
  reg [31:0] _RAND_1564;
  reg [31:0] _RAND_1565;
  reg [31:0] _RAND_1566;
  reg [31:0] _RAND_1567;
  reg [31:0] _RAND_1568;
  reg [31:0] _RAND_1569;
  reg [31:0] _RAND_1570;
  reg [31:0] _RAND_1571;
  reg [31:0] _RAND_1572;
  reg [31:0] _RAND_1573;
  reg [31:0] _RAND_1574;
  reg [31:0] _RAND_1575;
  reg [31:0] _RAND_1576;
  reg [31:0] _RAND_1577;
  reg [31:0] _RAND_1578;
  reg [31:0] _RAND_1579;
  reg [31:0] _RAND_1580;
  reg [31:0] _RAND_1581;
  reg [31:0] _RAND_1582;
  reg [31:0] _RAND_1583;
  reg [31:0] _RAND_1584;
  reg [31:0] _RAND_1585;
  reg [31:0] _RAND_1586;
  reg [31:0] _RAND_1587;
  reg [31:0] _RAND_1588;
  reg [31:0] _RAND_1589;
  reg [31:0] _RAND_1590;
  reg [31:0] _RAND_1591;
  reg [31:0] _RAND_1592;
  reg [31:0] _RAND_1593;
  reg [31:0] _RAND_1594;
  reg [31:0] _RAND_1595;
  reg [31:0] _RAND_1596;
  reg [31:0] _RAND_1597;
  reg [31:0] _RAND_1598;
  reg [31:0] _RAND_1599;
  reg [31:0] _RAND_1600;
  reg [31:0] _RAND_1601;
  reg [31:0] _RAND_1602;
  reg [31:0] _RAND_1603;
  reg [31:0] _RAND_1604;
  reg [31:0] _RAND_1605;
  reg [31:0] _RAND_1606;
  reg [31:0] _RAND_1607;
  reg [31:0] _RAND_1608;
  reg [31:0] _RAND_1609;
  reg [31:0] _RAND_1610;
  reg [31:0] _RAND_1611;
  reg [31:0] _RAND_1612;
  reg [31:0] _RAND_1613;
  reg [31:0] _RAND_1614;
  reg [31:0] _RAND_1615;
  reg [31:0] _RAND_1616;
  reg [31:0] _RAND_1617;
  reg [31:0] _RAND_1618;
  reg [31:0] _RAND_1619;
  reg [31:0] _RAND_1620;
  reg [31:0] _RAND_1621;
  reg [31:0] _RAND_1622;
  reg [31:0] _RAND_1623;
  reg [31:0] _RAND_1624;
  reg [31:0] _RAND_1625;
  reg [31:0] _RAND_1626;
  reg [31:0] _RAND_1627;
  reg [31:0] _RAND_1628;
  reg [31:0] _RAND_1629;
  reg [31:0] _RAND_1630;
  reg [31:0] _RAND_1631;
  reg [31:0] _RAND_1632;
  reg [31:0] _RAND_1633;
  reg [31:0] _RAND_1634;
  reg [31:0] _RAND_1635;
  reg [31:0] _RAND_1636;
  reg [31:0] _RAND_1637;
  reg [31:0] _RAND_1638;
  reg [31:0] _RAND_1639;
  reg [31:0] _RAND_1640;
  reg [31:0] _RAND_1641;
  reg [31:0] _RAND_1642;
  reg [31:0] _RAND_1643;
  reg [31:0] _RAND_1644;
  reg [31:0] _RAND_1645;
  reg [31:0] _RAND_1646;
  reg [31:0] _RAND_1647;
  reg [31:0] _RAND_1648;
  reg [31:0] _RAND_1649;
  reg [31:0] _RAND_1650;
  reg [31:0] _RAND_1651;
  reg [31:0] _RAND_1652;
  reg [31:0] _RAND_1653;
  reg [31:0] _RAND_1654;
  reg [31:0] _RAND_1655;
  reg [31:0] _RAND_1656;
  reg [31:0] _RAND_1657;
  reg [31:0] _RAND_1658;
  reg [31:0] _RAND_1659;
  reg [31:0] _RAND_1660;
  reg [31:0] _RAND_1661;
  reg [31:0] _RAND_1662;
  reg [31:0] _RAND_1663;
  reg [31:0] _RAND_1664;
  reg [31:0] _RAND_1665;
  reg [31:0] _RAND_1666;
  reg [31:0] _RAND_1667;
  reg [31:0] _RAND_1668;
  reg [31:0] _RAND_1669;
  reg [31:0] _RAND_1670;
  reg [31:0] _RAND_1671;
  reg [31:0] _RAND_1672;
  reg [31:0] _RAND_1673;
  reg [31:0] _RAND_1674;
  reg [31:0] _RAND_1675;
  reg [31:0] _RAND_1676;
  reg [31:0] _RAND_1677;
  reg [31:0] _RAND_1678;
  reg [31:0] _RAND_1679;
  reg [31:0] _RAND_1680;
  reg [31:0] _RAND_1681;
  reg [31:0] _RAND_1682;
  reg [31:0] _RAND_1683;
  reg [31:0] _RAND_1684;
  reg [31:0] _RAND_1685;
  reg [31:0] _RAND_1686;
  reg [31:0] _RAND_1687;
  reg [31:0] _RAND_1688;
  reg [31:0] _RAND_1689;
  reg [31:0] _RAND_1690;
  reg [31:0] _RAND_1691;
  reg [31:0] _RAND_1692;
  reg [31:0] _RAND_1693;
  reg [31:0] _RAND_1694;
  reg [31:0] _RAND_1695;
  reg [31:0] _RAND_1696;
  reg [31:0] _RAND_1697;
  reg [31:0] _RAND_1698;
  reg [31:0] _RAND_1699;
  reg [31:0] _RAND_1700;
  reg [31:0] _RAND_1701;
  reg [31:0] _RAND_1702;
  reg [31:0] _RAND_1703;
  reg [31:0] _RAND_1704;
  reg [31:0] _RAND_1705;
  reg [31:0] _RAND_1706;
  reg [31:0] _RAND_1707;
  reg [31:0] _RAND_1708;
  reg [31:0] _RAND_1709;
  reg [31:0] _RAND_1710;
  reg [31:0] _RAND_1711;
  reg [31:0] _RAND_1712;
  reg [31:0] _RAND_1713;
  reg [31:0] _RAND_1714;
  reg [31:0] _RAND_1715;
  reg [31:0] _RAND_1716;
  reg [31:0] _RAND_1717;
  reg [31:0] _RAND_1718;
  reg [31:0] _RAND_1719;
  reg [31:0] _RAND_1720;
  reg [31:0] _RAND_1721;
  reg [31:0] _RAND_1722;
  reg [31:0] _RAND_1723;
  reg [31:0] _RAND_1724;
  reg [31:0] _RAND_1725;
  reg [31:0] _RAND_1726;
  reg [31:0] _RAND_1727;
  reg [31:0] _RAND_1728;
  reg [31:0] _RAND_1729;
  reg [31:0] _RAND_1730;
  reg [31:0] _RAND_1731;
  reg [31:0] _RAND_1732;
  reg [31:0] _RAND_1733;
  reg [31:0] _RAND_1734;
  reg [31:0] _RAND_1735;
  reg [31:0] _RAND_1736;
  reg [31:0] _RAND_1737;
  reg [31:0] _RAND_1738;
  reg [31:0] _RAND_1739;
  reg [31:0] _RAND_1740;
  reg [31:0] _RAND_1741;
  reg [31:0] _RAND_1742;
  reg [31:0] _RAND_1743;
  reg [31:0] _RAND_1744;
  reg [31:0] _RAND_1745;
  reg [31:0] _RAND_1746;
  reg [31:0] _RAND_1747;
  reg [31:0] _RAND_1748;
  reg [31:0] _RAND_1749;
  reg [31:0] _RAND_1750;
  reg [31:0] _RAND_1751;
  reg [31:0] _RAND_1752;
  reg [31:0] _RAND_1753;
  reg [31:0] _RAND_1754;
  reg [31:0] _RAND_1755;
  reg [31:0] _RAND_1756;
  reg [31:0] _RAND_1757;
  reg [31:0] _RAND_1758;
  reg [31:0] _RAND_1759;
  reg [31:0] _RAND_1760;
  reg [31:0] _RAND_1761;
  reg [31:0] _RAND_1762;
  reg [31:0] _RAND_1763;
  reg [31:0] _RAND_1764;
  reg [31:0] _RAND_1765;
  reg [31:0] _RAND_1766;
  reg [31:0] _RAND_1767;
  reg [31:0] _RAND_1768;
  reg [31:0] _RAND_1769;
  reg [31:0] _RAND_1770;
  reg [31:0] _RAND_1771;
  reg [31:0] _RAND_1772;
  reg [31:0] _RAND_1773;
  reg [31:0] _RAND_1774;
  reg [31:0] _RAND_1775;
  reg [31:0] _RAND_1776;
  reg [31:0] _RAND_1777;
  reg [31:0] _RAND_1778;
  reg [31:0] _RAND_1779;
  reg [31:0] _RAND_1780;
  reg [31:0] _RAND_1781;
  reg [31:0] _RAND_1782;
  reg [31:0] _RAND_1783;
  reg [31:0] _RAND_1784;
  reg [31:0] _RAND_1785;
  reg [31:0] _RAND_1786;
  reg [31:0] _RAND_1787;
  reg [31:0] _RAND_1788;
  reg [31:0] _RAND_1789;
  reg [31:0] _RAND_1790;
  reg [31:0] _RAND_1791;
  reg [31:0] _RAND_1792;
  reg [31:0] _RAND_1793;
  reg [31:0] _RAND_1794;
  reg [31:0] _RAND_1795;
  reg [31:0] _RAND_1796;
  reg [31:0] _RAND_1797;
  reg [31:0] _RAND_1798;
  reg [31:0] _RAND_1799;
  reg [31:0] _RAND_1800;
  reg [31:0] _RAND_1801;
  reg [31:0] _RAND_1802;
  reg [31:0] _RAND_1803;
  reg [31:0] _RAND_1804;
  reg [31:0] _RAND_1805;
  reg [31:0] _RAND_1806;
  reg [31:0] _RAND_1807;
  reg [31:0] _RAND_1808;
  reg [31:0] _RAND_1809;
  reg [31:0] _RAND_1810;
  reg [31:0] _RAND_1811;
  reg [31:0] _RAND_1812;
  reg [31:0] _RAND_1813;
  reg [31:0] _RAND_1814;
  reg [31:0] _RAND_1815;
  reg [31:0] _RAND_1816;
  reg [31:0] _RAND_1817;
  reg [31:0] _RAND_1818;
  reg [31:0] _RAND_1819;
  reg [31:0] _RAND_1820;
  reg [31:0] _RAND_1821;
  reg [31:0] _RAND_1822;
  reg [31:0] _RAND_1823;
  reg [31:0] _RAND_1824;
  reg [31:0] _RAND_1825;
  reg [31:0] _RAND_1826;
  reg [31:0] _RAND_1827;
  reg [31:0] _RAND_1828;
  reg [31:0] _RAND_1829;
  reg [31:0] _RAND_1830;
  reg [31:0] _RAND_1831;
  reg [31:0] _RAND_1832;
  reg [31:0] _RAND_1833;
  reg [31:0] _RAND_1834;
  reg [31:0] _RAND_1835;
  reg [31:0] _RAND_1836;
  reg [31:0] _RAND_1837;
  reg [31:0] _RAND_1838;
  reg [31:0] _RAND_1839;
  reg [31:0] _RAND_1840;
  reg [31:0] _RAND_1841;
  reg [31:0] _RAND_1842;
  reg [31:0] _RAND_1843;
  reg [31:0] _RAND_1844;
  reg [31:0] _RAND_1845;
  reg [31:0] _RAND_1846;
  reg [31:0] _RAND_1847;
  reg [31:0] _RAND_1848;
  reg [31:0] _RAND_1849;
  reg [31:0] _RAND_1850;
  reg [31:0] _RAND_1851;
  reg [31:0] _RAND_1852;
  reg [31:0] _RAND_1853;
  reg [31:0] _RAND_1854;
  reg [31:0] _RAND_1855;
  reg [31:0] _RAND_1856;
  reg [31:0] _RAND_1857;
  reg [31:0] _RAND_1858;
  reg [31:0] _RAND_1859;
  reg [31:0] _RAND_1860;
  reg [31:0] _RAND_1861;
  reg [31:0] _RAND_1862;
  reg [31:0] _RAND_1863;
  reg [31:0] _RAND_1864;
  reg [31:0] _RAND_1865;
  reg [31:0] _RAND_1866;
  reg [31:0] _RAND_1867;
  reg [31:0] _RAND_1868;
  reg [31:0] _RAND_1869;
  reg [31:0] _RAND_1870;
  reg [31:0] _RAND_1871;
  reg [31:0] _RAND_1872;
  reg [31:0] _RAND_1873;
  reg [31:0] _RAND_1874;
  reg [31:0] _RAND_1875;
  reg [31:0] _RAND_1876;
  reg [31:0] _RAND_1877;
  reg [31:0] _RAND_1878;
  reg [31:0] _RAND_1879;
  reg [31:0] _RAND_1880;
  reg [31:0] _RAND_1881;
  reg [31:0] _RAND_1882;
  reg [31:0] _RAND_1883;
  reg [31:0] _RAND_1884;
  reg [31:0] _RAND_1885;
  reg [31:0] _RAND_1886;
  reg [31:0] _RAND_1887;
  reg [31:0] _RAND_1888;
  reg [31:0] _RAND_1889;
  reg [31:0] _RAND_1890;
  reg [31:0] _RAND_1891;
  reg [31:0] _RAND_1892;
  reg [31:0] _RAND_1893;
  reg [31:0] _RAND_1894;
  reg [31:0] _RAND_1895;
  reg [31:0] _RAND_1896;
  reg [31:0] _RAND_1897;
  reg [31:0] _RAND_1898;
  reg [31:0] _RAND_1899;
  reg [31:0] _RAND_1900;
  reg [31:0] _RAND_1901;
  reg [31:0] _RAND_1902;
  reg [31:0] _RAND_1903;
  reg [31:0] _RAND_1904;
  reg [31:0] _RAND_1905;
  reg [31:0] _RAND_1906;
  reg [31:0] _RAND_1907;
  reg [31:0] _RAND_1908;
  reg [31:0] _RAND_1909;
  reg [31:0] _RAND_1910;
  reg [31:0] _RAND_1911;
  reg [31:0] _RAND_1912;
  reg [31:0] _RAND_1913;
  reg [31:0] _RAND_1914;
  reg [31:0] _RAND_1915;
  reg [31:0] _RAND_1916;
  reg [31:0] _RAND_1917;
  reg [31:0] _RAND_1918;
  reg [31:0] _RAND_1919;
  reg [31:0] _RAND_1920;
  reg [31:0] _RAND_1921;
  reg [31:0] _RAND_1922;
  reg [31:0] _RAND_1923;
  reg [31:0] _RAND_1924;
  reg [31:0] _RAND_1925;
  reg [31:0] _RAND_1926;
  reg [31:0] _RAND_1927;
  reg [31:0] _RAND_1928;
  reg [31:0] _RAND_1929;
  reg [31:0] _RAND_1930;
  reg [31:0] _RAND_1931;
  reg [31:0] _RAND_1932;
  reg [31:0] _RAND_1933;
  reg [31:0] _RAND_1934;
  reg [31:0] _RAND_1935;
  reg [31:0] _RAND_1936;
  reg [31:0] _RAND_1937;
  reg [31:0] _RAND_1938;
  reg [31:0] _RAND_1939;
  reg [31:0] _RAND_1940;
  reg [31:0] _RAND_1941;
  reg [31:0] _RAND_1942;
  reg [31:0] _RAND_1943;
  reg [31:0] _RAND_1944;
  reg [31:0] _RAND_1945;
  reg [31:0] _RAND_1946;
  reg [31:0] _RAND_1947;
  reg [31:0] _RAND_1948;
  reg [31:0] _RAND_1949;
  reg [31:0] _RAND_1950;
  reg [31:0] _RAND_1951;
  reg [31:0] _RAND_1952;
  reg [31:0] _RAND_1953;
  reg [31:0] _RAND_1954;
  reg [31:0] _RAND_1955;
  reg [31:0] _RAND_1956;
  reg [31:0] _RAND_1957;
  reg [31:0] _RAND_1958;
  reg [31:0] _RAND_1959;
  reg [31:0] _RAND_1960;
  reg [31:0] _RAND_1961;
  reg [31:0] _RAND_1962;
  reg [31:0] _RAND_1963;
  reg [31:0] _RAND_1964;
  reg [31:0] _RAND_1965;
  reg [31:0] _RAND_1966;
  reg [31:0] _RAND_1967;
  reg [31:0] _RAND_1968;
  reg [31:0] _RAND_1969;
  reg [31:0] _RAND_1970;
  reg [31:0] _RAND_1971;
  reg [31:0] _RAND_1972;
  reg [31:0] _RAND_1973;
  reg [31:0] _RAND_1974;
  reg [31:0] _RAND_1975;
  reg [31:0] _RAND_1976;
  reg [31:0] _RAND_1977;
  reg [31:0] _RAND_1978;
  reg [31:0] _RAND_1979;
  reg [31:0] _RAND_1980;
  reg [31:0] _RAND_1981;
  reg [31:0] _RAND_1982;
  reg [31:0] _RAND_1983;
  reg [31:0] _RAND_1984;
  reg [31:0] _RAND_1985;
  reg [31:0] _RAND_1986;
  reg [31:0] _RAND_1987;
  reg [31:0] _RAND_1988;
  reg [31:0] _RAND_1989;
  reg [31:0] _RAND_1990;
  reg [31:0] _RAND_1991;
  reg [31:0] _RAND_1992;
  reg [31:0] _RAND_1993;
  reg [31:0] _RAND_1994;
  reg [31:0] _RAND_1995;
  reg [31:0] _RAND_1996;
  reg [31:0] _RAND_1997;
  reg [31:0] _RAND_1998;
  reg [31:0] _RAND_1999;
  reg [31:0] _RAND_2000;
  reg [31:0] _RAND_2001;
  reg [31:0] _RAND_2002;
  reg [31:0] _RAND_2003;
  reg [31:0] _RAND_2004;
  reg [31:0] _RAND_2005;
  reg [31:0] _RAND_2006;
  reg [31:0] _RAND_2007;
  reg [31:0] _RAND_2008;
  reg [31:0] _RAND_2009;
  reg [31:0] _RAND_2010;
  reg [31:0] _RAND_2011;
  reg [31:0] _RAND_2012;
  reg [31:0] _RAND_2013;
  reg [31:0] _RAND_2014;
  reg [31:0] _RAND_2015;
  reg [31:0] _RAND_2016;
  reg [31:0] _RAND_2017;
  reg [31:0] _RAND_2018;
  reg [31:0] _RAND_2019;
  reg [31:0] _RAND_2020;
  reg [31:0] _RAND_2021;
  reg [31:0] _RAND_2022;
  reg [31:0] _RAND_2023;
  reg [31:0] _RAND_2024;
  reg [31:0] _RAND_2025;
  reg [31:0] _RAND_2026;
  reg [31:0] _RAND_2027;
  reg [31:0] _RAND_2028;
  reg [31:0] _RAND_2029;
  reg [31:0] _RAND_2030;
  reg [31:0] _RAND_2031;
  reg [31:0] _RAND_2032;
  reg [31:0] _RAND_2033;
  reg [31:0] _RAND_2034;
  reg [31:0] _RAND_2035;
  reg [31:0] _RAND_2036;
  reg [31:0] _RAND_2037;
  reg [31:0] _RAND_2038;
  reg [31:0] _RAND_2039;
  reg [31:0] _RAND_2040;
  reg [31:0] _RAND_2041;
  reg [31:0] _RAND_2042;
  reg [31:0] _RAND_2043;
  reg [31:0] _RAND_2044;
  reg [31:0] _RAND_2045;
  reg [31:0] _RAND_2046;
  reg [31:0] _RAND_2047;
  reg [31:0] _RAND_2048;
  reg [31:0] _RAND_2049;
  reg [31:0] _RAND_2050;
  reg [31:0] _RAND_2051;
  reg [31:0] _RAND_2052;
  reg [31:0] _RAND_2053;
  reg [31:0] _RAND_2054;
  reg [31:0] _RAND_2055;
  reg [31:0] _RAND_2056;
  reg [31:0] _RAND_2057;
  reg [31:0] _RAND_2058;
  reg [31:0] _RAND_2059;
  reg [31:0] _RAND_2060;
  reg [31:0] _RAND_2061;
  reg [31:0] _RAND_2062;
  reg [31:0] _RAND_2063;
  reg [31:0] _RAND_2064;
  reg [31:0] _RAND_2065;
  reg [31:0] _RAND_2066;
  reg [31:0] _RAND_2067;
  reg [31:0] _RAND_2068;
  reg [31:0] _RAND_2069;
  reg [31:0] _RAND_2070;
  reg [31:0] _RAND_2071;
  reg [31:0] _RAND_2072;
  reg [31:0] _RAND_2073;
  reg [31:0] _RAND_2074;
  reg [31:0] _RAND_2075;
  reg [31:0] _RAND_2076;
  reg [31:0] _RAND_2077;
  reg [31:0] _RAND_2078;
  reg [31:0] _RAND_2079;
  reg [31:0] _RAND_2080;
  reg [31:0] _RAND_2081;
  reg [31:0] _RAND_2082;
  reg [31:0] _RAND_2083;
  reg [31:0] _RAND_2084;
  reg [31:0] _RAND_2085;
  reg [31:0] _RAND_2086;
  reg [31:0] _RAND_2087;
  reg [31:0] _RAND_2088;
  reg [31:0] _RAND_2089;
  reg [31:0] _RAND_2090;
  reg [31:0] _RAND_2091;
  reg [31:0] _RAND_2092;
  reg [31:0] _RAND_2093;
  reg [31:0] _RAND_2094;
  reg [31:0] _RAND_2095;
  reg [31:0] _RAND_2096;
  reg [31:0] _RAND_2097;
  reg [31:0] _RAND_2098;
  reg [31:0] _RAND_2099;
  reg [31:0] _RAND_2100;
  reg [31:0] _RAND_2101;
  reg [31:0] _RAND_2102;
  reg [31:0] _RAND_2103;
  reg [31:0] _RAND_2104;
  reg [31:0] _RAND_2105;
  reg [31:0] _RAND_2106;
  reg [31:0] _RAND_2107;
  reg [31:0] _RAND_2108;
  reg [31:0] _RAND_2109;
  reg [31:0] _RAND_2110;
  reg [31:0] _RAND_2111;
  reg [31:0] _RAND_2112;
  reg [31:0] _RAND_2113;
  reg [31:0] _RAND_2114;
  reg [31:0] _RAND_2115;
  reg [31:0] _RAND_2116;
  reg [31:0] _RAND_2117;
  reg [31:0] _RAND_2118;
  reg [31:0] _RAND_2119;
  reg [31:0] _RAND_2120;
  reg [31:0] _RAND_2121;
  reg [31:0] _RAND_2122;
  reg [31:0] _RAND_2123;
  reg [31:0] _RAND_2124;
  reg [31:0] _RAND_2125;
  reg [31:0] _RAND_2126;
  reg [31:0] _RAND_2127;
  reg [31:0] _RAND_2128;
  reg [31:0] _RAND_2129;
  reg [31:0] _RAND_2130;
  reg [31:0] _RAND_2131;
  reg [31:0] _RAND_2132;
  reg [31:0] _RAND_2133;
  reg [31:0] _RAND_2134;
  reg [31:0] _RAND_2135;
  reg [31:0] _RAND_2136;
  reg [31:0] _RAND_2137;
  reg [31:0] _RAND_2138;
  reg [31:0] _RAND_2139;
  reg [31:0] _RAND_2140;
  reg [31:0] _RAND_2141;
  reg [31:0] _RAND_2142;
  reg [31:0] _RAND_2143;
  reg [31:0] _RAND_2144;
  reg [31:0] _RAND_2145;
  reg [31:0] _RAND_2146;
  reg [31:0] _RAND_2147;
  reg [31:0] _RAND_2148;
  reg [31:0] _RAND_2149;
  reg [31:0] _RAND_2150;
  reg [31:0] _RAND_2151;
  reg [31:0] _RAND_2152;
  reg [31:0] _RAND_2153;
  reg [31:0] _RAND_2154;
  reg [31:0] _RAND_2155;
  reg [31:0] _RAND_2156;
  reg [31:0] _RAND_2157;
  reg [31:0] _RAND_2158;
  reg [31:0] _RAND_2159;
  reg [31:0] _RAND_2160;
  reg [31:0] _RAND_2161;
  reg [31:0] _RAND_2162;
  reg [31:0] _RAND_2163;
  reg [31:0] _RAND_2164;
  reg [31:0] _RAND_2165;
  reg [31:0] _RAND_2166;
  reg [31:0] _RAND_2167;
  reg [31:0] _RAND_2168;
  reg [31:0] _RAND_2169;
  reg [31:0] _RAND_2170;
  reg [31:0] _RAND_2171;
  reg [31:0] _RAND_2172;
  reg [31:0] _RAND_2173;
  reg [31:0] _RAND_2174;
  reg [31:0] _RAND_2175;
  reg [31:0] _RAND_2176;
  reg [31:0] _RAND_2177;
  reg [31:0] _RAND_2178;
  reg [31:0] _RAND_2179;
  reg [31:0] _RAND_2180;
  reg [31:0] _RAND_2181;
  reg [31:0] _RAND_2182;
  reg [31:0] _RAND_2183;
  reg [31:0] _RAND_2184;
  reg [31:0] _RAND_2185;
  reg [31:0] _RAND_2186;
  reg [31:0] _RAND_2187;
  reg [31:0] _RAND_2188;
  reg [31:0] _RAND_2189;
  reg [31:0] _RAND_2190;
  reg [31:0] _RAND_2191;
  reg [31:0] _RAND_2192;
  reg [31:0] _RAND_2193;
  reg [31:0] _RAND_2194;
  reg [31:0] _RAND_2195;
  reg [31:0] _RAND_2196;
  reg [31:0] _RAND_2197;
  reg [31:0] _RAND_2198;
  reg [31:0] _RAND_2199;
  reg [31:0] _RAND_2200;
  reg [31:0] _RAND_2201;
  reg [31:0] _RAND_2202;
  reg [31:0] _RAND_2203;
  reg [31:0] _RAND_2204;
  reg [31:0] _RAND_2205;
  reg [31:0] _RAND_2206;
  reg [31:0] _RAND_2207;
  reg [31:0] _RAND_2208;
  reg [31:0] _RAND_2209;
  reg [31:0] _RAND_2210;
  reg [31:0] _RAND_2211;
  reg [31:0] _RAND_2212;
  reg [31:0] _RAND_2213;
  reg [31:0] _RAND_2214;
  reg [31:0] _RAND_2215;
  reg [31:0] _RAND_2216;
  reg [31:0] _RAND_2217;
  reg [31:0] _RAND_2218;
  reg [31:0] _RAND_2219;
  reg [31:0] _RAND_2220;
  reg [31:0] _RAND_2221;
  reg [31:0] _RAND_2222;
  reg [31:0] _RAND_2223;
  reg [31:0] _RAND_2224;
  reg [31:0] _RAND_2225;
  reg [31:0] _RAND_2226;
  reg [31:0] _RAND_2227;
  reg [31:0] _RAND_2228;
  reg [31:0] _RAND_2229;
  reg [31:0] _RAND_2230;
  reg [31:0] _RAND_2231;
  reg [31:0] _RAND_2232;
  reg [31:0] _RAND_2233;
  reg [31:0] _RAND_2234;
  reg [31:0] _RAND_2235;
  reg [31:0] _RAND_2236;
  reg [31:0] _RAND_2237;
  reg [31:0] _RAND_2238;
  reg [31:0] _RAND_2239;
  reg [31:0] _RAND_2240;
  reg [31:0] _RAND_2241;
  reg [31:0] _RAND_2242;
  reg [31:0] _RAND_2243;
  reg [31:0] _RAND_2244;
  reg [31:0] _RAND_2245;
  reg [31:0] _RAND_2246;
  reg [31:0] _RAND_2247;
  reg [31:0] _RAND_2248;
  reg [31:0] _RAND_2249;
  reg [31:0] _RAND_2250;
  reg [31:0] _RAND_2251;
  reg [31:0] _RAND_2252;
  reg [31:0] _RAND_2253;
  reg [31:0] _RAND_2254;
  reg [31:0] _RAND_2255;
  reg [31:0] _RAND_2256;
  reg [31:0] _RAND_2257;
  reg [31:0] _RAND_2258;
  reg [31:0] _RAND_2259;
  reg [31:0] _RAND_2260;
  reg [31:0] _RAND_2261;
  reg [31:0] _RAND_2262;
  reg [31:0] _RAND_2263;
  reg [31:0] _RAND_2264;
  reg [31:0] _RAND_2265;
  reg [31:0] _RAND_2266;
  reg [31:0] _RAND_2267;
  reg [31:0] _RAND_2268;
  reg [31:0] _RAND_2269;
  reg [31:0] _RAND_2270;
  reg [31:0] _RAND_2271;
  reg [31:0] _RAND_2272;
  reg [31:0] _RAND_2273;
  reg [31:0] _RAND_2274;
  reg [31:0] _RAND_2275;
  reg [31:0] _RAND_2276;
  reg [31:0] _RAND_2277;
  reg [31:0] _RAND_2278;
  reg [31:0] _RAND_2279;
  reg [31:0] _RAND_2280;
  reg [31:0] _RAND_2281;
  reg [31:0] _RAND_2282;
  reg [31:0] _RAND_2283;
  reg [31:0] _RAND_2284;
  reg [31:0] _RAND_2285;
  reg [31:0] _RAND_2286;
  reg [31:0] _RAND_2287;
  reg [31:0] _RAND_2288;
  reg [31:0] _RAND_2289;
  reg [31:0] _RAND_2290;
  reg [31:0] _RAND_2291;
  reg [31:0] _RAND_2292;
  reg [31:0] _RAND_2293;
  reg [31:0] _RAND_2294;
  reg [31:0] _RAND_2295;
  reg [31:0] _RAND_2296;
  reg [31:0] _RAND_2297;
  reg [31:0] _RAND_2298;
  reg [31:0] _RAND_2299;
  reg [31:0] _RAND_2300;
  reg [31:0] _RAND_2301;
  reg [31:0] _RAND_2302;
  reg [31:0] _RAND_2303;
  reg [31:0] _RAND_2304;
  reg [31:0] _RAND_2305;
  reg [31:0] _RAND_2306;
  reg [31:0] _RAND_2307;
  reg [31:0] _RAND_2308;
  reg [31:0] _RAND_2309;
  reg [31:0] _RAND_2310;
  reg [31:0] _RAND_2311;
  reg [31:0] _RAND_2312;
  reg [31:0] _RAND_2313;
  reg [31:0] _RAND_2314;
  reg [31:0] _RAND_2315;
  reg [31:0] _RAND_2316;
  reg [31:0] _RAND_2317;
  reg [31:0] _RAND_2318;
  reg [31:0] _RAND_2319;
  reg [31:0] _RAND_2320;
  reg [31:0] _RAND_2321;
  reg [31:0] _RAND_2322;
  reg [31:0] _RAND_2323;
  reg [31:0] _RAND_2324;
  reg [31:0] _RAND_2325;
  reg [31:0] _RAND_2326;
  reg [31:0] _RAND_2327;
  reg [31:0] _RAND_2328;
  reg [31:0] _RAND_2329;
  reg [31:0] _RAND_2330;
  reg [31:0] _RAND_2331;
  reg [31:0] _RAND_2332;
  reg [31:0] _RAND_2333;
  reg [31:0] _RAND_2334;
  reg [31:0] _RAND_2335;
  reg [31:0] _RAND_2336;
  reg [31:0] _RAND_2337;
  reg [31:0] _RAND_2338;
  reg [31:0] _RAND_2339;
  reg [31:0] _RAND_2340;
  reg [31:0] _RAND_2341;
  reg [31:0] _RAND_2342;
  reg [31:0] _RAND_2343;
  reg [31:0] _RAND_2344;
  reg [31:0] _RAND_2345;
  reg [31:0] _RAND_2346;
  reg [31:0] _RAND_2347;
  reg [31:0] _RAND_2348;
  reg [31:0] _RAND_2349;
  reg [31:0] _RAND_2350;
  reg [31:0] _RAND_2351;
  reg [31:0] _RAND_2352;
  reg [31:0] _RAND_2353;
  reg [31:0] _RAND_2354;
  reg [31:0] _RAND_2355;
  reg [31:0] _RAND_2356;
  reg [31:0] _RAND_2357;
  reg [31:0] _RAND_2358;
  reg [31:0] _RAND_2359;
  reg [31:0] _RAND_2360;
  reg [31:0] _RAND_2361;
  reg [31:0] _RAND_2362;
  reg [31:0] _RAND_2363;
  reg [31:0] _RAND_2364;
  reg [31:0] _RAND_2365;
  reg [31:0] _RAND_2366;
  reg [31:0] _RAND_2367;
  reg [31:0] _RAND_2368;
  reg [31:0] _RAND_2369;
  reg [31:0] _RAND_2370;
  reg [31:0] _RAND_2371;
  reg [31:0] _RAND_2372;
  reg [31:0] _RAND_2373;
  reg [31:0] _RAND_2374;
  reg [31:0] _RAND_2375;
  reg [31:0] _RAND_2376;
  reg [31:0] _RAND_2377;
  reg [31:0] _RAND_2378;
  reg [31:0] _RAND_2379;
  reg [31:0] _RAND_2380;
  reg [31:0] _RAND_2381;
  reg [31:0] _RAND_2382;
  reg [31:0] _RAND_2383;
  reg [31:0] _RAND_2384;
  reg [31:0] _RAND_2385;
  reg [31:0] _RAND_2386;
  reg [31:0] _RAND_2387;
  reg [31:0] _RAND_2388;
  reg [31:0] _RAND_2389;
  reg [31:0] _RAND_2390;
  reg [31:0] _RAND_2391;
  reg [31:0] _RAND_2392;
  reg [31:0] _RAND_2393;
  reg [31:0] _RAND_2394;
  reg [31:0] _RAND_2395;
  reg [31:0] _RAND_2396;
  reg [31:0] _RAND_2397;
  reg [31:0] _RAND_2398;
  reg [31:0] _RAND_2399;
  reg [31:0] _RAND_2400;
  reg [31:0] _RAND_2401;
  reg [31:0] _RAND_2402;
  reg [31:0] _RAND_2403;
  reg [31:0] _RAND_2404;
  reg [31:0] _RAND_2405;
  reg [31:0] _RAND_2406;
  reg [31:0] _RAND_2407;
  reg [31:0] _RAND_2408;
  reg [31:0] _RAND_2409;
  reg [31:0] _RAND_2410;
  reg [31:0] _RAND_2411;
  reg [31:0] _RAND_2412;
  reg [31:0] _RAND_2413;
  reg [31:0] _RAND_2414;
  reg [31:0] _RAND_2415;
  reg [31:0] _RAND_2416;
  reg [31:0] _RAND_2417;
  reg [31:0] _RAND_2418;
  reg [31:0] _RAND_2419;
  reg [31:0] _RAND_2420;
  reg [31:0] _RAND_2421;
  reg [31:0] _RAND_2422;
  reg [31:0] _RAND_2423;
  reg [31:0] _RAND_2424;
  reg [31:0] _RAND_2425;
  reg [31:0] _RAND_2426;
  reg [31:0] _RAND_2427;
  reg [31:0] _RAND_2428;
  reg [31:0] _RAND_2429;
  reg [31:0] _RAND_2430;
  reg [31:0] _RAND_2431;
  reg [31:0] _RAND_2432;
  reg [31:0] _RAND_2433;
  reg [31:0] _RAND_2434;
  reg [31:0] _RAND_2435;
  reg [31:0] _RAND_2436;
  reg [31:0] _RAND_2437;
  reg [31:0] _RAND_2438;
  reg [31:0] _RAND_2439;
  reg [31:0] _RAND_2440;
  reg [31:0] _RAND_2441;
  reg [31:0] _RAND_2442;
  reg [31:0] _RAND_2443;
  reg [31:0] _RAND_2444;
  reg [31:0] _RAND_2445;
  reg [31:0] _RAND_2446;
  reg [31:0] _RAND_2447;
  reg [31:0] _RAND_2448;
  reg [31:0] _RAND_2449;
  reg [31:0] _RAND_2450;
  reg [31:0] _RAND_2451;
  reg [31:0] _RAND_2452;
  reg [31:0] _RAND_2453;
  reg [31:0] _RAND_2454;
  reg [31:0] _RAND_2455;
  reg [31:0] _RAND_2456;
  reg [31:0] _RAND_2457;
  reg [31:0] _RAND_2458;
  reg [31:0] _RAND_2459;
  reg [31:0] _RAND_2460;
  reg [31:0] _RAND_2461;
  reg [31:0] _RAND_2462;
  reg [31:0] _RAND_2463;
  reg [31:0] _RAND_2464;
  reg [31:0] _RAND_2465;
  reg [31:0] _RAND_2466;
  reg [31:0] _RAND_2467;
  reg [31:0] _RAND_2468;
  reg [31:0] _RAND_2469;
  reg [31:0] _RAND_2470;
  reg [31:0] _RAND_2471;
  reg [31:0] _RAND_2472;
  reg [31:0] _RAND_2473;
  reg [31:0] _RAND_2474;
  reg [31:0] _RAND_2475;
  reg [31:0] _RAND_2476;
  reg [31:0] _RAND_2477;
  reg [31:0] _RAND_2478;
  reg [31:0] _RAND_2479;
  reg [31:0] _RAND_2480;
  reg [31:0] _RAND_2481;
  reg [31:0] _RAND_2482;
  reg [31:0] _RAND_2483;
  reg [31:0] _RAND_2484;
  reg [31:0] _RAND_2485;
  reg [31:0] _RAND_2486;
  reg [31:0] _RAND_2487;
  reg [31:0] _RAND_2488;
  reg [31:0] _RAND_2489;
  reg [31:0] _RAND_2490;
  reg [31:0] _RAND_2491;
  reg [31:0] _RAND_2492;
  reg [31:0] _RAND_2493;
  reg [31:0] _RAND_2494;
  reg [31:0] _RAND_2495;
  reg [31:0] _RAND_2496;
  reg [31:0] _RAND_2497;
  reg [31:0] _RAND_2498;
  reg [31:0] _RAND_2499;
  reg [31:0] _RAND_2500;
  reg [31:0] _RAND_2501;
  reg [31:0] _RAND_2502;
  reg [31:0] _RAND_2503;
  reg [31:0] _RAND_2504;
  reg [31:0] _RAND_2505;
  reg [31:0] _RAND_2506;
  reg [31:0] _RAND_2507;
  reg [31:0] _RAND_2508;
  reg [31:0] _RAND_2509;
  reg [31:0] _RAND_2510;
  reg [31:0] _RAND_2511;
  reg [31:0] _RAND_2512;
  reg [31:0] _RAND_2513;
  reg [31:0] _RAND_2514;
  reg [31:0] _RAND_2515;
  reg [31:0] _RAND_2516;
  reg [31:0] _RAND_2517;
  reg [31:0] _RAND_2518;
  reg [31:0] _RAND_2519;
  reg [31:0] _RAND_2520;
  reg [31:0] _RAND_2521;
  reg [31:0] _RAND_2522;
  reg [31:0] _RAND_2523;
  reg [31:0] _RAND_2524;
  reg [31:0] _RAND_2525;
  reg [31:0] _RAND_2526;
  reg [31:0] _RAND_2527;
  reg [31:0] _RAND_2528;
  reg [31:0] _RAND_2529;
  reg [31:0] _RAND_2530;
  reg [31:0] _RAND_2531;
  reg [31:0] _RAND_2532;
  reg [31:0] _RAND_2533;
  reg [31:0] _RAND_2534;
  reg [31:0] _RAND_2535;
  reg [31:0] _RAND_2536;
  reg [31:0] _RAND_2537;
  reg [31:0] _RAND_2538;
  reg [31:0] _RAND_2539;
  reg [31:0] _RAND_2540;
  reg [31:0] _RAND_2541;
  reg [31:0] _RAND_2542;
  reg [31:0] _RAND_2543;
  reg [31:0] _RAND_2544;
  reg [31:0] _RAND_2545;
  reg [31:0] _RAND_2546;
  reg [31:0] _RAND_2547;
  reg [31:0] _RAND_2548;
  reg [31:0] _RAND_2549;
  reg [31:0] _RAND_2550;
`endif // RANDOMIZE_REG_INIT
  wire  KernelConvolution_clock; // @[Filter.scala 122:35]
  wire  KernelConvolution_reset; // @[Filter.scala 122:35]
  wire [4:0] KernelConvolution_io_kernelVal_in; // @[Filter.scala 122:35]
  wire [3:0] KernelConvolution_io_pixelVal_in_0; // @[Filter.scala 122:35]
  wire [3:0] KernelConvolution_io_pixelVal_in_1; // @[Filter.scala 122:35]
  wire [3:0] KernelConvolution_io_pixelVal_in_2; // @[Filter.scala 122:35]
  wire [3:0] KernelConvolution_io_pixelVal_in_3; // @[Filter.scala 122:35]
  wire [3:0] KernelConvolution_io_pixelVal_in_4; // @[Filter.scala 122:35]
  wire [3:0] KernelConvolution_io_pixelVal_in_5; // @[Filter.scala 122:35]
  wire [3:0] KernelConvolution_io_pixelVal_in_6; // @[Filter.scala 122:35]
  wire [3:0] KernelConvolution_io_pixelVal_in_7; // @[Filter.scala 122:35]
  wire [8:0] KernelConvolution_io_pixelVal_out_0; // @[Filter.scala 122:35]
  wire [8:0] KernelConvolution_io_pixelVal_out_1; // @[Filter.scala 122:35]
  wire [8:0] KernelConvolution_io_pixelVal_out_2; // @[Filter.scala 122:35]
  wire [8:0] KernelConvolution_io_pixelVal_out_3; // @[Filter.scala 122:35]
  wire [8:0] KernelConvolution_io_pixelVal_out_4; // @[Filter.scala 122:35]
  wire [8:0] KernelConvolution_io_pixelVal_out_5; // @[Filter.scala 122:35]
  wire [8:0] KernelConvolution_io_pixelVal_out_6; // @[Filter.scala 122:35]
  wire [8:0] KernelConvolution_io_pixelVal_out_7; // @[Filter.scala 122:35]
  wire  KernelConvolution_io_valid_out; // @[Filter.scala 122:35]
  reg [3:0] image_12; // @[Filter.scala 68:24]
  reg [3:0] image_14; // @[Filter.scala 68:24]
  reg [3:0] image_15; // @[Filter.scala 68:24]
  reg [3:0] image_16; // @[Filter.scala 68:24]
  reg [3:0] image_17; // @[Filter.scala 68:24]
  reg [3:0] image_18; // @[Filter.scala 68:24]
  reg [3:0] image_19; // @[Filter.scala 68:24]
  reg [3:0] image_20; // @[Filter.scala 68:24]
  reg [3:0] image_21; // @[Filter.scala 68:24]
  reg [3:0] image_22; // @[Filter.scala 68:24]
  reg [3:0] image_23; // @[Filter.scala 68:24]
  reg [3:0] image_35; // @[Filter.scala 68:24]
  reg [3:0] image_36; // @[Filter.scala 68:24]
  reg [3:0] image_37; // @[Filter.scala 68:24]
  reg [3:0] image_38; // @[Filter.scala 68:24]
  reg [3:0] image_39; // @[Filter.scala 68:24]
  reg [3:0] image_40; // @[Filter.scala 68:24]
  reg [3:0] image_41; // @[Filter.scala 68:24]
  reg [3:0] image_42; // @[Filter.scala 68:24]
  reg [3:0] image_75; // @[Filter.scala 68:24]
  reg [3:0] image_76; // @[Filter.scala 68:24]
  reg [3:0] image_77; // @[Filter.scala 68:24]
  reg [3:0] image_78; // @[Filter.scala 68:24]
  reg [3:0] image_79; // @[Filter.scala 68:24]
  reg [3:0] image_80; // @[Filter.scala 68:24]
  reg [3:0] image_81; // @[Filter.scala 68:24]
  reg [3:0] image_82; // @[Filter.scala 68:24]
  reg [3:0] image_83; // @[Filter.scala 68:24]
  reg [3:0] image_84; // @[Filter.scala 68:24]
  reg [3:0] image_85; // @[Filter.scala 68:24]
  reg [3:0] image_86; // @[Filter.scala 68:24]
  reg [3:0] image_87; // @[Filter.scala 68:24]
  reg [3:0] image_88; // @[Filter.scala 68:24]
  reg [3:0] image_89; // @[Filter.scala 68:24]
  reg [3:0] image_90; // @[Filter.scala 68:24]
  reg [3:0] image_93; // @[Filter.scala 68:24]
  reg [3:0] image_95; // @[Filter.scala 68:24]
  reg [3:0] image_96; // @[Filter.scala 68:24]
  reg [3:0] image_97; // @[Filter.scala 68:24]
  reg [3:0] image_98; // @[Filter.scala 68:24]
  reg [3:0] image_99; // @[Filter.scala 68:24]
  reg [3:0] image_100; // @[Filter.scala 68:24]
  reg [3:0] image_101; // @[Filter.scala 68:24]
  reg [3:0] image_102; // @[Filter.scala 68:24]
  reg [3:0] image_103; // @[Filter.scala 68:24]
  reg [3:0] image_104; // @[Filter.scala 68:24]
  reg [3:0] image_105; // @[Filter.scala 68:24]
  reg [3:0] image_106; // @[Filter.scala 68:24]
  reg [3:0] image_107; // @[Filter.scala 68:24]
  reg [3:0] image_108; // @[Filter.scala 68:24]
  reg [3:0] image_136; // @[Filter.scala 68:24]
  reg [3:0] image_137; // @[Filter.scala 68:24]
  reg [3:0] image_138; // @[Filter.scala 68:24]
  reg [3:0] image_139; // @[Filter.scala 68:24]
  reg [3:0] image_140; // @[Filter.scala 68:24]
  reg [3:0] image_141; // @[Filter.scala 68:24]
  reg [3:0] image_142; // @[Filter.scala 68:24]
  reg [3:0] image_143; // @[Filter.scala 68:24]
  reg [3:0] image_144; // @[Filter.scala 68:24]
  reg [3:0] image_145; // @[Filter.scala 68:24]
  reg [3:0] image_146; // @[Filter.scala 68:24]
  reg [3:0] image_147; // @[Filter.scala 68:24]
  reg [3:0] image_148; // @[Filter.scala 68:24]
  reg [3:0] image_149; // @[Filter.scala 68:24]
  reg [3:0] image_150; // @[Filter.scala 68:24]
  reg [3:0] image_151; // @[Filter.scala 68:24]
  reg [3:0] image_152; // @[Filter.scala 68:24]
  reg [3:0] image_153; // @[Filter.scala 68:24]
  reg [3:0] image_154; // @[Filter.scala 68:24]
  reg [3:0] image_155; // @[Filter.scala 68:24]
  reg [3:0] image_157; // @[Filter.scala 68:24]
  reg [3:0] image_158; // @[Filter.scala 68:24]
  reg [3:0] image_159; // @[Filter.scala 68:24]
  reg [3:0] image_160; // @[Filter.scala 68:24]
  reg [3:0] image_161; // @[Filter.scala 68:24]
  reg [3:0] image_162; // @[Filter.scala 68:24]
  reg [3:0] image_163; // @[Filter.scala 68:24]
  reg [3:0] image_164; // @[Filter.scala 68:24]
  reg [3:0] image_165; // @[Filter.scala 68:24]
  reg [3:0] image_166; // @[Filter.scala 68:24]
  reg [3:0] image_167; // @[Filter.scala 68:24]
  reg [3:0] image_168; // @[Filter.scala 68:24]
  reg [3:0] image_169; // @[Filter.scala 68:24]
  reg [3:0] image_170; // @[Filter.scala 68:24]
  reg [3:0] image_171; // @[Filter.scala 68:24]
  reg [3:0] image_172; // @[Filter.scala 68:24]
  reg [3:0] image_173; // @[Filter.scala 68:24]
  reg [3:0] image_174; // @[Filter.scala 68:24]
  reg [3:0] image_175; // @[Filter.scala 68:24]
  reg [3:0] image_176; // @[Filter.scala 68:24]
  reg [3:0] image_177; // @[Filter.scala 68:24]
  reg [3:0] image_178; // @[Filter.scala 68:24]
  reg [3:0] image_179; // @[Filter.scala 68:24]
  reg [3:0] image_199; // @[Filter.scala 68:24]
  reg [3:0] image_200; // @[Filter.scala 68:24]
  reg [3:0] image_201; // @[Filter.scala 68:24]
  reg [3:0] image_202; // @[Filter.scala 68:24]
  reg [3:0] image_203; // @[Filter.scala 68:24]
  reg [3:0] image_204; // @[Filter.scala 68:24]
  reg [3:0] image_205; // @[Filter.scala 68:24]
  reg [3:0] image_206; // @[Filter.scala 68:24]
  reg [3:0] image_207; // @[Filter.scala 68:24]
  reg [3:0] image_208; // @[Filter.scala 68:24]
  reg [3:0] image_209; // @[Filter.scala 68:24]
  reg [3:0] image_210; // @[Filter.scala 68:24]
  reg [3:0] image_211; // @[Filter.scala 68:24]
  reg [3:0] image_212; // @[Filter.scala 68:24]
  reg [3:0] image_213; // @[Filter.scala 68:24]
  reg [3:0] image_214; // @[Filter.scala 68:24]
  reg [3:0] image_215; // @[Filter.scala 68:24]
  reg [3:0] image_216; // @[Filter.scala 68:24]
  reg [3:0] image_217; // @[Filter.scala 68:24]
  reg [3:0] image_218; // @[Filter.scala 68:24]
  reg [3:0] image_219; // @[Filter.scala 68:24]
  reg [3:0] image_220; // @[Filter.scala 68:24]
  reg [3:0] image_221; // @[Filter.scala 68:24]
  reg [3:0] image_222; // @[Filter.scala 68:24]
  reg [3:0] image_223; // @[Filter.scala 68:24]
  reg [3:0] image_224; // @[Filter.scala 68:24]
  reg [3:0] image_225; // @[Filter.scala 68:24]
  reg [3:0] image_226; // @[Filter.scala 68:24]
  reg [3:0] image_227; // @[Filter.scala 68:24]
  reg [3:0] image_228; // @[Filter.scala 68:24]
  reg [3:0] image_229; // @[Filter.scala 68:24]
  reg [3:0] image_230; // @[Filter.scala 68:24]
  reg [3:0] image_231; // @[Filter.scala 68:24]
  reg [3:0] image_232; // @[Filter.scala 68:24]
  reg [3:0] image_233; // @[Filter.scala 68:24]
  reg [3:0] image_234; // @[Filter.scala 68:24]
  reg [3:0] image_235; // @[Filter.scala 68:24]
  reg [3:0] image_236; // @[Filter.scala 68:24]
  reg [3:0] image_237; // @[Filter.scala 68:24]
  reg [3:0] image_238; // @[Filter.scala 68:24]
  reg [3:0] image_239; // @[Filter.scala 68:24]
  reg [3:0] image_240; // @[Filter.scala 68:24]
  reg [3:0] image_241; // @[Filter.scala 68:24]
  reg [3:0] image_242; // @[Filter.scala 68:24]
  reg [3:0] image_243; // @[Filter.scala 68:24]
  reg [3:0] image_244; // @[Filter.scala 68:24]
  reg [3:0] image_245; // @[Filter.scala 68:24]
  reg [3:0] image_246; // @[Filter.scala 68:24]
  reg [3:0] image_262; // @[Filter.scala 68:24]
  reg [3:0] image_263; // @[Filter.scala 68:24]
  reg [3:0] image_264; // @[Filter.scala 68:24]
  reg [3:0] image_265; // @[Filter.scala 68:24]
  reg [3:0] image_266; // @[Filter.scala 68:24]
  reg [3:0] image_267; // @[Filter.scala 68:24]
  reg [3:0] image_268; // @[Filter.scala 68:24]
  reg [3:0] image_269; // @[Filter.scala 68:24]
  reg [3:0] image_270; // @[Filter.scala 68:24]
  reg [3:0] image_271; // @[Filter.scala 68:24]
  reg [3:0] image_272; // @[Filter.scala 68:24]
  reg [3:0] image_273; // @[Filter.scala 68:24]
  reg [3:0] image_274; // @[Filter.scala 68:24]
  reg [3:0] image_275; // @[Filter.scala 68:24]
  reg [3:0] image_276; // @[Filter.scala 68:24]
  reg [3:0] image_277; // @[Filter.scala 68:24]
  reg [3:0] image_278; // @[Filter.scala 68:24]
  reg [3:0] image_279; // @[Filter.scala 68:24]
  reg [3:0] image_280; // @[Filter.scala 68:24]
  reg [3:0] image_281; // @[Filter.scala 68:24]
  reg [3:0] image_282; // @[Filter.scala 68:24]
  reg [3:0] image_283; // @[Filter.scala 68:24]
  reg [3:0] image_284; // @[Filter.scala 68:24]
  reg [3:0] image_285; // @[Filter.scala 68:24]
  reg [3:0] image_286; // @[Filter.scala 68:24]
  reg [3:0] image_287; // @[Filter.scala 68:24]
  reg [3:0] image_288; // @[Filter.scala 68:24]
  reg [3:0] image_289; // @[Filter.scala 68:24]
  reg [3:0] image_290; // @[Filter.scala 68:24]
  reg [3:0] image_291; // @[Filter.scala 68:24]
  reg [3:0] image_292; // @[Filter.scala 68:24]
  reg [3:0] image_293; // @[Filter.scala 68:24]
  reg [3:0] image_294; // @[Filter.scala 68:24]
  reg [3:0] image_295; // @[Filter.scala 68:24]
  reg [3:0] image_296; // @[Filter.scala 68:24]
  reg [3:0] image_297; // @[Filter.scala 68:24]
  reg [3:0] image_298; // @[Filter.scala 68:24]
  reg [3:0] image_299; // @[Filter.scala 68:24]
  reg [3:0] image_300; // @[Filter.scala 68:24]
  reg [3:0] image_301; // @[Filter.scala 68:24]
  reg [3:0] image_302; // @[Filter.scala 68:24]
  reg [3:0] image_303; // @[Filter.scala 68:24]
  reg [3:0] image_304; // @[Filter.scala 68:24]
  reg [3:0] image_305; // @[Filter.scala 68:24]
  reg [3:0] image_306; // @[Filter.scala 68:24]
  reg [3:0] image_307; // @[Filter.scala 68:24]
  reg [3:0] image_308; // @[Filter.scala 68:24]
  reg [3:0] image_309; // @[Filter.scala 68:24]
  reg [3:0] image_310; // @[Filter.scala 68:24]
  reg [3:0] image_311; // @[Filter.scala 68:24]
  reg [3:0] image_312; // @[Filter.scala 68:24]
  reg [3:0] image_313; // @[Filter.scala 68:24]
  reg [3:0] image_314; // @[Filter.scala 68:24]
  reg [3:0] image_315; // @[Filter.scala 68:24]
  reg [3:0] image_325; // @[Filter.scala 68:24]
  reg [3:0] image_326; // @[Filter.scala 68:24]
  reg [3:0] image_327; // @[Filter.scala 68:24]
  reg [3:0] image_328; // @[Filter.scala 68:24]
  reg [3:0] image_329; // @[Filter.scala 68:24]
  reg [3:0] image_330; // @[Filter.scala 68:24]
  reg [3:0] image_331; // @[Filter.scala 68:24]
  reg [3:0] image_332; // @[Filter.scala 68:24]
  reg [3:0] image_333; // @[Filter.scala 68:24]
  reg [3:0] image_334; // @[Filter.scala 68:24]
  reg [3:0] image_335; // @[Filter.scala 68:24]
  reg [3:0] image_336; // @[Filter.scala 68:24]
  reg [3:0] image_337; // @[Filter.scala 68:24]
  reg [3:0] image_338; // @[Filter.scala 68:24]
  reg [3:0] image_339; // @[Filter.scala 68:24]
  reg [3:0] image_340; // @[Filter.scala 68:24]
  reg [3:0] image_341; // @[Filter.scala 68:24]
  reg [3:0] image_342; // @[Filter.scala 68:24]
  reg [3:0] image_343; // @[Filter.scala 68:24]
  reg [3:0] image_344; // @[Filter.scala 68:24]
  reg [3:0] image_345; // @[Filter.scala 68:24]
  reg [3:0] image_346; // @[Filter.scala 68:24]
  reg [3:0] image_347; // @[Filter.scala 68:24]
  reg [3:0] image_348; // @[Filter.scala 68:24]
  reg [3:0] image_349; // @[Filter.scala 68:24]
  reg [3:0] image_350; // @[Filter.scala 68:24]
  reg [3:0] image_351; // @[Filter.scala 68:24]
  reg [3:0] image_352; // @[Filter.scala 68:24]
  reg [3:0] image_353; // @[Filter.scala 68:24]
  reg [3:0] image_354; // @[Filter.scala 68:24]
  reg [3:0] image_355; // @[Filter.scala 68:24]
  reg [3:0] image_356; // @[Filter.scala 68:24]
  reg [3:0] image_357; // @[Filter.scala 68:24]
  reg [3:0] image_358; // @[Filter.scala 68:24]
  reg [3:0] image_359; // @[Filter.scala 68:24]
  reg [3:0] image_360; // @[Filter.scala 68:24]
  reg [3:0] image_361; // @[Filter.scala 68:24]
  reg [3:0] image_362; // @[Filter.scala 68:24]
  reg [3:0] image_363; // @[Filter.scala 68:24]
  reg [3:0] image_364; // @[Filter.scala 68:24]
  reg [3:0] image_365; // @[Filter.scala 68:24]
  reg [3:0] image_366; // @[Filter.scala 68:24]
  reg [3:0] image_367; // @[Filter.scala 68:24]
  reg [3:0] image_368; // @[Filter.scala 68:24]
  reg [3:0] image_369; // @[Filter.scala 68:24]
  reg [3:0] image_370; // @[Filter.scala 68:24]
  reg [3:0] image_371; // @[Filter.scala 68:24]
  reg [3:0] image_372; // @[Filter.scala 68:24]
  reg [3:0] image_373; // @[Filter.scala 68:24]
  reg [3:0] image_374; // @[Filter.scala 68:24]
  reg [3:0] image_375; // @[Filter.scala 68:24]
  reg [3:0] image_376; // @[Filter.scala 68:24]
  reg [3:0] image_377; // @[Filter.scala 68:24]
  reg [3:0] image_378; // @[Filter.scala 68:24]
  reg [3:0] image_379; // @[Filter.scala 68:24]
  reg [3:0] image_388; // @[Filter.scala 68:24]
  reg [3:0] image_389; // @[Filter.scala 68:24]
  reg [3:0] image_390; // @[Filter.scala 68:24]
  reg [3:0] image_391; // @[Filter.scala 68:24]
  reg [3:0] image_392; // @[Filter.scala 68:24]
  reg [3:0] image_393; // @[Filter.scala 68:24]
  reg [3:0] image_394; // @[Filter.scala 68:24]
  reg [3:0] image_395; // @[Filter.scala 68:24]
  reg [3:0] image_396; // @[Filter.scala 68:24]
  reg [3:0] image_397; // @[Filter.scala 68:24]
  reg [3:0] image_398; // @[Filter.scala 68:24]
  reg [3:0] image_399; // @[Filter.scala 68:24]
  reg [3:0] image_400; // @[Filter.scala 68:24]
  reg [3:0] image_401; // @[Filter.scala 68:24]
  reg [3:0] image_402; // @[Filter.scala 68:24]
  reg [3:0] image_403; // @[Filter.scala 68:24]
  reg [3:0] image_404; // @[Filter.scala 68:24]
  reg [3:0] image_405; // @[Filter.scala 68:24]
  reg [3:0] image_406; // @[Filter.scala 68:24]
  reg [3:0] image_407; // @[Filter.scala 68:24]
  reg [3:0] image_408; // @[Filter.scala 68:24]
  reg [3:0] image_409; // @[Filter.scala 68:24]
  reg [3:0] image_410; // @[Filter.scala 68:24]
  reg [3:0] image_411; // @[Filter.scala 68:24]
  reg [3:0] image_412; // @[Filter.scala 68:24]
  reg [3:0] image_413; // @[Filter.scala 68:24]
  reg [3:0] image_414; // @[Filter.scala 68:24]
  reg [3:0] image_415; // @[Filter.scala 68:24]
  reg [3:0] image_416; // @[Filter.scala 68:24]
  reg [3:0] image_417; // @[Filter.scala 68:24]
  reg [3:0] image_418; // @[Filter.scala 68:24]
  reg [3:0] image_419; // @[Filter.scala 68:24]
  reg [3:0] image_420; // @[Filter.scala 68:24]
  reg [3:0] image_421; // @[Filter.scala 68:24]
  reg [3:0] image_422; // @[Filter.scala 68:24]
  reg [3:0] image_423; // @[Filter.scala 68:24]
  reg [3:0] image_424; // @[Filter.scala 68:24]
  reg [3:0] image_425; // @[Filter.scala 68:24]
  reg [3:0] image_426; // @[Filter.scala 68:24]
  reg [3:0] image_427; // @[Filter.scala 68:24]
  reg [3:0] image_428; // @[Filter.scala 68:24]
  reg [3:0] image_429; // @[Filter.scala 68:24]
  reg [3:0] image_430; // @[Filter.scala 68:24]
  reg [3:0] image_431; // @[Filter.scala 68:24]
  reg [3:0] image_432; // @[Filter.scala 68:24]
  reg [3:0] image_433; // @[Filter.scala 68:24]
  reg [3:0] image_434; // @[Filter.scala 68:24]
  reg [3:0] image_435; // @[Filter.scala 68:24]
  reg [3:0] image_436; // @[Filter.scala 68:24]
  reg [3:0] image_437; // @[Filter.scala 68:24]
  reg [3:0] image_438; // @[Filter.scala 68:24]
  reg [3:0] image_439; // @[Filter.scala 68:24]
  reg [3:0] image_440; // @[Filter.scala 68:24]
  reg [3:0] image_441; // @[Filter.scala 68:24]
  reg [3:0] image_442; // @[Filter.scala 68:24]
  reg [3:0] image_443; // @[Filter.scala 68:24]
  reg [3:0] image_444; // @[Filter.scala 68:24]
  reg [3:0] image_451; // @[Filter.scala 68:24]
  reg [3:0] image_452; // @[Filter.scala 68:24]
  reg [3:0] image_453; // @[Filter.scala 68:24]
  reg [3:0] image_454; // @[Filter.scala 68:24]
  reg [3:0] image_455; // @[Filter.scala 68:24]
  reg [3:0] image_456; // @[Filter.scala 68:24]
  reg [3:0] image_457; // @[Filter.scala 68:24]
  reg [3:0] image_458; // @[Filter.scala 68:24]
  reg [3:0] image_459; // @[Filter.scala 68:24]
  reg [3:0] image_460; // @[Filter.scala 68:24]
  reg [3:0] image_461; // @[Filter.scala 68:24]
  reg [3:0] image_462; // @[Filter.scala 68:24]
  reg [3:0] image_463; // @[Filter.scala 68:24]
  reg [3:0] image_464; // @[Filter.scala 68:24]
  reg [3:0] image_465; // @[Filter.scala 68:24]
  reg [3:0] image_466; // @[Filter.scala 68:24]
  reg [3:0] image_467; // @[Filter.scala 68:24]
  reg [3:0] image_468; // @[Filter.scala 68:24]
  reg [3:0] image_469; // @[Filter.scala 68:24]
  reg [3:0] image_470; // @[Filter.scala 68:24]
  reg [3:0] image_471; // @[Filter.scala 68:24]
  reg [3:0] image_472; // @[Filter.scala 68:24]
  reg [3:0] image_473; // @[Filter.scala 68:24]
  reg [3:0] image_474; // @[Filter.scala 68:24]
  reg [3:0] image_475; // @[Filter.scala 68:24]
  reg [3:0] image_476; // @[Filter.scala 68:24]
  reg [3:0] image_477; // @[Filter.scala 68:24]
  reg [3:0] image_478; // @[Filter.scala 68:24]
  reg [3:0] image_479; // @[Filter.scala 68:24]
  reg [3:0] image_480; // @[Filter.scala 68:24]
  reg [3:0] image_481; // @[Filter.scala 68:24]
  reg [3:0] image_482; // @[Filter.scala 68:24]
  reg [3:0] image_483; // @[Filter.scala 68:24]
  reg [3:0] image_484; // @[Filter.scala 68:24]
  reg [3:0] image_485; // @[Filter.scala 68:24]
  reg [3:0] image_486; // @[Filter.scala 68:24]
  reg [3:0] image_487; // @[Filter.scala 68:24]
  reg [3:0] image_488; // @[Filter.scala 68:24]
  reg [3:0] image_489; // @[Filter.scala 68:24]
  reg [3:0] image_490; // @[Filter.scala 68:24]
  reg [3:0] image_491; // @[Filter.scala 68:24]
  reg [3:0] image_492; // @[Filter.scala 68:24]
  reg [3:0] image_493; // @[Filter.scala 68:24]
  reg [3:0] image_494; // @[Filter.scala 68:24]
  reg [3:0] image_495; // @[Filter.scala 68:24]
  reg [3:0] image_496; // @[Filter.scala 68:24]
  reg [3:0] image_497; // @[Filter.scala 68:24]
  reg [3:0] image_498; // @[Filter.scala 68:24]
  reg [3:0] image_499; // @[Filter.scala 68:24]
  reg [3:0] image_500; // @[Filter.scala 68:24]
  reg [3:0] image_501; // @[Filter.scala 68:24]
  reg [3:0] image_502; // @[Filter.scala 68:24]
  reg [3:0] image_503; // @[Filter.scala 68:24]
  reg [3:0] image_504; // @[Filter.scala 68:24]
  reg [3:0] image_505; // @[Filter.scala 68:24]
  reg [3:0] image_506; // @[Filter.scala 68:24]
  reg [3:0] image_507; // @[Filter.scala 68:24]
  reg [3:0] image_508; // @[Filter.scala 68:24]
  reg [3:0] image_509; // @[Filter.scala 68:24]
  reg [3:0] image_515; // @[Filter.scala 68:24]
  reg [3:0] image_516; // @[Filter.scala 68:24]
  reg [3:0] image_517; // @[Filter.scala 68:24]
  reg [3:0] image_518; // @[Filter.scala 68:24]
  reg [3:0] image_519; // @[Filter.scala 68:24]
  reg [3:0] image_520; // @[Filter.scala 68:24]
  reg [3:0] image_521; // @[Filter.scala 68:24]
  reg [3:0] image_522; // @[Filter.scala 68:24]
  reg [3:0] image_523; // @[Filter.scala 68:24]
  reg [3:0] image_524; // @[Filter.scala 68:24]
  reg [3:0] image_525; // @[Filter.scala 68:24]
  reg [3:0] image_526; // @[Filter.scala 68:24]
  reg [3:0] image_527; // @[Filter.scala 68:24]
  reg [3:0] image_528; // @[Filter.scala 68:24]
  reg [3:0] image_529; // @[Filter.scala 68:24]
  reg [3:0] image_530; // @[Filter.scala 68:24]
  reg [3:0] image_531; // @[Filter.scala 68:24]
  reg [3:0] image_532; // @[Filter.scala 68:24]
  reg [3:0] image_533; // @[Filter.scala 68:24]
  reg [3:0] image_534; // @[Filter.scala 68:24]
  reg [3:0] image_535; // @[Filter.scala 68:24]
  reg [3:0] image_536; // @[Filter.scala 68:24]
  reg [3:0] image_537; // @[Filter.scala 68:24]
  reg [3:0] image_538; // @[Filter.scala 68:24]
  reg [3:0] image_539; // @[Filter.scala 68:24]
  reg [3:0] image_540; // @[Filter.scala 68:24]
  reg [3:0] image_541; // @[Filter.scala 68:24]
  reg [3:0] image_542; // @[Filter.scala 68:24]
  reg [3:0] image_543; // @[Filter.scala 68:24]
  reg [3:0] image_544; // @[Filter.scala 68:24]
  reg [3:0] image_545; // @[Filter.scala 68:24]
  reg [3:0] image_546; // @[Filter.scala 68:24]
  reg [3:0] image_547; // @[Filter.scala 68:24]
  reg [3:0] image_548; // @[Filter.scala 68:24]
  reg [3:0] image_549; // @[Filter.scala 68:24]
  reg [3:0] image_550; // @[Filter.scala 68:24]
  reg [3:0] image_551; // @[Filter.scala 68:24]
  reg [3:0] image_552; // @[Filter.scala 68:24]
  reg [3:0] image_553; // @[Filter.scala 68:24]
  reg [3:0] image_554; // @[Filter.scala 68:24]
  reg [3:0] image_555; // @[Filter.scala 68:24]
  reg [3:0] image_556; // @[Filter.scala 68:24]
  reg [3:0] image_557; // @[Filter.scala 68:24]
  reg [3:0] image_558; // @[Filter.scala 68:24]
  reg [3:0] image_559; // @[Filter.scala 68:24]
  reg [3:0] image_560; // @[Filter.scala 68:24]
  reg [3:0] image_561; // @[Filter.scala 68:24]
  reg [3:0] image_562; // @[Filter.scala 68:24]
  reg [3:0] image_563; // @[Filter.scala 68:24]
  reg [3:0] image_564; // @[Filter.scala 68:24]
  reg [3:0] image_565; // @[Filter.scala 68:24]
  reg [3:0] image_566; // @[Filter.scala 68:24]
  reg [3:0] image_571; // @[Filter.scala 68:24]
  reg [3:0] image_572; // @[Filter.scala 68:24]
  reg [3:0] image_573; // @[Filter.scala 68:24]
  reg [3:0] image_574; // @[Filter.scala 68:24]
  reg [3:0] image_578; // @[Filter.scala 68:24]
  reg [3:0] image_579; // @[Filter.scala 68:24]
  reg [3:0] image_580; // @[Filter.scala 68:24]
  reg [3:0] image_581; // @[Filter.scala 68:24]
  reg [3:0] image_582; // @[Filter.scala 68:24]
  reg [3:0] image_583; // @[Filter.scala 68:24]
  reg [3:0] image_584; // @[Filter.scala 68:24]
  reg [3:0] image_585; // @[Filter.scala 68:24]
  reg [3:0] image_586; // @[Filter.scala 68:24]
  reg [3:0] image_587; // @[Filter.scala 68:24]
  reg [3:0] image_588; // @[Filter.scala 68:24]
  reg [3:0] image_589; // @[Filter.scala 68:24]
  reg [3:0] image_590; // @[Filter.scala 68:24]
  reg [3:0] image_591; // @[Filter.scala 68:24]
  reg [3:0] image_592; // @[Filter.scala 68:24]
  reg [3:0] image_593; // @[Filter.scala 68:24]
  reg [3:0] image_594; // @[Filter.scala 68:24]
  reg [3:0] image_595; // @[Filter.scala 68:24]
  reg [3:0] image_596; // @[Filter.scala 68:24]
  reg [3:0] image_597; // @[Filter.scala 68:24]
  reg [3:0] image_598; // @[Filter.scala 68:24]
  reg [3:0] image_599; // @[Filter.scala 68:24]
  reg [3:0] image_600; // @[Filter.scala 68:24]
  reg [3:0] image_601; // @[Filter.scala 68:24]
  reg [3:0] image_602; // @[Filter.scala 68:24]
  reg [3:0] image_603; // @[Filter.scala 68:24]
  reg [3:0] image_604; // @[Filter.scala 68:24]
  reg [3:0] image_605; // @[Filter.scala 68:24]
  reg [3:0] image_606; // @[Filter.scala 68:24]
  reg [3:0] image_607; // @[Filter.scala 68:24]
  reg [3:0] image_614; // @[Filter.scala 68:24]
  reg [3:0] image_615; // @[Filter.scala 68:24]
  reg [3:0] image_616; // @[Filter.scala 68:24]
  reg [3:0] image_617; // @[Filter.scala 68:24]
  reg [3:0] image_618; // @[Filter.scala 68:24]
  reg [3:0] image_619; // @[Filter.scala 68:24]
  reg [3:0] image_620; // @[Filter.scala 68:24]
  reg [3:0] image_621; // @[Filter.scala 68:24]
  reg [3:0] image_622; // @[Filter.scala 68:24]
  reg [3:0] image_623; // @[Filter.scala 68:24]
  reg [3:0] image_624; // @[Filter.scala 68:24]
  reg [3:0] image_625; // @[Filter.scala 68:24]
  reg [3:0] image_626; // @[Filter.scala 68:24]
  reg [3:0] image_627; // @[Filter.scala 68:24]
  reg [3:0] image_628; // @[Filter.scala 68:24]
  reg [3:0] image_636; // @[Filter.scala 68:24]
  reg [3:0] image_637; // @[Filter.scala 68:24]
  reg [3:0] image_638; // @[Filter.scala 68:24]
  reg [3:0] image_639; // @[Filter.scala 68:24]
  reg [3:0] image_642; // @[Filter.scala 68:24]
  reg [3:0] image_643; // @[Filter.scala 68:24]
  reg [3:0] image_644; // @[Filter.scala 68:24]
  reg [3:0] image_645; // @[Filter.scala 68:24]
  reg [3:0] image_646; // @[Filter.scala 68:24]
  reg [3:0] image_647; // @[Filter.scala 68:24]
  reg [3:0] image_648; // @[Filter.scala 68:24]
  reg [3:0] image_649; // @[Filter.scala 68:24]
  reg [3:0] image_650; // @[Filter.scala 68:24]
  reg [3:0] image_651; // @[Filter.scala 68:24]
  reg [3:0] image_652; // @[Filter.scala 68:24]
  reg [3:0] image_653; // @[Filter.scala 68:24]
  reg [3:0] image_654; // @[Filter.scala 68:24]
  reg [3:0] image_655; // @[Filter.scala 68:24]
  reg [3:0] image_656; // @[Filter.scala 68:24]
  reg [3:0] image_657; // @[Filter.scala 68:24]
  reg [3:0] image_658; // @[Filter.scala 68:24]
  reg [3:0] image_659; // @[Filter.scala 68:24]
  reg [3:0] image_660; // @[Filter.scala 68:24]
  reg [3:0] image_661; // @[Filter.scala 68:24]
  reg [3:0] image_662; // @[Filter.scala 68:24]
  reg [3:0] image_663; // @[Filter.scala 68:24]
  reg [3:0] image_664; // @[Filter.scala 68:24]
  reg [3:0] image_665; // @[Filter.scala 68:24]
  reg [3:0] image_666; // @[Filter.scala 68:24]
  reg [3:0] image_667; // @[Filter.scala 68:24]
  reg [3:0] image_668; // @[Filter.scala 68:24]
  reg [3:0] image_669; // @[Filter.scala 68:24]
  reg [3:0] image_670; // @[Filter.scala 68:24]
  reg [3:0] image_679; // @[Filter.scala 68:24]
  reg [3:0] image_680; // @[Filter.scala 68:24]
  reg [3:0] image_681; // @[Filter.scala 68:24]
  reg [3:0] image_682; // @[Filter.scala 68:24]
  reg [3:0] image_683; // @[Filter.scala 68:24]
  reg [3:0] image_684; // @[Filter.scala 68:24]
  reg [3:0] image_685; // @[Filter.scala 68:24]
  reg [3:0] image_686; // @[Filter.scala 68:24]
  reg [3:0] image_687; // @[Filter.scala 68:24]
  reg [3:0] image_688; // @[Filter.scala 68:24]
  reg [3:0] image_689; // @[Filter.scala 68:24]
  reg [3:0] image_690; // @[Filter.scala 68:24]
  reg [3:0] image_691; // @[Filter.scala 68:24]
  reg [3:0] image_692; // @[Filter.scala 68:24]
  reg [3:0] image_693; // @[Filter.scala 68:24]
  reg [3:0] image_694; // @[Filter.scala 68:24]
  reg [3:0] image_695; // @[Filter.scala 68:24]
  reg [3:0] image_696; // @[Filter.scala 68:24]
  reg [3:0] image_697; // @[Filter.scala 68:24]
  reg [3:0] image_698; // @[Filter.scala 68:24]
  reg [3:0] image_701; // @[Filter.scala 68:24]
  reg [3:0] image_702; // @[Filter.scala 68:24]
  reg [3:0] image_703; // @[Filter.scala 68:24]
  reg [3:0] image_705; // @[Filter.scala 68:24]
  reg [3:0] image_706; // @[Filter.scala 68:24]
  reg [3:0] image_707; // @[Filter.scala 68:24]
  reg [3:0] image_708; // @[Filter.scala 68:24]
  reg [3:0] image_709; // @[Filter.scala 68:24]
  reg [3:0] image_710; // @[Filter.scala 68:24]
  reg [3:0] image_711; // @[Filter.scala 68:24]
  reg [3:0] image_712; // @[Filter.scala 68:24]
  reg [3:0] image_713; // @[Filter.scala 68:24]
  reg [3:0] image_714; // @[Filter.scala 68:24]
  reg [3:0] image_715; // @[Filter.scala 68:24]
  reg [3:0] image_716; // @[Filter.scala 68:24]
  reg [3:0] image_717; // @[Filter.scala 68:24]
  reg [3:0] image_718; // @[Filter.scala 68:24]
  reg [3:0] image_719; // @[Filter.scala 68:24]
  reg [3:0] image_720; // @[Filter.scala 68:24]
  reg [3:0] image_721; // @[Filter.scala 68:24]
  reg [3:0] image_722; // @[Filter.scala 68:24]
  reg [3:0] image_723; // @[Filter.scala 68:24]
  reg [3:0] image_724; // @[Filter.scala 68:24]
  reg [3:0] image_725; // @[Filter.scala 68:24]
  reg [3:0] image_726; // @[Filter.scala 68:24]
  reg [3:0] image_727; // @[Filter.scala 68:24]
  reg [3:0] image_728; // @[Filter.scala 68:24]
  reg [3:0] image_729; // @[Filter.scala 68:24]
  reg [3:0] image_730; // @[Filter.scala 68:24]
  reg [3:0] image_731; // @[Filter.scala 68:24]
  reg [3:0] image_732; // @[Filter.scala 68:24]
  reg [3:0] image_733; // @[Filter.scala 68:24]
  reg [3:0] image_734; // @[Filter.scala 68:24]
  reg [3:0] image_736; // @[Filter.scala 68:24]
  reg [3:0] image_737; // @[Filter.scala 68:24]
  reg [3:0] image_739; // @[Filter.scala 68:24]
  reg [3:0] image_740; // @[Filter.scala 68:24]
  reg [3:0] image_741; // @[Filter.scala 68:24]
  reg [3:0] image_744; // @[Filter.scala 68:24]
  reg [3:0] image_745; // @[Filter.scala 68:24]
  reg [3:0] image_746; // @[Filter.scala 68:24]
  reg [3:0] image_747; // @[Filter.scala 68:24]
  reg [3:0] image_748; // @[Filter.scala 68:24]
  reg [3:0] image_749; // @[Filter.scala 68:24]
  reg [3:0] image_750; // @[Filter.scala 68:24]
  reg [3:0] image_751; // @[Filter.scala 68:24]
  reg [3:0] image_752; // @[Filter.scala 68:24]
  reg [3:0] image_753; // @[Filter.scala 68:24]
  reg [3:0] image_754; // @[Filter.scala 68:24]
  reg [3:0] image_755; // @[Filter.scala 68:24]
  reg [3:0] image_756; // @[Filter.scala 68:24]
  reg [3:0] image_758; // @[Filter.scala 68:24]
  reg [3:0] image_760; // @[Filter.scala 68:24]
  reg [3:0] image_761; // @[Filter.scala 68:24]
  reg [3:0] image_762; // @[Filter.scala 68:24]
  reg [3:0] image_763; // @[Filter.scala 68:24]
  reg [3:0] image_765; // @[Filter.scala 68:24]
  reg [3:0] image_766; // @[Filter.scala 68:24]
  reg [3:0] image_767; // @[Filter.scala 68:24]
  reg [3:0] image_768; // @[Filter.scala 68:24]
  reg [3:0] image_769; // @[Filter.scala 68:24]
  reg [3:0] image_770; // @[Filter.scala 68:24]
  reg [3:0] image_771; // @[Filter.scala 68:24]
  reg [3:0] image_772; // @[Filter.scala 68:24]
  reg [3:0] image_773; // @[Filter.scala 68:24]
  reg [3:0] image_774; // @[Filter.scala 68:24]
  reg [3:0] image_775; // @[Filter.scala 68:24]
  reg [3:0] image_776; // @[Filter.scala 68:24]
  reg [3:0] image_777; // @[Filter.scala 68:24]
  reg [3:0] image_778; // @[Filter.scala 68:24]
  reg [3:0] image_779; // @[Filter.scala 68:24]
  reg [3:0] image_780; // @[Filter.scala 68:24]
  reg [3:0] image_781; // @[Filter.scala 68:24]
  reg [3:0] image_782; // @[Filter.scala 68:24]
  reg [3:0] image_783; // @[Filter.scala 68:24]
  reg [3:0] image_784; // @[Filter.scala 68:24]
  reg [3:0] image_785; // @[Filter.scala 68:24]
  reg [3:0] image_786; // @[Filter.scala 68:24]
  reg [3:0] image_787; // @[Filter.scala 68:24]
  reg [3:0] image_788; // @[Filter.scala 68:24]
  reg [3:0] image_789; // @[Filter.scala 68:24]
  reg [3:0] image_790; // @[Filter.scala 68:24]
  reg [3:0] image_791; // @[Filter.scala 68:24]
  reg [3:0] image_792; // @[Filter.scala 68:24]
  reg [3:0] image_793; // @[Filter.scala 68:24]
  reg [3:0] image_794; // @[Filter.scala 68:24]
  reg [3:0] image_795; // @[Filter.scala 68:24]
  reg [3:0] image_796; // @[Filter.scala 68:24]
  reg [3:0] image_797; // @[Filter.scala 68:24]
  reg [3:0] image_800; // @[Filter.scala 68:24]
  reg [3:0] image_801; // @[Filter.scala 68:24]
  reg [3:0] image_802; // @[Filter.scala 68:24]
  reg [3:0] image_803; // @[Filter.scala 68:24]
  reg [3:0] image_804; // @[Filter.scala 68:24]
  reg [3:0] image_805; // @[Filter.scala 68:24]
  reg [3:0] image_806; // @[Filter.scala 68:24]
  reg [3:0] image_808; // @[Filter.scala 68:24]
  reg [3:0] image_809; // @[Filter.scala 68:24]
  reg [3:0] image_810; // @[Filter.scala 68:24]
  reg [3:0] image_811; // @[Filter.scala 68:24]
  reg [3:0] image_812; // @[Filter.scala 68:24]
  reg [3:0] image_813; // @[Filter.scala 68:24]
  reg [3:0] image_814; // @[Filter.scala 68:24]
  reg [3:0] image_815; // @[Filter.scala 68:24]
  reg [3:0] image_816; // @[Filter.scala 68:24]
  reg [3:0] image_817; // @[Filter.scala 68:24]
  reg [3:0] image_818; // @[Filter.scala 68:24]
  reg [3:0] image_819; // @[Filter.scala 68:24]
  reg [3:0] image_820; // @[Filter.scala 68:24]
  reg [3:0] image_822; // @[Filter.scala 68:24]
  reg [3:0] image_823; // @[Filter.scala 68:24]
  reg [3:0] image_824; // @[Filter.scala 68:24]
  reg [3:0] image_825; // @[Filter.scala 68:24]
  reg [3:0] image_826; // @[Filter.scala 68:24]
  reg [3:0] image_828; // @[Filter.scala 68:24]
  reg [3:0] image_829; // @[Filter.scala 68:24]
  reg [3:0] image_830; // @[Filter.scala 68:24]
  reg [3:0] image_831; // @[Filter.scala 68:24]
  reg [3:0] image_833; // @[Filter.scala 68:24]
  reg [3:0] image_834; // @[Filter.scala 68:24]
  reg [3:0] image_835; // @[Filter.scala 68:24]
  reg [3:0] image_836; // @[Filter.scala 68:24]
  reg [3:0] image_837; // @[Filter.scala 68:24]
  reg [3:0] image_838; // @[Filter.scala 68:24]
  reg [3:0] image_839; // @[Filter.scala 68:24]
  reg [3:0] image_840; // @[Filter.scala 68:24]
  reg [3:0] image_841; // @[Filter.scala 68:24]
  reg [3:0] image_842; // @[Filter.scala 68:24]
  reg [3:0] image_843; // @[Filter.scala 68:24]
  reg [3:0] image_844; // @[Filter.scala 68:24]
  reg [3:0] image_845; // @[Filter.scala 68:24]
  reg [3:0] image_846; // @[Filter.scala 68:24]
  reg [3:0] image_847; // @[Filter.scala 68:24]
  reg [3:0] image_848; // @[Filter.scala 68:24]
  reg [3:0] image_849; // @[Filter.scala 68:24]
  reg [3:0] image_850; // @[Filter.scala 68:24]
  reg [3:0] image_851; // @[Filter.scala 68:24]
  reg [3:0] image_852; // @[Filter.scala 68:24]
  reg [3:0] image_853; // @[Filter.scala 68:24]
  reg [3:0] image_854; // @[Filter.scala 68:24]
  reg [3:0] image_855; // @[Filter.scala 68:24]
  reg [3:0] image_856; // @[Filter.scala 68:24]
  reg [3:0] image_857; // @[Filter.scala 68:24]
  reg [3:0] image_858; // @[Filter.scala 68:24]
  reg [3:0] image_859; // @[Filter.scala 68:24]
  reg [3:0] image_860; // @[Filter.scala 68:24]
  reg [3:0] image_861; // @[Filter.scala 68:24]
  reg [3:0] image_862; // @[Filter.scala 68:24]
  reg [3:0] image_865; // @[Filter.scala 68:24]
  reg [3:0] image_866; // @[Filter.scala 68:24]
  reg [3:0] image_867; // @[Filter.scala 68:24]
  reg [3:0] image_868; // @[Filter.scala 68:24]
  reg [3:0] image_869; // @[Filter.scala 68:24]
  reg [3:0] image_872; // @[Filter.scala 68:24]
  reg [3:0] image_873; // @[Filter.scala 68:24]
  reg [3:0] image_874; // @[Filter.scala 68:24]
  reg [3:0] image_875; // @[Filter.scala 68:24]
  reg [3:0] image_876; // @[Filter.scala 68:24]
  reg [3:0] image_877; // @[Filter.scala 68:24]
  reg [3:0] image_878; // @[Filter.scala 68:24]
  reg [3:0] image_879; // @[Filter.scala 68:24]
  reg [3:0] image_880; // @[Filter.scala 68:24]
  reg [3:0] image_881; // @[Filter.scala 68:24]
  reg [3:0] image_882; // @[Filter.scala 68:24]
  reg [3:0] image_883; // @[Filter.scala 68:24]
  reg [3:0] image_884; // @[Filter.scala 68:24]
  reg [3:0] image_885; // @[Filter.scala 68:24]
  reg [3:0] image_891; // @[Filter.scala 68:24]
  reg [3:0] image_892; // @[Filter.scala 68:24]
  reg [3:0] image_893; // @[Filter.scala 68:24]
  reg [3:0] image_894; // @[Filter.scala 68:24]
  reg [3:0] image_895; // @[Filter.scala 68:24]
  reg [3:0] image_897; // @[Filter.scala 68:24]
  reg [3:0] image_898; // @[Filter.scala 68:24]
  reg [3:0] image_899; // @[Filter.scala 68:24]
  reg [3:0] image_900; // @[Filter.scala 68:24]
  reg [3:0] image_901; // @[Filter.scala 68:24]
  reg [3:0] image_902; // @[Filter.scala 68:24]
  reg [3:0] image_903; // @[Filter.scala 68:24]
  reg [3:0] image_904; // @[Filter.scala 68:24]
  reg [3:0] image_905; // @[Filter.scala 68:24]
  reg [3:0] image_906; // @[Filter.scala 68:24]
  reg [3:0] image_907; // @[Filter.scala 68:24]
  reg [3:0] image_908; // @[Filter.scala 68:24]
  reg [3:0] image_909; // @[Filter.scala 68:24]
  reg [3:0] image_910; // @[Filter.scala 68:24]
  reg [3:0] image_911; // @[Filter.scala 68:24]
  reg [3:0] image_912; // @[Filter.scala 68:24]
  reg [3:0] image_913; // @[Filter.scala 68:24]
  reg [3:0] image_914; // @[Filter.scala 68:24]
  reg [3:0] image_915; // @[Filter.scala 68:24]
  reg [3:0] image_916; // @[Filter.scala 68:24]
  reg [3:0] image_917; // @[Filter.scala 68:24]
  reg [3:0] image_918; // @[Filter.scala 68:24]
  reg [3:0] image_919; // @[Filter.scala 68:24]
  reg [3:0] image_920; // @[Filter.scala 68:24]
  reg [3:0] image_921; // @[Filter.scala 68:24]
  reg [3:0] image_922; // @[Filter.scala 68:24]
  reg [3:0] image_923; // @[Filter.scala 68:24]
  reg [3:0] image_924; // @[Filter.scala 68:24]
  reg [3:0] image_925; // @[Filter.scala 68:24]
  reg [3:0] image_926; // @[Filter.scala 68:24]
  reg [3:0] image_927; // @[Filter.scala 68:24]
  reg [3:0] image_929; // @[Filter.scala 68:24]
  reg [3:0] image_930; // @[Filter.scala 68:24]
  reg [3:0] image_935; // @[Filter.scala 68:24]
  reg [3:0] image_936; // @[Filter.scala 68:24]
  reg [3:0] image_937; // @[Filter.scala 68:24]
  reg [3:0] image_938; // @[Filter.scala 68:24]
  reg [3:0] image_939; // @[Filter.scala 68:24]
  reg [3:0] image_940; // @[Filter.scala 68:24]
  reg [3:0] image_941; // @[Filter.scala 68:24]
  reg [3:0] image_942; // @[Filter.scala 68:24]
  reg [3:0] image_943; // @[Filter.scala 68:24]
  reg [3:0] image_944; // @[Filter.scala 68:24]
  reg [3:0] image_945; // @[Filter.scala 68:24]
  reg [3:0] image_946; // @[Filter.scala 68:24]
  reg [3:0] image_947; // @[Filter.scala 68:24]
  reg [3:0] image_948; // @[Filter.scala 68:24]
  reg [3:0] image_949; // @[Filter.scala 68:24]
  reg [3:0] image_950; // @[Filter.scala 68:24]
  reg [3:0] image_951; // @[Filter.scala 68:24]
  reg [3:0] image_952; // @[Filter.scala 68:24]
  reg [3:0] image_953; // @[Filter.scala 68:24]
  reg [3:0] image_954; // @[Filter.scala 68:24]
  reg [3:0] image_955; // @[Filter.scala 68:24]
  reg [3:0] image_956; // @[Filter.scala 68:24]
  reg [3:0] image_957; // @[Filter.scala 68:24]
  reg [3:0] image_958; // @[Filter.scala 68:24]
  reg [3:0] image_959; // @[Filter.scala 68:24]
  reg [3:0] image_961; // @[Filter.scala 68:24]
  reg [3:0] image_962; // @[Filter.scala 68:24]
  reg [3:0] image_963; // @[Filter.scala 68:24]
  reg [3:0] image_964; // @[Filter.scala 68:24]
  reg [3:0] image_965; // @[Filter.scala 68:24]
  reg [3:0] image_966; // @[Filter.scala 68:24]
  reg [3:0] image_967; // @[Filter.scala 68:24]
  reg [3:0] image_968; // @[Filter.scala 68:24]
  reg [3:0] image_969; // @[Filter.scala 68:24]
  reg [3:0] image_970; // @[Filter.scala 68:24]
  reg [3:0] image_971; // @[Filter.scala 68:24]
  reg [3:0] image_972; // @[Filter.scala 68:24]
  reg [3:0] image_973; // @[Filter.scala 68:24]
  reg [3:0] image_974; // @[Filter.scala 68:24]
  reg [3:0] image_975; // @[Filter.scala 68:24]
  reg [3:0] image_976; // @[Filter.scala 68:24]
  reg [3:0] image_977; // @[Filter.scala 68:24]
  reg [3:0] image_978; // @[Filter.scala 68:24]
  reg [3:0] image_979; // @[Filter.scala 68:24]
  reg [3:0] image_980; // @[Filter.scala 68:24]
  reg [3:0] image_981; // @[Filter.scala 68:24]
  reg [3:0] image_982; // @[Filter.scala 68:24]
  reg [3:0] image_983; // @[Filter.scala 68:24]
  reg [3:0] image_984; // @[Filter.scala 68:24]
  reg [3:0] image_985; // @[Filter.scala 68:24]
  reg [3:0] image_986; // @[Filter.scala 68:24]
  reg [3:0] image_987; // @[Filter.scala 68:24]
  reg [3:0] image_988; // @[Filter.scala 68:24]
  reg [3:0] image_989; // @[Filter.scala 68:24]
  reg [3:0] image_990; // @[Filter.scala 68:24]
  reg [3:0] image_991; // @[Filter.scala 68:24]
  reg [3:0] image_992; // @[Filter.scala 68:24]
  reg [3:0] image_997; // @[Filter.scala 68:24]
  reg [3:0] image_998; // @[Filter.scala 68:24]
  reg [3:0] image_999; // @[Filter.scala 68:24]
  reg [3:0] image_1000; // @[Filter.scala 68:24]
  reg [3:0] image_1001; // @[Filter.scala 68:24]
  reg [3:0] image_1002; // @[Filter.scala 68:24]
  reg [3:0] image_1003; // @[Filter.scala 68:24]
  reg [3:0] image_1004; // @[Filter.scala 68:24]
  reg [3:0] image_1005; // @[Filter.scala 68:24]
  reg [3:0] image_1006; // @[Filter.scala 68:24]
  reg [3:0] image_1007; // @[Filter.scala 68:24]
  reg [3:0] image_1008; // @[Filter.scala 68:24]
  reg [3:0] image_1009; // @[Filter.scala 68:24]
  reg [3:0] image_1010; // @[Filter.scala 68:24]
  reg [3:0] image_1011; // @[Filter.scala 68:24]
  reg [3:0] image_1012; // @[Filter.scala 68:24]
  reg [3:0] image_1013; // @[Filter.scala 68:24]
  reg [3:0] image_1014; // @[Filter.scala 68:24]
  reg [3:0] image_1015; // @[Filter.scala 68:24]
  reg [3:0] image_1016; // @[Filter.scala 68:24]
  reg [3:0] image_1017; // @[Filter.scala 68:24]
  reg [3:0] image_1018; // @[Filter.scala 68:24]
  reg [3:0] image_1019; // @[Filter.scala 68:24]
  reg [3:0] image_1020; // @[Filter.scala 68:24]
  reg [3:0] image_1024; // @[Filter.scala 68:24]
  reg [3:0] image_1025; // @[Filter.scala 68:24]
  reg [3:0] image_1026; // @[Filter.scala 68:24]
  reg [3:0] image_1027; // @[Filter.scala 68:24]
  reg [3:0] image_1028; // @[Filter.scala 68:24]
  reg [3:0] image_1029; // @[Filter.scala 68:24]
  reg [3:0] image_1030; // @[Filter.scala 68:24]
  reg [3:0] image_1031; // @[Filter.scala 68:24]
  reg [3:0] image_1032; // @[Filter.scala 68:24]
  reg [3:0] image_1033; // @[Filter.scala 68:24]
  reg [3:0] image_1034; // @[Filter.scala 68:24]
  reg [3:0] image_1035; // @[Filter.scala 68:24]
  reg [3:0] image_1036; // @[Filter.scala 68:24]
  reg [3:0] image_1037; // @[Filter.scala 68:24]
  reg [3:0] image_1038; // @[Filter.scala 68:24]
  reg [3:0] image_1039; // @[Filter.scala 68:24]
  reg [3:0] image_1040; // @[Filter.scala 68:24]
  reg [3:0] image_1041; // @[Filter.scala 68:24]
  reg [3:0] image_1042; // @[Filter.scala 68:24]
  reg [3:0] image_1043; // @[Filter.scala 68:24]
  reg [3:0] image_1044; // @[Filter.scala 68:24]
  reg [3:0] image_1045; // @[Filter.scala 68:24]
  reg [3:0] image_1046; // @[Filter.scala 68:24]
  reg [3:0] image_1047; // @[Filter.scala 68:24]
  reg [3:0] image_1048; // @[Filter.scala 68:24]
  reg [3:0] image_1049; // @[Filter.scala 68:24]
  reg [3:0] image_1050; // @[Filter.scala 68:24]
  reg [3:0] image_1051; // @[Filter.scala 68:24]
  reg [3:0] image_1052; // @[Filter.scala 68:24]
  reg [3:0] image_1053; // @[Filter.scala 68:24]
  reg [3:0] image_1054; // @[Filter.scala 68:24]
  reg [3:0] image_1055; // @[Filter.scala 68:24]
  reg [3:0] image_1056; // @[Filter.scala 68:24]
  reg [3:0] image_1057; // @[Filter.scala 68:24]
  reg [3:0] image_1058; // @[Filter.scala 68:24]
  reg [3:0] image_1059; // @[Filter.scala 68:24]
  reg [3:0] image_1060; // @[Filter.scala 68:24]
  reg [3:0] image_1061; // @[Filter.scala 68:24]
  reg [3:0] image_1062; // @[Filter.scala 68:24]
  reg [3:0] image_1063; // @[Filter.scala 68:24]
  reg [3:0] image_1064; // @[Filter.scala 68:24]
  reg [3:0] image_1065; // @[Filter.scala 68:24]
  reg [3:0] image_1066; // @[Filter.scala 68:24]
  reg [3:0] image_1067; // @[Filter.scala 68:24]
  reg [3:0] image_1068; // @[Filter.scala 68:24]
  reg [3:0] image_1069; // @[Filter.scala 68:24]
  reg [3:0] image_1070; // @[Filter.scala 68:24]
  reg [3:0] image_1071; // @[Filter.scala 68:24]
  reg [3:0] image_1072; // @[Filter.scala 68:24]
  reg [3:0] image_1073; // @[Filter.scala 68:24]
  reg [3:0] image_1074; // @[Filter.scala 68:24]
  reg [3:0] image_1075; // @[Filter.scala 68:24]
  reg [3:0] image_1076; // @[Filter.scala 68:24]
  reg [3:0] image_1077; // @[Filter.scala 68:24]
  reg [3:0] image_1078; // @[Filter.scala 68:24]
  reg [3:0] image_1079; // @[Filter.scala 68:24]
  reg [3:0] image_1080; // @[Filter.scala 68:24]
  reg [3:0] image_1081; // @[Filter.scala 68:24]
  reg [3:0] image_1082; // @[Filter.scala 68:24]
  reg [3:0] image_1083; // @[Filter.scala 68:24]
  reg [3:0] image_1084; // @[Filter.scala 68:24]
  reg [3:0] image_1085; // @[Filter.scala 68:24]
  reg [3:0] image_1088; // @[Filter.scala 68:24]
  reg [3:0] image_1089; // @[Filter.scala 68:24]
  reg [3:0] image_1090; // @[Filter.scala 68:24]
  reg [3:0] image_1091; // @[Filter.scala 68:24]
  reg [3:0] image_1092; // @[Filter.scala 68:24]
  reg [3:0] image_1093; // @[Filter.scala 68:24]
  reg [3:0] image_1094; // @[Filter.scala 68:24]
  reg [3:0] image_1095; // @[Filter.scala 68:24]
  reg [3:0] image_1096; // @[Filter.scala 68:24]
  reg [3:0] image_1097; // @[Filter.scala 68:24]
  reg [3:0] image_1098; // @[Filter.scala 68:24]
  reg [3:0] image_1099; // @[Filter.scala 68:24]
  reg [3:0] image_1100; // @[Filter.scala 68:24]
  reg [3:0] image_1101; // @[Filter.scala 68:24]
  reg [3:0] image_1102; // @[Filter.scala 68:24]
  reg [3:0] image_1103; // @[Filter.scala 68:24]
  reg [3:0] image_1104; // @[Filter.scala 68:24]
  reg [3:0] image_1105; // @[Filter.scala 68:24]
  reg [3:0] image_1106; // @[Filter.scala 68:24]
  reg [3:0] image_1107; // @[Filter.scala 68:24]
  reg [3:0] image_1108; // @[Filter.scala 68:24]
  reg [3:0] image_1109; // @[Filter.scala 68:24]
  reg [3:0] image_1110; // @[Filter.scala 68:24]
  reg [3:0] image_1111; // @[Filter.scala 68:24]
  reg [3:0] image_1112; // @[Filter.scala 68:24]
  reg [3:0] image_1113; // @[Filter.scala 68:24]
  reg [3:0] image_1114; // @[Filter.scala 68:24]
  reg [3:0] image_1115; // @[Filter.scala 68:24]
  reg [3:0] image_1116; // @[Filter.scala 68:24]
  reg [3:0] image_1117; // @[Filter.scala 68:24]
  reg [3:0] image_1118; // @[Filter.scala 68:24]
  reg [3:0] image_1119; // @[Filter.scala 68:24]
  reg [3:0] image_1120; // @[Filter.scala 68:24]
  reg [3:0] image_1121; // @[Filter.scala 68:24]
  reg [3:0] image_1122; // @[Filter.scala 68:24]
  reg [3:0] image_1123; // @[Filter.scala 68:24]
  reg [3:0] image_1124; // @[Filter.scala 68:24]
  reg [3:0] image_1125; // @[Filter.scala 68:24]
  reg [3:0] image_1126; // @[Filter.scala 68:24]
  reg [3:0] image_1127; // @[Filter.scala 68:24]
  reg [3:0] image_1128; // @[Filter.scala 68:24]
  reg [3:0] image_1129; // @[Filter.scala 68:24]
  reg [3:0] image_1130; // @[Filter.scala 68:24]
  reg [3:0] image_1131; // @[Filter.scala 68:24]
  reg [3:0] image_1132; // @[Filter.scala 68:24]
  reg [3:0] image_1133; // @[Filter.scala 68:24]
  reg [3:0] image_1134; // @[Filter.scala 68:24]
  reg [3:0] image_1135; // @[Filter.scala 68:24]
  reg [3:0] image_1136; // @[Filter.scala 68:24]
  reg [3:0] image_1137; // @[Filter.scala 68:24]
  reg [3:0] image_1138; // @[Filter.scala 68:24]
  reg [3:0] image_1139; // @[Filter.scala 68:24]
  reg [3:0] image_1140; // @[Filter.scala 68:24]
  reg [3:0] image_1141; // @[Filter.scala 68:24]
  reg [3:0] image_1142; // @[Filter.scala 68:24]
  reg [3:0] image_1143; // @[Filter.scala 68:24]
  reg [3:0] image_1144; // @[Filter.scala 68:24]
  reg [3:0] image_1145; // @[Filter.scala 68:24]
  reg [3:0] image_1146; // @[Filter.scala 68:24]
  reg [3:0] image_1147; // @[Filter.scala 68:24]
  reg [3:0] image_1148; // @[Filter.scala 68:24]
  reg [3:0] image_1152; // @[Filter.scala 68:24]
  reg [3:0] image_1153; // @[Filter.scala 68:24]
  reg [3:0] image_1154; // @[Filter.scala 68:24]
  reg [3:0] image_1155; // @[Filter.scala 68:24]
  reg [3:0] image_1156; // @[Filter.scala 68:24]
  reg [3:0] image_1157; // @[Filter.scala 68:24]
  reg [3:0] image_1158; // @[Filter.scala 68:24]
  reg [3:0] image_1159; // @[Filter.scala 68:24]
  reg [3:0] image_1160; // @[Filter.scala 68:24]
  reg [3:0] image_1161; // @[Filter.scala 68:24]
  reg [3:0] image_1162; // @[Filter.scala 68:24]
  reg [3:0] image_1163; // @[Filter.scala 68:24]
  reg [3:0] image_1164; // @[Filter.scala 68:24]
  reg [3:0] image_1165; // @[Filter.scala 68:24]
  reg [3:0] image_1166; // @[Filter.scala 68:24]
  reg [3:0] image_1167; // @[Filter.scala 68:24]
  reg [3:0] image_1168; // @[Filter.scala 68:24]
  reg [3:0] image_1169; // @[Filter.scala 68:24]
  reg [3:0] image_1170; // @[Filter.scala 68:24]
  reg [3:0] image_1171; // @[Filter.scala 68:24]
  reg [3:0] image_1172; // @[Filter.scala 68:24]
  reg [3:0] image_1173; // @[Filter.scala 68:24]
  reg [3:0] image_1174; // @[Filter.scala 68:24]
  reg [3:0] image_1175; // @[Filter.scala 68:24]
  reg [3:0] image_1176; // @[Filter.scala 68:24]
  reg [3:0] image_1177; // @[Filter.scala 68:24]
  reg [3:0] image_1178; // @[Filter.scala 68:24]
  reg [3:0] image_1179; // @[Filter.scala 68:24]
  reg [3:0] image_1180; // @[Filter.scala 68:24]
  reg [3:0] image_1181; // @[Filter.scala 68:24]
  reg [3:0] image_1182; // @[Filter.scala 68:24]
  reg [3:0] image_1183; // @[Filter.scala 68:24]
  reg [3:0] image_1184; // @[Filter.scala 68:24]
  reg [3:0] image_1185; // @[Filter.scala 68:24]
  reg [3:0] image_1186; // @[Filter.scala 68:24]
  reg [3:0] image_1187; // @[Filter.scala 68:24]
  reg [3:0] image_1188; // @[Filter.scala 68:24]
  reg [3:0] image_1189; // @[Filter.scala 68:24]
  reg [3:0] image_1190; // @[Filter.scala 68:24]
  reg [3:0] image_1191; // @[Filter.scala 68:24]
  reg [3:0] image_1192; // @[Filter.scala 68:24]
  reg [3:0] image_1193; // @[Filter.scala 68:24]
  reg [3:0] image_1194; // @[Filter.scala 68:24]
  reg [3:0] image_1195; // @[Filter.scala 68:24]
  reg [3:0] image_1196; // @[Filter.scala 68:24]
  reg [3:0] image_1197; // @[Filter.scala 68:24]
  reg [3:0] image_1198; // @[Filter.scala 68:24]
  reg [3:0] image_1199; // @[Filter.scala 68:24]
  reg [3:0] image_1200; // @[Filter.scala 68:24]
  reg [3:0] image_1201; // @[Filter.scala 68:24]
  reg [3:0] image_1202; // @[Filter.scala 68:24]
  reg [3:0] image_1203; // @[Filter.scala 68:24]
  reg [3:0] image_1204; // @[Filter.scala 68:24]
  reg [3:0] image_1205; // @[Filter.scala 68:24]
  reg [3:0] image_1206; // @[Filter.scala 68:24]
  reg [3:0] image_1207; // @[Filter.scala 68:24]
  reg [3:0] image_1208; // @[Filter.scala 68:24]
  reg [3:0] image_1216; // @[Filter.scala 68:24]
  reg [3:0] image_1217; // @[Filter.scala 68:24]
  reg [3:0] image_1218; // @[Filter.scala 68:24]
  reg [3:0] image_1219; // @[Filter.scala 68:24]
  reg [3:0] image_1220; // @[Filter.scala 68:24]
  reg [3:0] image_1221; // @[Filter.scala 68:24]
  reg [3:0] image_1222; // @[Filter.scala 68:24]
  reg [3:0] image_1223; // @[Filter.scala 68:24]
  reg [3:0] image_1224; // @[Filter.scala 68:24]
  reg [3:0] image_1225; // @[Filter.scala 68:24]
  reg [3:0] image_1226; // @[Filter.scala 68:24]
  reg [3:0] image_1227; // @[Filter.scala 68:24]
  reg [3:0] image_1228; // @[Filter.scala 68:24]
  reg [3:0] image_1229; // @[Filter.scala 68:24]
  reg [3:0] image_1230; // @[Filter.scala 68:24]
  reg [3:0] image_1231; // @[Filter.scala 68:24]
  reg [3:0] image_1232; // @[Filter.scala 68:24]
  reg [3:0] image_1233; // @[Filter.scala 68:24]
  reg [3:0] image_1234; // @[Filter.scala 68:24]
  reg [3:0] image_1235; // @[Filter.scala 68:24]
  reg [3:0] image_1236; // @[Filter.scala 68:24]
  reg [3:0] image_1237; // @[Filter.scala 68:24]
  reg [3:0] image_1238; // @[Filter.scala 68:24]
  reg [3:0] image_1239; // @[Filter.scala 68:24]
  reg [3:0] image_1240; // @[Filter.scala 68:24]
  reg [3:0] image_1241; // @[Filter.scala 68:24]
  reg [3:0] image_1242; // @[Filter.scala 68:24]
  reg [3:0] image_1243; // @[Filter.scala 68:24]
  reg [3:0] image_1244; // @[Filter.scala 68:24]
  reg [3:0] image_1245; // @[Filter.scala 68:24]
  reg [3:0] image_1246; // @[Filter.scala 68:24]
  reg [3:0] image_1247; // @[Filter.scala 68:24]
  reg [3:0] image_1248; // @[Filter.scala 68:24]
  reg [3:0] image_1249; // @[Filter.scala 68:24]
  reg [3:0] image_1250; // @[Filter.scala 68:24]
  reg [3:0] image_1251; // @[Filter.scala 68:24]
  reg [3:0] image_1252; // @[Filter.scala 68:24]
  reg [3:0] image_1253; // @[Filter.scala 68:24]
  reg [3:0] image_1254; // @[Filter.scala 68:24]
  reg [3:0] image_1255; // @[Filter.scala 68:24]
  reg [3:0] image_1256; // @[Filter.scala 68:24]
  reg [3:0] image_1257; // @[Filter.scala 68:24]
  reg [3:0] image_1258; // @[Filter.scala 68:24]
  reg [3:0] image_1259; // @[Filter.scala 68:24]
  reg [3:0] image_1260; // @[Filter.scala 68:24]
  reg [3:0] image_1261; // @[Filter.scala 68:24]
  reg [3:0] image_1262; // @[Filter.scala 68:24]
  reg [3:0] image_1263; // @[Filter.scala 68:24]
  reg [3:0] image_1264; // @[Filter.scala 68:24]
  reg [3:0] image_1265; // @[Filter.scala 68:24]
  reg [3:0] image_1266; // @[Filter.scala 68:24]
  reg [3:0] image_1267; // @[Filter.scala 68:24]
  reg [3:0] image_1268; // @[Filter.scala 68:24]
  reg [3:0] image_1269; // @[Filter.scala 68:24]
  reg [3:0] image_1270; // @[Filter.scala 68:24]
  reg [3:0] image_1271; // @[Filter.scala 68:24]
  reg [3:0] image_1272; // @[Filter.scala 68:24]
  reg [3:0] image_1273; // @[Filter.scala 68:24]
  reg [3:0] image_1274; // @[Filter.scala 68:24]
  reg [3:0] image_1275; // @[Filter.scala 68:24]
  reg [3:0] image_1280; // @[Filter.scala 68:24]
  reg [3:0] image_1281; // @[Filter.scala 68:24]
  reg [3:0] image_1282; // @[Filter.scala 68:24]
  reg [3:0] image_1283; // @[Filter.scala 68:24]
  reg [3:0] image_1284; // @[Filter.scala 68:24]
  reg [3:0] image_1285; // @[Filter.scala 68:24]
  reg [3:0] image_1286; // @[Filter.scala 68:24]
  reg [3:0] image_1287; // @[Filter.scala 68:24]
  reg [3:0] image_1288; // @[Filter.scala 68:24]
  reg [3:0] image_1289; // @[Filter.scala 68:24]
  reg [3:0] image_1290; // @[Filter.scala 68:24]
  reg [3:0] image_1291; // @[Filter.scala 68:24]
  reg [3:0] image_1292; // @[Filter.scala 68:24]
  reg [3:0] image_1293; // @[Filter.scala 68:24]
  reg [3:0] image_1294; // @[Filter.scala 68:24]
  reg [3:0] image_1295; // @[Filter.scala 68:24]
  reg [3:0] image_1296; // @[Filter.scala 68:24]
  reg [3:0] image_1297; // @[Filter.scala 68:24]
  reg [3:0] image_1298; // @[Filter.scala 68:24]
  reg [3:0] image_1299; // @[Filter.scala 68:24]
  reg [3:0] image_1300; // @[Filter.scala 68:24]
  reg [3:0] image_1301; // @[Filter.scala 68:24]
  reg [3:0] image_1302; // @[Filter.scala 68:24]
  reg [3:0] image_1303; // @[Filter.scala 68:24]
  reg [3:0] image_1304; // @[Filter.scala 68:24]
  reg [3:0] image_1305; // @[Filter.scala 68:24]
  reg [3:0] image_1306; // @[Filter.scala 68:24]
  reg [3:0] image_1307; // @[Filter.scala 68:24]
  reg [3:0] image_1308; // @[Filter.scala 68:24]
  reg [3:0] image_1309; // @[Filter.scala 68:24]
  reg [3:0] image_1310; // @[Filter.scala 68:24]
  reg [3:0] image_1311; // @[Filter.scala 68:24]
  reg [3:0] image_1312; // @[Filter.scala 68:24]
  reg [3:0] image_1313; // @[Filter.scala 68:24]
  reg [3:0] image_1314; // @[Filter.scala 68:24]
  reg [3:0] image_1315; // @[Filter.scala 68:24]
  reg [3:0] image_1316; // @[Filter.scala 68:24]
  reg [3:0] image_1317; // @[Filter.scala 68:24]
  reg [3:0] image_1318; // @[Filter.scala 68:24]
  reg [3:0] image_1319; // @[Filter.scala 68:24]
  reg [3:0] image_1320; // @[Filter.scala 68:24]
  reg [3:0] image_1321; // @[Filter.scala 68:24]
  reg [3:0] image_1322; // @[Filter.scala 68:24]
  reg [3:0] image_1323; // @[Filter.scala 68:24]
  reg [3:0] image_1324; // @[Filter.scala 68:24]
  reg [3:0] image_1325; // @[Filter.scala 68:24]
  reg [3:0] image_1326; // @[Filter.scala 68:24]
  reg [3:0] image_1327; // @[Filter.scala 68:24]
  reg [3:0] image_1328; // @[Filter.scala 68:24]
  reg [3:0] image_1329; // @[Filter.scala 68:24]
  reg [3:0] image_1330; // @[Filter.scala 68:24]
  reg [3:0] image_1331; // @[Filter.scala 68:24]
  reg [3:0] image_1332; // @[Filter.scala 68:24]
  reg [3:0] image_1333; // @[Filter.scala 68:24]
  reg [3:0] image_1334; // @[Filter.scala 68:24]
  reg [3:0] image_1335; // @[Filter.scala 68:24]
  reg [3:0] image_1336; // @[Filter.scala 68:24]
  reg [3:0] image_1337; // @[Filter.scala 68:24]
  reg [3:0] image_1338; // @[Filter.scala 68:24]
  reg [3:0] image_1339; // @[Filter.scala 68:24]
  reg [3:0] image_1340; // @[Filter.scala 68:24]
  reg [3:0] image_1341; // @[Filter.scala 68:24]
  reg [3:0] image_1344; // @[Filter.scala 68:24]
  reg [3:0] image_1345; // @[Filter.scala 68:24]
  reg [3:0] image_1346; // @[Filter.scala 68:24]
  reg [3:0] image_1347; // @[Filter.scala 68:24]
  reg [3:0] image_1348; // @[Filter.scala 68:24]
  reg [3:0] image_1349; // @[Filter.scala 68:24]
  reg [3:0] image_1350; // @[Filter.scala 68:24]
  reg [3:0] image_1351; // @[Filter.scala 68:24]
  reg [3:0] image_1352; // @[Filter.scala 68:24]
  reg [3:0] image_1353; // @[Filter.scala 68:24]
  reg [3:0] image_1354; // @[Filter.scala 68:24]
  reg [3:0] image_1355; // @[Filter.scala 68:24]
  reg [3:0] image_1356; // @[Filter.scala 68:24]
  reg [3:0] image_1357; // @[Filter.scala 68:24]
  reg [3:0] image_1358; // @[Filter.scala 68:24]
  reg [3:0] image_1359; // @[Filter.scala 68:24]
  reg [3:0] image_1360; // @[Filter.scala 68:24]
  reg [3:0] image_1361; // @[Filter.scala 68:24]
  reg [3:0] image_1362; // @[Filter.scala 68:24]
  reg [3:0] image_1363; // @[Filter.scala 68:24]
  reg [3:0] image_1364; // @[Filter.scala 68:24]
  reg [3:0] image_1365; // @[Filter.scala 68:24]
  reg [3:0] image_1366; // @[Filter.scala 68:24]
  reg [3:0] image_1367; // @[Filter.scala 68:24]
  reg [3:0] image_1368; // @[Filter.scala 68:24]
  reg [3:0] image_1369; // @[Filter.scala 68:24]
  reg [3:0] image_1370; // @[Filter.scala 68:24]
  reg [3:0] image_1371; // @[Filter.scala 68:24]
  reg [3:0] image_1372; // @[Filter.scala 68:24]
  reg [3:0] image_1373; // @[Filter.scala 68:24]
  reg [3:0] image_1374; // @[Filter.scala 68:24]
  reg [3:0] image_1375; // @[Filter.scala 68:24]
  reg [3:0] image_1376; // @[Filter.scala 68:24]
  reg [3:0] image_1377; // @[Filter.scala 68:24]
  reg [3:0] image_1378; // @[Filter.scala 68:24]
  reg [3:0] image_1379; // @[Filter.scala 68:24]
  reg [3:0] image_1380; // @[Filter.scala 68:24]
  reg [3:0] image_1381; // @[Filter.scala 68:24]
  reg [3:0] image_1382; // @[Filter.scala 68:24]
  reg [3:0] image_1383; // @[Filter.scala 68:24]
  reg [3:0] image_1384; // @[Filter.scala 68:24]
  reg [3:0] image_1385; // @[Filter.scala 68:24]
  reg [3:0] image_1386; // @[Filter.scala 68:24]
  reg [3:0] image_1387; // @[Filter.scala 68:24]
  reg [3:0] image_1388; // @[Filter.scala 68:24]
  reg [3:0] image_1389; // @[Filter.scala 68:24]
  reg [3:0] image_1390; // @[Filter.scala 68:24]
  reg [3:0] image_1391; // @[Filter.scala 68:24]
  reg [3:0] image_1392; // @[Filter.scala 68:24]
  reg [3:0] image_1393; // @[Filter.scala 68:24]
  reg [3:0] image_1394; // @[Filter.scala 68:24]
  reg [3:0] image_1395; // @[Filter.scala 68:24]
  reg [3:0] image_1396; // @[Filter.scala 68:24]
  reg [3:0] image_1397; // @[Filter.scala 68:24]
  reg [3:0] image_1398; // @[Filter.scala 68:24]
  reg [3:0] image_1399; // @[Filter.scala 68:24]
  reg [3:0] image_1400; // @[Filter.scala 68:24]
  reg [3:0] image_1401; // @[Filter.scala 68:24]
  reg [3:0] image_1402; // @[Filter.scala 68:24]
  reg [3:0] image_1403; // @[Filter.scala 68:24]
  reg [3:0] image_1404; // @[Filter.scala 68:24]
  reg [3:0] image_1405; // @[Filter.scala 68:24]
  reg [3:0] image_1408; // @[Filter.scala 68:24]
  reg [3:0] image_1409; // @[Filter.scala 68:24]
  reg [3:0] image_1410; // @[Filter.scala 68:24]
  reg [3:0] image_1411; // @[Filter.scala 68:24]
  reg [3:0] image_1412; // @[Filter.scala 68:24]
  reg [3:0] image_1413; // @[Filter.scala 68:24]
  reg [3:0] image_1414; // @[Filter.scala 68:24]
  reg [3:0] image_1415; // @[Filter.scala 68:24]
  reg [3:0] image_1416; // @[Filter.scala 68:24]
  reg [3:0] image_1417; // @[Filter.scala 68:24]
  reg [3:0] image_1418; // @[Filter.scala 68:24]
  reg [3:0] image_1419; // @[Filter.scala 68:24]
  reg [3:0] image_1420; // @[Filter.scala 68:24]
  reg [3:0] image_1421; // @[Filter.scala 68:24]
  reg [3:0] image_1422; // @[Filter.scala 68:24]
  reg [3:0] image_1423; // @[Filter.scala 68:24]
  reg [3:0] image_1424; // @[Filter.scala 68:24]
  reg [3:0] image_1425; // @[Filter.scala 68:24]
  reg [3:0] image_1426; // @[Filter.scala 68:24]
  reg [3:0] image_1427; // @[Filter.scala 68:24]
  reg [3:0] image_1428; // @[Filter.scala 68:24]
  reg [3:0] image_1429; // @[Filter.scala 68:24]
  reg [3:0] image_1430; // @[Filter.scala 68:24]
  reg [3:0] image_1431; // @[Filter.scala 68:24]
  reg [3:0] image_1432; // @[Filter.scala 68:24]
  reg [3:0] image_1433; // @[Filter.scala 68:24]
  reg [3:0] image_1434; // @[Filter.scala 68:24]
  reg [3:0] image_1435; // @[Filter.scala 68:24]
  reg [3:0] image_1436; // @[Filter.scala 68:24]
  reg [3:0] image_1437; // @[Filter.scala 68:24]
  reg [3:0] image_1438; // @[Filter.scala 68:24]
  reg [3:0] image_1439; // @[Filter.scala 68:24]
  reg [3:0] image_1440; // @[Filter.scala 68:24]
  reg [3:0] image_1441; // @[Filter.scala 68:24]
  reg [3:0] image_1442; // @[Filter.scala 68:24]
  reg [3:0] image_1443; // @[Filter.scala 68:24]
  reg [3:0] image_1444; // @[Filter.scala 68:24]
  reg [3:0] image_1445; // @[Filter.scala 68:24]
  reg [3:0] image_1446; // @[Filter.scala 68:24]
  reg [3:0] image_1447; // @[Filter.scala 68:24]
  reg [3:0] image_1448; // @[Filter.scala 68:24]
  reg [3:0] image_1449; // @[Filter.scala 68:24]
  reg [3:0] image_1450; // @[Filter.scala 68:24]
  reg [3:0] image_1451; // @[Filter.scala 68:24]
  reg [3:0] image_1452; // @[Filter.scala 68:24]
  reg [3:0] image_1453; // @[Filter.scala 68:24]
  reg [3:0] image_1454; // @[Filter.scala 68:24]
  reg [3:0] image_1455; // @[Filter.scala 68:24]
  reg [3:0] image_1456; // @[Filter.scala 68:24]
  reg [3:0] image_1457; // @[Filter.scala 68:24]
  reg [3:0] image_1458; // @[Filter.scala 68:24]
  reg [3:0] image_1459; // @[Filter.scala 68:24]
  reg [3:0] image_1460; // @[Filter.scala 68:24]
  reg [3:0] image_1461; // @[Filter.scala 68:24]
  reg [3:0] image_1462; // @[Filter.scala 68:24]
  reg [3:0] image_1463; // @[Filter.scala 68:24]
  reg [3:0] image_1464; // @[Filter.scala 68:24]
  reg [3:0] image_1465; // @[Filter.scala 68:24]
  reg [3:0] image_1466; // @[Filter.scala 68:24]
  reg [3:0] image_1467; // @[Filter.scala 68:24]
  reg [3:0] image_1468; // @[Filter.scala 68:24]
  reg [3:0] image_1469; // @[Filter.scala 68:24]
  reg [3:0] image_1472; // @[Filter.scala 68:24]
  reg [3:0] image_1473; // @[Filter.scala 68:24]
  reg [3:0] image_1474; // @[Filter.scala 68:24]
  reg [3:0] image_1475; // @[Filter.scala 68:24]
  reg [3:0] image_1476; // @[Filter.scala 68:24]
  reg [3:0] image_1477; // @[Filter.scala 68:24]
  reg [3:0] image_1478; // @[Filter.scala 68:24]
  reg [3:0] image_1479; // @[Filter.scala 68:24]
  reg [3:0] image_1480; // @[Filter.scala 68:24]
  reg [3:0] image_1481; // @[Filter.scala 68:24]
  reg [3:0] image_1482; // @[Filter.scala 68:24]
  reg [3:0] image_1483; // @[Filter.scala 68:24]
  reg [3:0] image_1484; // @[Filter.scala 68:24]
  reg [3:0] image_1485; // @[Filter.scala 68:24]
  reg [3:0] image_1486; // @[Filter.scala 68:24]
  reg [3:0] image_1487; // @[Filter.scala 68:24]
  reg [3:0] image_1488; // @[Filter.scala 68:24]
  reg [3:0] image_1489; // @[Filter.scala 68:24]
  reg [3:0] image_1490; // @[Filter.scala 68:24]
  reg [3:0] image_1491; // @[Filter.scala 68:24]
  reg [3:0] image_1492; // @[Filter.scala 68:24]
  reg [3:0] image_1493; // @[Filter.scala 68:24]
  reg [3:0] image_1494; // @[Filter.scala 68:24]
  reg [3:0] image_1495; // @[Filter.scala 68:24]
  reg [3:0] image_1496; // @[Filter.scala 68:24]
  reg [3:0] image_1497; // @[Filter.scala 68:24]
  reg [3:0] image_1498; // @[Filter.scala 68:24]
  reg [3:0] image_1499; // @[Filter.scala 68:24]
  reg [3:0] image_1500; // @[Filter.scala 68:24]
  reg [3:0] image_1501; // @[Filter.scala 68:24]
  reg [3:0] image_1502; // @[Filter.scala 68:24]
  reg [3:0] image_1503; // @[Filter.scala 68:24]
  reg [3:0] image_1504; // @[Filter.scala 68:24]
  reg [3:0] image_1505; // @[Filter.scala 68:24]
  reg [3:0] image_1506; // @[Filter.scala 68:24]
  reg [3:0] image_1507; // @[Filter.scala 68:24]
  reg [3:0] image_1508; // @[Filter.scala 68:24]
  reg [3:0] image_1509; // @[Filter.scala 68:24]
  reg [3:0] image_1510; // @[Filter.scala 68:24]
  reg [3:0] image_1511; // @[Filter.scala 68:24]
  reg [3:0] image_1512; // @[Filter.scala 68:24]
  reg [3:0] image_1513; // @[Filter.scala 68:24]
  reg [3:0] image_1514; // @[Filter.scala 68:24]
  reg [3:0] image_1515; // @[Filter.scala 68:24]
  reg [3:0] image_1516; // @[Filter.scala 68:24]
  reg [3:0] image_1517; // @[Filter.scala 68:24]
  reg [3:0] image_1518; // @[Filter.scala 68:24]
  reg [3:0] image_1519; // @[Filter.scala 68:24]
  reg [3:0] image_1520; // @[Filter.scala 68:24]
  reg [3:0] image_1521; // @[Filter.scala 68:24]
  reg [3:0] image_1522; // @[Filter.scala 68:24]
  reg [3:0] image_1523; // @[Filter.scala 68:24]
  reg [3:0] image_1524; // @[Filter.scala 68:24]
  reg [3:0] image_1525; // @[Filter.scala 68:24]
  reg [3:0] image_1526; // @[Filter.scala 68:24]
  reg [3:0] image_1527; // @[Filter.scala 68:24]
  reg [3:0] image_1528; // @[Filter.scala 68:24]
  reg [3:0] image_1529; // @[Filter.scala 68:24]
  reg [3:0] image_1530; // @[Filter.scala 68:24]
  reg [3:0] image_1531; // @[Filter.scala 68:24]
  reg [3:0] image_1532; // @[Filter.scala 68:24]
  reg [3:0] image_1533; // @[Filter.scala 68:24]
  reg [3:0] image_1536; // @[Filter.scala 68:24]
  reg [3:0] image_1537; // @[Filter.scala 68:24]
  reg [3:0] image_1538; // @[Filter.scala 68:24]
  reg [3:0] image_1539; // @[Filter.scala 68:24]
  reg [3:0] image_1540; // @[Filter.scala 68:24]
  reg [3:0] image_1541; // @[Filter.scala 68:24]
  reg [3:0] image_1542; // @[Filter.scala 68:24]
  reg [3:0] image_1543; // @[Filter.scala 68:24]
  reg [3:0] image_1544; // @[Filter.scala 68:24]
  reg [3:0] image_1545; // @[Filter.scala 68:24]
  reg [3:0] image_1546; // @[Filter.scala 68:24]
  reg [3:0] image_1547; // @[Filter.scala 68:24]
  reg [3:0] image_1548; // @[Filter.scala 68:24]
  reg [3:0] image_1549; // @[Filter.scala 68:24]
  reg [3:0] image_1550; // @[Filter.scala 68:24]
  reg [3:0] image_1551; // @[Filter.scala 68:24]
  reg [3:0] image_1552; // @[Filter.scala 68:24]
  reg [3:0] image_1553; // @[Filter.scala 68:24]
  reg [3:0] image_1554; // @[Filter.scala 68:24]
  reg [3:0] image_1555; // @[Filter.scala 68:24]
  reg [3:0] image_1556; // @[Filter.scala 68:24]
  reg [3:0] image_1557; // @[Filter.scala 68:24]
  reg [3:0] image_1558; // @[Filter.scala 68:24]
  reg [3:0] image_1559; // @[Filter.scala 68:24]
  reg [3:0] image_1560; // @[Filter.scala 68:24]
  reg [3:0] image_1561; // @[Filter.scala 68:24]
  reg [3:0] image_1562; // @[Filter.scala 68:24]
  reg [3:0] image_1563; // @[Filter.scala 68:24]
  reg [3:0] image_1564; // @[Filter.scala 68:24]
  reg [3:0] image_1565; // @[Filter.scala 68:24]
  reg [3:0] image_1566; // @[Filter.scala 68:24]
  reg [3:0] image_1567; // @[Filter.scala 68:24]
  reg [3:0] image_1568; // @[Filter.scala 68:24]
  reg [3:0] image_1569; // @[Filter.scala 68:24]
  reg [3:0] image_1570; // @[Filter.scala 68:24]
  reg [3:0] image_1571; // @[Filter.scala 68:24]
  reg [3:0] image_1572; // @[Filter.scala 68:24]
  reg [3:0] image_1573; // @[Filter.scala 68:24]
  reg [3:0] image_1574; // @[Filter.scala 68:24]
  reg [3:0] image_1575; // @[Filter.scala 68:24]
  reg [3:0] image_1576; // @[Filter.scala 68:24]
  reg [3:0] image_1577; // @[Filter.scala 68:24]
  reg [3:0] image_1578; // @[Filter.scala 68:24]
  reg [3:0] image_1579; // @[Filter.scala 68:24]
  reg [3:0] image_1580; // @[Filter.scala 68:24]
  reg [3:0] image_1581; // @[Filter.scala 68:24]
  reg [3:0] image_1582; // @[Filter.scala 68:24]
  reg [3:0] image_1583; // @[Filter.scala 68:24]
  reg [3:0] image_1584; // @[Filter.scala 68:24]
  reg [3:0] image_1585; // @[Filter.scala 68:24]
  reg [3:0] image_1586; // @[Filter.scala 68:24]
  reg [3:0] image_1587; // @[Filter.scala 68:24]
  reg [3:0] image_1588; // @[Filter.scala 68:24]
  reg [3:0] image_1589; // @[Filter.scala 68:24]
  reg [3:0] image_1590; // @[Filter.scala 68:24]
  reg [3:0] image_1591; // @[Filter.scala 68:24]
  reg [3:0] image_1592; // @[Filter.scala 68:24]
  reg [3:0] image_1593; // @[Filter.scala 68:24]
  reg [3:0] image_1594; // @[Filter.scala 68:24]
  reg [3:0] image_1595; // @[Filter.scala 68:24]
  reg [3:0] image_1596; // @[Filter.scala 68:24]
  reg [3:0] image_1597; // @[Filter.scala 68:24]
  reg [3:0] image_1600; // @[Filter.scala 68:24]
  reg [3:0] image_1601; // @[Filter.scala 68:24]
  reg [3:0] image_1602; // @[Filter.scala 68:24]
  reg [3:0] image_1603; // @[Filter.scala 68:24]
  reg [3:0] image_1604; // @[Filter.scala 68:24]
  reg [3:0] image_1605; // @[Filter.scala 68:24]
  reg [3:0] image_1606; // @[Filter.scala 68:24]
  reg [3:0] image_1607; // @[Filter.scala 68:24]
  reg [3:0] image_1608; // @[Filter.scala 68:24]
  reg [3:0] image_1609; // @[Filter.scala 68:24]
  reg [3:0] image_1610; // @[Filter.scala 68:24]
  reg [3:0] image_1611; // @[Filter.scala 68:24]
  reg [3:0] image_1612; // @[Filter.scala 68:24]
  reg [3:0] image_1613; // @[Filter.scala 68:24]
  reg [3:0] image_1614; // @[Filter.scala 68:24]
  reg [3:0] image_1615; // @[Filter.scala 68:24]
  reg [3:0] image_1616; // @[Filter.scala 68:24]
  reg [3:0] image_1617; // @[Filter.scala 68:24]
  reg [3:0] image_1618; // @[Filter.scala 68:24]
  reg [3:0] image_1619; // @[Filter.scala 68:24]
  reg [3:0] image_1620; // @[Filter.scala 68:24]
  reg [3:0] image_1621; // @[Filter.scala 68:24]
  reg [3:0] image_1622; // @[Filter.scala 68:24]
  reg [3:0] image_1623; // @[Filter.scala 68:24]
  reg [3:0] image_1624; // @[Filter.scala 68:24]
  reg [3:0] image_1625; // @[Filter.scala 68:24]
  reg [3:0] image_1626; // @[Filter.scala 68:24]
  reg [3:0] image_1627; // @[Filter.scala 68:24]
  reg [3:0] image_1628; // @[Filter.scala 68:24]
  reg [3:0] image_1629; // @[Filter.scala 68:24]
  reg [3:0] image_1630; // @[Filter.scala 68:24]
  reg [3:0] image_1631; // @[Filter.scala 68:24]
  reg [3:0] image_1632; // @[Filter.scala 68:24]
  reg [3:0] image_1633; // @[Filter.scala 68:24]
  reg [3:0] image_1634; // @[Filter.scala 68:24]
  reg [3:0] image_1635; // @[Filter.scala 68:24]
  reg [3:0] image_1636; // @[Filter.scala 68:24]
  reg [3:0] image_1637; // @[Filter.scala 68:24]
  reg [3:0] image_1638; // @[Filter.scala 68:24]
  reg [3:0] image_1639; // @[Filter.scala 68:24]
  reg [3:0] image_1640; // @[Filter.scala 68:24]
  reg [3:0] image_1641; // @[Filter.scala 68:24]
  reg [3:0] image_1642; // @[Filter.scala 68:24]
  reg [3:0] image_1643; // @[Filter.scala 68:24]
  reg [3:0] image_1644; // @[Filter.scala 68:24]
  reg [3:0] image_1645; // @[Filter.scala 68:24]
  reg [3:0] image_1646; // @[Filter.scala 68:24]
  reg [3:0] image_1647; // @[Filter.scala 68:24]
  reg [3:0] image_1648; // @[Filter.scala 68:24]
  reg [3:0] image_1649; // @[Filter.scala 68:24]
  reg [3:0] image_1650; // @[Filter.scala 68:24]
  reg [3:0] image_1651; // @[Filter.scala 68:24]
  reg [3:0] image_1652; // @[Filter.scala 68:24]
  reg [3:0] image_1653; // @[Filter.scala 68:24]
  reg [3:0] image_1654; // @[Filter.scala 68:24]
  reg [3:0] image_1655; // @[Filter.scala 68:24]
  reg [3:0] image_1656; // @[Filter.scala 68:24]
  reg [3:0] image_1657; // @[Filter.scala 68:24]
  reg [3:0] image_1658; // @[Filter.scala 68:24]
  reg [3:0] image_1659; // @[Filter.scala 68:24]
  reg [3:0] image_1660; // @[Filter.scala 68:24]
  reg [3:0] image_1664; // @[Filter.scala 68:24]
  reg [3:0] image_1665; // @[Filter.scala 68:24]
  reg [3:0] image_1666; // @[Filter.scala 68:24]
  reg [3:0] image_1667; // @[Filter.scala 68:24]
  reg [3:0] image_1668; // @[Filter.scala 68:24]
  reg [3:0] image_1669; // @[Filter.scala 68:24]
  reg [3:0] image_1670; // @[Filter.scala 68:24]
  reg [3:0] image_1671; // @[Filter.scala 68:24]
  reg [3:0] image_1672; // @[Filter.scala 68:24]
  reg [3:0] image_1673; // @[Filter.scala 68:24]
  reg [3:0] image_1674; // @[Filter.scala 68:24]
  reg [3:0] image_1675; // @[Filter.scala 68:24]
  reg [3:0] image_1676; // @[Filter.scala 68:24]
  reg [3:0] image_1677; // @[Filter.scala 68:24]
  reg [3:0] image_1678; // @[Filter.scala 68:24]
  reg [3:0] image_1679; // @[Filter.scala 68:24]
  reg [3:0] image_1680; // @[Filter.scala 68:24]
  reg [3:0] image_1681; // @[Filter.scala 68:24]
  reg [3:0] image_1682; // @[Filter.scala 68:24]
  reg [3:0] image_1683; // @[Filter.scala 68:24]
  reg [3:0] image_1684; // @[Filter.scala 68:24]
  reg [3:0] image_1685; // @[Filter.scala 68:24]
  reg [3:0] image_1686; // @[Filter.scala 68:24]
  reg [3:0] image_1687; // @[Filter.scala 68:24]
  reg [3:0] image_1688; // @[Filter.scala 68:24]
  reg [3:0] image_1689; // @[Filter.scala 68:24]
  reg [3:0] image_1690; // @[Filter.scala 68:24]
  reg [3:0] image_1691; // @[Filter.scala 68:24]
  reg [3:0] image_1692; // @[Filter.scala 68:24]
  reg [3:0] image_1693; // @[Filter.scala 68:24]
  reg [3:0] image_1694; // @[Filter.scala 68:24]
  reg [3:0] image_1695; // @[Filter.scala 68:24]
  reg [3:0] image_1696; // @[Filter.scala 68:24]
  reg [3:0] image_1697; // @[Filter.scala 68:24]
  reg [3:0] image_1698; // @[Filter.scala 68:24]
  reg [3:0] image_1699; // @[Filter.scala 68:24]
  reg [3:0] image_1700; // @[Filter.scala 68:24]
  reg [3:0] image_1701; // @[Filter.scala 68:24]
  reg [3:0] image_1702; // @[Filter.scala 68:24]
  reg [3:0] image_1703; // @[Filter.scala 68:24]
  reg [3:0] image_1704; // @[Filter.scala 68:24]
  reg [3:0] image_1705; // @[Filter.scala 68:24]
  reg [3:0] image_1706; // @[Filter.scala 68:24]
  reg [3:0] image_1707; // @[Filter.scala 68:24]
  reg [3:0] image_1708; // @[Filter.scala 68:24]
  reg [3:0] image_1709; // @[Filter.scala 68:24]
  reg [3:0] image_1710; // @[Filter.scala 68:24]
  reg [3:0] image_1711; // @[Filter.scala 68:24]
  reg [3:0] image_1712; // @[Filter.scala 68:24]
  reg [3:0] image_1713; // @[Filter.scala 68:24]
  reg [3:0] image_1714; // @[Filter.scala 68:24]
  reg [3:0] image_1715; // @[Filter.scala 68:24]
  reg [3:0] image_1716; // @[Filter.scala 68:24]
  reg [3:0] image_1717; // @[Filter.scala 68:24]
  reg [3:0] image_1718; // @[Filter.scala 68:24]
  reg [3:0] image_1719; // @[Filter.scala 68:24]
  reg [3:0] image_1720; // @[Filter.scala 68:24]
  reg [3:0] image_1721; // @[Filter.scala 68:24]
  reg [3:0] image_1722; // @[Filter.scala 68:24]
  reg [3:0] image_1723; // @[Filter.scala 68:24]
  reg [3:0] image_1728; // @[Filter.scala 68:24]
  reg [3:0] image_1729; // @[Filter.scala 68:24]
  reg [3:0] image_1730; // @[Filter.scala 68:24]
  reg [3:0] image_1731; // @[Filter.scala 68:24]
  reg [3:0] image_1732; // @[Filter.scala 68:24]
  reg [3:0] image_1733; // @[Filter.scala 68:24]
  reg [3:0] image_1734; // @[Filter.scala 68:24]
  reg [3:0] image_1735; // @[Filter.scala 68:24]
  reg [3:0] image_1736; // @[Filter.scala 68:24]
  reg [3:0] image_1737; // @[Filter.scala 68:24]
  reg [3:0] image_1738; // @[Filter.scala 68:24]
  reg [3:0] image_1739; // @[Filter.scala 68:24]
  reg [3:0] image_1740; // @[Filter.scala 68:24]
  reg [3:0] image_1741; // @[Filter.scala 68:24]
  reg [3:0] image_1742; // @[Filter.scala 68:24]
  reg [3:0] image_1743; // @[Filter.scala 68:24]
  reg [3:0] image_1744; // @[Filter.scala 68:24]
  reg [3:0] image_1745; // @[Filter.scala 68:24]
  reg [3:0] image_1746; // @[Filter.scala 68:24]
  reg [3:0] image_1747; // @[Filter.scala 68:24]
  reg [3:0] image_1748; // @[Filter.scala 68:24]
  reg [3:0] image_1749; // @[Filter.scala 68:24]
  reg [3:0] image_1750; // @[Filter.scala 68:24]
  reg [3:0] image_1751; // @[Filter.scala 68:24]
  reg [3:0] image_1752; // @[Filter.scala 68:24]
  reg [3:0] image_1753; // @[Filter.scala 68:24]
  reg [3:0] image_1754; // @[Filter.scala 68:24]
  reg [3:0] image_1755; // @[Filter.scala 68:24]
  reg [3:0] image_1756; // @[Filter.scala 68:24]
  reg [3:0] image_1757; // @[Filter.scala 68:24]
  reg [3:0] image_1758; // @[Filter.scala 68:24]
  reg [3:0] image_1759; // @[Filter.scala 68:24]
  reg [3:0] image_1760; // @[Filter.scala 68:24]
  reg [3:0] image_1761; // @[Filter.scala 68:24]
  reg [3:0] image_1762; // @[Filter.scala 68:24]
  reg [3:0] image_1763; // @[Filter.scala 68:24]
  reg [3:0] image_1764; // @[Filter.scala 68:24]
  reg [3:0] image_1765; // @[Filter.scala 68:24]
  reg [3:0] image_1766; // @[Filter.scala 68:24]
  reg [3:0] image_1767; // @[Filter.scala 68:24]
  reg [3:0] image_1768; // @[Filter.scala 68:24]
  reg [3:0] image_1769; // @[Filter.scala 68:24]
  reg [3:0] image_1770; // @[Filter.scala 68:24]
  reg [3:0] image_1771; // @[Filter.scala 68:24]
  reg [3:0] image_1772; // @[Filter.scala 68:24]
  reg [3:0] image_1773; // @[Filter.scala 68:24]
  reg [3:0] image_1774; // @[Filter.scala 68:24]
  reg [3:0] image_1775; // @[Filter.scala 68:24]
  reg [3:0] image_1776; // @[Filter.scala 68:24]
  reg [3:0] image_1777; // @[Filter.scala 68:24]
  reg [3:0] image_1778; // @[Filter.scala 68:24]
  reg [3:0] image_1779; // @[Filter.scala 68:24]
  reg [3:0] image_1780; // @[Filter.scala 68:24]
  reg [3:0] image_1781; // @[Filter.scala 68:24]
  reg [3:0] image_1782; // @[Filter.scala 68:24]
  reg [3:0] image_1783; // @[Filter.scala 68:24]
  reg [3:0] image_1784; // @[Filter.scala 68:24]
  reg [3:0] image_1785; // @[Filter.scala 68:24]
  reg [3:0] image_1786; // @[Filter.scala 68:24]
  reg [3:0] image_1793; // @[Filter.scala 68:24]
  reg [3:0] image_1794; // @[Filter.scala 68:24]
  reg [3:0] image_1795; // @[Filter.scala 68:24]
  reg [3:0] image_1796; // @[Filter.scala 68:24]
  reg [3:0] image_1797; // @[Filter.scala 68:24]
  reg [3:0] image_1798; // @[Filter.scala 68:24]
  reg [3:0] image_1799; // @[Filter.scala 68:24]
  reg [3:0] image_1800; // @[Filter.scala 68:24]
  reg [3:0] image_1801; // @[Filter.scala 68:24]
  reg [3:0] image_1802; // @[Filter.scala 68:24]
  reg [3:0] image_1803; // @[Filter.scala 68:24]
  reg [3:0] image_1804; // @[Filter.scala 68:24]
  reg [3:0] image_1805; // @[Filter.scala 68:24]
  reg [3:0] image_1806; // @[Filter.scala 68:24]
  reg [3:0] image_1807; // @[Filter.scala 68:24]
  reg [3:0] image_1808; // @[Filter.scala 68:24]
  reg [3:0] image_1809; // @[Filter.scala 68:24]
  reg [3:0] image_1810; // @[Filter.scala 68:24]
  reg [3:0] image_1811; // @[Filter.scala 68:24]
  reg [3:0] image_1812; // @[Filter.scala 68:24]
  reg [3:0] image_1813; // @[Filter.scala 68:24]
  reg [3:0] image_1814; // @[Filter.scala 68:24]
  reg [3:0] image_1815; // @[Filter.scala 68:24]
  reg [3:0] image_1816; // @[Filter.scala 68:24]
  reg [3:0] image_1817; // @[Filter.scala 68:24]
  reg [3:0] image_1818; // @[Filter.scala 68:24]
  reg [3:0] image_1819; // @[Filter.scala 68:24]
  reg [3:0] image_1820; // @[Filter.scala 68:24]
  reg [3:0] image_1821; // @[Filter.scala 68:24]
  reg [3:0] image_1822; // @[Filter.scala 68:24]
  reg [3:0] image_1823; // @[Filter.scala 68:24]
  reg [3:0] image_1824; // @[Filter.scala 68:24]
  reg [3:0] image_1825; // @[Filter.scala 68:24]
  reg [3:0] image_1826; // @[Filter.scala 68:24]
  reg [3:0] image_1827; // @[Filter.scala 68:24]
  reg [3:0] image_1828; // @[Filter.scala 68:24]
  reg [3:0] image_1829; // @[Filter.scala 68:24]
  reg [3:0] image_1830; // @[Filter.scala 68:24]
  reg [3:0] image_1831; // @[Filter.scala 68:24]
  reg [3:0] image_1832; // @[Filter.scala 68:24]
  reg [3:0] image_1833; // @[Filter.scala 68:24]
  reg [3:0] image_1834; // @[Filter.scala 68:24]
  reg [3:0] image_1835; // @[Filter.scala 68:24]
  reg [3:0] image_1836; // @[Filter.scala 68:24]
  reg [3:0] image_1837; // @[Filter.scala 68:24]
  reg [3:0] image_1838; // @[Filter.scala 68:24]
  reg [3:0] image_1839; // @[Filter.scala 68:24]
  reg [3:0] image_1840; // @[Filter.scala 68:24]
  reg [3:0] image_1841; // @[Filter.scala 68:24]
  reg [3:0] image_1842; // @[Filter.scala 68:24]
  reg [3:0] image_1843; // @[Filter.scala 68:24]
  reg [3:0] image_1844; // @[Filter.scala 68:24]
  reg [3:0] image_1845; // @[Filter.scala 68:24]
  reg [3:0] image_1846; // @[Filter.scala 68:24]
  reg [3:0] image_1847; // @[Filter.scala 68:24]
  reg [3:0] image_1848; // @[Filter.scala 68:24]
  reg [3:0] image_1849; // @[Filter.scala 68:24]
  reg [3:0] image_1857; // @[Filter.scala 68:24]
  reg [3:0] image_1858; // @[Filter.scala 68:24]
  reg [3:0] image_1859; // @[Filter.scala 68:24]
  reg [3:0] image_1860; // @[Filter.scala 68:24]
  reg [3:0] image_1861; // @[Filter.scala 68:24]
  reg [3:0] image_1862; // @[Filter.scala 68:24]
  reg [3:0] image_1863; // @[Filter.scala 68:24]
  reg [3:0] image_1864; // @[Filter.scala 68:24]
  reg [3:0] image_1865; // @[Filter.scala 68:24]
  reg [3:0] image_1866; // @[Filter.scala 68:24]
  reg [3:0] image_1867; // @[Filter.scala 68:24]
  reg [3:0] image_1868; // @[Filter.scala 68:24]
  reg [3:0] image_1869; // @[Filter.scala 68:24]
  reg [3:0] image_1870; // @[Filter.scala 68:24]
  reg [3:0] image_1871; // @[Filter.scala 68:24]
  reg [3:0] image_1872; // @[Filter.scala 68:24]
  reg [3:0] image_1873; // @[Filter.scala 68:24]
  reg [3:0] image_1874; // @[Filter.scala 68:24]
  reg [3:0] image_1875; // @[Filter.scala 68:24]
  reg [3:0] image_1876; // @[Filter.scala 68:24]
  reg [3:0] image_1877; // @[Filter.scala 68:24]
  reg [3:0] image_1878; // @[Filter.scala 68:24]
  reg [3:0] image_1879; // @[Filter.scala 68:24]
  reg [3:0] image_1880; // @[Filter.scala 68:24]
  reg [3:0] image_1881; // @[Filter.scala 68:24]
  reg [3:0] image_1882; // @[Filter.scala 68:24]
  reg [3:0] image_1883; // @[Filter.scala 68:24]
  reg [3:0] image_1884; // @[Filter.scala 68:24]
  reg [3:0] image_1885; // @[Filter.scala 68:24]
  reg [3:0] image_1886; // @[Filter.scala 68:24]
  reg [3:0] image_1887; // @[Filter.scala 68:24]
  reg [3:0] image_1888; // @[Filter.scala 68:24]
  reg [3:0] image_1889; // @[Filter.scala 68:24]
  reg [3:0] image_1890; // @[Filter.scala 68:24]
  reg [3:0] image_1891; // @[Filter.scala 68:24]
  reg [3:0] image_1892; // @[Filter.scala 68:24]
  reg [3:0] image_1893; // @[Filter.scala 68:24]
  reg [3:0] image_1894; // @[Filter.scala 68:24]
  reg [3:0] image_1895; // @[Filter.scala 68:24]
  reg [3:0] image_1896; // @[Filter.scala 68:24]
  reg [3:0] image_1897; // @[Filter.scala 68:24]
  reg [3:0] image_1898; // @[Filter.scala 68:24]
  reg [3:0] image_1899; // @[Filter.scala 68:24]
  reg [3:0] image_1900; // @[Filter.scala 68:24]
  reg [3:0] image_1901; // @[Filter.scala 68:24]
  reg [3:0] image_1902; // @[Filter.scala 68:24]
  reg [3:0] image_1903; // @[Filter.scala 68:24]
  reg [3:0] image_1904; // @[Filter.scala 68:24]
  reg [3:0] image_1905; // @[Filter.scala 68:24]
  reg [3:0] image_1906; // @[Filter.scala 68:24]
  reg [3:0] image_1907; // @[Filter.scala 68:24]
  reg [3:0] image_1908; // @[Filter.scala 68:24]
  reg [3:0] image_1909; // @[Filter.scala 68:24]
  reg [3:0] image_1910; // @[Filter.scala 68:24]
  reg [3:0] image_1911; // @[Filter.scala 68:24]
  reg [3:0] image_1912; // @[Filter.scala 68:24]
  reg [3:0] image_1913; // @[Filter.scala 68:24]
  reg [3:0] image_1921; // @[Filter.scala 68:24]
  reg [3:0] image_1922; // @[Filter.scala 68:24]
  reg [3:0] image_1923; // @[Filter.scala 68:24]
  reg [3:0] image_1924; // @[Filter.scala 68:24]
  reg [3:0] image_1925; // @[Filter.scala 68:24]
  reg [3:0] image_1926; // @[Filter.scala 68:24]
  reg [3:0] image_1927; // @[Filter.scala 68:24]
  reg [3:0] image_1928; // @[Filter.scala 68:24]
  reg [3:0] image_1929; // @[Filter.scala 68:24]
  reg [3:0] image_1930; // @[Filter.scala 68:24]
  reg [3:0] image_1931; // @[Filter.scala 68:24]
  reg [3:0] image_1932; // @[Filter.scala 68:24]
  reg [3:0] image_1933; // @[Filter.scala 68:24]
  reg [3:0] image_1934; // @[Filter.scala 68:24]
  reg [3:0] image_1935; // @[Filter.scala 68:24]
  reg [3:0] image_1936; // @[Filter.scala 68:24]
  reg [3:0] image_1937; // @[Filter.scala 68:24]
  reg [3:0] image_1938; // @[Filter.scala 68:24]
  reg [3:0] image_1939; // @[Filter.scala 68:24]
  reg [3:0] image_1940; // @[Filter.scala 68:24]
  reg [3:0] image_1941; // @[Filter.scala 68:24]
  reg [3:0] image_1942; // @[Filter.scala 68:24]
  reg [3:0] image_1943; // @[Filter.scala 68:24]
  reg [3:0] image_1944; // @[Filter.scala 68:24]
  reg [3:0] image_1945; // @[Filter.scala 68:24]
  reg [3:0] image_1946; // @[Filter.scala 68:24]
  reg [3:0] image_1947; // @[Filter.scala 68:24]
  reg [3:0] image_1948; // @[Filter.scala 68:24]
  reg [3:0] image_1949; // @[Filter.scala 68:24]
  reg [3:0] image_1950; // @[Filter.scala 68:24]
  reg [3:0] image_1951; // @[Filter.scala 68:24]
  reg [3:0] image_1952; // @[Filter.scala 68:24]
  reg [3:0] image_1953; // @[Filter.scala 68:24]
  reg [3:0] image_1954; // @[Filter.scala 68:24]
  reg [3:0] image_1955; // @[Filter.scala 68:24]
  reg [3:0] image_1956; // @[Filter.scala 68:24]
  reg [3:0] image_1957; // @[Filter.scala 68:24]
  reg [3:0] image_1958; // @[Filter.scala 68:24]
  reg [3:0] image_1959; // @[Filter.scala 68:24]
  reg [3:0] image_1960; // @[Filter.scala 68:24]
  reg [3:0] image_1961; // @[Filter.scala 68:24]
  reg [3:0] image_1962; // @[Filter.scala 68:24]
  reg [3:0] image_1963; // @[Filter.scala 68:24]
  reg [3:0] image_1964; // @[Filter.scala 68:24]
  reg [3:0] image_1965; // @[Filter.scala 68:24]
  reg [3:0] image_1966; // @[Filter.scala 68:24]
  reg [3:0] image_1967; // @[Filter.scala 68:24]
  reg [3:0] image_1968; // @[Filter.scala 68:24]
  reg [3:0] image_1969; // @[Filter.scala 68:24]
  reg [3:0] image_1970; // @[Filter.scala 68:24]
  reg [3:0] image_1971; // @[Filter.scala 68:24]
  reg [3:0] image_1972; // @[Filter.scala 68:24]
  reg [3:0] image_1973; // @[Filter.scala 68:24]
  reg [3:0] image_1974; // @[Filter.scala 68:24]
  reg [3:0] image_1975; // @[Filter.scala 68:24]
  reg [3:0] image_1976; // @[Filter.scala 68:24]
  reg [3:0] image_1977; // @[Filter.scala 68:24]
  reg [3:0] image_1985; // @[Filter.scala 68:24]
  reg [3:0] image_1986; // @[Filter.scala 68:24]
  reg [3:0] image_1987; // @[Filter.scala 68:24]
  reg [3:0] image_1988; // @[Filter.scala 68:24]
  reg [3:0] image_1989; // @[Filter.scala 68:24]
  reg [3:0] image_1990; // @[Filter.scala 68:24]
  reg [3:0] image_1991; // @[Filter.scala 68:24]
  reg [3:0] image_1992; // @[Filter.scala 68:24]
  reg [3:0] image_1993; // @[Filter.scala 68:24]
  reg [3:0] image_1994; // @[Filter.scala 68:24]
  reg [3:0] image_1995; // @[Filter.scala 68:24]
  reg [3:0] image_1996; // @[Filter.scala 68:24]
  reg [3:0] image_1997; // @[Filter.scala 68:24]
  reg [3:0] image_1998; // @[Filter.scala 68:24]
  reg [3:0] image_1999; // @[Filter.scala 68:24]
  reg [3:0] image_2000; // @[Filter.scala 68:24]
  reg [3:0] image_2001; // @[Filter.scala 68:24]
  reg [3:0] image_2002; // @[Filter.scala 68:24]
  reg [3:0] image_2003; // @[Filter.scala 68:24]
  reg [3:0] image_2004; // @[Filter.scala 68:24]
  reg [3:0] image_2005; // @[Filter.scala 68:24]
  reg [3:0] image_2006; // @[Filter.scala 68:24]
  reg [3:0] image_2007; // @[Filter.scala 68:24]
  reg [3:0] image_2008; // @[Filter.scala 68:24]
  reg [3:0] image_2009; // @[Filter.scala 68:24]
  reg [3:0] image_2010; // @[Filter.scala 68:24]
  reg [3:0] image_2011; // @[Filter.scala 68:24]
  reg [3:0] image_2012; // @[Filter.scala 68:24]
  reg [3:0] image_2013; // @[Filter.scala 68:24]
  reg [3:0] image_2014; // @[Filter.scala 68:24]
  reg [3:0] image_2015; // @[Filter.scala 68:24]
  reg [3:0] image_2016; // @[Filter.scala 68:24]
  reg [3:0] image_2017; // @[Filter.scala 68:24]
  reg [3:0] image_2018; // @[Filter.scala 68:24]
  reg [3:0] image_2019; // @[Filter.scala 68:24]
  reg [3:0] image_2020; // @[Filter.scala 68:24]
  reg [3:0] image_2021; // @[Filter.scala 68:24]
  reg [3:0] image_2022; // @[Filter.scala 68:24]
  reg [3:0] image_2023; // @[Filter.scala 68:24]
  reg [3:0] image_2024; // @[Filter.scala 68:24]
  reg [3:0] image_2025; // @[Filter.scala 68:24]
  reg [3:0] image_2026; // @[Filter.scala 68:24]
  reg [3:0] image_2027; // @[Filter.scala 68:24]
  reg [3:0] image_2028; // @[Filter.scala 68:24]
  reg [3:0] image_2029; // @[Filter.scala 68:24]
  reg [3:0] image_2030; // @[Filter.scala 68:24]
  reg [3:0] image_2031; // @[Filter.scala 68:24]
  reg [3:0] image_2032; // @[Filter.scala 68:24]
  reg [3:0] image_2033; // @[Filter.scala 68:24]
  reg [3:0] image_2034; // @[Filter.scala 68:24]
  reg [3:0] image_2035; // @[Filter.scala 68:24]
  reg [3:0] image_2036; // @[Filter.scala 68:24]
  reg [3:0] image_2037; // @[Filter.scala 68:24]
  reg [3:0] image_2038; // @[Filter.scala 68:24]
  reg [3:0] image_2039; // @[Filter.scala 68:24]
  reg [3:0] image_2040; // @[Filter.scala 68:24]
  reg [3:0] image_2041; // @[Filter.scala 68:24]
  reg [3:0] image_2049; // @[Filter.scala 68:24]
  reg [3:0] image_2050; // @[Filter.scala 68:24]
  reg [3:0] image_2051; // @[Filter.scala 68:24]
  reg [3:0] image_2052; // @[Filter.scala 68:24]
  reg [3:0] image_2053; // @[Filter.scala 68:24]
  reg [3:0] image_2054; // @[Filter.scala 68:24]
  reg [3:0] image_2055; // @[Filter.scala 68:24]
  reg [3:0] image_2056; // @[Filter.scala 68:24]
  reg [3:0] image_2057; // @[Filter.scala 68:24]
  reg [3:0] image_2058; // @[Filter.scala 68:24]
  reg [3:0] image_2059; // @[Filter.scala 68:24]
  reg [3:0] image_2060; // @[Filter.scala 68:24]
  reg [3:0] image_2061; // @[Filter.scala 68:24]
  reg [3:0] image_2062; // @[Filter.scala 68:24]
  reg [3:0] image_2063; // @[Filter.scala 68:24]
  reg [3:0] image_2064; // @[Filter.scala 68:24]
  reg [3:0] image_2065; // @[Filter.scala 68:24]
  reg [3:0] image_2066; // @[Filter.scala 68:24]
  reg [3:0] image_2067; // @[Filter.scala 68:24]
  reg [3:0] image_2068; // @[Filter.scala 68:24]
  reg [3:0] image_2069; // @[Filter.scala 68:24]
  reg [3:0] image_2070; // @[Filter.scala 68:24]
  reg [3:0] image_2071; // @[Filter.scala 68:24]
  reg [3:0] image_2072; // @[Filter.scala 68:24]
  reg [3:0] image_2073; // @[Filter.scala 68:24]
  reg [3:0] image_2074; // @[Filter.scala 68:24]
  reg [3:0] image_2075; // @[Filter.scala 68:24]
  reg [3:0] image_2076; // @[Filter.scala 68:24]
  reg [3:0] image_2077; // @[Filter.scala 68:24]
  reg [3:0] image_2078; // @[Filter.scala 68:24]
  reg [3:0] image_2079; // @[Filter.scala 68:24]
  reg [3:0] image_2080; // @[Filter.scala 68:24]
  reg [3:0] image_2081; // @[Filter.scala 68:24]
  reg [3:0] image_2082; // @[Filter.scala 68:24]
  reg [3:0] image_2083; // @[Filter.scala 68:24]
  reg [3:0] image_2084; // @[Filter.scala 68:24]
  reg [3:0] image_2085; // @[Filter.scala 68:24]
  reg [3:0] image_2086; // @[Filter.scala 68:24]
  reg [3:0] image_2087; // @[Filter.scala 68:24]
  reg [3:0] image_2088; // @[Filter.scala 68:24]
  reg [3:0] image_2089; // @[Filter.scala 68:24]
  reg [3:0] image_2090; // @[Filter.scala 68:24]
  reg [3:0] image_2091; // @[Filter.scala 68:24]
  reg [3:0] image_2092; // @[Filter.scala 68:24]
  reg [3:0] image_2093; // @[Filter.scala 68:24]
  reg [3:0] image_2094; // @[Filter.scala 68:24]
  reg [3:0] image_2095; // @[Filter.scala 68:24]
  reg [3:0] image_2096; // @[Filter.scala 68:24]
  reg [3:0] image_2097; // @[Filter.scala 68:24]
  reg [3:0] image_2098; // @[Filter.scala 68:24]
  reg [3:0] image_2099; // @[Filter.scala 68:24]
  reg [3:0] image_2100; // @[Filter.scala 68:24]
  reg [3:0] image_2101; // @[Filter.scala 68:24]
  reg [3:0] image_2102; // @[Filter.scala 68:24]
  reg [3:0] image_2103; // @[Filter.scala 68:24]
  reg [3:0] image_2104; // @[Filter.scala 68:24]
  reg [3:0] image_2105; // @[Filter.scala 68:24]
  reg [3:0] image_2106; // @[Filter.scala 68:24]
  reg [3:0] image_2114; // @[Filter.scala 68:24]
  reg [3:0] image_2115; // @[Filter.scala 68:24]
  reg [3:0] image_2116; // @[Filter.scala 68:24]
  reg [3:0] image_2117; // @[Filter.scala 68:24]
  reg [3:0] image_2118; // @[Filter.scala 68:24]
  reg [3:0] image_2119; // @[Filter.scala 68:24]
  reg [3:0] image_2120; // @[Filter.scala 68:24]
  reg [3:0] image_2121; // @[Filter.scala 68:24]
  reg [3:0] image_2122; // @[Filter.scala 68:24]
  reg [3:0] image_2123; // @[Filter.scala 68:24]
  reg [3:0] image_2124; // @[Filter.scala 68:24]
  reg [3:0] image_2125; // @[Filter.scala 68:24]
  reg [3:0] image_2126; // @[Filter.scala 68:24]
  reg [3:0] image_2127; // @[Filter.scala 68:24]
  reg [3:0] image_2128; // @[Filter.scala 68:24]
  reg [3:0] image_2129; // @[Filter.scala 68:24]
  reg [3:0] image_2130; // @[Filter.scala 68:24]
  reg [3:0] image_2131; // @[Filter.scala 68:24]
  reg [3:0] image_2132; // @[Filter.scala 68:24]
  reg [3:0] image_2133; // @[Filter.scala 68:24]
  reg [3:0] image_2134; // @[Filter.scala 68:24]
  reg [3:0] image_2135; // @[Filter.scala 68:24]
  reg [3:0] image_2136; // @[Filter.scala 68:24]
  reg [3:0] image_2137; // @[Filter.scala 68:24]
  reg [3:0] image_2138; // @[Filter.scala 68:24]
  reg [3:0] image_2139; // @[Filter.scala 68:24]
  reg [3:0] image_2140; // @[Filter.scala 68:24]
  reg [3:0] image_2141; // @[Filter.scala 68:24]
  reg [3:0] image_2142; // @[Filter.scala 68:24]
  reg [3:0] image_2143; // @[Filter.scala 68:24]
  reg [3:0] image_2144; // @[Filter.scala 68:24]
  reg [3:0] image_2145; // @[Filter.scala 68:24]
  reg [3:0] image_2146; // @[Filter.scala 68:24]
  reg [3:0] image_2147; // @[Filter.scala 68:24]
  reg [3:0] image_2148; // @[Filter.scala 68:24]
  reg [3:0] image_2149; // @[Filter.scala 68:24]
  reg [3:0] image_2150; // @[Filter.scala 68:24]
  reg [3:0] image_2151; // @[Filter.scala 68:24]
  reg [3:0] image_2152; // @[Filter.scala 68:24]
  reg [3:0] image_2153; // @[Filter.scala 68:24]
  reg [3:0] image_2154; // @[Filter.scala 68:24]
  reg [3:0] image_2155; // @[Filter.scala 68:24]
  reg [3:0] image_2156; // @[Filter.scala 68:24]
  reg [3:0] image_2157; // @[Filter.scala 68:24]
  reg [3:0] image_2158; // @[Filter.scala 68:24]
  reg [3:0] image_2159; // @[Filter.scala 68:24]
  reg [3:0] image_2160; // @[Filter.scala 68:24]
  reg [3:0] image_2161; // @[Filter.scala 68:24]
  reg [3:0] image_2162; // @[Filter.scala 68:24]
  reg [3:0] image_2163; // @[Filter.scala 68:24]
  reg [3:0] image_2164; // @[Filter.scala 68:24]
  reg [3:0] image_2165; // @[Filter.scala 68:24]
  reg [3:0] image_2166; // @[Filter.scala 68:24]
  reg [3:0] image_2167; // @[Filter.scala 68:24]
  reg [3:0] image_2168; // @[Filter.scala 68:24]
  reg [3:0] image_2169; // @[Filter.scala 68:24]
  reg [3:0] image_2170; // @[Filter.scala 68:24]
  reg [3:0] image_2177; // @[Filter.scala 68:24]
  reg [3:0] image_2178; // @[Filter.scala 68:24]
  reg [3:0] image_2179; // @[Filter.scala 68:24]
  reg [3:0] image_2180; // @[Filter.scala 68:24]
  reg [3:0] image_2181; // @[Filter.scala 68:24]
  reg [3:0] image_2182; // @[Filter.scala 68:24]
  reg [3:0] image_2183; // @[Filter.scala 68:24]
  reg [3:0] image_2184; // @[Filter.scala 68:24]
  reg [3:0] image_2185; // @[Filter.scala 68:24]
  reg [3:0] image_2186; // @[Filter.scala 68:24]
  reg [3:0] image_2187; // @[Filter.scala 68:24]
  reg [3:0] image_2188; // @[Filter.scala 68:24]
  reg [3:0] image_2189; // @[Filter.scala 68:24]
  reg [3:0] image_2190; // @[Filter.scala 68:24]
  reg [3:0] image_2191; // @[Filter.scala 68:24]
  reg [3:0] image_2192; // @[Filter.scala 68:24]
  reg [3:0] image_2193; // @[Filter.scala 68:24]
  reg [3:0] image_2194; // @[Filter.scala 68:24]
  reg [3:0] image_2195; // @[Filter.scala 68:24]
  reg [3:0] image_2196; // @[Filter.scala 68:24]
  reg [3:0] image_2197; // @[Filter.scala 68:24]
  reg [3:0] image_2198; // @[Filter.scala 68:24]
  reg [3:0] image_2199; // @[Filter.scala 68:24]
  reg [3:0] image_2200; // @[Filter.scala 68:24]
  reg [3:0] image_2201; // @[Filter.scala 68:24]
  reg [3:0] image_2202; // @[Filter.scala 68:24]
  reg [3:0] image_2203; // @[Filter.scala 68:24]
  reg [3:0] image_2204; // @[Filter.scala 68:24]
  reg [3:0] image_2205; // @[Filter.scala 68:24]
  reg [3:0] image_2206; // @[Filter.scala 68:24]
  reg [3:0] image_2207; // @[Filter.scala 68:24]
  reg [3:0] image_2208; // @[Filter.scala 68:24]
  reg [3:0] image_2209; // @[Filter.scala 68:24]
  reg [3:0] image_2210; // @[Filter.scala 68:24]
  reg [3:0] image_2211; // @[Filter.scala 68:24]
  reg [3:0] image_2212; // @[Filter.scala 68:24]
  reg [3:0] image_2213; // @[Filter.scala 68:24]
  reg [3:0] image_2214; // @[Filter.scala 68:24]
  reg [3:0] image_2215; // @[Filter.scala 68:24]
  reg [3:0] image_2216; // @[Filter.scala 68:24]
  reg [3:0] image_2217; // @[Filter.scala 68:24]
  reg [3:0] image_2218; // @[Filter.scala 68:24]
  reg [3:0] image_2219; // @[Filter.scala 68:24]
  reg [3:0] image_2220; // @[Filter.scala 68:24]
  reg [3:0] image_2221; // @[Filter.scala 68:24]
  reg [3:0] image_2222; // @[Filter.scala 68:24]
  reg [3:0] image_2223; // @[Filter.scala 68:24]
  reg [3:0] image_2224; // @[Filter.scala 68:24]
  reg [3:0] image_2225; // @[Filter.scala 68:24]
  reg [3:0] image_2226; // @[Filter.scala 68:24]
  reg [3:0] image_2227; // @[Filter.scala 68:24]
  reg [3:0] image_2228; // @[Filter.scala 68:24]
  reg [3:0] image_2229; // @[Filter.scala 68:24]
  reg [3:0] image_2230; // @[Filter.scala 68:24]
  reg [3:0] image_2231; // @[Filter.scala 68:24]
  reg [3:0] image_2232; // @[Filter.scala 68:24]
  reg [3:0] image_2233; // @[Filter.scala 68:24]
  reg [3:0] image_2234; // @[Filter.scala 68:24]
  reg [3:0] image_2243; // @[Filter.scala 68:24]
  reg [3:0] image_2244; // @[Filter.scala 68:24]
  reg [3:0] image_2245; // @[Filter.scala 68:24]
  reg [3:0] image_2246; // @[Filter.scala 68:24]
  reg [3:0] image_2247; // @[Filter.scala 68:24]
  reg [3:0] image_2248; // @[Filter.scala 68:24]
  reg [3:0] image_2249; // @[Filter.scala 68:24]
  reg [3:0] image_2250; // @[Filter.scala 68:24]
  reg [3:0] image_2251; // @[Filter.scala 68:24]
  reg [3:0] image_2252; // @[Filter.scala 68:24]
  reg [3:0] image_2253; // @[Filter.scala 68:24]
  reg [3:0] image_2254; // @[Filter.scala 68:24]
  reg [3:0] image_2255; // @[Filter.scala 68:24]
  reg [3:0] image_2256; // @[Filter.scala 68:24]
  reg [3:0] image_2257; // @[Filter.scala 68:24]
  reg [3:0] image_2258; // @[Filter.scala 68:24]
  reg [3:0] image_2259; // @[Filter.scala 68:24]
  reg [3:0] image_2260; // @[Filter.scala 68:24]
  reg [3:0] image_2261; // @[Filter.scala 68:24]
  reg [3:0] image_2262; // @[Filter.scala 68:24]
  reg [3:0] image_2263; // @[Filter.scala 68:24]
  reg [3:0] image_2264; // @[Filter.scala 68:24]
  reg [3:0] image_2265; // @[Filter.scala 68:24]
  reg [3:0] image_2266; // @[Filter.scala 68:24]
  reg [3:0] image_2267; // @[Filter.scala 68:24]
  reg [3:0] image_2268; // @[Filter.scala 68:24]
  reg [3:0] image_2269; // @[Filter.scala 68:24]
  reg [3:0] image_2270; // @[Filter.scala 68:24]
  reg [3:0] image_2271; // @[Filter.scala 68:24]
  reg [3:0] image_2272; // @[Filter.scala 68:24]
  reg [3:0] image_2273; // @[Filter.scala 68:24]
  reg [3:0] image_2274; // @[Filter.scala 68:24]
  reg [3:0] image_2275; // @[Filter.scala 68:24]
  reg [3:0] image_2276; // @[Filter.scala 68:24]
  reg [3:0] image_2277; // @[Filter.scala 68:24]
  reg [3:0] image_2278; // @[Filter.scala 68:24]
  reg [3:0] image_2279; // @[Filter.scala 68:24]
  reg [3:0] image_2280; // @[Filter.scala 68:24]
  reg [3:0] image_2281; // @[Filter.scala 68:24]
  reg [3:0] image_2282; // @[Filter.scala 68:24]
  reg [3:0] image_2283; // @[Filter.scala 68:24]
  reg [3:0] image_2284; // @[Filter.scala 68:24]
  reg [3:0] image_2285; // @[Filter.scala 68:24]
  reg [3:0] image_2286; // @[Filter.scala 68:24]
  reg [3:0] image_2287; // @[Filter.scala 68:24]
  reg [3:0] image_2288; // @[Filter.scala 68:24]
  reg [3:0] image_2289; // @[Filter.scala 68:24]
  reg [3:0] image_2290; // @[Filter.scala 68:24]
  reg [3:0] image_2291; // @[Filter.scala 68:24]
  reg [3:0] image_2292; // @[Filter.scala 68:24]
  reg [3:0] image_2293; // @[Filter.scala 68:24]
  reg [3:0] image_2294; // @[Filter.scala 68:24]
  reg [3:0] image_2295; // @[Filter.scala 68:24]
  reg [3:0] image_2296; // @[Filter.scala 68:24]
  reg [3:0] image_2297; // @[Filter.scala 68:24]
  reg [3:0] image_2298; // @[Filter.scala 68:24]
  reg [3:0] image_2307; // @[Filter.scala 68:24]
  reg [3:0] image_2308; // @[Filter.scala 68:24]
  reg [3:0] image_2309; // @[Filter.scala 68:24]
  reg [3:0] image_2310; // @[Filter.scala 68:24]
  reg [3:0] image_2311; // @[Filter.scala 68:24]
  reg [3:0] image_2312; // @[Filter.scala 68:24]
  reg [3:0] image_2313; // @[Filter.scala 68:24]
  reg [3:0] image_2314; // @[Filter.scala 68:24]
  reg [3:0] image_2315; // @[Filter.scala 68:24]
  reg [3:0] image_2316; // @[Filter.scala 68:24]
  reg [3:0] image_2317; // @[Filter.scala 68:24]
  reg [3:0] image_2318; // @[Filter.scala 68:24]
  reg [3:0] image_2319; // @[Filter.scala 68:24]
  reg [3:0] image_2320; // @[Filter.scala 68:24]
  reg [3:0] image_2321; // @[Filter.scala 68:24]
  reg [3:0] image_2322; // @[Filter.scala 68:24]
  reg [3:0] image_2323; // @[Filter.scala 68:24]
  reg [3:0] image_2324; // @[Filter.scala 68:24]
  reg [3:0] image_2325; // @[Filter.scala 68:24]
  reg [3:0] image_2326; // @[Filter.scala 68:24]
  reg [3:0] image_2327; // @[Filter.scala 68:24]
  reg [3:0] image_2328; // @[Filter.scala 68:24]
  reg [3:0] image_2329; // @[Filter.scala 68:24]
  reg [3:0] image_2330; // @[Filter.scala 68:24]
  reg [3:0] image_2331; // @[Filter.scala 68:24]
  reg [3:0] image_2332; // @[Filter.scala 68:24]
  reg [3:0] image_2333; // @[Filter.scala 68:24]
  reg [3:0] image_2334; // @[Filter.scala 68:24]
  reg [3:0] image_2335; // @[Filter.scala 68:24]
  reg [3:0] image_2336; // @[Filter.scala 68:24]
  reg [3:0] image_2337; // @[Filter.scala 68:24]
  reg [3:0] image_2338; // @[Filter.scala 68:24]
  reg [3:0] image_2339; // @[Filter.scala 68:24]
  reg [3:0] image_2340; // @[Filter.scala 68:24]
  reg [3:0] image_2341; // @[Filter.scala 68:24]
  reg [3:0] image_2342; // @[Filter.scala 68:24]
  reg [3:0] image_2343; // @[Filter.scala 68:24]
  reg [3:0] image_2344; // @[Filter.scala 68:24]
  reg [3:0] image_2345; // @[Filter.scala 68:24]
  reg [3:0] image_2346; // @[Filter.scala 68:24]
  reg [3:0] image_2347; // @[Filter.scala 68:24]
  reg [3:0] image_2348; // @[Filter.scala 68:24]
  reg [3:0] image_2349; // @[Filter.scala 68:24]
  reg [3:0] image_2350; // @[Filter.scala 68:24]
  reg [3:0] image_2351; // @[Filter.scala 68:24]
  reg [3:0] image_2352; // @[Filter.scala 68:24]
  reg [3:0] image_2353; // @[Filter.scala 68:24]
  reg [3:0] image_2354; // @[Filter.scala 68:24]
  reg [3:0] image_2355; // @[Filter.scala 68:24]
  reg [3:0] image_2356; // @[Filter.scala 68:24]
  reg [3:0] image_2357; // @[Filter.scala 68:24]
  reg [3:0] image_2358; // @[Filter.scala 68:24]
  reg [3:0] image_2359; // @[Filter.scala 68:24]
  reg [3:0] image_2360; // @[Filter.scala 68:24]
  reg [3:0] image_2361; // @[Filter.scala 68:24]
  reg [3:0] image_2362; // @[Filter.scala 68:24]
  reg [3:0] image_2372; // @[Filter.scala 68:24]
  reg [3:0] image_2373; // @[Filter.scala 68:24]
  reg [3:0] image_2374; // @[Filter.scala 68:24]
  reg [3:0] image_2375; // @[Filter.scala 68:24]
  reg [3:0] image_2376; // @[Filter.scala 68:24]
  reg [3:0] image_2377; // @[Filter.scala 68:24]
  reg [3:0] image_2378; // @[Filter.scala 68:24]
  reg [3:0] image_2379; // @[Filter.scala 68:24]
  reg [3:0] image_2380; // @[Filter.scala 68:24]
  reg [3:0] image_2381; // @[Filter.scala 68:24]
  reg [3:0] image_2382; // @[Filter.scala 68:24]
  reg [3:0] image_2383; // @[Filter.scala 68:24]
  reg [3:0] image_2384; // @[Filter.scala 68:24]
  reg [3:0] image_2385; // @[Filter.scala 68:24]
  reg [3:0] image_2386; // @[Filter.scala 68:24]
  reg [3:0] image_2387; // @[Filter.scala 68:24]
  reg [3:0] image_2388; // @[Filter.scala 68:24]
  reg [3:0] image_2389; // @[Filter.scala 68:24]
  reg [3:0] image_2390; // @[Filter.scala 68:24]
  reg [3:0] image_2391; // @[Filter.scala 68:24]
  reg [3:0] image_2392; // @[Filter.scala 68:24]
  reg [3:0] image_2393; // @[Filter.scala 68:24]
  reg [3:0] image_2394; // @[Filter.scala 68:24]
  reg [3:0] image_2395; // @[Filter.scala 68:24]
  reg [3:0] image_2396; // @[Filter.scala 68:24]
  reg [3:0] image_2397; // @[Filter.scala 68:24]
  reg [3:0] image_2398; // @[Filter.scala 68:24]
  reg [3:0] image_2399; // @[Filter.scala 68:24]
  reg [3:0] image_2400; // @[Filter.scala 68:24]
  reg [3:0] image_2401; // @[Filter.scala 68:24]
  reg [3:0] image_2402; // @[Filter.scala 68:24]
  reg [3:0] image_2403; // @[Filter.scala 68:24]
  reg [3:0] image_2404; // @[Filter.scala 68:24]
  reg [3:0] image_2405; // @[Filter.scala 68:24]
  reg [3:0] image_2406; // @[Filter.scala 68:24]
  reg [3:0] image_2407; // @[Filter.scala 68:24]
  reg [3:0] image_2408; // @[Filter.scala 68:24]
  reg [3:0] image_2409; // @[Filter.scala 68:24]
  reg [3:0] image_2410; // @[Filter.scala 68:24]
  reg [3:0] image_2411; // @[Filter.scala 68:24]
  reg [3:0] image_2412; // @[Filter.scala 68:24]
  reg [3:0] image_2413; // @[Filter.scala 68:24]
  reg [3:0] image_2414; // @[Filter.scala 68:24]
  reg [3:0] image_2415; // @[Filter.scala 68:24]
  reg [3:0] image_2416; // @[Filter.scala 68:24]
  reg [3:0] image_2417; // @[Filter.scala 68:24]
  reg [3:0] image_2418; // @[Filter.scala 68:24]
  reg [3:0] image_2419; // @[Filter.scala 68:24]
  reg [3:0] image_2420; // @[Filter.scala 68:24]
  reg [3:0] image_2421; // @[Filter.scala 68:24]
  reg [3:0] image_2422; // @[Filter.scala 68:24]
  reg [3:0] image_2423; // @[Filter.scala 68:24]
  reg [3:0] image_2424; // @[Filter.scala 68:24]
  reg [3:0] image_2425; // @[Filter.scala 68:24]
  reg [3:0] image_2426; // @[Filter.scala 68:24]
  reg [3:0] image_2437; // @[Filter.scala 68:24]
  reg [3:0] image_2438; // @[Filter.scala 68:24]
  reg [3:0] image_2439; // @[Filter.scala 68:24]
  reg [3:0] image_2440; // @[Filter.scala 68:24]
  reg [3:0] image_2441; // @[Filter.scala 68:24]
  reg [3:0] image_2442; // @[Filter.scala 68:24]
  reg [3:0] image_2443; // @[Filter.scala 68:24]
  reg [3:0] image_2444; // @[Filter.scala 68:24]
  reg [3:0] image_2445; // @[Filter.scala 68:24]
  reg [3:0] image_2446; // @[Filter.scala 68:24]
  reg [3:0] image_2447; // @[Filter.scala 68:24]
  reg [3:0] image_2448; // @[Filter.scala 68:24]
  reg [3:0] image_2449; // @[Filter.scala 68:24]
  reg [3:0] image_2450; // @[Filter.scala 68:24]
  reg [3:0] image_2451; // @[Filter.scala 68:24]
  reg [3:0] image_2452; // @[Filter.scala 68:24]
  reg [3:0] image_2453; // @[Filter.scala 68:24]
  reg [3:0] image_2454; // @[Filter.scala 68:24]
  reg [3:0] image_2455; // @[Filter.scala 68:24]
  reg [3:0] image_2456; // @[Filter.scala 68:24]
  reg [3:0] image_2457; // @[Filter.scala 68:24]
  reg [3:0] image_2458; // @[Filter.scala 68:24]
  reg [3:0] image_2459; // @[Filter.scala 68:24]
  reg [3:0] image_2460; // @[Filter.scala 68:24]
  reg [3:0] image_2461; // @[Filter.scala 68:24]
  reg [3:0] image_2462; // @[Filter.scala 68:24]
  reg [3:0] image_2463; // @[Filter.scala 68:24]
  reg [3:0] image_2464; // @[Filter.scala 68:24]
  reg [3:0] image_2465; // @[Filter.scala 68:24]
  reg [3:0] image_2466; // @[Filter.scala 68:24]
  reg [3:0] image_2467; // @[Filter.scala 68:24]
  reg [3:0] image_2468; // @[Filter.scala 68:24]
  reg [3:0] image_2469; // @[Filter.scala 68:24]
  reg [3:0] image_2470; // @[Filter.scala 68:24]
  reg [3:0] image_2471; // @[Filter.scala 68:24]
  reg [3:0] image_2472; // @[Filter.scala 68:24]
  reg [3:0] image_2473; // @[Filter.scala 68:24]
  reg [3:0] image_2474; // @[Filter.scala 68:24]
  reg [3:0] image_2475; // @[Filter.scala 68:24]
  reg [3:0] image_2476; // @[Filter.scala 68:24]
  reg [3:0] image_2477; // @[Filter.scala 68:24]
  reg [3:0] image_2478; // @[Filter.scala 68:24]
  reg [3:0] image_2479; // @[Filter.scala 68:24]
  reg [3:0] image_2480; // @[Filter.scala 68:24]
  reg [3:0] image_2481; // @[Filter.scala 68:24]
  reg [3:0] image_2482; // @[Filter.scala 68:24]
  reg [3:0] image_2483; // @[Filter.scala 68:24]
  reg [3:0] image_2484; // @[Filter.scala 68:24]
  reg [3:0] image_2485; // @[Filter.scala 68:24]
  reg [3:0] image_2486; // @[Filter.scala 68:24]
  reg [3:0] image_2487; // @[Filter.scala 68:24]
  reg [3:0] image_2488; // @[Filter.scala 68:24]
  reg [3:0] image_2489; // @[Filter.scala 68:24]
  reg [3:0] image_2490; // @[Filter.scala 68:24]
  reg [3:0] image_2502; // @[Filter.scala 68:24]
  reg [3:0] image_2503; // @[Filter.scala 68:24]
  reg [3:0] image_2504; // @[Filter.scala 68:24]
  reg [3:0] image_2505; // @[Filter.scala 68:24]
  reg [3:0] image_2506; // @[Filter.scala 68:24]
  reg [3:0] image_2507; // @[Filter.scala 68:24]
  reg [3:0] image_2508; // @[Filter.scala 68:24]
  reg [3:0] image_2509; // @[Filter.scala 68:24]
  reg [3:0] image_2510; // @[Filter.scala 68:24]
  reg [3:0] image_2511; // @[Filter.scala 68:24]
  reg [3:0] image_2512; // @[Filter.scala 68:24]
  reg [3:0] image_2513; // @[Filter.scala 68:24]
  reg [3:0] image_2514; // @[Filter.scala 68:24]
  reg [3:0] image_2515; // @[Filter.scala 68:24]
  reg [3:0] image_2516; // @[Filter.scala 68:24]
  reg [3:0] image_2517; // @[Filter.scala 68:24]
  reg [3:0] image_2518; // @[Filter.scala 68:24]
  reg [3:0] image_2519; // @[Filter.scala 68:24]
  reg [3:0] image_2520; // @[Filter.scala 68:24]
  reg [3:0] image_2521; // @[Filter.scala 68:24]
  reg [3:0] image_2522; // @[Filter.scala 68:24]
  reg [3:0] image_2523; // @[Filter.scala 68:24]
  reg [3:0] image_2524; // @[Filter.scala 68:24]
  reg [3:0] image_2525; // @[Filter.scala 68:24]
  reg [3:0] image_2526; // @[Filter.scala 68:24]
  reg [3:0] image_2527; // @[Filter.scala 68:24]
  reg [3:0] image_2528; // @[Filter.scala 68:24]
  reg [3:0] image_2529; // @[Filter.scala 68:24]
  reg [3:0] image_2530; // @[Filter.scala 68:24]
  reg [3:0] image_2531; // @[Filter.scala 68:24]
  reg [3:0] image_2532; // @[Filter.scala 68:24]
  reg [3:0] image_2533; // @[Filter.scala 68:24]
  reg [3:0] image_2534; // @[Filter.scala 68:24]
  reg [3:0] image_2535; // @[Filter.scala 68:24]
  reg [3:0] image_2536; // @[Filter.scala 68:24]
  reg [3:0] image_2537; // @[Filter.scala 68:24]
  reg [3:0] image_2538; // @[Filter.scala 68:24]
  reg [3:0] image_2539; // @[Filter.scala 68:24]
  reg [3:0] image_2540; // @[Filter.scala 68:24]
  reg [3:0] image_2541; // @[Filter.scala 68:24]
  reg [3:0] image_2542; // @[Filter.scala 68:24]
  reg [3:0] image_2543; // @[Filter.scala 68:24]
  reg [3:0] image_2544; // @[Filter.scala 68:24]
  reg [3:0] image_2545; // @[Filter.scala 68:24]
  reg [3:0] image_2546; // @[Filter.scala 68:24]
  reg [3:0] image_2547; // @[Filter.scala 68:24]
  reg [3:0] image_2548; // @[Filter.scala 68:24]
  reg [3:0] image_2549; // @[Filter.scala 68:24]
  reg [3:0] image_2550; // @[Filter.scala 68:24]
  reg [3:0] image_2551; // @[Filter.scala 68:24]
  reg [3:0] image_2552; // @[Filter.scala 68:24]
  reg [3:0] image_2553; // @[Filter.scala 68:24]
  reg [3:0] image_2554; // @[Filter.scala 68:24]
  reg [3:0] image_2567; // @[Filter.scala 68:24]
  reg [3:0] image_2568; // @[Filter.scala 68:24]
  reg [3:0] image_2569; // @[Filter.scala 68:24]
  reg [3:0] image_2570; // @[Filter.scala 68:24]
  reg [3:0] image_2571; // @[Filter.scala 68:24]
  reg [3:0] image_2572; // @[Filter.scala 68:24]
  reg [3:0] image_2573; // @[Filter.scala 68:24]
  reg [3:0] image_2574; // @[Filter.scala 68:24]
  reg [3:0] image_2575; // @[Filter.scala 68:24]
  reg [3:0] image_2576; // @[Filter.scala 68:24]
  reg [3:0] image_2577; // @[Filter.scala 68:24]
  reg [3:0] image_2578; // @[Filter.scala 68:24]
  reg [3:0] image_2579; // @[Filter.scala 68:24]
  reg [3:0] image_2580; // @[Filter.scala 68:24]
  reg [3:0] image_2581; // @[Filter.scala 68:24]
  reg [3:0] image_2582; // @[Filter.scala 68:24]
  reg [3:0] image_2583; // @[Filter.scala 68:24]
  reg [3:0] image_2584; // @[Filter.scala 68:24]
  reg [3:0] image_2585; // @[Filter.scala 68:24]
  reg [3:0] image_2586; // @[Filter.scala 68:24]
  reg [3:0] image_2587; // @[Filter.scala 68:24]
  reg [3:0] image_2588; // @[Filter.scala 68:24]
  reg [3:0] image_2589; // @[Filter.scala 68:24]
  reg [3:0] image_2590; // @[Filter.scala 68:24]
  reg [3:0] image_2591; // @[Filter.scala 68:24]
  reg [3:0] image_2592; // @[Filter.scala 68:24]
  reg [3:0] image_2593; // @[Filter.scala 68:24]
  reg [3:0] image_2594; // @[Filter.scala 68:24]
  reg [3:0] image_2595; // @[Filter.scala 68:24]
  reg [3:0] image_2596; // @[Filter.scala 68:24]
  reg [3:0] image_2597; // @[Filter.scala 68:24]
  reg [3:0] image_2598; // @[Filter.scala 68:24]
  reg [3:0] image_2599; // @[Filter.scala 68:24]
  reg [3:0] image_2600; // @[Filter.scala 68:24]
  reg [3:0] image_2601; // @[Filter.scala 68:24]
  reg [3:0] image_2602; // @[Filter.scala 68:24]
  reg [3:0] image_2603; // @[Filter.scala 68:24]
  reg [3:0] image_2604; // @[Filter.scala 68:24]
  reg [3:0] image_2605; // @[Filter.scala 68:24]
  reg [3:0] image_2606; // @[Filter.scala 68:24]
  reg [3:0] image_2607; // @[Filter.scala 68:24]
  reg [3:0] image_2608; // @[Filter.scala 68:24]
  reg [3:0] image_2609; // @[Filter.scala 68:24]
  reg [3:0] image_2610; // @[Filter.scala 68:24]
  reg [3:0] image_2611; // @[Filter.scala 68:24]
  reg [3:0] image_2612; // @[Filter.scala 68:24]
  reg [3:0] image_2613; // @[Filter.scala 68:24]
  reg [3:0] image_2614; // @[Filter.scala 68:24]
  reg [3:0] image_2615; // @[Filter.scala 68:24]
  reg [3:0] image_2616; // @[Filter.scala 68:24]
  reg [3:0] image_2617; // @[Filter.scala 68:24]
  reg [3:0] image_2618; // @[Filter.scala 68:24]
  reg [3:0] image_2632; // @[Filter.scala 68:24]
  reg [3:0] image_2633; // @[Filter.scala 68:24]
  reg [3:0] image_2634; // @[Filter.scala 68:24]
  reg [3:0] image_2635; // @[Filter.scala 68:24]
  reg [3:0] image_2636; // @[Filter.scala 68:24]
  reg [3:0] image_2637; // @[Filter.scala 68:24]
  reg [3:0] image_2638; // @[Filter.scala 68:24]
  reg [3:0] image_2639; // @[Filter.scala 68:24]
  reg [3:0] image_2640; // @[Filter.scala 68:24]
  reg [3:0] image_2641; // @[Filter.scala 68:24]
  reg [3:0] image_2642; // @[Filter.scala 68:24]
  reg [3:0] image_2643; // @[Filter.scala 68:24]
  reg [3:0] image_2644; // @[Filter.scala 68:24]
  reg [3:0] image_2645; // @[Filter.scala 68:24]
  reg [3:0] image_2646; // @[Filter.scala 68:24]
  reg [3:0] image_2647; // @[Filter.scala 68:24]
  reg [3:0] image_2648; // @[Filter.scala 68:24]
  reg [3:0] image_2649; // @[Filter.scala 68:24]
  reg [3:0] image_2650; // @[Filter.scala 68:24]
  reg [3:0] image_2651; // @[Filter.scala 68:24]
  reg [3:0] image_2652; // @[Filter.scala 68:24]
  reg [3:0] image_2653; // @[Filter.scala 68:24]
  reg [3:0] image_2654; // @[Filter.scala 68:24]
  reg [3:0] image_2655; // @[Filter.scala 68:24]
  reg [3:0] image_2656; // @[Filter.scala 68:24]
  reg [3:0] image_2657; // @[Filter.scala 68:24]
  reg [3:0] image_2658; // @[Filter.scala 68:24]
  reg [3:0] image_2659; // @[Filter.scala 68:24]
  reg [3:0] image_2660; // @[Filter.scala 68:24]
  reg [3:0] image_2661; // @[Filter.scala 68:24]
  reg [3:0] image_2662; // @[Filter.scala 68:24]
  reg [3:0] image_2663; // @[Filter.scala 68:24]
  reg [3:0] image_2664; // @[Filter.scala 68:24]
  reg [3:0] image_2665; // @[Filter.scala 68:24]
  reg [3:0] image_2666; // @[Filter.scala 68:24]
  reg [3:0] image_2667; // @[Filter.scala 68:24]
  reg [3:0] image_2668; // @[Filter.scala 68:24]
  reg [3:0] image_2669; // @[Filter.scala 68:24]
  reg [3:0] image_2670; // @[Filter.scala 68:24]
  reg [3:0] image_2671; // @[Filter.scala 68:24]
  reg [3:0] image_2672; // @[Filter.scala 68:24]
  reg [3:0] image_2673; // @[Filter.scala 68:24]
  reg [3:0] image_2674; // @[Filter.scala 68:24]
  reg [3:0] image_2675; // @[Filter.scala 68:24]
  reg [3:0] image_2676; // @[Filter.scala 68:24]
  reg [3:0] image_2677; // @[Filter.scala 68:24]
  reg [3:0] image_2678; // @[Filter.scala 68:24]
  reg [3:0] image_2679; // @[Filter.scala 68:24]
  reg [3:0] image_2680; // @[Filter.scala 68:24]
  reg [3:0] image_2681; // @[Filter.scala 68:24]
  reg [3:0] image_2682; // @[Filter.scala 68:24]
  reg [3:0] image_2697; // @[Filter.scala 68:24]
  reg [3:0] image_2698; // @[Filter.scala 68:24]
  reg [3:0] image_2699; // @[Filter.scala 68:24]
  reg [3:0] image_2700; // @[Filter.scala 68:24]
  reg [3:0] image_2701; // @[Filter.scala 68:24]
  reg [3:0] image_2702; // @[Filter.scala 68:24]
  reg [3:0] image_2703; // @[Filter.scala 68:24]
  reg [3:0] image_2704; // @[Filter.scala 68:24]
  reg [3:0] image_2705; // @[Filter.scala 68:24]
  reg [3:0] image_2706; // @[Filter.scala 68:24]
  reg [3:0] image_2707; // @[Filter.scala 68:24]
  reg [3:0] image_2708; // @[Filter.scala 68:24]
  reg [3:0] image_2709; // @[Filter.scala 68:24]
  reg [3:0] image_2710; // @[Filter.scala 68:24]
  reg [3:0] image_2711; // @[Filter.scala 68:24]
  reg [3:0] image_2712; // @[Filter.scala 68:24]
  reg [3:0] image_2713; // @[Filter.scala 68:24]
  reg [3:0] image_2714; // @[Filter.scala 68:24]
  reg [3:0] image_2715; // @[Filter.scala 68:24]
  reg [3:0] image_2716; // @[Filter.scala 68:24]
  reg [3:0] image_2717; // @[Filter.scala 68:24]
  reg [3:0] image_2718; // @[Filter.scala 68:24]
  reg [3:0] image_2719; // @[Filter.scala 68:24]
  reg [3:0] image_2720; // @[Filter.scala 68:24]
  reg [3:0] image_2721; // @[Filter.scala 68:24]
  reg [3:0] image_2722; // @[Filter.scala 68:24]
  reg [3:0] image_2723; // @[Filter.scala 68:24]
  reg [3:0] image_2724; // @[Filter.scala 68:24]
  reg [3:0] image_2725; // @[Filter.scala 68:24]
  reg [3:0] image_2726; // @[Filter.scala 68:24]
  reg [3:0] image_2727; // @[Filter.scala 68:24]
  reg [3:0] image_2728; // @[Filter.scala 68:24]
  reg [3:0] image_2729; // @[Filter.scala 68:24]
  reg [3:0] image_2730; // @[Filter.scala 68:24]
  reg [3:0] image_2731; // @[Filter.scala 68:24]
  reg [3:0] image_2732; // @[Filter.scala 68:24]
  reg [3:0] image_2733; // @[Filter.scala 68:24]
  reg [3:0] image_2734; // @[Filter.scala 68:24]
  reg [3:0] image_2735; // @[Filter.scala 68:24]
  reg [3:0] image_2736; // @[Filter.scala 68:24]
  reg [3:0] image_2737; // @[Filter.scala 68:24]
  reg [3:0] image_2738; // @[Filter.scala 68:24]
  reg [3:0] image_2739; // @[Filter.scala 68:24]
  reg [3:0] image_2740; // @[Filter.scala 68:24]
  reg [3:0] image_2741; // @[Filter.scala 68:24]
  reg [3:0] image_2742; // @[Filter.scala 68:24]
  reg [3:0] image_2743; // @[Filter.scala 68:24]
  reg [3:0] image_2744; // @[Filter.scala 68:24]
  reg [3:0] image_2745; // @[Filter.scala 68:24]
  reg [3:0] image_2763; // @[Filter.scala 68:24]
  reg [3:0] image_2764; // @[Filter.scala 68:24]
  reg [3:0] image_2765; // @[Filter.scala 68:24]
  reg [3:0] image_2766; // @[Filter.scala 68:24]
  reg [3:0] image_2767; // @[Filter.scala 68:24]
  reg [3:0] image_2768; // @[Filter.scala 68:24]
  reg [3:0] image_2769; // @[Filter.scala 68:24]
  reg [3:0] image_2770; // @[Filter.scala 68:24]
  reg [3:0] image_2771; // @[Filter.scala 68:24]
  reg [3:0] image_2772; // @[Filter.scala 68:24]
  reg [3:0] image_2773; // @[Filter.scala 68:24]
  reg [3:0] image_2774; // @[Filter.scala 68:24]
  reg [3:0] image_2775; // @[Filter.scala 68:24]
  reg [3:0] image_2776; // @[Filter.scala 68:24]
  reg [3:0] image_2777; // @[Filter.scala 68:24]
  reg [3:0] image_2778; // @[Filter.scala 68:24]
  reg [3:0] image_2779; // @[Filter.scala 68:24]
  reg [3:0] image_2780; // @[Filter.scala 68:24]
  reg [3:0] image_2781; // @[Filter.scala 68:24]
  reg [3:0] image_2782; // @[Filter.scala 68:24]
  reg [3:0] image_2783; // @[Filter.scala 68:24]
  reg [3:0] image_2784; // @[Filter.scala 68:24]
  reg [3:0] image_2785; // @[Filter.scala 68:24]
  reg [3:0] image_2786; // @[Filter.scala 68:24]
  reg [3:0] image_2787; // @[Filter.scala 68:24]
  reg [3:0] image_2788; // @[Filter.scala 68:24]
  reg [3:0] image_2789; // @[Filter.scala 68:24]
  reg [3:0] image_2790; // @[Filter.scala 68:24]
  reg [3:0] image_2791; // @[Filter.scala 68:24]
  reg [3:0] image_2792; // @[Filter.scala 68:24]
  reg [3:0] image_2793; // @[Filter.scala 68:24]
  reg [3:0] image_2794; // @[Filter.scala 68:24]
  reg [3:0] image_2795; // @[Filter.scala 68:24]
  reg [3:0] image_2796; // @[Filter.scala 68:24]
  reg [3:0] image_2797; // @[Filter.scala 68:24]
  reg [3:0] image_2798; // @[Filter.scala 68:24]
  reg [3:0] image_2799; // @[Filter.scala 68:24]
  reg [3:0] image_2800; // @[Filter.scala 68:24]
  reg [3:0] image_2801; // @[Filter.scala 68:24]
  reg [3:0] image_2802; // @[Filter.scala 68:24]
  reg [3:0] image_2803; // @[Filter.scala 68:24]
  reg [3:0] image_2804; // @[Filter.scala 68:24]
  reg [3:0] image_2805; // @[Filter.scala 68:24]
  reg [3:0] image_2806; // @[Filter.scala 68:24]
  reg [3:0] image_2807; // @[Filter.scala 68:24]
  reg [3:0] image_2808; // @[Filter.scala 68:24]
  reg [3:0] image_2828; // @[Filter.scala 68:24]
  reg [3:0] image_2829; // @[Filter.scala 68:24]
  reg [3:0] image_2830; // @[Filter.scala 68:24]
  reg [3:0] image_2831; // @[Filter.scala 68:24]
  reg [3:0] image_2832; // @[Filter.scala 68:24]
  reg [3:0] image_2833; // @[Filter.scala 68:24]
  reg [3:0] image_2834; // @[Filter.scala 68:24]
  reg [3:0] image_2835; // @[Filter.scala 68:24]
  reg [3:0] image_2836; // @[Filter.scala 68:24]
  reg [3:0] image_2837; // @[Filter.scala 68:24]
  reg [3:0] image_2838; // @[Filter.scala 68:24]
  reg [3:0] image_2839; // @[Filter.scala 68:24]
  reg [3:0] image_2840; // @[Filter.scala 68:24]
  reg [3:0] image_2841; // @[Filter.scala 68:24]
  reg [3:0] image_2842; // @[Filter.scala 68:24]
  reg [3:0] image_2843; // @[Filter.scala 68:24]
  reg [3:0] image_2844; // @[Filter.scala 68:24]
  reg [3:0] image_2845; // @[Filter.scala 68:24]
  reg [3:0] image_2846; // @[Filter.scala 68:24]
  reg [3:0] image_2847; // @[Filter.scala 68:24]
  reg [3:0] image_2848; // @[Filter.scala 68:24]
  reg [3:0] image_2849; // @[Filter.scala 68:24]
  reg [3:0] image_2850; // @[Filter.scala 68:24]
  reg [3:0] image_2851; // @[Filter.scala 68:24]
  reg [3:0] image_2852; // @[Filter.scala 68:24]
  reg [3:0] image_2853; // @[Filter.scala 68:24]
  reg [3:0] image_2854; // @[Filter.scala 68:24]
  reg [3:0] image_2855; // @[Filter.scala 68:24]
  reg [3:0] image_2856; // @[Filter.scala 68:24]
  reg [3:0] image_2857; // @[Filter.scala 68:24]
  reg [3:0] image_2858; // @[Filter.scala 68:24]
  reg [3:0] image_2859; // @[Filter.scala 68:24]
  reg [3:0] image_2860; // @[Filter.scala 68:24]
  reg [3:0] image_2861; // @[Filter.scala 68:24]
  reg [3:0] image_2862; // @[Filter.scala 68:24]
  reg [3:0] image_2863; // @[Filter.scala 68:24]
  reg [3:0] image_2864; // @[Filter.scala 68:24]
  reg [3:0] image_2865; // @[Filter.scala 68:24]
  reg [3:0] image_2866; // @[Filter.scala 68:24]
  reg [3:0] image_2867; // @[Filter.scala 68:24]
  reg [3:0] image_2868; // @[Filter.scala 68:24]
  reg [3:0] image_2869; // @[Filter.scala 68:24]
  reg [3:0] image_2870; // @[Filter.scala 68:24]
  reg [3:0] image_2871; // @[Filter.scala 68:24]
  reg [3:0] image_2895; // @[Filter.scala 68:24]
  reg [3:0] image_2896; // @[Filter.scala 68:24]
  reg [3:0] image_2897; // @[Filter.scala 68:24]
  reg [3:0] image_2898; // @[Filter.scala 68:24]
  reg [3:0] image_2899; // @[Filter.scala 68:24]
  reg [3:0] image_2900; // @[Filter.scala 68:24]
  reg [3:0] image_2901; // @[Filter.scala 68:24]
  reg [3:0] image_2902; // @[Filter.scala 68:24]
  reg [3:0] image_2903; // @[Filter.scala 68:24]
  reg [3:0] image_2904; // @[Filter.scala 68:24]
  reg [3:0] image_2905; // @[Filter.scala 68:24]
  reg [3:0] image_2906; // @[Filter.scala 68:24]
  reg [3:0] image_2907; // @[Filter.scala 68:24]
  reg [3:0] image_2908; // @[Filter.scala 68:24]
  reg [3:0] image_2909; // @[Filter.scala 68:24]
  reg [3:0] image_2910; // @[Filter.scala 68:24]
  reg [3:0] image_2911; // @[Filter.scala 68:24]
  reg [3:0] image_2912; // @[Filter.scala 68:24]
  reg [3:0] image_2913; // @[Filter.scala 68:24]
  reg [3:0] image_2914; // @[Filter.scala 68:24]
  reg [3:0] image_2915; // @[Filter.scala 68:24]
  reg [3:0] image_2916; // @[Filter.scala 68:24]
  reg [3:0] image_2917; // @[Filter.scala 68:24]
  reg [3:0] image_2918; // @[Filter.scala 68:24]
  reg [3:0] image_2919; // @[Filter.scala 68:24]
  reg [3:0] image_2920; // @[Filter.scala 68:24]
  reg [3:0] image_2921; // @[Filter.scala 68:24]
  reg [3:0] image_2922; // @[Filter.scala 68:24]
  reg [3:0] image_2923; // @[Filter.scala 68:24]
  reg [3:0] image_2924; // @[Filter.scala 68:24]
  reg [3:0] image_2925; // @[Filter.scala 68:24]
  reg [3:0] image_2926; // @[Filter.scala 68:24]
  reg [3:0] image_2927; // @[Filter.scala 68:24]
  reg [3:0] image_2928; // @[Filter.scala 68:24]
  reg [3:0] image_2929; // @[Filter.scala 68:24]
  reg [3:0] image_2930; // @[Filter.scala 68:24]
  reg [3:0] image_2931; // @[Filter.scala 68:24]
  reg [3:0] image_2932; // @[Filter.scala 68:24]
  reg [3:0] image_2933; // @[Filter.scala 68:24]
  reg [3:0] image_2934; // @[Filter.scala 68:24]
  reg [3:0] image_2965; // @[Filter.scala 68:24]
  reg [3:0] image_2966; // @[Filter.scala 68:24]
  reg [3:0] image_2967; // @[Filter.scala 68:24]
  reg [3:0] image_2968; // @[Filter.scala 68:24]
  reg [3:0] image_2969; // @[Filter.scala 68:24]
  reg [3:0] image_2970; // @[Filter.scala 68:24]
  reg [3:0] image_2971; // @[Filter.scala 68:24]
  reg [3:0] image_2972; // @[Filter.scala 68:24]
  reg [3:0] image_2973; // @[Filter.scala 68:24]
  reg [3:0] image_2974; // @[Filter.scala 68:24]
  reg [3:0] image_2975; // @[Filter.scala 68:24]
  reg [3:0] image_2976; // @[Filter.scala 68:24]
  reg [3:0] image_2977; // @[Filter.scala 68:24]
  reg [3:0] image_2978; // @[Filter.scala 68:24]
  reg [3:0] image_2979; // @[Filter.scala 68:24]
  reg [3:0] image_2980; // @[Filter.scala 68:24]
  reg [3:0] image_2981; // @[Filter.scala 68:24]
  reg [3:0] image_2982; // @[Filter.scala 68:24]
  reg [3:0] image_2983; // @[Filter.scala 68:24]
  reg [3:0] image_2984; // @[Filter.scala 68:24]
  reg [3:0] image_2985; // @[Filter.scala 68:24]
  reg [3:0] image_2986; // @[Filter.scala 68:24]
  reg [3:0] image_2987; // @[Filter.scala 68:24]
  reg [3:0] image_2988; // @[Filter.scala 68:24]
  reg [3:0] image_2989; // @[Filter.scala 68:24]
  reg [3:0] image_2990; // @[Filter.scala 68:24]
  reg [3:0] image_2991; // @[Filter.scala 68:24]
  reg [3:0] image_2992; // @[Filter.scala 68:24]
  reg [3:0] image_2993; // @[Filter.scala 68:24]
  reg [3:0] image_2994; // @[Filter.scala 68:24]
  reg [3:0] image_2995; // @[Filter.scala 68:24]
  reg [3:0] image_2996; // @[Filter.scala 68:24]
  reg [3:0] image_3035; // @[Filter.scala 68:24]
  reg [3:0] image_3036; // @[Filter.scala 68:24]
  reg [3:0] image_3037; // @[Filter.scala 68:24]
  reg [3:0] image_3038; // @[Filter.scala 68:24]
  reg [3:0] image_3039; // @[Filter.scala 68:24]
  reg [3:0] image_3040; // @[Filter.scala 68:24]
  reg [3:0] image_3041; // @[Filter.scala 68:24]
  reg [3:0] image_3042; // @[Filter.scala 68:24]
  reg [3:0] image_3043; // @[Filter.scala 68:24]
  reg [3:0] image_3044; // @[Filter.scala 68:24]
  reg [3:0] image_3045; // @[Filter.scala 68:24]
  reg [3:0] image_3046; // @[Filter.scala 68:24]
  reg [3:0] image_3047; // @[Filter.scala 68:24]
  reg [3:0] image_3048; // @[Filter.scala 68:24]
  reg [3:0] image_3049; // @[Filter.scala 68:24]
  reg [3:0] image_3050; // @[Filter.scala 68:24]
  reg [3:0] image_3051; // @[Filter.scala 68:24]
  reg [3:0] image_3052; // @[Filter.scala 68:24]
  reg [3:0] image_3053; // @[Filter.scala 68:24]
  reg [3:0] image_3054; // @[Filter.scala 68:24]
  reg [3:0] image_3055; // @[Filter.scala 68:24]
  reg [3:0] image_3056; // @[Filter.scala 68:24]
  reg [3:0] kernelCounter; // @[Counter.scala 29:33]
  wire  kernelCountReset = kernelCounter == 4'h8; // @[Counter.scala 38:24]
  wire [3:0] _T_15 = kernelCounter + 4'h1; // @[Counter.scala 39:22]
  wire  _GEN_24705 = 3'h0 == io_SPI_filterIndex[2:0]; // @[Filter.scala 125:36]
  wire  _GEN_24706 = 4'h4 == kernelCounter; // @[Filter.scala 125:36]
  wire [4:0] _GEN_7 = _GEN_24705 & _GEN_24706 ? $signed(5'sh1) : $signed(5'sh0); // @[Filter.scala 125:36]
  wire  _GEN_24708 = 4'h5 == kernelCounter; // @[Filter.scala 125:36]
  wire [4:0] _GEN_8 = _GEN_24705 & _GEN_24708 ? $signed(5'sh0) : $signed(_GEN_7); // @[Filter.scala 125:36]
  wire  _GEN_24710 = 4'h6 == kernelCounter; // @[Filter.scala 125:36]
  wire [4:0] _GEN_9 = _GEN_24705 & _GEN_24710 ? $signed(5'sh0) : $signed(_GEN_8); // @[Filter.scala 125:36]
  wire  _GEN_24712 = 4'h7 == kernelCounter; // @[Filter.scala 125:36]
  wire [4:0] _GEN_10 = _GEN_24705 & _GEN_24712 ? $signed(5'sh0) : $signed(_GEN_9); // @[Filter.scala 125:36]
  wire  _GEN_24714 = 4'h8 == kernelCounter; // @[Filter.scala 125:36]
  wire [4:0] _GEN_11 = _GEN_24705 & _GEN_24714 ? $signed(5'sh0) : $signed(_GEN_10); // @[Filter.scala 125:36]
  wire  _GEN_24715 = 3'h1 == io_SPI_filterIndex[2:0]; // @[Filter.scala 125:36]
  wire  _GEN_24716 = 4'h0 == kernelCounter; // @[Filter.scala 125:36]
  wire [4:0] _GEN_12 = _GEN_24715 & _GEN_24716 ? $signed(5'sh1) : $signed(_GEN_11); // @[Filter.scala 125:36]
  wire  _GEN_24718 = 4'h1 == kernelCounter; // @[Filter.scala 125:36]
  wire [4:0] _GEN_13 = _GEN_24715 & _GEN_24718 ? $signed(5'sh1) : $signed(_GEN_12); // @[Filter.scala 125:36]
  wire  _GEN_24720 = 4'h2 == kernelCounter; // @[Filter.scala 125:36]
  wire [4:0] _GEN_14 = _GEN_24715 & _GEN_24720 ? $signed(5'sh1) : $signed(_GEN_13); // @[Filter.scala 125:36]
  wire  _GEN_24722 = 4'h3 == kernelCounter; // @[Filter.scala 125:36]
  wire [4:0] _GEN_15 = _GEN_24715 & _GEN_24722 ? $signed(5'sh1) : $signed(_GEN_14); // @[Filter.scala 125:36]
  wire [4:0] _GEN_16 = _GEN_24715 & _GEN_24706 ? $signed(5'sh1) : $signed(_GEN_15); // @[Filter.scala 125:36]
  wire [4:0] _GEN_17 = _GEN_24715 & _GEN_24708 ? $signed(5'sh1) : $signed(_GEN_16); // @[Filter.scala 125:36]
  wire [4:0] _GEN_18 = _GEN_24715 & _GEN_24710 ? $signed(5'sh1) : $signed(_GEN_17); // @[Filter.scala 125:36]
  wire [4:0] _GEN_19 = _GEN_24715 & _GEN_24712 ? $signed(5'sh1) : $signed(_GEN_18); // @[Filter.scala 125:36]
  wire [4:0] _GEN_20 = _GEN_24715 & _GEN_24714 ? $signed(5'sh1) : $signed(_GEN_19); // @[Filter.scala 125:36]
  wire  _GEN_24733 = 3'h2 == io_SPI_filterIndex[2:0]; // @[Filter.scala 125:36]
  wire [4:0] _GEN_21 = _GEN_24733 & _GEN_24716 ? $signed(5'sh1) : $signed(_GEN_20); // @[Filter.scala 125:36]
  wire [4:0] _GEN_22 = _GEN_24733 & _GEN_24718 ? $signed(5'sh2) : $signed(_GEN_21); // @[Filter.scala 125:36]
  wire [4:0] _GEN_23 = _GEN_24733 & _GEN_24720 ? $signed(5'sh1) : $signed(_GEN_22); // @[Filter.scala 125:36]
  wire [4:0] _GEN_24 = _GEN_24733 & _GEN_24722 ? $signed(5'sh2) : $signed(_GEN_23); // @[Filter.scala 125:36]
  wire [4:0] _GEN_25 = _GEN_24733 & _GEN_24706 ? $signed(5'sh4) : $signed(_GEN_24); // @[Filter.scala 125:36]
  wire [4:0] _GEN_26 = _GEN_24733 & _GEN_24708 ? $signed(5'sh2) : $signed(_GEN_25); // @[Filter.scala 125:36]
  wire [4:0] _GEN_27 = _GEN_24733 & _GEN_24710 ? $signed(5'sh1) : $signed(_GEN_26); // @[Filter.scala 125:36]
  wire [4:0] _GEN_28 = _GEN_24733 & _GEN_24712 ? $signed(5'sh2) : $signed(_GEN_27); // @[Filter.scala 125:36]
  wire [4:0] _GEN_29 = _GEN_24733 & _GEN_24714 ? $signed(5'sh1) : $signed(_GEN_28); // @[Filter.scala 125:36]
  wire  _GEN_24751 = 3'h3 == io_SPI_filterIndex[2:0]; // @[Filter.scala 125:36]
  wire [4:0] _GEN_30 = _GEN_24751 & _GEN_24716 ? $signed(5'sh0) : $signed(_GEN_29); // @[Filter.scala 125:36]
  wire [4:0] _GEN_31 = _GEN_24751 & _GEN_24718 ? $signed(-5'sh1) : $signed(_GEN_30); // @[Filter.scala 125:36]
  wire [4:0] _GEN_32 = _GEN_24751 & _GEN_24720 ? $signed(5'sh0) : $signed(_GEN_31); // @[Filter.scala 125:36]
  wire [4:0] _GEN_33 = _GEN_24751 & _GEN_24722 ? $signed(-5'sh1) : $signed(_GEN_32); // @[Filter.scala 125:36]
  wire [4:0] _GEN_34 = _GEN_24751 & _GEN_24706 ? $signed(5'sh4) : $signed(_GEN_33); // @[Filter.scala 125:36]
  wire [4:0] _GEN_35 = _GEN_24751 & _GEN_24708 ? $signed(-5'sh1) : $signed(_GEN_34); // @[Filter.scala 125:36]
  wire [4:0] _GEN_36 = _GEN_24751 & _GEN_24710 ? $signed(5'sh0) : $signed(_GEN_35); // @[Filter.scala 125:36]
  wire [4:0] _GEN_37 = _GEN_24751 & _GEN_24712 ? $signed(-5'sh1) : $signed(_GEN_36); // @[Filter.scala 125:36]
  wire [4:0] _GEN_38 = _GEN_24751 & _GEN_24714 ? $signed(5'sh0) : $signed(_GEN_37); // @[Filter.scala 125:36]
  wire  _GEN_24769 = 3'h4 == io_SPI_filterIndex[2:0]; // @[Filter.scala 125:36]
  wire [4:0] _GEN_39 = _GEN_24769 & _GEN_24716 ? $signed(-5'sh1) : $signed(_GEN_38); // @[Filter.scala 125:36]
  wire [4:0] _GEN_40 = _GEN_24769 & _GEN_24718 ? $signed(-5'sh1) : $signed(_GEN_39); // @[Filter.scala 125:36]
  wire [4:0] _GEN_41 = _GEN_24769 & _GEN_24720 ? $signed(-5'sh1) : $signed(_GEN_40); // @[Filter.scala 125:36]
  wire [4:0] _GEN_42 = _GEN_24769 & _GEN_24722 ? $signed(-5'sh1) : $signed(_GEN_41); // @[Filter.scala 125:36]
  wire [4:0] _GEN_43 = _GEN_24769 & _GEN_24706 ? $signed(5'sh8) : $signed(_GEN_42); // @[Filter.scala 125:36]
  wire [4:0] _GEN_44 = _GEN_24769 & _GEN_24708 ? $signed(-5'sh1) : $signed(_GEN_43); // @[Filter.scala 125:36]
  wire [4:0] _GEN_45 = _GEN_24769 & _GEN_24710 ? $signed(-5'sh1) : $signed(_GEN_44); // @[Filter.scala 125:36]
  wire [4:0] _GEN_46 = _GEN_24769 & _GEN_24712 ? $signed(-5'sh1) : $signed(_GEN_45); // @[Filter.scala 125:36]
  wire [4:0] _GEN_47 = _GEN_24769 & _GEN_24714 ? $signed(-5'sh1) : $signed(_GEN_46); // @[Filter.scala 125:36]
  wire  _GEN_24787 = 3'h5 == io_SPI_filterIndex[2:0]; // @[Filter.scala 125:36]
  wire [4:0] _GEN_48 = _GEN_24787 & _GEN_24716 ? $signed(5'sh0) : $signed(_GEN_47); // @[Filter.scala 125:36]
  wire [4:0] _GEN_49 = _GEN_24787 & _GEN_24718 ? $signed(-5'sh1) : $signed(_GEN_48); // @[Filter.scala 125:36]
  wire [4:0] _GEN_50 = _GEN_24787 & _GEN_24720 ? $signed(5'sh0) : $signed(_GEN_49); // @[Filter.scala 125:36]
  wire [4:0] _GEN_51 = _GEN_24787 & _GEN_24722 ? $signed(-5'sh1) : $signed(_GEN_50); // @[Filter.scala 125:36]
  wire [4:0] _GEN_52 = _GEN_24787 & _GEN_24706 ? $signed(5'sh5) : $signed(_GEN_51); // @[Filter.scala 125:36]
  wire [4:0] _GEN_53 = _GEN_24787 & _GEN_24708 ? $signed(-5'sh1) : $signed(_GEN_52); // @[Filter.scala 125:36]
  wire [4:0] _GEN_54 = _GEN_24787 & _GEN_24710 ? $signed(5'sh0) : $signed(_GEN_53); // @[Filter.scala 125:36]
  wire [4:0] _GEN_55 = _GEN_24787 & _GEN_24712 ? $signed(-5'sh1) : $signed(_GEN_54); // @[Filter.scala 125:36]
  reg [1:0] imageCounterX; // @[Counter.scala 29:33]
  wire  imageCounterXReset = imageCounterX == 2'h2; // @[Counter.scala 38:24]
  wire [1:0] _T_19 = imageCounterX + 2'h1; // @[Counter.scala 39:22]
  reg [1:0] imageCounterY; // @[Counter.scala 29:33]
  wire  _T_20 = imageCounterY == 2'h2; // @[Counter.scala 38:24]
  wire [1:0] _T_22 = imageCounterY + 2'h1; // @[Counter.scala 39:22]
  reg [31:0] pixelIndex; // @[Filter.scala 130:29]
  wire [32:0] _T_23 = {{1'd0}, pixelIndex}; // @[Filter.scala 133:29]
  wire [31:0] _T_25 = _T_23[31:0] / 32'h40; // @[Filter.scala 133:36]
  wire [31:0] _GEN_24805 = {{30'd0}, imageCounterX}; // @[Filter.scala 133:51]
  wire [31:0] _T_27 = _T_25 + _GEN_24805; // @[Filter.scala 133:51]
  wire [31:0] _T_29 = _T_27 - 32'h1; // @[Filter.scala 133:67]
  wire [31:0] _GEN_0 = _T_23[31:0] % 32'h40; // @[Filter.scala 134:36]
  wire [6:0] _T_32 = _GEN_0[6:0]; // @[Filter.scala 134:36]
  wire [6:0] _GEN_24806 = {{5'd0}, imageCounterY}; // @[Filter.scala 134:51]
  wire [6:0] _T_34 = _T_32 + _GEN_24806; // @[Filter.scala 134:51]
  wire [6:0] _T_36 = _T_34 - 7'h1; // @[Filter.scala 134:67]
  wire  _T_38 = _T_29 >= 32'h40; // @[Filter.scala 135:27]
  wire  _T_42 = _T_36 >= 7'h30; // @[Filter.scala 135:59]
  wire  _T_43 = _T_38 | _T_42; // @[Filter.scala 135:54]
  wire [13:0] _T_44 = _T_36 * 7'h40; // @[Filter.scala 138:57]
  wire [31:0] _GEN_24807 = {{18'd0}, _T_44}; // @[Filter.scala 138:72]
  wire [31:0] _T_46 = _GEN_24807 + _T_29; // @[Filter.scala 138:72]
  wire [3:0] _GEN_75 = 12'hc == _T_46[11:0] ? image_12 : 4'h0; // @[Filter.scala 138:46]
  wire [3:0] _GEN_76 = 12'hd == _T_46[11:0] ? 4'h0 : _GEN_75; // @[Filter.scala 138:46]
  wire [3:0] _GEN_77 = 12'he == _T_46[11:0] ? image_14 : _GEN_76; // @[Filter.scala 138:46]
  wire [3:0] _GEN_78 = 12'hf == _T_46[11:0] ? image_15 : _GEN_77; // @[Filter.scala 138:46]
  wire [3:0] _GEN_79 = 12'h10 == _T_46[11:0] ? image_16 : _GEN_78; // @[Filter.scala 138:46]
  wire [3:0] _GEN_80 = 12'h11 == _T_46[11:0] ? image_17 : _GEN_79; // @[Filter.scala 138:46]
  wire [3:0] _GEN_81 = 12'h12 == _T_46[11:0] ? image_18 : _GEN_80; // @[Filter.scala 138:46]
  wire [3:0] _GEN_82 = 12'h13 == _T_46[11:0] ? image_19 : _GEN_81; // @[Filter.scala 138:46]
  wire [3:0] _GEN_83 = 12'h14 == _T_46[11:0] ? image_20 : _GEN_82; // @[Filter.scala 138:46]
  wire [3:0] _GEN_84 = 12'h15 == _T_46[11:0] ? image_21 : _GEN_83; // @[Filter.scala 138:46]
  wire [3:0] _GEN_85 = 12'h16 == _T_46[11:0] ? image_22 : _GEN_84; // @[Filter.scala 138:46]
  wire [3:0] _GEN_86 = 12'h17 == _T_46[11:0] ? image_23 : _GEN_85; // @[Filter.scala 138:46]
  wire [3:0] _GEN_87 = 12'h18 == _T_46[11:0] ? 4'h0 : _GEN_86; // @[Filter.scala 138:46]
  wire [3:0] _GEN_88 = 12'h19 == _T_46[11:0] ? 4'h0 : _GEN_87; // @[Filter.scala 138:46]
  wire [3:0] _GEN_89 = 12'h1a == _T_46[11:0] ? 4'h0 : _GEN_88; // @[Filter.scala 138:46]
  wire [3:0] _GEN_90 = 12'h1b == _T_46[11:0] ? 4'h0 : _GEN_89; // @[Filter.scala 138:46]
  wire [3:0] _GEN_91 = 12'h1c == _T_46[11:0] ? 4'h0 : _GEN_90; // @[Filter.scala 138:46]
  wire [3:0] _GEN_92 = 12'h1d == _T_46[11:0] ? 4'h0 : _GEN_91; // @[Filter.scala 138:46]
  wire [3:0] _GEN_93 = 12'h1e == _T_46[11:0] ? 4'h0 : _GEN_92; // @[Filter.scala 138:46]
  wire [3:0] _GEN_94 = 12'h1f == _T_46[11:0] ? 4'h0 : _GEN_93; // @[Filter.scala 138:46]
  wire [3:0] _GEN_95 = 12'h20 == _T_46[11:0] ? 4'h0 : _GEN_94; // @[Filter.scala 138:46]
  wire [3:0] _GEN_96 = 12'h21 == _T_46[11:0] ? 4'h0 : _GEN_95; // @[Filter.scala 138:46]
  wire [3:0] _GEN_97 = 12'h22 == _T_46[11:0] ? 4'h0 : _GEN_96; // @[Filter.scala 138:46]
  wire [3:0] _GEN_98 = 12'h23 == _T_46[11:0] ? image_35 : _GEN_97; // @[Filter.scala 138:46]
  wire [3:0] _GEN_99 = 12'h24 == _T_46[11:0] ? image_36 : _GEN_98; // @[Filter.scala 138:46]
  wire [3:0] _GEN_100 = 12'h25 == _T_46[11:0] ? image_37 : _GEN_99; // @[Filter.scala 138:46]
  wire [3:0] _GEN_101 = 12'h26 == _T_46[11:0] ? image_38 : _GEN_100; // @[Filter.scala 138:46]
  wire [3:0] _GEN_102 = 12'h27 == _T_46[11:0] ? image_39 : _GEN_101; // @[Filter.scala 138:46]
  wire [3:0] _GEN_103 = 12'h28 == _T_46[11:0] ? image_40 : _GEN_102; // @[Filter.scala 138:46]
  wire [3:0] _GEN_104 = 12'h29 == _T_46[11:0] ? image_41 : _GEN_103; // @[Filter.scala 138:46]
  wire [3:0] _GEN_105 = 12'h2a == _T_46[11:0] ? image_42 : _GEN_104; // @[Filter.scala 138:46]
  wire [3:0] _GEN_106 = 12'h2b == _T_46[11:0] ? 4'h0 : _GEN_105; // @[Filter.scala 138:46]
  wire [3:0] _GEN_107 = 12'h2c == _T_46[11:0] ? 4'h0 : _GEN_106; // @[Filter.scala 138:46]
  wire [3:0] _GEN_108 = 12'h2d == _T_46[11:0] ? 4'h0 : _GEN_107; // @[Filter.scala 138:46]
  wire [3:0] _GEN_109 = 12'h2e == _T_46[11:0] ? 4'h0 : _GEN_108; // @[Filter.scala 138:46]
  wire [3:0] _GEN_110 = 12'h2f == _T_46[11:0] ? 4'h0 : _GEN_109; // @[Filter.scala 138:46]
  wire [3:0] _GEN_111 = 12'h30 == _T_46[11:0] ? 4'h0 : _GEN_110; // @[Filter.scala 138:46]
  wire [3:0] _GEN_112 = 12'h31 == _T_46[11:0] ? 4'h0 : _GEN_111; // @[Filter.scala 138:46]
  wire [3:0] _GEN_113 = 12'h32 == _T_46[11:0] ? 4'h0 : _GEN_112; // @[Filter.scala 138:46]
  wire [3:0] _GEN_114 = 12'h33 == _T_46[11:0] ? 4'h0 : _GEN_113; // @[Filter.scala 138:46]
  wire [3:0] _GEN_115 = 12'h34 == _T_46[11:0] ? 4'h0 : _GEN_114; // @[Filter.scala 138:46]
  wire [3:0] _GEN_116 = 12'h35 == _T_46[11:0] ? 4'h0 : _GEN_115; // @[Filter.scala 138:46]
  wire [3:0] _GEN_117 = 12'h36 == _T_46[11:0] ? 4'h0 : _GEN_116; // @[Filter.scala 138:46]
  wire [3:0] _GEN_118 = 12'h37 == _T_46[11:0] ? 4'h0 : _GEN_117; // @[Filter.scala 138:46]
  wire [3:0] _GEN_119 = 12'h38 == _T_46[11:0] ? 4'h0 : _GEN_118; // @[Filter.scala 138:46]
  wire [3:0] _GEN_120 = 12'h39 == _T_46[11:0] ? 4'h0 : _GEN_119; // @[Filter.scala 138:46]
  wire [3:0] _GEN_121 = 12'h3a == _T_46[11:0] ? 4'h0 : _GEN_120; // @[Filter.scala 138:46]
  wire [3:0] _GEN_122 = 12'h3b == _T_46[11:0] ? 4'h0 : _GEN_121; // @[Filter.scala 138:46]
  wire [3:0] _GEN_123 = 12'h3c == _T_46[11:0] ? 4'h0 : _GEN_122; // @[Filter.scala 138:46]
  wire [3:0] _GEN_124 = 12'h3d == _T_46[11:0] ? 4'h0 : _GEN_123; // @[Filter.scala 138:46]
  wire [3:0] _GEN_125 = 12'h3e == _T_46[11:0] ? 4'h0 : _GEN_124; // @[Filter.scala 138:46]
  wire [3:0] _GEN_126 = 12'h3f == _T_46[11:0] ? 4'h0 : _GEN_125; // @[Filter.scala 138:46]
  wire [3:0] _GEN_127 = 12'h40 == _T_46[11:0] ? 4'h0 : _GEN_126; // @[Filter.scala 138:46]
  wire [3:0] _GEN_128 = 12'h41 == _T_46[11:0] ? 4'h0 : _GEN_127; // @[Filter.scala 138:46]
  wire [3:0] _GEN_129 = 12'h42 == _T_46[11:0] ? 4'h0 : _GEN_128; // @[Filter.scala 138:46]
  wire [3:0] _GEN_130 = 12'h43 == _T_46[11:0] ? 4'h0 : _GEN_129; // @[Filter.scala 138:46]
  wire [3:0] _GEN_131 = 12'h44 == _T_46[11:0] ? 4'h0 : _GEN_130; // @[Filter.scala 138:46]
  wire [3:0] _GEN_132 = 12'h45 == _T_46[11:0] ? 4'h0 : _GEN_131; // @[Filter.scala 138:46]
  wire [3:0] _GEN_133 = 12'h46 == _T_46[11:0] ? 4'h0 : _GEN_132; // @[Filter.scala 138:46]
  wire [3:0] _GEN_134 = 12'h47 == _T_46[11:0] ? 4'h0 : _GEN_133; // @[Filter.scala 138:46]
  wire [3:0] _GEN_135 = 12'h48 == _T_46[11:0] ? 4'h0 : _GEN_134; // @[Filter.scala 138:46]
  wire [3:0] _GEN_136 = 12'h49 == _T_46[11:0] ? 4'h0 : _GEN_135; // @[Filter.scala 138:46]
  wire [3:0] _GEN_137 = 12'h4a == _T_46[11:0] ? 4'h0 : _GEN_136; // @[Filter.scala 138:46]
  wire [3:0] _GEN_138 = 12'h4b == _T_46[11:0] ? image_75 : _GEN_137; // @[Filter.scala 138:46]
  wire [3:0] _GEN_139 = 12'h4c == _T_46[11:0] ? image_76 : _GEN_138; // @[Filter.scala 138:46]
  wire [3:0] _GEN_140 = 12'h4d == _T_46[11:0] ? image_77 : _GEN_139; // @[Filter.scala 138:46]
  wire [3:0] _GEN_141 = 12'h4e == _T_46[11:0] ? image_78 : _GEN_140; // @[Filter.scala 138:46]
  wire [3:0] _GEN_142 = 12'h4f == _T_46[11:0] ? image_79 : _GEN_141; // @[Filter.scala 138:46]
  wire [3:0] _GEN_143 = 12'h50 == _T_46[11:0] ? image_80 : _GEN_142; // @[Filter.scala 138:46]
  wire [3:0] _GEN_144 = 12'h51 == _T_46[11:0] ? image_81 : _GEN_143; // @[Filter.scala 138:46]
  wire [3:0] _GEN_145 = 12'h52 == _T_46[11:0] ? image_82 : _GEN_144; // @[Filter.scala 138:46]
  wire [3:0] _GEN_146 = 12'h53 == _T_46[11:0] ? image_83 : _GEN_145; // @[Filter.scala 138:46]
  wire [3:0] _GEN_147 = 12'h54 == _T_46[11:0] ? image_84 : _GEN_146; // @[Filter.scala 138:46]
  wire [3:0] _GEN_148 = 12'h55 == _T_46[11:0] ? image_85 : _GEN_147; // @[Filter.scala 138:46]
  wire [3:0] _GEN_149 = 12'h56 == _T_46[11:0] ? image_86 : _GEN_148; // @[Filter.scala 138:46]
  wire [3:0] _GEN_150 = 12'h57 == _T_46[11:0] ? image_87 : _GEN_149; // @[Filter.scala 138:46]
  wire [3:0] _GEN_151 = 12'h58 == _T_46[11:0] ? image_88 : _GEN_150; // @[Filter.scala 138:46]
  wire [3:0] _GEN_152 = 12'h59 == _T_46[11:0] ? image_89 : _GEN_151; // @[Filter.scala 138:46]
  wire [3:0] _GEN_153 = 12'h5a == _T_46[11:0] ? image_90 : _GEN_152; // @[Filter.scala 138:46]
  wire [3:0] _GEN_154 = 12'h5b == _T_46[11:0] ? 4'h0 : _GEN_153; // @[Filter.scala 138:46]
  wire [3:0] _GEN_155 = 12'h5c == _T_46[11:0] ? 4'h0 : _GEN_154; // @[Filter.scala 138:46]
  wire [3:0] _GEN_156 = 12'h5d == _T_46[11:0] ? image_93 : _GEN_155; // @[Filter.scala 138:46]
  wire [3:0] _GEN_157 = 12'h5e == _T_46[11:0] ? 4'h0 : _GEN_156; // @[Filter.scala 138:46]
  wire [3:0] _GEN_158 = 12'h5f == _T_46[11:0] ? image_95 : _GEN_157; // @[Filter.scala 138:46]
  wire [3:0] _GEN_159 = 12'h60 == _T_46[11:0] ? image_96 : _GEN_158; // @[Filter.scala 138:46]
  wire [3:0] _GEN_160 = 12'h61 == _T_46[11:0] ? image_97 : _GEN_159; // @[Filter.scala 138:46]
  wire [3:0] _GEN_161 = 12'h62 == _T_46[11:0] ? image_98 : _GEN_160; // @[Filter.scala 138:46]
  wire [3:0] _GEN_162 = 12'h63 == _T_46[11:0] ? image_99 : _GEN_161; // @[Filter.scala 138:46]
  wire [3:0] _GEN_163 = 12'h64 == _T_46[11:0] ? image_100 : _GEN_162; // @[Filter.scala 138:46]
  wire [3:0] _GEN_164 = 12'h65 == _T_46[11:0] ? image_101 : _GEN_163; // @[Filter.scala 138:46]
  wire [3:0] _GEN_165 = 12'h66 == _T_46[11:0] ? image_102 : _GEN_164; // @[Filter.scala 138:46]
  wire [3:0] _GEN_166 = 12'h67 == _T_46[11:0] ? image_103 : _GEN_165; // @[Filter.scala 138:46]
  wire [3:0] _GEN_167 = 12'h68 == _T_46[11:0] ? image_104 : _GEN_166; // @[Filter.scala 138:46]
  wire [3:0] _GEN_168 = 12'h69 == _T_46[11:0] ? image_105 : _GEN_167; // @[Filter.scala 138:46]
  wire [3:0] _GEN_169 = 12'h6a == _T_46[11:0] ? image_106 : _GEN_168; // @[Filter.scala 138:46]
  wire [3:0] _GEN_170 = 12'h6b == _T_46[11:0] ? image_107 : _GEN_169; // @[Filter.scala 138:46]
  wire [3:0] _GEN_171 = 12'h6c == _T_46[11:0] ? image_108 : _GEN_170; // @[Filter.scala 138:46]
  wire [3:0] _GEN_172 = 12'h6d == _T_46[11:0] ? 4'h0 : _GEN_171; // @[Filter.scala 138:46]
  wire [3:0] _GEN_173 = 12'h6e == _T_46[11:0] ? 4'h0 : _GEN_172; // @[Filter.scala 138:46]
  wire [3:0] _GEN_174 = 12'h6f == _T_46[11:0] ? 4'h0 : _GEN_173; // @[Filter.scala 138:46]
  wire [3:0] _GEN_175 = 12'h70 == _T_46[11:0] ? 4'h0 : _GEN_174; // @[Filter.scala 138:46]
  wire [3:0] _GEN_176 = 12'h71 == _T_46[11:0] ? 4'h0 : _GEN_175; // @[Filter.scala 138:46]
  wire [3:0] _GEN_177 = 12'h72 == _T_46[11:0] ? 4'h0 : _GEN_176; // @[Filter.scala 138:46]
  wire [3:0] _GEN_178 = 12'h73 == _T_46[11:0] ? 4'h0 : _GEN_177; // @[Filter.scala 138:46]
  wire [3:0] _GEN_179 = 12'h74 == _T_46[11:0] ? 4'h0 : _GEN_178; // @[Filter.scala 138:46]
  wire [3:0] _GEN_180 = 12'h75 == _T_46[11:0] ? 4'h0 : _GEN_179; // @[Filter.scala 138:46]
  wire [3:0] _GEN_181 = 12'h76 == _T_46[11:0] ? 4'h0 : _GEN_180; // @[Filter.scala 138:46]
  wire [3:0] _GEN_182 = 12'h77 == _T_46[11:0] ? 4'h0 : _GEN_181; // @[Filter.scala 138:46]
  wire [3:0] _GEN_183 = 12'h78 == _T_46[11:0] ? 4'h0 : _GEN_182; // @[Filter.scala 138:46]
  wire [3:0] _GEN_184 = 12'h79 == _T_46[11:0] ? 4'h0 : _GEN_183; // @[Filter.scala 138:46]
  wire [3:0] _GEN_185 = 12'h7a == _T_46[11:0] ? 4'h0 : _GEN_184; // @[Filter.scala 138:46]
  wire [3:0] _GEN_186 = 12'h7b == _T_46[11:0] ? 4'h0 : _GEN_185; // @[Filter.scala 138:46]
  wire [3:0] _GEN_187 = 12'h7c == _T_46[11:0] ? 4'h0 : _GEN_186; // @[Filter.scala 138:46]
  wire [3:0] _GEN_188 = 12'h7d == _T_46[11:0] ? 4'h0 : _GEN_187; // @[Filter.scala 138:46]
  wire [3:0] _GEN_189 = 12'h7e == _T_46[11:0] ? 4'h0 : _GEN_188; // @[Filter.scala 138:46]
  wire [3:0] _GEN_190 = 12'h7f == _T_46[11:0] ? 4'h0 : _GEN_189; // @[Filter.scala 138:46]
  wire [3:0] _GEN_191 = 12'h80 == _T_46[11:0] ? 4'h0 : _GEN_190; // @[Filter.scala 138:46]
  wire [3:0] _GEN_192 = 12'h81 == _T_46[11:0] ? 4'h0 : _GEN_191; // @[Filter.scala 138:46]
  wire [3:0] _GEN_193 = 12'h82 == _T_46[11:0] ? 4'h0 : _GEN_192; // @[Filter.scala 138:46]
  wire [3:0] _GEN_194 = 12'h83 == _T_46[11:0] ? 4'h0 : _GEN_193; // @[Filter.scala 138:46]
  wire [3:0] _GEN_195 = 12'h84 == _T_46[11:0] ? 4'h0 : _GEN_194; // @[Filter.scala 138:46]
  wire [3:0] _GEN_196 = 12'h85 == _T_46[11:0] ? 4'h0 : _GEN_195; // @[Filter.scala 138:46]
  wire [3:0] _GEN_197 = 12'h86 == _T_46[11:0] ? 4'h0 : _GEN_196; // @[Filter.scala 138:46]
  wire [3:0] _GEN_198 = 12'h87 == _T_46[11:0] ? 4'h0 : _GEN_197; // @[Filter.scala 138:46]
  wire [3:0] _GEN_199 = 12'h88 == _T_46[11:0] ? image_136 : _GEN_198; // @[Filter.scala 138:46]
  wire [3:0] _GEN_200 = 12'h89 == _T_46[11:0] ? image_137 : _GEN_199; // @[Filter.scala 138:46]
  wire [3:0] _GEN_201 = 12'h8a == _T_46[11:0] ? image_138 : _GEN_200; // @[Filter.scala 138:46]
  wire [3:0] _GEN_202 = 12'h8b == _T_46[11:0] ? image_139 : _GEN_201; // @[Filter.scala 138:46]
  wire [3:0] _GEN_203 = 12'h8c == _T_46[11:0] ? image_140 : _GEN_202; // @[Filter.scala 138:46]
  wire [3:0] _GEN_204 = 12'h8d == _T_46[11:0] ? image_141 : _GEN_203; // @[Filter.scala 138:46]
  wire [3:0] _GEN_205 = 12'h8e == _T_46[11:0] ? image_142 : _GEN_204; // @[Filter.scala 138:46]
  wire [3:0] _GEN_206 = 12'h8f == _T_46[11:0] ? image_143 : _GEN_205; // @[Filter.scala 138:46]
  wire [3:0] _GEN_207 = 12'h90 == _T_46[11:0] ? image_144 : _GEN_206; // @[Filter.scala 138:46]
  wire [3:0] _GEN_208 = 12'h91 == _T_46[11:0] ? image_145 : _GEN_207; // @[Filter.scala 138:46]
  wire [3:0] _GEN_209 = 12'h92 == _T_46[11:0] ? image_146 : _GEN_208; // @[Filter.scala 138:46]
  wire [3:0] _GEN_210 = 12'h93 == _T_46[11:0] ? image_147 : _GEN_209; // @[Filter.scala 138:46]
  wire [3:0] _GEN_211 = 12'h94 == _T_46[11:0] ? image_148 : _GEN_210; // @[Filter.scala 138:46]
  wire [3:0] _GEN_212 = 12'h95 == _T_46[11:0] ? image_149 : _GEN_211; // @[Filter.scala 138:46]
  wire [3:0] _GEN_213 = 12'h96 == _T_46[11:0] ? image_150 : _GEN_212; // @[Filter.scala 138:46]
  wire [3:0] _GEN_214 = 12'h97 == _T_46[11:0] ? image_151 : _GEN_213; // @[Filter.scala 138:46]
  wire [3:0] _GEN_215 = 12'h98 == _T_46[11:0] ? image_152 : _GEN_214; // @[Filter.scala 138:46]
  wire [3:0] _GEN_216 = 12'h99 == _T_46[11:0] ? image_153 : _GEN_215; // @[Filter.scala 138:46]
  wire [3:0] _GEN_217 = 12'h9a == _T_46[11:0] ? image_154 : _GEN_216; // @[Filter.scala 138:46]
  wire [3:0] _GEN_218 = 12'h9b == _T_46[11:0] ? image_155 : _GEN_217; // @[Filter.scala 138:46]
  wire [3:0] _GEN_219 = 12'h9c == _T_46[11:0] ? 4'h0 : _GEN_218; // @[Filter.scala 138:46]
  wire [3:0] _GEN_220 = 12'h9d == _T_46[11:0] ? image_157 : _GEN_219; // @[Filter.scala 138:46]
  wire [3:0] _GEN_221 = 12'h9e == _T_46[11:0] ? image_158 : _GEN_220; // @[Filter.scala 138:46]
  wire [3:0] _GEN_222 = 12'h9f == _T_46[11:0] ? image_159 : _GEN_221; // @[Filter.scala 138:46]
  wire [3:0] _GEN_223 = 12'ha0 == _T_46[11:0] ? image_160 : _GEN_222; // @[Filter.scala 138:46]
  wire [3:0] _GEN_224 = 12'ha1 == _T_46[11:0] ? image_161 : _GEN_223; // @[Filter.scala 138:46]
  wire [3:0] _GEN_225 = 12'ha2 == _T_46[11:0] ? image_162 : _GEN_224; // @[Filter.scala 138:46]
  wire [3:0] _GEN_226 = 12'ha3 == _T_46[11:0] ? image_163 : _GEN_225; // @[Filter.scala 138:46]
  wire [3:0] _GEN_227 = 12'ha4 == _T_46[11:0] ? image_164 : _GEN_226; // @[Filter.scala 138:46]
  wire [3:0] _GEN_228 = 12'ha5 == _T_46[11:0] ? image_165 : _GEN_227; // @[Filter.scala 138:46]
  wire [3:0] _GEN_229 = 12'ha6 == _T_46[11:0] ? image_166 : _GEN_228; // @[Filter.scala 138:46]
  wire [3:0] _GEN_230 = 12'ha7 == _T_46[11:0] ? image_167 : _GEN_229; // @[Filter.scala 138:46]
  wire [3:0] _GEN_231 = 12'ha8 == _T_46[11:0] ? image_168 : _GEN_230; // @[Filter.scala 138:46]
  wire [3:0] _GEN_232 = 12'ha9 == _T_46[11:0] ? image_169 : _GEN_231; // @[Filter.scala 138:46]
  wire [3:0] _GEN_233 = 12'haa == _T_46[11:0] ? image_170 : _GEN_232; // @[Filter.scala 138:46]
  wire [3:0] _GEN_234 = 12'hab == _T_46[11:0] ? image_171 : _GEN_233; // @[Filter.scala 138:46]
  wire [3:0] _GEN_235 = 12'hac == _T_46[11:0] ? image_172 : _GEN_234; // @[Filter.scala 138:46]
  wire [3:0] _GEN_236 = 12'had == _T_46[11:0] ? image_173 : _GEN_235; // @[Filter.scala 138:46]
  wire [3:0] _GEN_237 = 12'hae == _T_46[11:0] ? image_174 : _GEN_236; // @[Filter.scala 138:46]
  wire [3:0] _GEN_238 = 12'haf == _T_46[11:0] ? image_175 : _GEN_237; // @[Filter.scala 138:46]
  wire [3:0] _GEN_239 = 12'hb0 == _T_46[11:0] ? image_176 : _GEN_238; // @[Filter.scala 138:46]
  wire [3:0] _GEN_240 = 12'hb1 == _T_46[11:0] ? image_177 : _GEN_239; // @[Filter.scala 138:46]
  wire [3:0] _GEN_241 = 12'hb2 == _T_46[11:0] ? image_178 : _GEN_240; // @[Filter.scala 138:46]
  wire [3:0] _GEN_242 = 12'hb3 == _T_46[11:0] ? image_179 : _GEN_241; // @[Filter.scala 138:46]
  wire [3:0] _GEN_243 = 12'hb4 == _T_46[11:0] ? 4'h0 : _GEN_242; // @[Filter.scala 138:46]
  wire [3:0] _GEN_244 = 12'hb5 == _T_46[11:0] ? 4'h0 : _GEN_243; // @[Filter.scala 138:46]
  wire [3:0] _GEN_245 = 12'hb6 == _T_46[11:0] ? 4'h0 : _GEN_244; // @[Filter.scala 138:46]
  wire [3:0] _GEN_246 = 12'hb7 == _T_46[11:0] ? 4'h0 : _GEN_245; // @[Filter.scala 138:46]
  wire [3:0] _GEN_247 = 12'hb8 == _T_46[11:0] ? 4'h0 : _GEN_246; // @[Filter.scala 138:46]
  wire [3:0] _GEN_248 = 12'hb9 == _T_46[11:0] ? 4'h0 : _GEN_247; // @[Filter.scala 138:46]
  wire [3:0] _GEN_249 = 12'hba == _T_46[11:0] ? 4'h0 : _GEN_248; // @[Filter.scala 138:46]
  wire [3:0] _GEN_250 = 12'hbb == _T_46[11:0] ? 4'h0 : _GEN_249; // @[Filter.scala 138:46]
  wire [3:0] _GEN_251 = 12'hbc == _T_46[11:0] ? 4'h0 : _GEN_250; // @[Filter.scala 138:46]
  wire [3:0] _GEN_252 = 12'hbd == _T_46[11:0] ? 4'h0 : _GEN_251; // @[Filter.scala 138:46]
  wire [3:0] _GEN_253 = 12'hbe == _T_46[11:0] ? 4'h0 : _GEN_252; // @[Filter.scala 138:46]
  wire [3:0] _GEN_254 = 12'hbf == _T_46[11:0] ? 4'h0 : _GEN_253; // @[Filter.scala 138:46]
  wire [3:0] _GEN_255 = 12'hc0 == _T_46[11:0] ? 4'h0 : _GEN_254; // @[Filter.scala 138:46]
  wire [3:0] _GEN_256 = 12'hc1 == _T_46[11:0] ? 4'h0 : _GEN_255; // @[Filter.scala 138:46]
  wire [3:0] _GEN_257 = 12'hc2 == _T_46[11:0] ? 4'h0 : _GEN_256; // @[Filter.scala 138:46]
  wire [3:0] _GEN_258 = 12'hc3 == _T_46[11:0] ? 4'h0 : _GEN_257; // @[Filter.scala 138:46]
  wire [3:0] _GEN_259 = 12'hc4 == _T_46[11:0] ? 4'h0 : _GEN_258; // @[Filter.scala 138:46]
  wire [3:0] _GEN_260 = 12'hc5 == _T_46[11:0] ? 4'h0 : _GEN_259; // @[Filter.scala 138:46]
  wire [3:0] _GEN_261 = 12'hc6 == _T_46[11:0] ? 4'h0 : _GEN_260; // @[Filter.scala 138:46]
  wire [3:0] _GEN_262 = 12'hc7 == _T_46[11:0] ? image_199 : _GEN_261; // @[Filter.scala 138:46]
  wire [3:0] _GEN_263 = 12'hc8 == _T_46[11:0] ? image_200 : _GEN_262; // @[Filter.scala 138:46]
  wire [3:0] _GEN_264 = 12'hc9 == _T_46[11:0] ? image_201 : _GEN_263; // @[Filter.scala 138:46]
  wire [3:0] _GEN_265 = 12'hca == _T_46[11:0] ? image_202 : _GEN_264; // @[Filter.scala 138:46]
  wire [3:0] _GEN_266 = 12'hcb == _T_46[11:0] ? image_203 : _GEN_265; // @[Filter.scala 138:46]
  wire [3:0] _GEN_267 = 12'hcc == _T_46[11:0] ? image_204 : _GEN_266; // @[Filter.scala 138:46]
  wire [3:0] _GEN_268 = 12'hcd == _T_46[11:0] ? image_205 : _GEN_267; // @[Filter.scala 138:46]
  wire [3:0] _GEN_269 = 12'hce == _T_46[11:0] ? image_206 : _GEN_268; // @[Filter.scala 138:46]
  wire [3:0] _GEN_270 = 12'hcf == _T_46[11:0] ? image_207 : _GEN_269; // @[Filter.scala 138:46]
  wire [3:0] _GEN_271 = 12'hd0 == _T_46[11:0] ? image_208 : _GEN_270; // @[Filter.scala 138:46]
  wire [3:0] _GEN_272 = 12'hd1 == _T_46[11:0] ? image_209 : _GEN_271; // @[Filter.scala 138:46]
  wire [3:0] _GEN_273 = 12'hd2 == _T_46[11:0] ? image_210 : _GEN_272; // @[Filter.scala 138:46]
  wire [3:0] _GEN_274 = 12'hd3 == _T_46[11:0] ? image_211 : _GEN_273; // @[Filter.scala 138:46]
  wire [3:0] _GEN_275 = 12'hd4 == _T_46[11:0] ? image_212 : _GEN_274; // @[Filter.scala 138:46]
  wire [3:0] _GEN_276 = 12'hd5 == _T_46[11:0] ? image_213 : _GEN_275; // @[Filter.scala 138:46]
  wire [3:0] _GEN_277 = 12'hd6 == _T_46[11:0] ? image_214 : _GEN_276; // @[Filter.scala 138:46]
  wire [3:0] _GEN_278 = 12'hd7 == _T_46[11:0] ? image_215 : _GEN_277; // @[Filter.scala 138:46]
  wire [3:0] _GEN_279 = 12'hd8 == _T_46[11:0] ? image_216 : _GEN_278; // @[Filter.scala 138:46]
  wire [3:0] _GEN_280 = 12'hd9 == _T_46[11:0] ? image_217 : _GEN_279; // @[Filter.scala 138:46]
  wire [3:0] _GEN_281 = 12'hda == _T_46[11:0] ? image_218 : _GEN_280; // @[Filter.scala 138:46]
  wire [3:0] _GEN_282 = 12'hdb == _T_46[11:0] ? image_219 : _GEN_281; // @[Filter.scala 138:46]
  wire [3:0] _GEN_283 = 12'hdc == _T_46[11:0] ? image_220 : _GEN_282; // @[Filter.scala 138:46]
  wire [3:0] _GEN_284 = 12'hdd == _T_46[11:0] ? image_221 : _GEN_283; // @[Filter.scala 138:46]
  wire [3:0] _GEN_285 = 12'hde == _T_46[11:0] ? image_222 : _GEN_284; // @[Filter.scala 138:46]
  wire [3:0] _GEN_286 = 12'hdf == _T_46[11:0] ? image_223 : _GEN_285; // @[Filter.scala 138:46]
  wire [3:0] _GEN_287 = 12'he0 == _T_46[11:0] ? image_224 : _GEN_286; // @[Filter.scala 138:46]
  wire [3:0] _GEN_288 = 12'he1 == _T_46[11:0] ? image_225 : _GEN_287; // @[Filter.scala 138:46]
  wire [3:0] _GEN_289 = 12'he2 == _T_46[11:0] ? image_226 : _GEN_288; // @[Filter.scala 138:46]
  wire [3:0] _GEN_290 = 12'he3 == _T_46[11:0] ? image_227 : _GEN_289; // @[Filter.scala 138:46]
  wire [3:0] _GEN_291 = 12'he4 == _T_46[11:0] ? image_228 : _GEN_290; // @[Filter.scala 138:46]
  wire [3:0] _GEN_292 = 12'he5 == _T_46[11:0] ? image_229 : _GEN_291; // @[Filter.scala 138:46]
  wire [3:0] _GEN_293 = 12'he6 == _T_46[11:0] ? image_230 : _GEN_292; // @[Filter.scala 138:46]
  wire [3:0] _GEN_294 = 12'he7 == _T_46[11:0] ? image_231 : _GEN_293; // @[Filter.scala 138:46]
  wire [3:0] _GEN_295 = 12'he8 == _T_46[11:0] ? image_232 : _GEN_294; // @[Filter.scala 138:46]
  wire [3:0] _GEN_296 = 12'he9 == _T_46[11:0] ? image_233 : _GEN_295; // @[Filter.scala 138:46]
  wire [3:0] _GEN_297 = 12'hea == _T_46[11:0] ? image_234 : _GEN_296; // @[Filter.scala 138:46]
  wire [3:0] _GEN_298 = 12'heb == _T_46[11:0] ? image_235 : _GEN_297; // @[Filter.scala 138:46]
  wire [3:0] _GEN_299 = 12'hec == _T_46[11:0] ? image_236 : _GEN_298; // @[Filter.scala 138:46]
  wire [3:0] _GEN_300 = 12'hed == _T_46[11:0] ? image_237 : _GEN_299; // @[Filter.scala 138:46]
  wire [3:0] _GEN_301 = 12'hee == _T_46[11:0] ? image_238 : _GEN_300; // @[Filter.scala 138:46]
  wire [3:0] _GEN_302 = 12'hef == _T_46[11:0] ? image_239 : _GEN_301; // @[Filter.scala 138:46]
  wire [3:0] _GEN_303 = 12'hf0 == _T_46[11:0] ? image_240 : _GEN_302; // @[Filter.scala 138:46]
  wire [3:0] _GEN_304 = 12'hf1 == _T_46[11:0] ? image_241 : _GEN_303; // @[Filter.scala 138:46]
  wire [3:0] _GEN_305 = 12'hf2 == _T_46[11:0] ? image_242 : _GEN_304; // @[Filter.scala 138:46]
  wire [3:0] _GEN_306 = 12'hf3 == _T_46[11:0] ? image_243 : _GEN_305; // @[Filter.scala 138:46]
  wire [3:0] _GEN_307 = 12'hf4 == _T_46[11:0] ? image_244 : _GEN_306; // @[Filter.scala 138:46]
  wire [3:0] _GEN_308 = 12'hf5 == _T_46[11:0] ? image_245 : _GEN_307; // @[Filter.scala 138:46]
  wire [3:0] _GEN_309 = 12'hf6 == _T_46[11:0] ? image_246 : _GEN_308; // @[Filter.scala 138:46]
  wire [3:0] _GEN_310 = 12'hf7 == _T_46[11:0] ? 4'h0 : _GEN_309; // @[Filter.scala 138:46]
  wire [3:0] _GEN_311 = 12'hf8 == _T_46[11:0] ? 4'h0 : _GEN_310; // @[Filter.scala 138:46]
  wire [3:0] _GEN_312 = 12'hf9 == _T_46[11:0] ? 4'h0 : _GEN_311; // @[Filter.scala 138:46]
  wire [3:0] _GEN_313 = 12'hfa == _T_46[11:0] ? 4'h0 : _GEN_312; // @[Filter.scala 138:46]
  wire [3:0] _GEN_314 = 12'hfb == _T_46[11:0] ? 4'h0 : _GEN_313; // @[Filter.scala 138:46]
  wire [3:0] _GEN_315 = 12'hfc == _T_46[11:0] ? 4'h0 : _GEN_314; // @[Filter.scala 138:46]
  wire [3:0] _GEN_316 = 12'hfd == _T_46[11:0] ? 4'h0 : _GEN_315; // @[Filter.scala 138:46]
  wire [3:0] _GEN_317 = 12'hfe == _T_46[11:0] ? 4'h0 : _GEN_316; // @[Filter.scala 138:46]
  wire [3:0] _GEN_318 = 12'hff == _T_46[11:0] ? 4'h0 : _GEN_317; // @[Filter.scala 138:46]
  wire [3:0] _GEN_319 = 12'h100 == _T_46[11:0] ? 4'h0 : _GEN_318; // @[Filter.scala 138:46]
  wire [3:0] _GEN_320 = 12'h101 == _T_46[11:0] ? 4'h0 : _GEN_319; // @[Filter.scala 138:46]
  wire [3:0] _GEN_321 = 12'h102 == _T_46[11:0] ? 4'h0 : _GEN_320; // @[Filter.scala 138:46]
  wire [3:0] _GEN_322 = 12'h103 == _T_46[11:0] ? 4'h0 : _GEN_321; // @[Filter.scala 138:46]
  wire [3:0] _GEN_323 = 12'h104 == _T_46[11:0] ? 4'h0 : _GEN_322; // @[Filter.scala 138:46]
  wire [3:0] _GEN_324 = 12'h105 == _T_46[11:0] ? 4'h0 : _GEN_323; // @[Filter.scala 138:46]
  wire [3:0] _GEN_325 = 12'h106 == _T_46[11:0] ? image_262 : _GEN_324; // @[Filter.scala 138:46]
  wire [3:0] _GEN_326 = 12'h107 == _T_46[11:0] ? image_263 : _GEN_325; // @[Filter.scala 138:46]
  wire [3:0] _GEN_327 = 12'h108 == _T_46[11:0] ? image_264 : _GEN_326; // @[Filter.scala 138:46]
  wire [3:0] _GEN_328 = 12'h109 == _T_46[11:0] ? image_265 : _GEN_327; // @[Filter.scala 138:46]
  wire [3:0] _GEN_329 = 12'h10a == _T_46[11:0] ? image_266 : _GEN_328; // @[Filter.scala 138:46]
  wire [3:0] _GEN_330 = 12'h10b == _T_46[11:0] ? image_267 : _GEN_329; // @[Filter.scala 138:46]
  wire [3:0] _GEN_331 = 12'h10c == _T_46[11:0] ? image_268 : _GEN_330; // @[Filter.scala 138:46]
  wire [3:0] _GEN_332 = 12'h10d == _T_46[11:0] ? image_269 : _GEN_331; // @[Filter.scala 138:46]
  wire [3:0] _GEN_333 = 12'h10e == _T_46[11:0] ? image_270 : _GEN_332; // @[Filter.scala 138:46]
  wire [3:0] _GEN_334 = 12'h10f == _T_46[11:0] ? image_271 : _GEN_333; // @[Filter.scala 138:46]
  wire [3:0] _GEN_335 = 12'h110 == _T_46[11:0] ? image_272 : _GEN_334; // @[Filter.scala 138:46]
  wire [3:0] _GEN_336 = 12'h111 == _T_46[11:0] ? image_273 : _GEN_335; // @[Filter.scala 138:46]
  wire [3:0] _GEN_337 = 12'h112 == _T_46[11:0] ? image_274 : _GEN_336; // @[Filter.scala 138:46]
  wire [3:0] _GEN_338 = 12'h113 == _T_46[11:0] ? image_275 : _GEN_337; // @[Filter.scala 138:46]
  wire [3:0] _GEN_339 = 12'h114 == _T_46[11:0] ? image_276 : _GEN_338; // @[Filter.scala 138:46]
  wire [3:0] _GEN_340 = 12'h115 == _T_46[11:0] ? image_277 : _GEN_339; // @[Filter.scala 138:46]
  wire [3:0] _GEN_341 = 12'h116 == _T_46[11:0] ? image_278 : _GEN_340; // @[Filter.scala 138:46]
  wire [3:0] _GEN_342 = 12'h117 == _T_46[11:0] ? image_279 : _GEN_341; // @[Filter.scala 138:46]
  wire [3:0] _GEN_343 = 12'h118 == _T_46[11:0] ? image_280 : _GEN_342; // @[Filter.scala 138:46]
  wire [3:0] _GEN_344 = 12'h119 == _T_46[11:0] ? image_281 : _GEN_343; // @[Filter.scala 138:46]
  wire [3:0] _GEN_345 = 12'h11a == _T_46[11:0] ? image_282 : _GEN_344; // @[Filter.scala 138:46]
  wire [3:0] _GEN_346 = 12'h11b == _T_46[11:0] ? image_283 : _GEN_345; // @[Filter.scala 138:46]
  wire [3:0] _GEN_347 = 12'h11c == _T_46[11:0] ? image_284 : _GEN_346; // @[Filter.scala 138:46]
  wire [3:0] _GEN_348 = 12'h11d == _T_46[11:0] ? image_285 : _GEN_347; // @[Filter.scala 138:46]
  wire [3:0] _GEN_349 = 12'h11e == _T_46[11:0] ? image_286 : _GEN_348; // @[Filter.scala 138:46]
  wire [3:0] _GEN_350 = 12'h11f == _T_46[11:0] ? image_287 : _GEN_349; // @[Filter.scala 138:46]
  wire [3:0] _GEN_351 = 12'h120 == _T_46[11:0] ? image_288 : _GEN_350; // @[Filter.scala 138:46]
  wire [3:0] _GEN_352 = 12'h121 == _T_46[11:0] ? image_289 : _GEN_351; // @[Filter.scala 138:46]
  wire [3:0] _GEN_353 = 12'h122 == _T_46[11:0] ? image_290 : _GEN_352; // @[Filter.scala 138:46]
  wire [3:0] _GEN_354 = 12'h123 == _T_46[11:0] ? image_291 : _GEN_353; // @[Filter.scala 138:46]
  wire [3:0] _GEN_355 = 12'h124 == _T_46[11:0] ? image_292 : _GEN_354; // @[Filter.scala 138:46]
  wire [3:0] _GEN_356 = 12'h125 == _T_46[11:0] ? image_293 : _GEN_355; // @[Filter.scala 138:46]
  wire [3:0] _GEN_357 = 12'h126 == _T_46[11:0] ? image_294 : _GEN_356; // @[Filter.scala 138:46]
  wire [3:0] _GEN_358 = 12'h127 == _T_46[11:0] ? image_295 : _GEN_357; // @[Filter.scala 138:46]
  wire [3:0] _GEN_359 = 12'h128 == _T_46[11:0] ? image_296 : _GEN_358; // @[Filter.scala 138:46]
  wire [3:0] _GEN_360 = 12'h129 == _T_46[11:0] ? image_297 : _GEN_359; // @[Filter.scala 138:46]
  wire [3:0] _GEN_361 = 12'h12a == _T_46[11:0] ? image_298 : _GEN_360; // @[Filter.scala 138:46]
  wire [3:0] _GEN_362 = 12'h12b == _T_46[11:0] ? image_299 : _GEN_361; // @[Filter.scala 138:46]
  wire [3:0] _GEN_363 = 12'h12c == _T_46[11:0] ? image_300 : _GEN_362; // @[Filter.scala 138:46]
  wire [3:0] _GEN_364 = 12'h12d == _T_46[11:0] ? image_301 : _GEN_363; // @[Filter.scala 138:46]
  wire [3:0] _GEN_365 = 12'h12e == _T_46[11:0] ? image_302 : _GEN_364; // @[Filter.scala 138:46]
  wire [3:0] _GEN_366 = 12'h12f == _T_46[11:0] ? image_303 : _GEN_365; // @[Filter.scala 138:46]
  wire [3:0] _GEN_367 = 12'h130 == _T_46[11:0] ? image_304 : _GEN_366; // @[Filter.scala 138:46]
  wire [3:0] _GEN_368 = 12'h131 == _T_46[11:0] ? image_305 : _GEN_367; // @[Filter.scala 138:46]
  wire [3:0] _GEN_369 = 12'h132 == _T_46[11:0] ? image_306 : _GEN_368; // @[Filter.scala 138:46]
  wire [3:0] _GEN_370 = 12'h133 == _T_46[11:0] ? image_307 : _GEN_369; // @[Filter.scala 138:46]
  wire [3:0] _GEN_371 = 12'h134 == _T_46[11:0] ? image_308 : _GEN_370; // @[Filter.scala 138:46]
  wire [3:0] _GEN_372 = 12'h135 == _T_46[11:0] ? image_309 : _GEN_371; // @[Filter.scala 138:46]
  wire [3:0] _GEN_373 = 12'h136 == _T_46[11:0] ? image_310 : _GEN_372; // @[Filter.scala 138:46]
  wire [3:0] _GEN_374 = 12'h137 == _T_46[11:0] ? image_311 : _GEN_373; // @[Filter.scala 138:46]
  wire [3:0] _GEN_375 = 12'h138 == _T_46[11:0] ? image_312 : _GEN_374; // @[Filter.scala 138:46]
  wire [3:0] _GEN_376 = 12'h139 == _T_46[11:0] ? image_313 : _GEN_375; // @[Filter.scala 138:46]
  wire [3:0] _GEN_377 = 12'h13a == _T_46[11:0] ? image_314 : _GEN_376; // @[Filter.scala 138:46]
  wire [3:0] _GEN_378 = 12'h13b == _T_46[11:0] ? image_315 : _GEN_377; // @[Filter.scala 138:46]
  wire [3:0] _GEN_379 = 12'h13c == _T_46[11:0] ? 4'h0 : _GEN_378; // @[Filter.scala 138:46]
  wire [3:0] _GEN_380 = 12'h13d == _T_46[11:0] ? 4'h0 : _GEN_379; // @[Filter.scala 138:46]
  wire [3:0] _GEN_381 = 12'h13e == _T_46[11:0] ? 4'h0 : _GEN_380; // @[Filter.scala 138:46]
  wire [3:0] _GEN_382 = 12'h13f == _T_46[11:0] ? 4'h0 : _GEN_381; // @[Filter.scala 138:46]
  wire [3:0] _GEN_383 = 12'h140 == _T_46[11:0] ? 4'h0 : _GEN_382; // @[Filter.scala 138:46]
  wire [3:0] _GEN_384 = 12'h141 == _T_46[11:0] ? 4'h0 : _GEN_383; // @[Filter.scala 138:46]
  wire [3:0] _GEN_385 = 12'h142 == _T_46[11:0] ? 4'h0 : _GEN_384; // @[Filter.scala 138:46]
  wire [3:0] _GEN_386 = 12'h143 == _T_46[11:0] ? 4'h0 : _GEN_385; // @[Filter.scala 138:46]
  wire [3:0] _GEN_387 = 12'h144 == _T_46[11:0] ? 4'h0 : _GEN_386; // @[Filter.scala 138:46]
  wire [3:0] _GEN_388 = 12'h145 == _T_46[11:0] ? image_325 : _GEN_387; // @[Filter.scala 138:46]
  wire [3:0] _GEN_389 = 12'h146 == _T_46[11:0] ? image_326 : _GEN_388; // @[Filter.scala 138:46]
  wire [3:0] _GEN_390 = 12'h147 == _T_46[11:0] ? image_327 : _GEN_389; // @[Filter.scala 138:46]
  wire [3:0] _GEN_391 = 12'h148 == _T_46[11:0] ? image_328 : _GEN_390; // @[Filter.scala 138:46]
  wire [3:0] _GEN_392 = 12'h149 == _T_46[11:0] ? image_329 : _GEN_391; // @[Filter.scala 138:46]
  wire [3:0] _GEN_393 = 12'h14a == _T_46[11:0] ? image_330 : _GEN_392; // @[Filter.scala 138:46]
  wire [3:0] _GEN_394 = 12'h14b == _T_46[11:0] ? image_331 : _GEN_393; // @[Filter.scala 138:46]
  wire [3:0] _GEN_395 = 12'h14c == _T_46[11:0] ? image_332 : _GEN_394; // @[Filter.scala 138:46]
  wire [3:0] _GEN_396 = 12'h14d == _T_46[11:0] ? image_333 : _GEN_395; // @[Filter.scala 138:46]
  wire [3:0] _GEN_397 = 12'h14e == _T_46[11:0] ? image_334 : _GEN_396; // @[Filter.scala 138:46]
  wire [3:0] _GEN_398 = 12'h14f == _T_46[11:0] ? image_335 : _GEN_397; // @[Filter.scala 138:46]
  wire [3:0] _GEN_399 = 12'h150 == _T_46[11:0] ? image_336 : _GEN_398; // @[Filter.scala 138:46]
  wire [3:0] _GEN_400 = 12'h151 == _T_46[11:0] ? image_337 : _GEN_399; // @[Filter.scala 138:46]
  wire [3:0] _GEN_401 = 12'h152 == _T_46[11:0] ? image_338 : _GEN_400; // @[Filter.scala 138:46]
  wire [3:0] _GEN_402 = 12'h153 == _T_46[11:0] ? image_339 : _GEN_401; // @[Filter.scala 138:46]
  wire [3:0] _GEN_403 = 12'h154 == _T_46[11:0] ? image_340 : _GEN_402; // @[Filter.scala 138:46]
  wire [3:0] _GEN_404 = 12'h155 == _T_46[11:0] ? image_341 : _GEN_403; // @[Filter.scala 138:46]
  wire [3:0] _GEN_405 = 12'h156 == _T_46[11:0] ? image_342 : _GEN_404; // @[Filter.scala 138:46]
  wire [3:0] _GEN_406 = 12'h157 == _T_46[11:0] ? image_343 : _GEN_405; // @[Filter.scala 138:46]
  wire [3:0] _GEN_407 = 12'h158 == _T_46[11:0] ? image_344 : _GEN_406; // @[Filter.scala 138:46]
  wire [3:0] _GEN_408 = 12'h159 == _T_46[11:0] ? image_345 : _GEN_407; // @[Filter.scala 138:46]
  wire [3:0] _GEN_409 = 12'h15a == _T_46[11:0] ? image_346 : _GEN_408; // @[Filter.scala 138:46]
  wire [3:0] _GEN_410 = 12'h15b == _T_46[11:0] ? image_347 : _GEN_409; // @[Filter.scala 138:46]
  wire [3:0] _GEN_411 = 12'h15c == _T_46[11:0] ? image_348 : _GEN_410; // @[Filter.scala 138:46]
  wire [3:0] _GEN_412 = 12'h15d == _T_46[11:0] ? image_349 : _GEN_411; // @[Filter.scala 138:46]
  wire [3:0] _GEN_413 = 12'h15e == _T_46[11:0] ? image_350 : _GEN_412; // @[Filter.scala 138:46]
  wire [3:0] _GEN_414 = 12'h15f == _T_46[11:0] ? image_351 : _GEN_413; // @[Filter.scala 138:46]
  wire [3:0] _GEN_415 = 12'h160 == _T_46[11:0] ? image_352 : _GEN_414; // @[Filter.scala 138:46]
  wire [3:0] _GEN_416 = 12'h161 == _T_46[11:0] ? image_353 : _GEN_415; // @[Filter.scala 138:46]
  wire [3:0] _GEN_417 = 12'h162 == _T_46[11:0] ? image_354 : _GEN_416; // @[Filter.scala 138:46]
  wire [3:0] _GEN_418 = 12'h163 == _T_46[11:0] ? image_355 : _GEN_417; // @[Filter.scala 138:46]
  wire [3:0] _GEN_419 = 12'h164 == _T_46[11:0] ? image_356 : _GEN_418; // @[Filter.scala 138:46]
  wire [3:0] _GEN_420 = 12'h165 == _T_46[11:0] ? image_357 : _GEN_419; // @[Filter.scala 138:46]
  wire [3:0] _GEN_421 = 12'h166 == _T_46[11:0] ? image_358 : _GEN_420; // @[Filter.scala 138:46]
  wire [3:0] _GEN_422 = 12'h167 == _T_46[11:0] ? image_359 : _GEN_421; // @[Filter.scala 138:46]
  wire [3:0] _GEN_423 = 12'h168 == _T_46[11:0] ? image_360 : _GEN_422; // @[Filter.scala 138:46]
  wire [3:0] _GEN_424 = 12'h169 == _T_46[11:0] ? image_361 : _GEN_423; // @[Filter.scala 138:46]
  wire [3:0] _GEN_425 = 12'h16a == _T_46[11:0] ? image_362 : _GEN_424; // @[Filter.scala 138:46]
  wire [3:0] _GEN_426 = 12'h16b == _T_46[11:0] ? image_363 : _GEN_425; // @[Filter.scala 138:46]
  wire [3:0] _GEN_427 = 12'h16c == _T_46[11:0] ? image_364 : _GEN_426; // @[Filter.scala 138:46]
  wire [3:0] _GEN_428 = 12'h16d == _T_46[11:0] ? image_365 : _GEN_427; // @[Filter.scala 138:46]
  wire [3:0] _GEN_429 = 12'h16e == _T_46[11:0] ? image_366 : _GEN_428; // @[Filter.scala 138:46]
  wire [3:0] _GEN_430 = 12'h16f == _T_46[11:0] ? image_367 : _GEN_429; // @[Filter.scala 138:46]
  wire [3:0] _GEN_431 = 12'h170 == _T_46[11:0] ? image_368 : _GEN_430; // @[Filter.scala 138:46]
  wire [3:0] _GEN_432 = 12'h171 == _T_46[11:0] ? image_369 : _GEN_431; // @[Filter.scala 138:46]
  wire [3:0] _GEN_433 = 12'h172 == _T_46[11:0] ? image_370 : _GEN_432; // @[Filter.scala 138:46]
  wire [3:0] _GEN_434 = 12'h173 == _T_46[11:0] ? image_371 : _GEN_433; // @[Filter.scala 138:46]
  wire [3:0] _GEN_435 = 12'h174 == _T_46[11:0] ? image_372 : _GEN_434; // @[Filter.scala 138:46]
  wire [3:0] _GEN_436 = 12'h175 == _T_46[11:0] ? image_373 : _GEN_435; // @[Filter.scala 138:46]
  wire [3:0] _GEN_437 = 12'h176 == _T_46[11:0] ? image_374 : _GEN_436; // @[Filter.scala 138:46]
  wire [3:0] _GEN_438 = 12'h177 == _T_46[11:0] ? image_375 : _GEN_437; // @[Filter.scala 138:46]
  wire [3:0] _GEN_439 = 12'h178 == _T_46[11:0] ? image_376 : _GEN_438; // @[Filter.scala 138:46]
  wire [3:0] _GEN_440 = 12'h179 == _T_46[11:0] ? image_377 : _GEN_439; // @[Filter.scala 138:46]
  wire [3:0] _GEN_441 = 12'h17a == _T_46[11:0] ? image_378 : _GEN_440; // @[Filter.scala 138:46]
  wire [3:0] _GEN_442 = 12'h17b == _T_46[11:0] ? image_379 : _GEN_441; // @[Filter.scala 138:46]
  wire [3:0] _GEN_443 = 12'h17c == _T_46[11:0] ? 4'h0 : _GEN_442; // @[Filter.scala 138:46]
  wire [3:0] _GEN_444 = 12'h17d == _T_46[11:0] ? 4'h0 : _GEN_443; // @[Filter.scala 138:46]
  wire [3:0] _GEN_445 = 12'h17e == _T_46[11:0] ? 4'h0 : _GEN_444; // @[Filter.scala 138:46]
  wire [3:0] _GEN_446 = 12'h17f == _T_46[11:0] ? 4'h0 : _GEN_445; // @[Filter.scala 138:46]
  wire [3:0] _GEN_447 = 12'h180 == _T_46[11:0] ? 4'h0 : _GEN_446; // @[Filter.scala 138:46]
  wire [3:0] _GEN_448 = 12'h181 == _T_46[11:0] ? 4'h0 : _GEN_447; // @[Filter.scala 138:46]
  wire [3:0] _GEN_449 = 12'h182 == _T_46[11:0] ? 4'h0 : _GEN_448; // @[Filter.scala 138:46]
  wire [3:0] _GEN_450 = 12'h183 == _T_46[11:0] ? 4'h0 : _GEN_449; // @[Filter.scala 138:46]
  wire [3:0] _GEN_451 = 12'h184 == _T_46[11:0] ? image_388 : _GEN_450; // @[Filter.scala 138:46]
  wire [3:0] _GEN_452 = 12'h185 == _T_46[11:0] ? image_389 : _GEN_451; // @[Filter.scala 138:46]
  wire [3:0] _GEN_453 = 12'h186 == _T_46[11:0] ? image_390 : _GEN_452; // @[Filter.scala 138:46]
  wire [3:0] _GEN_454 = 12'h187 == _T_46[11:0] ? image_391 : _GEN_453; // @[Filter.scala 138:46]
  wire [3:0] _GEN_455 = 12'h188 == _T_46[11:0] ? image_392 : _GEN_454; // @[Filter.scala 138:46]
  wire [3:0] _GEN_456 = 12'h189 == _T_46[11:0] ? image_393 : _GEN_455; // @[Filter.scala 138:46]
  wire [3:0] _GEN_457 = 12'h18a == _T_46[11:0] ? image_394 : _GEN_456; // @[Filter.scala 138:46]
  wire [3:0] _GEN_458 = 12'h18b == _T_46[11:0] ? image_395 : _GEN_457; // @[Filter.scala 138:46]
  wire [3:0] _GEN_459 = 12'h18c == _T_46[11:0] ? image_396 : _GEN_458; // @[Filter.scala 138:46]
  wire [3:0] _GEN_460 = 12'h18d == _T_46[11:0] ? image_397 : _GEN_459; // @[Filter.scala 138:46]
  wire [3:0] _GEN_461 = 12'h18e == _T_46[11:0] ? image_398 : _GEN_460; // @[Filter.scala 138:46]
  wire [3:0] _GEN_462 = 12'h18f == _T_46[11:0] ? image_399 : _GEN_461; // @[Filter.scala 138:46]
  wire [3:0] _GEN_463 = 12'h190 == _T_46[11:0] ? image_400 : _GEN_462; // @[Filter.scala 138:46]
  wire [3:0] _GEN_464 = 12'h191 == _T_46[11:0] ? image_401 : _GEN_463; // @[Filter.scala 138:46]
  wire [3:0] _GEN_465 = 12'h192 == _T_46[11:0] ? image_402 : _GEN_464; // @[Filter.scala 138:46]
  wire [3:0] _GEN_466 = 12'h193 == _T_46[11:0] ? image_403 : _GEN_465; // @[Filter.scala 138:46]
  wire [3:0] _GEN_467 = 12'h194 == _T_46[11:0] ? image_404 : _GEN_466; // @[Filter.scala 138:46]
  wire [3:0] _GEN_468 = 12'h195 == _T_46[11:0] ? image_405 : _GEN_467; // @[Filter.scala 138:46]
  wire [3:0] _GEN_469 = 12'h196 == _T_46[11:0] ? image_406 : _GEN_468; // @[Filter.scala 138:46]
  wire [3:0] _GEN_470 = 12'h197 == _T_46[11:0] ? image_407 : _GEN_469; // @[Filter.scala 138:46]
  wire [3:0] _GEN_471 = 12'h198 == _T_46[11:0] ? image_408 : _GEN_470; // @[Filter.scala 138:46]
  wire [3:0] _GEN_472 = 12'h199 == _T_46[11:0] ? image_409 : _GEN_471; // @[Filter.scala 138:46]
  wire [3:0] _GEN_473 = 12'h19a == _T_46[11:0] ? image_410 : _GEN_472; // @[Filter.scala 138:46]
  wire [3:0] _GEN_474 = 12'h19b == _T_46[11:0] ? image_411 : _GEN_473; // @[Filter.scala 138:46]
  wire [3:0] _GEN_475 = 12'h19c == _T_46[11:0] ? image_412 : _GEN_474; // @[Filter.scala 138:46]
  wire [3:0] _GEN_476 = 12'h19d == _T_46[11:0] ? image_413 : _GEN_475; // @[Filter.scala 138:46]
  wire [3:0] _GEN_477 = 12'h19e == _T_46[11:0] ? image_414 : _GEN_476; // @[Filter.scala 138:46]
  wire [3:0] _GEN_478 = 12'h19f == _T_46[11:0] ? image_415 : _GEN_477; // @[Filter.scala 138:46]
  wire [3:0] _GEN_479 = 12'h1a0 == _T_46[11:0] ? image_416 : _GEN_478; // @[Filter.scala 138:46]
  wire [3:0] _GEN_480 = 12'h1a1 == _T_46[11:0] ? image_417 : _GEN_479; // @[Filter.scala 138:46]
  wire [3:0] _GEN_481 = 12'h1a2 == _T_46[11:0] ? image_418 : _GEN_480; // @[Filter.scala 138:46]
  wire [3:0] _GEN_482 = 12'h1a3 == _T_46[11:0] ? image_419 : _GEN_481; // @[Filter.scala 138:46]
  wire [3:0] _GEN_483 = 12'h1a4 == _T_46[11:0] ? image_420 : _GEN_482; // @[Filter.scala 138:46]
  wire [3:0] _GEN_484 = 12'h1a5 == _T_46[11:0] ? image_421 : _GEN_483; // @[Filter.scala 138:46]
  wire [3:0] _GEN_485 = 12'h1a6 == _T_46[11:0] ? image_422 : _GEN_484; // @[Filter.scala 138:46]
  wire [3:0] _GEN_486 = 12'h1a7 == _T_46[11:0] ? image_423 : _GEN_485; // @[Filter.scala 138:46]
  wire [3:0] _GEN_487 = 12'h1a8 == _T_46[11:0] ? image_424 : _GEN_486; // @[Filter.scala 138:46]
  wire [3:0] _GEN_488 = 12'h1a9 == _T_46[11:0] ? image_425 : _GEN_487; // @[Filter.scala 138:46]
  wire [3:0] _GEN_489 = 12'h1aa == _T_46[11:0] ? image_426 : _GEN_488; // @[Filter.scala 138:46]
  wire [3:0] _GEN_490 = 12'h1ab == _T_46[11:0] ? image_427 : _GEN_489; // @[Filter.scala 138:46]
  wire [3:0] _GEN_491 = 12'h1ac == _T_46[11:0] ? image_428 : _GEN_490; // @[Filter.scala 138:46]
  wire [3:0] _GEN_492 = 12'h1ad == _T_46[11:0] ? image_429 : _GEN_491; // @[Filter.scala 138:46]
  wire [3:0] _GEN_493 = 12'h1ae == _T_46[11:0] ? image_430 : _GEN_492; // @[Filter.scala 138:46]
  wire [3:0] _GEN_494 = 12'h1af == _T_46[11:0] ? image_431 : _GEN_493; // @[Filter.scala 138:46]
  wire [3:0] _GEN_495 = 12'h1b0 == _T_46[11:0] ? image_432 : _GEN_494; // @[Filter.scala 138:46]
  wire [3:0] _GEN_496 = 12'h1b1 == _T_46[11:0] ? image_433 : _GEN_495; // @[Filter.scala 138:46]
  wire [3:0] _GEN_497 = 12'h1b2 == _T_46[11:0] ? image_434 : _GEN_496; // @[Filter.scala 138:46]
  wire [3:0] _GEN_498 = 12'h1b3 == _T_46[11:0] ? image_435 : _GEN_497; // @[Filter.scala 138:46]
  wire [3:0] _GEN_499 = 12'h1b4 == _T_46[11:0] ? image_436 : _GEN_498; // @[Filter.scala 138:46]
  wire [3:0] _GEN_500 = 12'h1b5 == _T_46[11:0] ? image_437 : _GEN_499; // @[Filter.scala 138:46]
  wire [3:0] _GEN_501 = 12'h1b6 == _T_46[11:0] ? image_438 : _GEN_500; // @[Filter.scala 138:46]
  wire [3:0] _GEN_502 = 12'h1b7 == _T_46[11:0] ? image_439 : _GEN_501; // @[Filter.scala 138:46]
  wire [3:0] _GEN_503 = 12'h1b8 == _T_46[11:0] ? image_440 : _GEN_502; // @[Filter.scala 138:46]
  wire [3:0] _GEN_504 = 12'h1b9 == _T_46[11:0] ? image_441 : _GEN_503; // @[Filter.scala 138:46]
  wire [3:0] _GEN_505 = 12'h1ba == _T_46[11:0] ? image_442 : _GEN_504; // @[Filter.scala 138:46]
  wire [3:0] _GEN_506 = 12'h1bb == _T_46[11:0] ? image_443 : _GEN_505; // @[Filter.scala 138:46]
  wire [3:0] _GEN_507 = 12'h1bc == _T_46[11:0] ? image_444 : _GEN_506; // @[Filter.scala 138:46]
  wire [3:0] _GEN_508 = 12'h1bd == _T_46[11:0] ? 4'h0 : _GEN_507; // @[Filter.scala 138:46]
  wire [3:0] _GEN_509 = 12'h1be == _T_46[11:0] ? 4'h0 : _GEN_508; // @[Filter.scala 138:46]
  wire [3:0] _GEN_510 = 12'h1bf == _T_46[11:0] ? 4'h0 : _GEN_509; // @[Filter.scala 138:46]
  wire [3:0] _GEN_511 = 12'h1c0 == _T_46[11:0] ? 4'h0 : _GEN_510; // @[Filter.scala 138:46]
  wire [3:0] _GEN_512 = 12'h1c1 == _T_46[11:0] ? 4'h0 : _GEN_511; // @[Filter.scala 138:46]
  wire [3:0] _GEN_513 = 12'h1c2 == _T_46[11:0] ? 4'h0 : _GEN_512; // @[Filter.scala 138:46]
  wire [3:0] _GEN_514 = 12'h1c3 == _T_46[11:0] ? image_451 : _GEN_513; // @[Filter.scala 138:46]
  wire [3:0] _GEN_515 = 12'h1c4 == _T_46[11:0] ? image_452 : _GEN_514; // @[Filter.scala 138:46]
  wire [3:0] _GEN_516 = 12'h1c5 == _T_46[11:0] ? image_453 : _GEN_515; // @[Filter.scala 138:46]
  wire [3:0] _GEN_517 = 12'h1c6 == _T_46[11:0] ? image_454 : _GEN_516; // @[Filter.scala 138:46]
  wire [3:0] _GEN_518 = 12'h1c7 == _T_46[11:0] ? image_455 : _GEN_517; // @[Filter.scala 138:46]
  wire [3:0] _GEN_519 = 12'h1c8 == _T_46[11:0] ? image_456 : _GEN_518; // @[Filter.scala 138:46]
  wire [3:0] _GEN_520 = 12'h1c9 == _T_46[11:0] ? image_457 : _GEN_519; // @[Filter.scala 138:46]
  wire [3:0] _GEN_521 = 12'h1ca == _T_46[11:0] ? image_458 : _GEN_520; // @[Filter.scala 138:46]
  wire [3:0] _GEN_522 = 12'h1cb == _T_46[11:0] ? image_459 : _GEN_521; // @[Filter.scala 138:46]
  wire [3:0] _GEN_523 = 12'h1cc == _T_46[11:0] ? image_460 : _GEN_522; // @[Filter.scala 138:46]
  wire [3:0] _GEN_524 = 12'h1cd == _T_46[11:0] ? image_461 : _GEN_523; // @[Filter.scala 138:46]
  wire [3:0] _GEN_525 = 12'h1ce == _T_46[11:0] ? image_462 : _GEN_524; // @[Filter.scala 138:46]
  wire [3:0] _GEN_526 = 12'h1cf == _T_46[11:0] ? image_463 : _GEN_525; // @[Filter.scala 138:46]
  wire [3:0] _GEN_527 = 12'h1d0 == _T_46[11:0] ? image_464 : _GEN_526; // @[Filter.scala 138:46]
  wire [3:0] _GEN_528 = 12'h1d1 == _T_46[11:0] ? image_465 : _GEN_527; // @[Filter.scala 138:46]
  wire [3:0] _GEN_529 = 12'h1d2 == _T_46[11:0] ? image_466 : _GEN_528; // @[Filter.scala 138:46]
  wire [3:0] _GEN_530 = 12'h1d3 == _T_46[11:0] ? image_467 : _GEN_529; // @[Filter.scala 138:46]
  wire [3:0] _GEN_531 = 12'h1d4 == _T_46[11:0] ? image_468 : _GEN_530; // @[Filter.scala 138:46]
  wire [3:0] _GEN_532 = 12'h1d5 == _T_46[11:0] ? image_469 : _GEN_531; // @[Filter.scala 138:46]
  wire [3:0] _GEN_533 = 12'h1d6 == _T_46[11:0] ? image_470 : _GEN_532; // @[Filter.scala 138:46]
  wire [3:0] _GEN_534 = 12'h1d7 == _T_46[11:0] ? image_471 : _GEN_533; // @[Filter.scala 138:46]
  wire [3:0] _GEN_535 = 12'h1d8 == _T_46[11:0] ? image_472 : _GEN_534; // @[Filter.scala 138:46]
  wire [3:0] _GEN_536 = 12'h1d9 == _T_46[11:0] ? image_473 : _GEN_535; // @[Filter.scala 138:46]
  wire [3:0] _GEN_537 = 12'h1da == _T_46[11:0] ? image_474 : _GEN_536; // @[Filter.scala 138:46]
  wire [3:0] _GEN_538 = 12'h1db == _T_46[11:0] ? image_475 : _GEN_537; // @[Filter.scala 138:46]
  wire [3:0] _GEN_539 = 12'h1dc == _T_46[11:0] ? image_476 : _GEN_538; // @[Filter.scala 138:46]
  wire [3:0] _GEN_540 = 12'h1dd == _T_46[11:0] ? image_477 : _GEN_539; // @[Filter.scala 138:46]
  wire [3:0] _GEN_541 = 12'h1de == _T_46[11:0] ? image_478 : _GEN_540; // @[Filter.scala 138:46]
  wire [3:0] _GEN_542 = 12'h1df == _T_46[11:0] ? image_479 : _GEN_541; // @[Filter.scala 138:46]
  wire [3:0] _GEN_543 = 12'h1e0 == _T_46[11:0] ? image_480 : _GEN_542; // @[Filter.scala 138:46]
  wire [3:0] _GEN_544 = 12'h1e1 == _T_46[11:0] ? image_481 : _GEN_543; // @[Filter.scala 138:46]
  wire [3:0] _GEN_545 = 12'h1e2 == _T_46[11:0] ? image_482 : _GEN_544; // @[Filter.scala 138:46]
  wire [3:0] _GEN_546 = 12'h1e3 == _T_46[11:0] ? image_483 : _GEN_545; // @[Filter.scala 138:46]
  wire [3:0] _GEN_547 = 12'h1e4 == _T_46[11:0] ? image_484 : _GEN_546; // @[Filter.scala 138:46]
  wire [3:0] _GEN_548 = 12'h1e5 == _T_46[11:0] ? image_485 : _GEN_547; // @[Filter.scala 138:46]
  wire [3:0] _GEN_549 = 12'h1e6 == _T_46[11:0] ? image_486 : _GEN_548; // @[Filter.scala 138:46]
  wire [3:0] _GEN_550 = 12'h1e7 == _T_46[11:0] ? image_487 : _GEN_549; // @[Filter.scala 138:46]
  wire [3:0] _GEN_551 = 12'h1e8 == _T_46[11:0] ? image_488 : _GEN_550; // @[Filter.scala 138:46]
  wire [3:0] _GEN_552 = 12'h1e9 == _T_46[11:0] ? image_489 : _GEN_551; // @[Filter.scala 138:46]
  wire [3:0] _GEN_553 = 12'h1ea == _T_46[11:0] ? image_490 : _GEN_552; // @[Filter.scala 138:46]
  wire [3:0] _GEN_554 = 12'h1eb == _T_46[11:0] ? image_491 : _GEN_553; // @[Filter.scala 138:46]
  wire [3:0] _GEN_555 = 12'h1ec == _T_46[11:0] ? image_492 : _GEN_554; // @[Filter.scala 138:46]
  wire [3:0] _GEN_556 = 12'h1ed == _T_46[11:0] ? image_493 : _GEN_555; // @[Filter.scala 138:46]
  wire [3:0] _GEN_557 = 12'h1ee == _T_46[11:0] ? image_494 : _GEN_556; // @[Filter.scala 138:46]
  wire [3:0] _GEN_558 = 12'h1ef == _T_46[11:0] ? image_495 : _GEN_557; // @[Filter.scala 138:46]
  wire [3:0] _GEN_559 = 12'h1f0 == _T_46[11:0] ? image_496 : _GEN_558; // @[Filter.scala 138:46]
  wire [3:0] _GEN_560 = 12'h1f1 == _T_46[11:0] ? image_497 : _GEN_559; // @[Filter.scala 138:46]
  wire [3:0] _GEN_561 = 12'h1f2 == _T_46[11:0] ? image_498 : _GEN_560; // @[Filter.scala 138:46]
  wire [3:0] _GEN_562 = 12'h1f3 == _T_46[11:0] ? image_499 : _GEN_561; // @[Filter.scala 138:46]
  wire [3:0] _GEN_563 = 12'h1f4 == _T_46[11:0] ? image_500 : _GEN_562; // @[Filter.scala 138:46]
  wire [3:0] _GEN_564 = 12'h1f5 == _T_46[11:0] ? image_501 : _GEN_563; // @[Filter.scala 138:46]
  wire [3:0] _GEN_565 = 12'h1f6 == _T_46[11:0] ? image_502 : _GEN_564; // @[Filter.scala 138:46]
  wire [3:0] _GEN_566 = 12'h1f7 == _T_46[11:0] ? image_503 : _GEN_565; // @[Filter.scala 138:46]
  wire [3:0] _GEN_567 = 12'h1f8 == _T_46[11:0] ? image_504 : _GEN_566; // @[Filter.scala 138:46]
  wire [3:0] _GEN_568 = 12'h1f9 == _T_46[11:0] ? image_505 : _GEN_567; // @[Filter.scala 138:46]
  wire [3:0] _GEN_569 = 12'h1fa == _T_46[11:0] ? image_506 : _GEN_568; // @[Filter.scala 138:46]
  wire [3:0] _GEN_570 = 12'h1fb == _T_46[11:0] ? image_507 : _GEN_569; // @[Filter.scala 138:46]
  wire [3:0] _GEN_571 = 12'h1fc == _T_46[11:0] ? image_508 : _GEN_570; // @[Filter.scala 138:46]
  wire [3:0] _GEN_572 = 12'h1fd == _T_46[11:0] ? image_509 : _GEN_571; // @[Filter.scala 138:46]
  wire [3:0] _GEN_573 = 12'h1fe == _T_46[11:0] ? 4'h0 : _GEN_572; // @[Filter.scala 138:46]
  wire [3:0] _GEN_574 = 12'h1ff == _T_46[11:0] ? 4'h0 : _GEN_573; // @[Filter.scala 138:46]
  wire [3:0] _GEN_575 = 12'h200 == _T_46[11:0] ? 4'h0 : _GEN_574; // @[Filter.scala 138:46]
  wire [3:0] _GEN_576 = 12'h201 == _T_46[11:0] ? 4'h0 : _GEN_575; // @[Filter.scala 138:46]
  wire [3:0] _GEN_577 = 12'h202 == _T_46[11:0] ? 4'h0 : _GEN_576; // @[Filter.scala 138:46]
  wire [3:0] _GEN_578 = 12'h203 == _T_46[11:0] ? image_515 : _GEN_577; // @[Filter.scala 138:46]
  wire [3:0] _GEN_579 = 12'h204 == _T_46[11:0] ? image_516 : _GEN_578; // @[Filter.scala 138:46]
  wire [3:0] _GEN_580 = 12'h205 == _T_46[11:0] ? image_517 : _GEN_579; // @[Filter.scala 138:46]
  wire [3:0] _GEN_581 = 12'h206 == _T_46[11:0] ? image_518 : _GEN_580; // @[Filter.scala 138:46]
  wire [3:0] _GEN_582 = 12'h207 == _T_46[11:0] ? image_519 : _GEN_581; // @[Filter.scala 138:46]
  wire [3:0] _GEN_583 = 12'h208 == _T_46[11:0] ? image_520 : _GEN_582; // @[Filter.scala 138:46]
  wire [3:0] _GEN_584 = 12'h209 == _T_46[11:0] ? image_521 : _GEN_583; // @[Filter.scala 138:46]
  wire [3:0] _GEN_585 = 12'h20a == _T_46[11:0] ? image_522 : _GEN_584; // @[Filter.scala 138:46]
  wire [3:0] _GEN_586 = 12'h20b == _T_46[11:0] ? image_523 : _GEN_585; // @[Filter.scala 138:46]
  wire [3:0] _GEN_587 = 12'h20c == _T_46[11:0] ? image_524 : _GEN_586; // @[Filter.scala 138:46]
  wire [3:0] _GEN_588 = 12'h20d == _T_46[11:0] ? image_525 : _GEN_587; // @[Filter.scala 138:46]
  wire [3:0] _GEN_589 = 12'h20e == _T_46[11:0] ? image_526 : _GEN_588; // @[Filter.scala 138:46]
  wire [3:0] _GEN_590 = 12'h20f == _T_46[11:0] ? image_527 : _GEN_589; // @[Filter.scala 138:46]
  wire [3:0] _GEN_591 = 12'h210 == _T_46[11:0] ? image_528 : _GEN_590; // @[Filter.scala 138:46]
  wire [3:0] _GEN_592 = 12'h211 == _T_46[11:0] ? image_529 : _GEN_591; // @[Filter.scala 138:46]
  wire [3:0] _GEN_593 = 12'h212 == _T_46[11:0] ? image_530 : _GEN_592; // @[Filter.scala 138:46]
  wire [3:0] _GEN_594 = 12'h213 == _T_46[11:0] ? image_531 : _GEN_593; // @[Filter.scala 138:46]
  wire [3:0] _GEN_595 = 12'h214 == _T_46[11:0] ? image_532 : _GEN_594; // @[Filter.scala 138:46]
  wire [3:0] _GEN_596 = 12'h215 == _T_46[11:0] ? image_533 : _GEN_595; // @[Filter.scala 138:46]
  wire [3:0] _GEN_597 = 12'h216 == _T_46[11:0] ? image_534 : _GEN_596; // @[Filter.scala 138:46]
  wire [3:0] _GEN_598 = 12'h217 == _T_46[11:0] ? image_535 : _GEN_597; // @[Filter.scala 138:46]
  wire [3:0] _GEN_599 = 12'h218 == _T_46[11:0] ? image_536 : _GEN_598; // @[Filter.scala 138:46]
  wire [3:0] _GEN_600 = 12'h219 == _T_46[11:0] ? image_537 : _GEN_599; // @[Filter.scala 138:46]
  wire [3:0] _GEN_601 = 12'h21a == _T_46[11:0] ? image_538 : _GEN_600; // @[Filter.scala 138:46]
  wire [3:0] _GEN_602 = 12'h21b == _T_46[11:0] ? image_539 : _GEN_601; // @[Filter.scala 138:46]
  wire [3:0] _GEN_603 = 12'h21c == _T_46[11:0] ? image_540 : _GEN_602; // @[Filter.scala 138:46]
  wire [3:0] _GEN_604 = 12'h21d == _T_46[11:0] ? image_541 : _GEN_603; // @[Filter.scala 138:46]
  wire [3:0] _GEN_605 = 12'h21e == _T_46[11:0] ? image_542 : _GEN_604; // @[Filter.scala 138:46]
  wire [3:0] _GEN_606 = 12'h21f == _T_46[11:0] ? image_543 : _GEN_605; // @[Filter.scala 138:46]
  wire [3:0] _GEN_607 = 12'h220 == _T_46[11:0] ? image_544 : _GEN_606; // @[Filter.scala 138:46]
  wire [3:0] _GEN_608 = 12'h221 == _T_46[11:0] ? image_545 : _GEN_607; // @[Filter.scala 138:46]
  wire [3:0] _GEN_609 = 12'h222 == _T_46[11:0] ? image_546 : _GEN_608; // @[Filter.scala 138:46]
  wire [3:0] _GEN_610 = 12'h223 == _T_46[11:0] ? image_547 : _GEN_609; // @[Filter.scala 138:46]
  wire [3:0] _GEN_611 = 12'h224 == _T_46[11:0] ? image_548 : _GEN_610; // @[Filter.scala 138:46]
  wire [3:0] _GEN_612 = 12'h225 == _T_46[11:0] ? image_549 : _GEN_611; // @[Filter.scala 138:46]
  wire [3:0] _GEN_613 = 12'h226 == _T_46[11:0] ? image_550 : _GEN_612; // @[Filter.scala 138:46]
  wire [3:0] _GEN_614 = 12'h227 == _T_46[11:0] ? image_551 : _GEN_613; // @[Filter.scala 138:46]
  wire [3:0] _GEN_615 = 12'h228 == _T_46[11:0] ? image_552 : _GEN_614; // @[Filter.scala 138:46]
  wire [3:0] _GEN_616 = 12'h229 == _T_46[11:0] ? image_553 : _GEN_615; // @[Filter.scala 138:46]
  wire [3:0] _GEN_617 = 12'h22a == _T_46[11:0] ? image_554 : _GEN_616; // @[Filter.scala 138:46]
  wire [3:0] _GEN_618 = 12'h22b == _T_46[11:0] ? image_555 : _GEN_617; // @[Filter.scala 138:46]
  wire [3:0] _GEN_619 = 12'h22c == _T_46[11:0] ? image_556 : _GEN_618; // @[Filter.scala 138:46]
  wire [3:0] _GEN_620 = 12'h22d == _T_46[11:0] ? image_557 : _GEN_619; // @[Filter.scala 138:46]
  wire [3:0] _GEN_621 = 12'h22e == _T_46[11:0] ? image_558 : _GEN_620; // @[Filter.scala 138:46]
  wire [3:0] _GEN_622 = 12'h22f == _T_46[11:0] ? image_559 : _GEN_621; // @[Filter.scala 138:46]
  wire [3:0] _GEN_623 = 12'h230 == _T_46[11:0] ? image_560 : _GEN_622; // @[Filter.scala 138:46]
  wire [3:0] _GEN_624 = 12'h231 == _T_46[11:0] ? image_561 : _GEN_623; // @[Filter.scala 138:46]
  wire [3:0] _GEN_625 = 12'h232 == _T_46[11:0] ? image_562 : _GEN_624; // @[Filter.scala 138:46]
  wire [3:0] _GEN_626 = 12'h233 == _T_46[11:0] ? image_563 : _GEN_625; // @[Filter.scala 138:46]
  wire [3:0] _GEN_627 = 12'h234 == _T_46[11:0] ? image_564 : _GEN_626; // @[Filter.scala 138:46]
  wire [3:0] _GEN_628 = 12'h235 == _T_46[11:0] ? image_565 : _GEN_627; // @[Filter.scala 138:46]
  wire [3:0] _GEN_629 = 12'h236 == _T_46[11:0] ? image_566 : _GEN_628; // @[Filter.scala 138:46]
  wire [3:0] _GEN_630 = 12'h237 == _T_46[11:0] ? 4'h0 : _GEN_629; // @[Filter.scala 138:46]
  wire [3:0] _GEN_631 = 12'h238 == _T_46[11:0] ? 4'h0 : _GEN_630; // @[Filter.scala 138:46]
  wire [3:0] _GEN_632 = 12'h239 == _T_46[11:0] ? 4'h0 : _GEN_631; // @[Filter.scala 138:46]
  wire [3:0] _GEN_633 = 12'h23a == _T_46[11:0] ? 4'h0 : _GEN_632; // @[Filter.scala 138:46]
  wire [3:0] _GEN_634 = 12'h23b == _T_46[11:0] ? image_571 : _GEN_633; // @[Filter.scala 138:46]
  wire [3:0] _GEN_635 = 12'h23c == _T_46[11:0] ? image_572 : _GEN_634; // @[Filter.scala 138:46]
  wire [3:0] _GEN_636 = 12'h23d == _T_46[11:0] ? image_573 : _GEN_635; // @[Filter.scala 138:46]
  wire [3:0] _GEN_637 = 12'h23e == _T_46[11:0] ? image_574 : _GEN_636; // @[Filter.scala 138:46]
  wire [3:0] _GEN_638 = 12'h23f == _T_46[11:0] ? 4'h0 : _GEN_637; // @[Filter.scala 138:46]
  wire [3:0] _GEN_639 = 12'h240 == _T_46[11:0] ? 4'h0 : _GEN_638; // @[Filter.scala 138:46]
  wire [3:0] _GEN_640 = 12'h241 == _T_46[11:0] ? 4'h0 : _GEN_639; // @[Filter.scala 138:46]
  wire [3:0] _GEN_641 = 12'h242 == _T_46[11:0] ? image_578 : _GEN_640; // @[Filter.scala 138:46]
  wire [3:0] _GEN_642 = 12'h243 == _T_46[11:0] ? image_579 : _GEN_641; // @[Filter.scala 138:46]
  wire [3:0] _GEN_643 = 12'h244 == _T_46[11:0] ? image_580 : _GEN_642; // @[Filter.scala 138:46]
  wire [3:0] _GEN_644 = 12'h245 == _T_46[11:0] ? image_581 : _GEN_643; // @[Filter.scala 138:46]
  wire [3:0] _GEN_645 = 12'h246 == _T_46[11:0] ? image_582 : _GEN_644; // @[Filter.scala 138:46]
  wire [3:0] _GEN_646 = 12'h247 == _T_46[11:0] ? image_583 : _GEN_645; // @[Filter.scala 138:46]
  wire [3:0] _GEN_647 = 12'h248 == _T_46[11:0] ? image_584 : _GEN_646; // @[Filter.scala 138:46]
  wire [3:0] _GEN_648 = 12'h249 == _T_46[11:0] ? image_585 : _GEN_647; // @[Filter.scala 138:46]
  wire [3:0] _GEN_649 = 12'h24a == _T_46[11:0] ? image_586 : _GEN_648; // @[Filter.scala 138:46]
  wire [3:0] _GEN_650 = 12'h24b == _T_46[11:0] ? image_587 : _GEN_649; // @[Filter.scala 138:46]
  wire [3:0] _GEN_651 = 12'h24c == _T_46[11:0] ? image_588 : _GEN_650; // @[Filter.scala 138:46]
  wire [3:0] _GEN_652 = 12'h24d == _T_46[11:0] ? image_589 : _GEN_651; // @[Filter.scala 138:46]
  wire [3:0] _GEN_653 = 12'h24e == _T_46[11:0] ? image_590 : _GEN_652; // @[Filter.scala 138:46]
  wire [3:0] _GEN_654 = 12'h24f == _T_46[11:0] ? image_591 : _GEN_653; // @[Filter.scala 138:46]
  wire [3:0] _GEN_655 = 12'h250 == _T_46[11:0] ? image_592 : _GEN_654; // @[Filter.scala 138:46]
  wire [3:0] _GEN_656 = 12'h251 == _T_46[11:0] ? image_593 : _GEN_655; // @[Filter.scala 138:46]
  wire [3:0] _GEN_657 = 12'h252 == _T_46[11:0] ? image_594 : _GEN_656; // @[Filter.scala 138:46]
  wire [3:0] _GEN_658 = 12'h253 == _T_46[11:0] ? image_595 : _GEN_657; // @[Filter.scala 138:46]
  wire [3:0] _GEN_659 = 12'h254 == _T_46[11:0] ? image_596 : _GEN_658; // @[Filter.scala 138:46]
  wire [3:0] _GEN_660 = 12'h255 == _T_46[11:0] ? image_597 : _GEN_659; // @[Filter.scala 138:46]
  wire [3:0] _GEN_661 = 12'h256 == _T_46[11:0] ? image_598 : _GEN_660; // @[Filter.scala 138:46]
  wire [3:0] _GEN_662 = 12'h257 == _T_46[11:0] ? image_599 : _GEN_661; // @[Filter.scala 138:46]
  wire [3:0] _GEN_663 = 12'h258 == _T_46[11:0] ? image_600 : _GEN_662; // @[Filter.scala 138:46]
  wire [3:0] _GEN_664 = 12'h259 == _T_46[11:0] ? image_601 : _GEN_663; // @[Filter.scala 138:46]
  wire [3:0] _GEN_665 = 12'h25a == _T_46[11:0] ? image_602 : _GEN_664; // @[Filter.scala 138:46]
  wire [3:0] _GEN_666 = 12'h25b == _T_46[11:0] ? image_603 : _GEN_665; // @[Filter.scala 138:46]
  wire [3:0] _GEN_667 = 12'h25c == _T_46[11:0] ? image_604 : _GEN_666; // @[Filter.scala 138:46]
  wire [3:0] _GEN_668 = 12'h25d == _T_46[11:0] ? image_605 : _GEN_667; // @[Filter.scala 138:46]
  wire [3:0] _GEN_669 = 12'h25e == _T_46[11:0] ? image_606 : _GEN_668; // @[Filter.scala 138:46]
  wire [3:0] _GEN_670 = 12'h25f == _T_46[11:0] ? image_607 : _GEN_669; // @[Filter.scala 138:46]
  wire [3:0] _GEN_671 = 12'h260 == _T_46[11:0] ? 4'h0 : _GEN_670; // @[Filter.scala 138:46]
  wire [3:0] _GEN_672 = 12'h261 == _T_46[11:0] ? 4'h0 : _GEN_671; // @[Filter.scala 138:46]
  wire [3:0] _GEN_673 = 12'h262 == _T_46[11:0] ? 4'h0 : _GEN_672; // @[Filter.scala 138:46]
  wire [3:0] _GEN_674 = 12'h263 == _T_46[11:0] ? 4'h0 : _GEN_673; // @[Filter.scala 138:46]
  wire [3:0] _GEN_675 = 12'h264 == _T_46[11:0] ? 4'h0 : _GEN_674; // @[Filter.scala 138:46]
  wire [3:0] _GEN_676 = 12'h265 == _T_46[11:0] ? 4'h0 : _GEN_675; // @[Filter.scala 138:46]
  wire [3:0] _GEN_677 = 12'h266 == _T_46[11:0] ? image_614 : _GEN_676; // @[Filter.scala 138:46]
  wire [3:0] _GEN_678 = 12'h267 == _T_46[11:0] ? image_615 : _GEN_677; // @[Filter.scala 138:46]
  wire [3:0] _GEN_679 = 12'h268 == _T_46[11:0] ? image_616 : _GEN_678; // @[Filter.scala 138:46]
  wire [3:0] _GEN_680 = 12'h269 == _T_46[11:0] ? image_617 : _GEN_679; // @[Filter.scala 138:46]
  wire [3:0] _GEN_681 = 12'h26a == _T_46[11:0] ? image_618 : _GEN_680; // @[Filter.scala 138:46]
  wire [3:0] _GEN_682 = 12'h26b == _T_46[11:0] ? image_619 : _GEN_681; // @[Filter.scala 138:46]
  wire [3:0] _GEN_683 = 12'h26c == _T_46[11:0] ? image_620 : _GEN_682; // @[Filter.scala 138:46]
  wire [3:0] _GEN_684 = 12'h26d == _T_46[11:0] ? image_621 : _GEN_683; // @[Filter.scala 138:46]
  wire [3:0] _GEN_685 = 12'h26e == _T_46[11:0] ? image_622 : _GEN_684; // @[Filter.scala 138:46]
  wire [3:0] _GEN_686 = 12'h26f == _T_46[11:0] ? image_623 : _GEN_685; // @[Filter.scala 138:46]
  wire [3:0] _GEN_687 = 12'h270 == _T_46[11:0] ? image_624 : _GEN_686; // @[Filter.scala 138:46]
  wire [3:0] _GEN_688 = 12'h271 == _T_46[11:0] ? image_625 : _GEN_687; // @[Filter.scala 138:46]
  wire [3:0] _GEN_689 = 12'h272 == _T_46[11:0] ? image_626 : _GEN_688; // @[Filter.scala 138:46]
  wire [3:0] _GEN_690 = 12'h273 == _T_46[11:0] ? image_627 : _GEN_689; // @[Filter.scala 138:46]
  wire [3:0] _GEN_691 = 12'h274 == _T_46[11:0] ? image_628 : _GEN_690; // @[Filter.scala 138:46]
  wire [3:0] _GEN_692 = 12'h275 == _T_46[11:0] ? 4'h0 : _GEN_691; // @[Filter.scala 138:46]
  wire [3:0] _GEN_693 = 12'h276 == _T_46[11:0] ? 4'h0 : _GEN_692; // @[Filter.scala 138:46]
  wire [3:0] _GEN_694 = 12'h277 == _T_46[11:0] ? 4'h0 : _GEN_693; // @[Filter.scala 138:46]
  wire [3:0] _GEN_695 = 12'h278 == _T_46[11:0] ? 4'h0 : _GEN_694; // @[Filter.scala 138:46]
  wire [3:0] _GEN_696 = 12'h279 == _T_46[11:0] ? 4'h0 : _GEN_695; // @[Filter.scala 138:46]
  wire [3:0] _GEN_697 = 12'h27a == _T_46[11:0] ? 4'h0 : _GEN_696; // @[Filter.scala 138:46]
  wire [3:0] _GEN_698 = 12'h27b == _T_46[11:0] ? 4'h0 : _GEN_697; // @[Filter.scala 138:46]
  wire [3:0] _GEN_699 = 12'h27c == _T_46[11:0] ? image_636 : _GEN_698; // @[Filter.scala 138:46]
  wire [3:0] _GEN_700 = 12'h27d == _T_46[11:0] ? image_637 : _GEN_699; // @[Filter.scala 138:46]
  wire [3:0] _GEN_701 = 12'h27e == _T_46[11:0] ? image_638 : _GEN_700; // @[Filter.scala 138:46]
  wire [3:0] _GEN_702 = 12'h27f == _T_46[11:0] ? image_639 : _GEN_701; // @[Filter.scala 138:46]
  wire [3:0] _GEN_703 = 12'h280 == _T_46[11:0] ? 4'h0 : _GEN_702; // @[Filter.scala 138:46]
  wire [3:0] _GEN_704 = 12'h281 == _T_46[11:0] ? 4'h0 : _GEN_703; // @[Filter.scala 138:46]
  wire [3:0] _GEN_705 = 12'h282 == _T_46[11:0] ? image_642 : _GEN_704; // @[Filter.scala 138:46]
  wire [3:0] _GEN_706 = 12'h283 == _T_46[11:0] ? image_643 : _GEN_705; // @[Filter.scala 138:46]
  wire [3:0] _GEN_707 = 12'h284 == _T_46[11:0] ? image_644 : _GEN_706; // @[Filter.scala 138:46]
  wire [3:0] _GEN_708 = 12'h285 == _T_46[11:0] ? image_645 : _GEN_707; // @[Filter.scala 138:46]
  wire [3:0] _GEN_709 = 12'h286 == _T_46[11:0] ? image_646 : _GEN_708; // @[Filter.scala 138:46]
  wire [3:0] _GEN_710 = 12'h287 == _T_46[11:0] ? image_647 : _GEN_709; // @[Filter.scala 138:46]
  wire [3:0] _GEN_711 = 12'h288 == _T_46[11:0] ? image_648 : _GEN_710; // @[Filter.scala 138:46]
  wire [3:0] _GEN_712 = 12'h289 == _T_46[11:0] ? image_649 : _GEN_711; // @[Filter.scala 138:46]
  wire [3:0] _GEN_713 = 12'h28a == _T_46[11:0] ? image_650 : _GEN_712; // @[Filter.scala 138:46]
  wire [3:0] _GEN_714 = 12'h28b == _T_46[11:0] ? image_651 : _GEN_713; // @[Filter.scala 138:46]
  wire [3:0] _GEN_715 = 12'h28c == _T_46[11:0] ? image_652 : _GEN_714; // @[Filter.scala 138:46]
  wire [3:0] _GEN_716 = 12'h28d == _T_46[11:0] ? image_653 : _GEN_715; // @[Filter.scala 138:46]
  wire [3:0] _GEN_717 = 12'h28e == _T_46[11:0] ? image_654 : _GEN_716; // @[Filter.scala 138:46]
  wire [3:0] _GEN_718 = 12'h28f == _T_46[11:0] ? image_655 : _GEN_717; // @[Filter.scala 138:46]
  wire [3:0] _GEN_719 = 12'h290 == _T_46[11:0] ? image_656 : _GEN_718; // @[Filter.scala 138:46]
  wire [3:0] _GEN_720 = 12'h291 == _T_46[11:0] ? image_657 : _GEN_719; // @[Filter.scala 138:46]
  wire [3:0] _GEN_721 = 12'h292 == _T_46[11:0] ? image_658 : _GEN_720; // @[Filter.scala 138:46]
  wire [3:0] _GEN_722 = 12'h293 == _T_46[11:0] ? image_659 : _GEN_721; // @[Filter.scala 138:46]
  wire [3:0] _GEN_723 = 12'h294 == _T_46[11:0] ? image_660 : _GEN_722; // @[Filter.scala 138:46]
  wire [3:0] _GEN_724 = 12'h295 == _T_46[11:0] ? image_661 : _GEN_723; // @[Filter.scala 138:46]
  wire [3:0] _GEN_725 = 12'h296 == _T_46[11:0] ? image_662 : _GEN_724; // @[Filter.scala 138:46]
  wire [3:0] _GEN_726 = 12'h297 == _T_46[11:0] ? image_663 : _GEN_725; // @[Filter.scala 138:46]
  wire [3:0] _GEN_727 = 12'h298 == _T_46[11:0] ? image_664 : _GEN_726; // @[Filter.scala 138:46]
  wire [3:0] _GEN_728 = 12'h299 == _T_46[11:0] ? image_665 : _GEN_727; // @[Filter.scala 138:46]
  wire [3:0] _GEN_729 = 12'h29a == _T_46[11:0] ? image_666 : _GEN_728; // @[Filter.scala 138:46]
  wire [3:0] _GEN_730 = 12'h29b == _T_46[11:0] ? image_667 : _GEN_729; // @[Filter.scala 138:46]
  wire [3:0] _GEN_731 = 12'h29c == _T_46[11:0] ? image_668 : _GEN_730; // @[Filter.scala 138:46]
  wire [3:0] _GEN_732 = 12'h29d == _T_46[11:0] ? image_669 : _GEN_731; // @[Filter.scala 138:46]
  wire [3:0] _GEN_733 = 12'h29e == _T_46[11:0] ? image_670 : _GEN_732; // @[Filter.scala 138:46]
  wire [3:0] _GEN_734 = 12'h29f == _T_46[11:0] ? 4'h0 : _GEN_733; // @[Filter.scala 138:46]
  wire [3:0] _GEN_735 = 12'h2a0 == _T_46[11:0] ? 4'h0 : _GEN_734; // @[Filter.scala 138:46]
  wire [3:0] _GEN_736 = 12'h2a1 == _T_46[11:0] ? 4'h0 : _GEN_735; // @[Filter.scala 138:46]
  wire [3:0] _GEN_737 = 12'h2a2 == _T_46[11:0] ? 4'h0 : _GEN_736; // @[Filter.scala 138:46]
  wire [3:0] _GEN_738 = 12'h2a3 == _T_46[11:0] ? 4'h0 : _GEN_737; // @[Filter.scala 138:46]
  wire [3:0] _GEN_739 = 12'h2a4 == _T_46[11:0] ? 4'h0 : _GEN_738; // @[Filter.scala 138:46]
  wire [3:0] _GEN_740 = 12'h2a5 == _T_46[11:0] ? 4'h0 : _GEN_739; // @[Filter.scala 138:46]
  wire [3:0] _GEN_741 = 12'h2a6 == _T_46[11:0] ? 4'h0 : _GEN_740; // @[Filter.scala 138:46]
  wire [3:0] _GEN_742 = 12'h2a7 == _T_46[11:0] ? image_679 : _GEN_741; // @[Filter.scala 138:46]
  wire [3:0] _GEN_743 = 12'h2a8 == _T_46[11:0] ? image_680 : _GEN_742; // @[Filter.scala 138:46]
  wire [3:0] _GEN_744 = 12'h2a9 == _T_46[11:0] ? image_681 : _GEN_743; // @[Filter.scala 138:46]
  wire [3:0] _GEN_745 = 12'h2aa == _T_46[11:0] ? image_682 : _GEN_744; // @[Filter.scala 138:46]
  wire [3:0] _GEN_746 = 12'h2ab == _T_46[11:0] ? image_683 : _GEN_745; // @[Filter.scala 138:46]
  wire [3:0] _GEN_747 = 12'h2ac == _T_46[11:0] ? image_684 : _GEN_746; // @[Filter.scala 138:46]
  wire [3:0] _GEN_748 = 12'h2ad == _T_46[11:0] ? image_685 : _GEN_747; // @[Filter.scala 138:46]
  wire [3:0] _GEN_749 = 12'h2ae == _T_46[11:0] ? image_686 : _GEN_748; // @[Filter.scala 138:46]
  wire [3:0] _GEN_750 = 12'h2af == _T_46[11:0] ? image_687 : _GEN_749; // @[Filter.scala 138:46]
  wire [3:0] _GEN_751 = 12'h2b0 == _T_46[11:0] ? image_688 : _GEN_750; // @[Filter.scala 138:46]
  wire [3:0] _GEN_752 = 12'h2b1 == _T_46[11:0] ? image_689 : _GEN_751; // @[Filter.scala 138:46]
  wire [3:0] _GEN_753 = 12'h2b2 == _T_46[11:0] ? image_690 : _GEN_752; // @[Filter.scala 138:46]
  wire [3:0] _GEN_754 = 12'h2b3 == _T_46[11:0] ? image_691 : _GEN_753; // @[Filter.scala 138:46]
  wire [3:0] _GEN_755 = 12'h2b4 == _T_46[11:0] ? image_692 : _GEN_754; // @[Filter.scala 138:46]
  wire [3:0] _GEN_756 = 12'h2b5 == _T_46[11:0] ? image_693 : _GEN_755; // @[Filter.scala 138:46]
  wire [3:0] _GEN_757 = 12'h2b6 == _T_46[11:0] ? image_694 : _GEN_756; // @[Filter.scala 138:46]
  wire [3:0] _GEN_758 = 12'h2b7 == _T_46[11:0] ? image_695 : _GEN_757; // @[Filter.scala 138:46]
  wire [3:0] _GEN_759 = 12'h2b8 == _T_46[11:0] ? image_696 : _GEN_758; // @[Filter.scala 138:46]
  wire [3:0] _GEN_760 = 12'h2b9 == _T_46[11:0] ? image_697 : _GEN_759; // @[Filter.scala 138:46]
  wire [3:0] _GEN_761 = 12'h2ba == _T_46[11:0] ? image_698 : _GEN_760; // @[Filter.scala 138:46]
  wire [3:0] _GEN_762 = 12'h2bb == _T_46[11:0] ? 4'h0 : _GEN_761; // @[Filter.scala 138:46]
  wire [3:0] _GEN_763 = 12'h2bc == _T_46[11:0] ? 4'h0 : _GEN_762; // @[Filter.scala 138:46]
  wire [3:0] _GEN_764 = 12'h2bd == _T_46[11:0] ? image_701 : _GEN_763; // @[Filter.scala 138:46]
  wire [3:0] _GEN_765 = 12'h2be == _T_46[11:0] ? image_702 : _GEN_764; // @[Filter.scala 138:46]
  wire [3:0] _GEN_766 = 12'h2bf == _T_46[11:0] ? image_703 : _GEN_765; // @[Filter.scala 138:46]
  wire [3:0] _GEN_767 = 12'h2c0 == _T_46[11:0] ? 4'h0 : _GEN_766; // @[Filter.scala 138:46]
  wire [3:0] _GEN_768 = 12'h2c1 == _T_46[11:0] ? image_705 : _GEN_767; // @[Filter.scala 138:46]
  wire [3:0] _GEN_769 = 12'h2c2 == _T_46[11:0] ? image_706 : _GEN_768; // @[Filter.scala 138:46]
  wire [3:0] _GEN_770 = 12'h2c3 == _T_46[11:0] ? image_707 : _GEN_769; // @[Filter.scala 138:46]
  wire [3:0] _GEN_771 = 12'h2c4 == _T_46[11:0] ? image_708 : _GEN_770; // @[Filter.scala 138:46]
  wire [3:0] _GEN_772 = 12'h2c5 == _T_46[11:0] ? image_709 : _GEN_771; // @[Filter.scala 138:46]
  wire [3:0] _GEN_773 = 12'h2c6 == _T_46[11:0] ? image_710 : _GEN_772; // @[Filter.scala 138:46]
  wire [3:0] _GEN_774 = 12'h2c7 == _T_46[11:0] ? image_711 : _GEN_773; // @[Filter.scala 138:46]
  wire [3:0] _GEN_775 = 12'h2c8 == _T_46[11:0] ? image_712 : _GEN_774; // @[Filter.scala 138:46]
  wire [3:0] _GEN_776 = 12'h2c9 == _T_46[11:0] ? image_713 : _GEN_775; // @[Filter.scala 138:46]
  wire [3:0] _GEN_777 = 12'h2ca == _T_46[11:0] ? image_714 : _GEN_776; // @[Filter.scala 138:46]
  wire [3:0] _GEN_778 = 12'h2cb == _T_46[11:0] ? image_715 : _GEN_777; // @[Filter.scala 138:46]
  wire [3:0] _GEN_779 = 12'h2cc == _T_46[11:0] ? image_716 : _GEN_778; // @[Filter.scala 138:46]
  wire [3:0] _GEN_780 = 12'h2cd == _T_46[11:0] ? image_717 : _GEN_779; // @[Filter.scala 138:46]
  wire [3:0] _GEN_781 = 12'h2ce == _T_46[11:0] ? image_718 : _GEN_780; // @[Filter.scala 138:46]
  wire [3:0] _GEN_782 = 12'h2cf == _T_46[11:0] ? image_719 : _GEN_781; // @[Filter.scala 138:46]
  wire [3:0] _GEN_783 = 12'h2d0 == _T_46[11:0] ? image_720 : _GEN_782; // @[Filter.scala 138:46]
  wire [3:0] _GEN_784 = 12'h2d1 == _T_46[11:0] ? image_721 : _GEN_783; // @[Filter.scala 138:46]
  wire [3:0] _GEN_785 = 12'h2d2 == _T_46[11:0] ? image_722 : _GEN_784; // @[Filter.scala 138:46]
  wire [3:0] _GEN_786 = 12'h2d3 == _T_46[11:0] ? image_723 : _GEN_785; // @[Filter.scala 138:46]
  wire [3:0] _GEN_787 = 12'h2d4 == _T_46[11:0] ? image_724 : _GEN_786; // @[Filter.scala 138:46]
  wire [3:0] _GEN_788 = 12'h2d5 == _T_46[11:0] ? image_725 : _GEN_787; // @[Filter.scala 138:46]
  wire [3:0] _GEN_789 = 12'h2d6 == _T_46[11:0] ? image_726 : _GEN_788; // @[Filter.scala 138:46]
  wire [3:0] _GEN_790 = 12'h2d7 == _T_46[11:0] ? image_727 : _GEN_789; // @[Filter.scala 138:46]
  wire [3:0] _GEN_791 = 12'h2d8 == _T_46[11:0] ? image_728 : _GEN_790; // @[Filter.scala 138:46]
  wire [3:0] _GEN_792 = 12'h2d9 == _T_46[11:0] ? image_729 : _GEN_791; // @[Filter.scala 138:46]
  wire [3:0] _GEN_793 = 12'h2da == _T_46[11:0] ? image_730 : _GEN_792; // @[Filter.scala 138:46]
  wire [3:0] _GEN_794 = 12'h2db == _T_46[11:0] ? image_731 : _GEN_793; // @[Filter.scala 138:46]
  wire [3:0] _GEN_795 = 12'h2dc == _T_46[11:0] ? image_732 : _GEN_794; // @[Filter.scala 138:46]
  wire [3:0] _GEN_796 = 12'h2dd == _T_46[11:0] ? image_733 : _GEN_795; // @[Filter.scala 138:46]
  wire [3:0] _GEN_797 = 12'h2de == _T_46[11:0] ? image_734 : _GEN_796; // @[Filter.scala 138:46]
  wire [3:0] _GEN_798 = 12'h2df == _T_46[11:0] ? 4'h0 : _GEN_797; // @[Filter.scala 138:46]
  wire [3:0] _GEN_799 = 12'h2e0 == _T_46[11:0] ? image_736 : _GEN_798; // @[Filter.scala 138:46]
  wire [3:0] _GEN_800 = 12'h2e1 == _T_46[11:0] ? image_737 : _GEN_799; // @[Filter.scala 138:46]
  wire [3:0] _GEN_801 = 12'h2e2 == _T_46[11:0] ? 4'h0 : _GEN_800; // @[Filter.scala 138:46]
  wire [3:0] _GEN_802 = 12'h2e3 == _T_46[11:0] ? image_739 : _GEN_801; // @[Filter.scala 138:46]
  wire [3:0] _GEN_803 = 12'h2e4 == _T_46[11:0] ? image_740 : _GEN_802; // @[Filter.scala 138:46]
  wire [3:0] _GEN_804 = 12'h2e5 == _T_46[11:0] ? image_741 : _GEN_803; // @[Filter.scala 138:46]
  wire [3:0] _GEN_805 = 12'h2e6 == _T_46[11:0] ? 4'h0 : _GEN_804; // @[Filter.scala 138:46]
  wire [3:0] _GEN_806 = 12'h2e7 == _T_46[11:0] ? 4'h0 : _GEN_805; // @[Filter.scala 138:46]
  wire [3:0] _GEN_807 = 12'h2e8 == _T_46[11:0] ? image_744 : _GEN_806; // @[Filter.scala 138:46]
  wire [3:0] _GEN_808 = 12'h2e9 == _T_46[11:0] ? image_745 : _GEN_807; // @[Filter.scala 138:46]
  wire [3:0] _GEN_809 = 12'h2ea == _T_46[11:0] ? image_746 : _GEN_808; // @[Filter.scala 138:46]
  wire [3:0] _GEN_810 = 12'h2eb == _T_46[11:0] ? image_747 : _GEN_809; // @[Filter.scala 138:46]
  wire [3:0] _GEN_811 = 12'h2ec == _T_46[11:0] ? image_748 : _GEN_810; // @[Filter.scala 138:46]
  wire [3:0] _GEN_812 = 12'h2ed == _T_46[11:0] ? image_749 : _GEN_811; // @[Filter.scala 138:46]
  wire [3:0] _GEN_813 = 12'h2ee == _T_46[11:0] ? image_750 : _GEN_812; // @[Filter.scala 138:46]
  wire [3:0] _GEN_814 = 12'h2ef == _T_46[11:0] ? image_751 : _GEN_813; // @[Filter.scala 138:46]
  wire [3:0] _GEN_815 = 12'h2f0 == _T_46[11:0] ? image_752 : _GEN_814; // @[Filter.scala 138:46]
  wire [3:0] _GEN_816 = 12'h2f1 == _T_46[11:0] ? image_753 : _GEN_815; // @[Filter.scala 138:46]
  wire [3:0] _GEN_817 = 12'h2f2 == _T_46[11:0] ? image_754 : _GEN_816; // @[Filter.scala 138:46]
  wire [3:0] _GEN_818 = 12'h2f3 == _T_46[11:0] ? image_755 : _GEN_817; // @[Filter.scala 138:46]
  wire [3:0] _GEN_819 = 12'h2f4 == _T_46[11:0] ? image_756 : _GEN_818; // @[Filter.scala 138:46]
  wire [3:0] _GEN_820 = 12'h2f5 == _T_46[11:0] ? 4'h0 : _GEN_819; // @[Filter.scala 138:46]
  wire [3:0] _GEN_821 = 12'h2f6 == _T_46[11:0] ? image_758 : _GEN_820; // @[Filter.scala 138:46]
  wire [3:0] _GEN_822 = 12'h2f7 == _T_46[11:0] ? 4'h0 : _GEN_821; // @[Filter.scala 138:46]
  wire [3:0] _GEN_823 = 12'h2f8 == _T_46[11:0] ? image_760 : _GEN_822; // @[Filter.scala 138:46]
  wire [3:0] _GEN_824 = 12'h2f9 == _T_46[11:0] ? image_761 : _GEN_823; // @[Filter.scala 138:46]
  wire [3:0] _GEN_825 = 12'h2fa == _T_46[11:0] ? image_762 : _GEN_824; // @[Filter.scala 138:46]
  wire [3:0] _GEN_826 = 12'h2fb == _T_46[11:0] ? image_763 : _GEN_825; // @[Filter.scala 138:46]
  wire [3:0] _GEN_827 = 12'h2fc == _T_46[11:0] ? 4'h0 : _GEN_826; // @[Filter.scala 138:46]
  wire [3:0] _GEN_828 = 12'h2fd == _T_46[11:0] ? image_765 : _GEN_827; // @[Filter.scala 138:46]
  wire [3:0] _GEN_829 = 12'h2fe == _T_46[11:0] ? image_766 : _GEN_828; // @[Filter.scala 138:46]
  wire [3:0] _GEN_830 = 12'h2ff == _T_46[11:0] ? image_767 : _GEN_829; // @[Filter.scala 138:46]
  wire [3:0] _GEN_831 = 12'h300 == _T_46[11:0] ? image_768 : _GEN_830; // @[Filter.scala 138:46]
  wire [3:0] _GEN_832 = 12'h301 == _T_46[11:0] ? image_769 : _GEN_831; // @[Filter.scala 138:46]
  wire [3:0] _GEN_833 = 12'h302 == _T_46[11:0] ? image_770 : _GEN_832; // @[Filter.scala 138:46]
  wire [3:0] _GEN_834 = 12'h303 == _T_46[11:0] ? image_771 : _GEN_833; // @[Filter.scala 138:46]
  wire [3:0] _GEN_835 = 12'h304 == _T_46[11:0] ? image_772 : _GEN_834; // @[Filter.scala 138:46]
  wire [3:0] _GEN_836 = 12'h305 == _T_46[11:0] ? image_773 : _GEN_835; // @[Filter.scala 138:46]
  wire [3:0] _GEN_837 = 12'h306 == _T_46[11:0] ? image_774 : _GEN_836; // @[Filter.scala 138:46]
  wire [3:0] _GEN_838 = 12'h307 == _T_46[11:0] ? image_775 : _GEN_837; // @[Filter.scala 138:46]
  wire [3:0] _GEN_839 = 12'h308 == _T_46[11:0] ? image_776 : _GEN_838; // @[Filter.scala 138:46]
  wire [3:0] _GEN_840 = 12'h309 == _T_46[11:0] ? image_777 : _GEN_839; // @[Filter.scala 138:46]
  wire [3:0] _GEN_841 = 12'h30a == _T_46[11:0] ? image_778 : _GEN_840; // @[Filter.scala 138:46]
  wire [3:0] _GEN_842 = 12'h30b == _T_46[11:0] ? image_779 : _GEN_841; // @[Filter.scala 138:46]
  wire [3:0] _GEN_843 = 12'h30c == _T_46[11:0] ? image_780 : _GEN_842; // @[Filter.scala 138:46]
  wire [3:0] _GEN_844 = 12'h30d == _T_46[11:0] ? image_781 : _GEN_843; // @[Filter.scala 138:46]
  wire [3:0] _GEN_845 = 12'h30e == _T_46[11:0] ? image_782 : _GEN_844; // @[Filter.scala 138:46]
  wire [3:0] _GEN_846 = 12'h30f == _T_46[11:0] ? image_783 : _GEN_845; // @[Filter.scala 138:46]
  wire [3:0] _GEN_847 = 12'h310 == _T_46[11:0] ? image_784 : _GEN_846; // @[Filter.scala 138:46]
  wire [3:0] _GEN_848 = 12'h311 == _T_46[11:0] ? image_785 : _GEN_847; // @[Filter.scala 138:46]
  wire [3:0] _GEN_849 = 12'h312 == _T_46[11:0] ? image_786 : _GEN_848; // @[Filter.scala 138:46]
  wire [3:0] _GEN_850 = 12'h313 == _T_46[11:0] ? image_787 : _GEN_849; // @[Filter.scala 138:46]
  wire [3:0] _GEN_851 = 12'h314 == _T_46[11:0] ? image_788 : _GEN_850; // @[Filter.scala 138:46]
  wire [3:0] _GEN_852 = 12'h315 == _T_46[11:0] ? image_789 : _GEN_851; // @[Filter.scala 138:46]
  wire [3:0] _GEN_853 = 12'h316 == _T_46[11:0] ? image_790 : _GEN_852; // @[Filter.scala 138:46]
  wire [3:0] _GEN_854 = 12'h317 == _T_46[11:0] ? image_791 : _GEN_853; // @[Filter.scala 138:46]
  wire [3:0] _GEN_855 = 12'h318 == _T_46[11:0] ? image_792 : _GEN_854; // @[Filter.scala 138:46]
  wire [3:0] _GEN_856 = 12'h319 == _T_46[11:0] ? image_793 : _GEN_855; // @[Filter.scala 138:46]
  wire [3:0] _GEN_857 = 12'h31a == _T_46[11:0] ? image_794 : _GEN_856; // @[Filter.scala 138:46]
  wire [3:0] _GEN_858 = 12'h31b == _T_46[11:0] ? image_795 : _GEN_857; // @[Filter.scala 138:46]
  wire [3:0] _GEN_859 = 12'h31c == _T_46[11:0] ? image_796 : _GEN_858; // @[Filter.scala 138:46]
  wire [3:0] _GEN_860 = 12'h31d == _T_46[11:0] ? image_797 : _GEN_859; // @[Filter.scala 138:46]
  wire [3:0] _GEN_861 = 12'h31e == _T_46[11:0] ? 4'h0 : _GEN_860; // @[Filter.scala 138:46]
  wire [3:0] _GEN_862 = 12'h31f == _T_46[11:0] ? 4'h0 : _GEN_861; // @[Filter.scala 138:46]
  wire [3:0] _GEN_863 = 12'h320 == _T_46[11:0] ? image_800 : _GEN_862; // @[Filter.scala 138:46]
  wire [3:0] _GEN_864 = 12'h321 == _T_46[11:0] ? image_801 : _GEN_863; // @[Filter.scala 138:46]
  wire [3:0] _GEN_865 = 12'h322 == _T_46[11:0] ? image_802 : _GEN_864; // @[Filter.scala 138:46]
  wire [3:0] _GEN_866 = 12'h323 == _T_46[11:0] ? image_803 : _GEN_865; // @[Filter.scala 138:46]
  wire [3:0] _GEN_867 = 12'h324 == _T_46[11:0] ? image_804 : _GEN_866; // @[Filter.scala 138:46]
  wire [3:0] _GEN_868 = 12'h325 == _T_46[11:0] ? image_805 : _GEN_867; // @[Filter.scala 138:46]
  wire [3:0] _GEN_869 = 12'h326 == _T_46[11:0] ? image_806 : _GEN_868; // @[Filter.scala 138:46]
  wire [3:0] _GEN_870 = 12'h327 == _T_46[11:0] ? 4'h0 : _GEN_869; // @[Filter.scala 138:46]
  wire [3:0] _GEN_871 = 12'h328 == _T_46[11:0] ? image_808 : _GEN_870; // @[Filter.scala 138:46]
  wire [3:0] _GEN_872 = 12'h329 == _T_46[11:0] ? image_809 : _GEN_871; // @[Filter.scala 138:46]
  wire [3:0] _GEN_873 = 12'h32a == _T_46[11:0] ? image_810 : _GEN_872; // @[Filter.scala 138:46]
  wire [3:0] _GEN_874 = 12'h32b == _T_46[11:0] ? image_811 : _GEN_873; // @[Filter.scala 138:46]
  wire [3:0] _GEN_875 = 12'h32c == _T_46[11:0] ? image_812 : _GEN_874; // @[Filter.scala 138:46]
  wire [3:0] _GEN_876 = 12'h32d == _T_46[11:0] ? image_813 : _GEN_875; // @[Filter.scala 138:46]
  wire [3:0] _GEN_877 = 12'h32e == _T_46[11:0] ? image_814 : _GEN_876; // @[Filter.scala 138:46]
  wire [3:0] _GEN_878 = 12'h32f == _T_46[11:0] ? image_815 : _GEN_877; // @[Filter.scala 138:46]
  wire [3:0] _GEN_879 = 12'h330 == _T_46[11:0] ? image_816 : _GEN_878; // @[Filter.scala 138:46]
  wire [3:0] _GEN_880 = 12'h331 == _T_46[11:0] ? image_817 : _GEN_879; // @[Filter.scala 138:46]
  wire [3:0] _GEN_881 = 12'h332 == _T_46[11:0] ? image_818 : _GEN_880; // @[Filter.scala 138:46]
  wire [3:0] _GEN_882 = 12'h333 == _T_46[11:0] ? image_819 : _GEN_881; // @[Filter.scala 138:46]
  wire [3:0] _GEN_883 = 12'h334 == _T_46[11:0] ? image_820 : _GEN_882; // @[Filter.scala 138:46]
  wire [3:0] _GEN_884 = 12'h335 == _T_46[11:0] ? 4'h0 : _GEN_883; // @[Filter.scala 138:46]
  wire [3:0] _GEN_885 = 12'h336 == _T_46[11:0] ? image_822 : _GEN_884; // @[Filter.scala 138:46]
  wire [3:0] _GEN_886 = 12'h337 == _T_46[11:0] ? image_823 : _GEN_885; // @[Filter.scala 138:46]
  wire [3:0] _GEN_887 = 12'h338 == _T_46[11:0] ? image_824 : _GEN_886; // @[Filter.scala 138:46]
  wire [3:0] _GEN_888 = 12'h339 == _T_46[11:0] ? image_825 : _GEN_887; // @[Filter.scala 138:46]
  wire [3:0] _GEN_889 = 12'h33a == _T_46[11:0] ? image_826 : _GEN_888; // @[Filter.scala 138:46]
  wire [3:0] _GEN_890 = 12'h33b == _T_46[11:0] ? 4'h0 : _GEN_889; // @[Filter.scala 138:46]
  wire [3:0] _GEN_891 = 12'h33c == _T_46[11:0] ? image_828 : _GEN_890; // @[Filter.scala 138:46]
  wire [3:0] _GEN_892 = 12'h33d == _T_46[11:0] ? image_829 : _GEN_891; // @[Filter.scala 138:46]
  wire [3:0] _GEN_893 = 12'h33e == _T_46[11:0] ? image_830 : _GEN_892; // @[Filter.scala 138:46]
  wire [3:0] _GEN_894 = 12'h33f == _T_46[11:0] ? image_831 : _GEN_893; // @[Filter.scala 138:46]
  wire [3:0] _GEN_895 = 12'h340 == _T_46[11:0] ? 4'h0 : _GEN_894; // @[Filter.scala 138:46]
  wire [3:0] _GEN_896 = 12'h341 == _T_46[11:0] ? image_833 : _GEN_895; // @[Filter.scala 138:46]
  wire [3:0] _GEN_897 = 12'h342 == _T_46[11:0] ? image_834 : _GEN_896; // @[Filter.scala 138:46]
  wire [3:0] _GEN_898 = 12'h343 == _T_46[11:0] ? image_835 : _GEN_897; // @[Filter.scala 138:46]
  wire [3:0] _GEN_899 = 12'h344 == _T_46[11:0] ? image_836 : _GEN_898; // @[Filter.scala 138:46]
  wire [3:0] _GEN_900 = 12'h345 == _T_46[11:0] ? image_837 : _GEN_899; // @[Filter.scala 138:46]
  wire [3:0] _GEN_901 = 12'h346 == _T_46[11:0] ? image_838 : _GEN_900; // @[Filter.scala 138:46]
  wire [3:0] _GEN_902 = 12'h347 == _T_46[11:0] ? image_839 : _GEN_901; // @[Filter.scala 138:46]
  wire [3:0] _GEN_903 = 12'h348 == _T_46[11:0] ? image_840 : _GEN_902; // @[Filter.scala 138:46]
  wire [3:0] _GEN_904 = 12'h349 == _T_46[11:0] ? image_841 : _GEN_903; // @[Filter.scala 138:46]
  wire [3:0] _GEN_905 = 12'h34a == _T_46[11:0] ? image_842 : _GEN_904; // @[Filter.scala 138:46]
  wire [3:0] _GEN_906 = 12'h34b == _T_46[11:0] ? image_843 : _GEN_905; // @[Filter.scala 138:46]
  wire [3:0] _GEN_907 = 12'h34c == _T_46[11:0] ? image_844 : _GEN_906; // @[Filter.scala 138:46]
  wire [3:0] _GEN_908 = 12'h34d == _T_46[11:0] ? image_845 : _GEN_907; // @[Filter.scala 138:46]
  wire [3:0] _GEN_909 = 12'h34e == _T_46[11:0] ? image_846 : _GEN_908; // @[Filter.scala 138:46]
  wire [3:0] _GEN_910 = 12'h34f == _T_46[11:0] ? image_847 : _GEN_909; // @[Filter.scala 138:46]
  wire [3:0] _GEN_911 = 12'h350 == _T_46[11:0] ? image_848 : _GEN_910; // @[Filter.scala 138:46]
  wire [3:0] _GEN_912 = 12'h351 == _T_46[11:0] ? image_849 : _GEN_911; // @[Filter.scala 138:46]
  wire [3:0] _GEN_913 = 12'h352 == _T_46[11:0] ? image_850 : _GEN_912; // @[Filter.scala 138:46]
  wire [3:0] _GEN_914 = 12'h353 == _T_46[11:0] ? image_851 : _GEN_913; // @[Filter.scala 138:46]
  wire [3:0] _GEN_915 = 12'h354 == _T_46[11:0] ? image_852 : _GEN_914; // @[Filter.scala 138:46]
  wire [3:0] _GEN_916 = 12'h355 == _T_46[11:0] ? image_853 : _GEN_915; // @[Filter.scala 138:46]
  wire [3:0] _GEN_917 = 12'h356 == _T_46[11:0] ? image_854 : _GEN_916; // @[Filter.scala 138:46]
  wire [3:0] _GEN_918 = 12'h357 == _T_46[11:0] ? image_855 : _GEN_917; // @[Filter.scala 138:46]
  wire [3:0] _GEN_919 = 12'h358 == _T_46[11:0] ? image_856 : _GEN_918; // @[Filter.scala 138:46]
  wire [3:0] _GEN_920 = 12'h359 == _T_46[11:0] ? image_857 : _GEN_919; // @[Filter.scala 138:46]
  wire [3:0] _GEN_921 = 12'h35a == _T_46[11:0] ? image_858 : _GEN_920; // @[Filter.scala 138:46]
  wire [3:0] _GEN_922 = 12'h35b == _T_46[11:0] ? image_859 : _GEN_921; // @[Filter.scala 138:46]
  wire [3:0] _GEN_923 = 12'h35c == _T_46[11:0] ? image_860 : _GEN_922; // @[Filter.scala 138:46]
  wire [3:0] _GEN_924 = 12'h35d == _T_46[11:0] ? image_861 : _GEN_923; // @[Filter.scala 138:46]
  wire [3:0] _GEN_925 = 12'h35e == _T_46[11:0] ? image_862 : _GEN_924; // @[Filter.scala 138:46]
  wire [3:0] _GEN_926 = 12'h35f == _T_46[11:0] ? 4'h0 : _GEN_925; // @[Filter.scala 138:46]
  wire [3:0] _GEN_927 = 12'h360 == _T_46[11:0] ? 4'h0 : _GEN_926; // @[Filter.scala 138:46]
  wire [3:0] _GEN_928 = 12'h361 == _T_46[11:0] ? image_865 : _GEN_927; // @[Filter.scala 138:46]
  wire [3:0] _GEN_929 = 12'h362 == _T_46[11:0] ? image_866 : _GEN_928; // @[Filter.scala 138:46]
  wire [3:0] _GEN_930 = 12'h363 == _T_46[11:0] ? image_867 : _GEN_929; // @[Filter.scala 138:46]
  wire [3:0] _GEN_931 = 12'h364 == _T_46[11:0] ? image_868 : _GEN_930; // @[Filter.scala 138:46]
  wire [3:0] _GEN_932 = 12'h365 == _T_46[11:0] ? image_869 : _GEN_931; // @[Filter.scala 138:46]
  wire [3:0] _GEN_933 = 12'h366 == _T_46[11:0] ? 4'h0 : _GEN_932; // @[Filter.scala 138:46]
  wire [3:0] _GEN_934 = 12'h367 == _T_46[11:0] ? 4'h0 : _GEN_933; // @[Filter.scala 138:46]
  wire [3:0] _GEN_935 = 12'h368 == _T_46[11:0] ? image_872 : _GEN_934; // @[Filter.scala 138:46]
  wire [3:0] _GEN_936 = 12'h369 == _T_46[11:0] ? image_873 : _GEN_935; // @[Filter.scala 138:46]
  wire [3:0] _GEN_937 = 12'h36a == _T_46[11:0] ? image_874 : _GEN_936; // @[Filter.scala 138:46]
  wire [3:0] _GEN_938 = 12'h36b == _T_46[11:0] ? image_875 : _GEN_937; // @[Filter.scala 138:46]
  wire [3:0] _GEN_939 = 12'h36c == _T_46[11:0] ? image_876 : _GEN_938; // @[Filter.scala 138:46]
  wire [3:0] _GEN_940 = 12'h36d == _T_46[11:0] ? image_877 : _GEN_939; // @[Filter.scala 138:46]
  wire [3:0] _GEN_941 = 12'h36e == _T_46[11:0] ? image_878 : _GEN_940; // @[Filter.scala 138:46]
  wire [3:0] _GEN_942 = 12'h36f == _T_46[11:0] ? image_879 : _GEN_941; // @[Filter.scala 138:46]
  wire [3:0] _GEN_943 = 12'h370 == _T_46[11:0] ? image_880 : _GEN_942; // @[Filter.scala 138:46]
  wire [3:0] _GEN_944 = 12'h371 == _T_46[11:0] ? image_881 : _GEN_943; // @[Filter.scala 138:46]
  wire [3:0] _GEN_945 = 12'h372 == _T_46[11:0] ? image_882 : _GEN_944; // @[Filter.scala 138:46]
  wire [3:0] _GEN_946 = 12'h373 == _T_46[11:0] ? image_883 : _GEN_945; // @[Filter.scala 138:46]
  wire [3:0] _GEN_947 = 12'h374 == _T_46[11:0] ? image_884 : _GEN_946; // @[Filter.scala 138:46]
  wire [3:0] _GEN_948 = 12'h375 == _T_46[11:0] ? image_885 : _GEN_947; // @[Filter.scala 138:46]
  wire [3:0] _GEN_949 = 12'h376 == _T_46[11:0] ? 4'h0 : _GEN_948; // @[Filter.scala 138:46]
  wire [3:0] _GEN_950 = 12'h377 == _T_46[11:0] ? 4'h0 : _GEN_949; // @[Filter.scala 138:46]
  wire [3:0] _GEN_951 = 12'h378 == _T_46[11:0] ? 4'h0 : _GEN_950; // @[Filter.scala 138:46]
  wire [3:0] _GEN_952 = 12'h379 == _T_46[11:0] ? 4'h0 : _GEN_951; // @[Filter.scala 138:46]
  wire [3:0] _GEN_953 = 12'h37a == _T_46[11:0] ? 4'h0 : _GEN_952; // @[Filter.scala 138:46]
  wire [3:0] _GEN_954 = 12'h37b == _T_46[11:0] ? image_891 : _GEN_953; // @[Filter.scala 138:46]
  wire [3:0] _GEN_955 = 12'h37c == _T_46[11:0] ? image_892 : _GEN_954; // @[Filter.scala 138:46]
  wire [3:0] _GEN_956 = 12'h37d == _T_46[11:0] ? image_893 : _GEN_955; // @[Filter.scala 138:46]
  wire [3:0] _GEN_957 = 12'h37e == _T_46[11:0] ? image_894 : _GEN_956; // @[Filter.scala 138:46]
  wire [3:0] _GEN_958 = 12'h37f == _T_46[11:0] ? image_895 : _GEN_957; // @[Filter.scala 138:46]
  wire [3:0] _GEN_959 = 12'h380 == _T_46[11:0] ? 4'h0 : _GEN_958; // @[Filter.scala 138:46]
  wire [3:0] _GEN_960 = 12'h381 == _T_46[11:0] ? image_897 : _GEN_959; // @[Filter.scala 138:46]
  wire [3:0] _GEN_961 = 12'h382 == _T_46[11:0] ? image_898 : _GEN_960; // @[Filter.scala 138:46]
  wire [3:0] _GEN_962 = 12'h383 == _T_46[11:0] ? image_899 : _GEN_961; // @[Filter.scala 138:46]
  wire [3:0] _GEN_963 = 12'h384 == _T_46[11:0] ? image_900 : _GEN_962; // @[Filter.scala 138:46]
  wire [3:0] _GEN_964 = 12'h385 == _T_46[11:0] ? image_901 : _GEN_963; // @[Filter.scala 138:46]
  wire [3:0] _GEN_965 = 12'h386 == _T_46[11:0] ? image_902 : _GEN_964; // @[Filter.scala 138:46]
  wire [3:0] _GEN_966 = 12'h387 == _T_46[11:0] ? image_903 : _GEN_965; // @[Filter.scala 138:46]
  wire [3:0] _GEN_967 = 12'h388 == _T_46[11:0] ? image_904 : _GEN_966; // @[Filter.scala 138:46]
  wire [3:0] _GEN_968 = 12'h389 == _T_46[11:0] ? image_905 : _GEN_967; // @[Filter.scala 138:46]
  wire [3:0] _GEN_969 = 12'h38a == _T_46[11:0] ? image_906 : _GEN_968; // @[Filter.scala 138:46]
  wire [3:0] _GEN_970 = 12'h38b == _T_46[11:0] ? image_907 : _GEN_969; // @[Filter.scala 138:46]
  wire [3:0] _GEN_971 = 12'h38c == _T_46[11:0] ? image_908 : _GEN_970; // @[Filter.scala 138:46]
  wire [3:0] _GEN_972 = 12'h38d == _T_46[11:0] ? image_909 : _GEN_971; // @[Filter.scala 138:46]
  wire [3:0] _GEN_973 = 12'h38e == _T_46[11:0] ? image_910 : _GEN_972; // @[Filter.scala 138:46]
  wire [3:0] _GEN_974 = 12'h38f == _T_46[11:0] ? image_911 : _GEN_973; // @[Filter.scala 138:46]
  wire [3:0] _GEN_975 = 12'h390 == _T_46[11:0] ? image_912 : _GEN_974; // @[Filter.scala 138:46]
  wire [3:0] _GEN_976 = 12'h391 == _T_46[11:0] ? image_913 : _GEN_975; // @[Filter.scala 138:46]
  wire [3:0] _GEN_977 = 12'h392 == _T_46[11:0] ? image_914 : _GEN_976; // @[Filter.scala 138:46]
  wire [3:0] _GEN_978 = 12'h393 == _T_46[11:0] ? image_915 : _GEN_977; // @[Filter.scala 138:46]
  wire [3:0] _GEN_979 = 12'h394 == _T_46[11:0] ? image_916 : _GEN_978; // @[Filter.scala 138:46]
  wire [3:0] _GEN_980 = 12'h395 == _T_46[11:0] ? image_917 : _GEN_979; // @[Filter.scala 138:46]
  wire [3:0] _GEN_981 = 12'h396 == _T_46[11:0] ? image_918 : _GEN_980; // @[Filter.scala 138:46]
  wire [3:0] _GEN_982 = 12'h397 == _T_46[11:0] ? image_919 : _GEN_981; // @[Filter.scala 138:46]
  wire [3:0] _GEN_983 = 12'h398 == _T_46[11:0] ? image_920 : _GEN_982; // @[Filter.scala 138:46]
  wire [3:0] _GEN_984 = 12'h399 == _T_46[11:0] ? image_921 : _GEN_983; // @[Filter.scala 138:46]
  wire [3:0] _GEN_985 = 12'h39a == _T_46[11:0] ? image_922 : _GEN_984; // @[Filter.scala 138:46]
  wire [3:0] _GEN_986 = 12'h39b == _T_46[11:0] ? image_923 : _GEN_985; // @[Filter.scala 138:46]
  wire [3:0] _GEN_987 = 12'h39c == _T_46[11:0] ? image_924 : _GEN_986; // @[Filter.scala 138:46]
  wire [3:0] _GEN_988 = 12'h39d == _T_46[11:0] ? image_925 : _GEN_987; // @[Filter.scala 138:46]
  wire [3:0] _GEN_989 = 12'h39e == _T_46[11:0] ? image_926 : _GEN_988; // @[Filter.scala 138:46]
  wire [3:0] _GEN_990 = 12'h39f == _T_46[11:0] ? image_927 : _GEN_989; // @[Filter.scala 138:46]
  wire [3:0] _GEN_991 = 12'h3a0 == _T_46[11:0] ? 4'h0 : _GEN_990; // @[Filter.scala 138:46]
  wire [3:0] _GEN_992 = 12'h3a1 == _T_46[11:0] ? image_929 : _GEN_991; // @[Filter.scala 138:46]
  wire [3:0] _GEN_993 = 12'h3a2 == _T_46[11:0] ? image_930 : _GEN_992; // @[Filter.scala 138:46]
  wire [3:0] _GEN_994 = 12'h3a3 == _T_46[11:0] ? 4'h0 : _GEN_993; // @[Filter.scala 138:46]
  wire [3:0] _GEN_995 = 12'h3a4 == _T_46[11:0] ? 4'h0 : _GEN_994; // @[Filter.scala 138:46]
  wire [3:0] _GEN_996 = 12'h3a5 == _T_46[11:0] ? 4'h0 : _GEN_995; // @[Filter.scala 138:46]
  wire [3:0] _GEN_997 = 12'h3a6 == _T_46[11:0] ? 4'h0 : _GEN_996; // @[Filter.scala 138:46]
  wire [3:0] _GEN_998 = 12'h3a7 == _T_46[11:0] ? image_935 : _GEN_997; // @[Filter.scala 138:46]
  wire [3:0] _GEN_999 = 12'h3a8 == _T_46[11:0] ? image_936 : _GEN_998; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1000 = 12'h3a9 == _T_46[11:0] ? image_937 : _GEN_999; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1001 = 12'h3aa == _T_46[11:0] ? image_938 : _GEN_1000; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1002 = 12'h3ab == _T_46[11:0] ? image_939 : _GEN_1001; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1003 = 12'h3ac == _T_46[11:0] ? image_940 : _GEN_1002; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1004 = 12'h3ad == _T_46[11:0] ? image_941 : _GEN_1003; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1005 = 12'h3ae == _T_46[11:0] ? image_942 : _GEN_1004; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1006 = 12'h3af == _T_46[11:0] ? image_943 : _GEN_1005; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1007 = 12'h3b0 == _T_46[11:0] ? image_944 : _GEN_1006; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1008 = 12'h3b1 == _T_46[11:0] ? image_945 : _GEN_1007; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1009 = 12'h3b2 == _T_46[11:0] ? image_946 : _GEN_1008; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1010 = 12'h3b3 == _T_46[11:0] ? image_947 : _GEN_1009; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1011 = 12'h3b4 == _T_46[11:0] ? image_948 : _GEN_1010; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1012 = 12'h3b5 == _T_46[11:0] ? image_949 : _GEN_1011; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1013 = 12'h3b6 == _T_46[11:0] ? image_950 : _GEN_1012; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1014 = 12'h3b7 == _T_46[11:0] ? image_951 : _GEN_1013; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1015 = 12'h3b8 == _T_46[11:0] ? image_952 : _GEN_1014; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1016 = 12'h3b9 == _T_46[11:0] ? image_953 : _GEN_1015; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1017 = 12'h3ba == _T_46[11:0] ? image_954 : _GEN_1016; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1018 = 12'h3bb == _T_46[11:0] ? image_955 : _GEN_1017; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1019 = 12'h3bc == _T_46[11:0] ? image_956 : _GEN_1018; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1020 = 12'h3bd == _T_46[11:0] ? image_957 : _GEN_1019; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1021 = 12'h3be == _T_46[11:0] ? image_958 : _GEN_1020; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1022 = 12'h3bf == _T_46[11:0] ? image_959 : _GEN_1021; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1023 = 12'h3c0 == _T_46[11:0] ? 4'h0 : _GEN_1022; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1024 = 12'h3c1 == _T_46[11:0] ? image_961 : _GEN_1023; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1025 = 12'h3c2 == _T_46[11:0] ? image_962 : _GEN_1024; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1026 = 12'h3c3 == _T_46[11:0] ? image_963 : _GEN_1025; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1027 = 12'h3c4 == _T_46[11:0] ? image_964 : _GEN_1026; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1028 = 12'h3c5 == _T_46[11:0] ? image_965 : _GEN_1027; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1029 = 12'h3c6 == _T_46[11:0] ? image_966 : _GEN_1028; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1030 = 12'h3c7 == _T_46[11:0] ? image_967 : _GEN_1029; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1031 = 12'h3c8 == _T_46[11:0] ? image_968 : _GEN_1030; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1032 = 12'h3c9 == _T_46[11:0] ? image_969 : _GEN_1031; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1033 = 12'h3ca == _T_46[11:0] ? image_970 : _GEN_1032; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1034 = 12'h3cb == _T_46[11:0] ? image_971 : _GEN_1033; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1035 = 12'h3cc == _T_46[11:0] ? image_972 : _GEN_1034; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1036 = 12'h3cd == _T_46[11:0] ? image_973 : _GEN_1035; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1037 = 12'h3ce == _T_46[11:0] ? image_974 : _GEN_1036; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1038 = 12'h3cf == _T_46[11:0] ? image_975 : _GEN_1037; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1039 = 12'h3d0 == _T_46[11:0] ? image_976 : _GEN_1038; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1040 = 12'h3d1 == _T_46[11:0] ? image_977 : _GEN_1039; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1041 = 12'h3d2 == _T_46[11:0] ? image_978 : _GEN_1040; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1042 = 12'h3d3 == _T_46[11:0] ? image_979 : _GEN_1041; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1043 = 12'h3d4 == _T_46[11:0] ? image_980 : _GEN_1042; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1044 = 12'h3d5 == _T_46[11:0] ? image_981 : _GEN_1043; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1045 = 12'h3d6 == _T_46[11:0] ? image_982 : _GEN_1044; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1046 = 12'h3d7 == _T_46[11:0] ? image_983 : _GEN_1045; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1047 = 12'h3d8 == _T_46[11:0] ? image_984 : _GEN_1046; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1048 = 12'h3d9 == _T_46[11:0] ? image_985 : _GEN_1047; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1049 = 12'h3da == _T_46[11:0] ? image_986 : _GEN_1048; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1050 = 12'h3db == _T_46[11:0] ? image_987 : _GEN_1049; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1051 = 12'h3dc == _T_46[11:0] ? image_988 : _GEN_1050; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1052 = 12'h3dd == _T_46[11:0] ? image_989 : _GEN_1051; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1053 = 12'h3de == _T_46[11:0] ? image_990 : _GEN_1052; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1054 = 12'h3df == _T_46[11:0] ? image_991 : _GEN_1053; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1055 = 12'h3e0 == _T_46[11:0] ? image_992 : _GEN_1054; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1056 = 12'h3e1 == _T_46[11:0] ? 4'h0 : _GEN_1055; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1057 = 12'h3e2 == _T_46[11:0] ? 4'h0 : _GEN_1056; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1058 = 12'h3e3 == _T_46[11:0] ? 4'h0 : _GEN_1057; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1059 = 12'h3e4 == _T_46[11:0] ? 4'h0 : _GEN_1058; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1060 = 12'h3e5 == _T_46[11:0] ? image_997 : _GEN_1059; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1061 = 12'h3e6 == _T_46[11:0] ? image_998 : _GEN_1060; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1062 = 12'h3e7 == _T_46[11:0] ? image_999 : _GEN_1061; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1063 = 12'h3e8 == _T_46[11:0] ? image_1000 : _GEN_1062; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1064 = 12'h3e9 == _T_46[11:0] ? image_1001 : _GEN_1063; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1065 = 12'h3ea == _T_46[11:0] ? image_1002 : _GEN_1064; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1066 = 12'h3eb == _T_46[11:0] ? image_1003 : _GEN_1065; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1067 = 12'h3ec == _T_46[11:0] ? image_1004 : _GEN_1066; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1068 = 12'h3ed == _T_46[11:0] ? image_1005 : _GEN_1067; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1069 = 12'h3ee == _T_46[11:0] ? image_1006 : _GEN_1068; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1070 = 12'h3ef == _T_46[11:0] ? image_1007 : _GEN_1069; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1071 = 12'h3f0 == _T_46[11:0] ? image_1008 : _GEN_1070; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1072 = 12'h3f1 == _T_46[11:0] ? image_1009 : _GEN_1071; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1073 = 12'h3f2 == _T_46[11:0] ? image_1010 : _GEN_1072; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1074 = 12'h3f3 == _T_46[11:0] ? image_1011 : _GEN_1073; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1075 = 12'h3f4 == _T_46[11:0] ? image_1012 : _GEN_1074; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1076 = 12'h3f5 == _T_46[11:0] ? image_1013 : _GEN_1075; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1077 = 12'h3f6 == _T_46[11:0] ? image_1014 : _GEN_1076; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1078 = 12'h3f7 == _T_46[11:0] ? image_1015 : _GEN_1077; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1079 = 12'h3f8 == _T_46[11:0] ? image_1016 : _GEN_1078; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1080 = 12'h3f9 == _T_46[11:0] ? image_1017 : _GEN_1079; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1081 = 12'h3fa == _T_46[11:0] ? image_1018 : _GEN_1080; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1082 = 12'h3fb == _T_46[11:0] ? image_1019 : _GEN_1081; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1083 = 12'h3fc == _T_46[11:0] ? image_1020 : _GEN_1082; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1084 = 12'h3fd == _T_46[11:0] ? 4'h0 : _GEN_1083; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1085 = 12'h3fe == _T_46[11:0] ? 4'h0 : _GEN_1084; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1086 = 12'h3ff == _T_46[11:0] ? 4'h0 : _GEN_1085; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1087 = 12'h400 == _T_46[11:0] ? image_1024 : _GEN_1086; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1088 = 12'h401 == _T_46[11:0] ? image_1025 : _GEN_1087; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1089 = 12'h402 == _T_46[11:0] ? image_1026 : _GEN_1088; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1090 = 12'h403 == _T_46[11:0] ? image_1027 : _GEN_1089; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1091 = 12'h404 == _T_46[11:0] ? image_1028 : _GEN_1090; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1092 = 12'h405 == _T_46[11:0] ? image_1029 : _GEN_1091; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1093 = 12'h406 == _T_46[11:0] ? image_1030 : _GEN_1092; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1094 = 12'h407 == _T_46[11:0] ? image_1031 : _GEN_1093; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1095 = 12'h408 == _T_46[11:0] ? image_1032 : _GEN_1094; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1096 = 12'h409 == _T_46[11:0] ? image_1033 : _GEN_1095; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1097 = 12'h40a == _T_46[11:0] ? image_1034 : _GEN_1096; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1098 = 12'h40b == _T_46[11:0] ? image_1035 : _GEN_1097; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1099 = 12'h40c == _T_46[11:0] ? image_1036 : _GEN_1098; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1100 = 12'h40d == _T_46[11:0] ? image_1037 : _GEN_1099; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1101 = 12'h40e == _T_46[11:0] ? image_1038 : _GEN_1100; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1102 = 12'h40f == _T_46[11:0] ? image_1039 : _GEN_1101; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1103 = 12'h410 == _T_46[11:0] ? image_1040 : _GEN_1102; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1104 = 12'h411 == _T_46[11:0] ? image_1041 : _GEN_1103; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1105 = 12'h412 == _T_46[11:0] ? image_1042 : _GEN_1104; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1106 = 12'h413 == _T_46[11:0] ? image_1043 : _GEN_1105; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1107 = 12'h414 == _T_46[11:0] ? image_1044 : _GEN_1106; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1108 = 12'h415 == _T_46[11:0] ? image_1045 : _GEN_1107; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1109 = 12'h416 == _T_46[11:0] ? image_1046 : _GEN_1108; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1110 = 12'h417 == _T_46[11:0] ? image_1047 : _GEN_1109; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1111 = 12'h418 == _T_46[11:0] ? image_1048 : _GEN_1110; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1112 = 12'h419 == _T_46[11:0] ? image_1049 : _GEN_1111; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1113 = 12'h41a == _T_46[11:0] ? image_1050 : _GEN_1112; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1114 = 12'h41b == _T_46[11:0] ? image_1051 : _GEN_1113; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1115 = 12'h41c == _T_46[11:0] ? image_1052 : _GEN_1114; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1116 = 12'h41d == _T_46[11:0] ? image_1053 : _GEN_1115; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1117 = 12'h41e == _T_46[11:0] ? image_1054 : _GEN_1116; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1118 = 12'h41f == _T_46[11:0] ? image_1055 : _GEN_1117; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1119 = 12'h420 == _T_46[11:0] ? image_1056 : _GEN_1118; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1120 = 12'h421 == _T_46[11:0] ? image_1057 : _GEN_1119; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1121 = 12'h422 == _T_46[11:0] ? image_1058 : _GEN_1120; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1122 = 12'h423 == _T_46[11:0] ? image_1059 : _GEN_1121; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1123 = 12'h424 == _T_46[11:0] ? image_1060 : _GEN_1122; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1124 = 12'h425 == _T_46[11:0] ? image_1061 : _GEN_1123; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1125 = 12'h426 == _T_46[11:0] ? image_1062 : _GEN_1124; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1126 = 12'h427 == _T_46[11:0] ? image_1063 : _GEN_1125; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1127 = 12'h428 == _T_46[11:0] ? image_1064 : _GEN_1126; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1128 = 12'h429 == _T_46[11:0] ? image_1065 : _GEN_1127; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1129 = 12'h42a == _T_46[11:0] ? image_1066 : _GEN_1128; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1130 = 12'h42b == _T_46[11:0] ? image_1067 : _GEN_1129; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1131 = 12'h42c == _T_46[11:0] ? image_1068 : _GEN_1130; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1132 = 12'h42d == _T_46[11:0] ? image_1069 : _GEN_1131; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1133 = 12'h42e == _T_46[11:0] ? image_1070 : _GEN_1132; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1134 = 12'h42f == _T_46[11:0] ? image_1071 : _GEN_1133; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1135 = 12'h430 == _T_46[11:0] ? image_1072 : _GEN_1134; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1136 = 12'h431 == _T_46[11:0] ? image_1073 : _GEN_1135; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1137 = 12'h432 == _T_46[11:0] ? image_1074 : _GEN_1136; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1138 = 12'h433 == _T_46[11:0] ? image_1075 : _GEN_1137; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1139 = 12'h434 == _T_46[11:0] ? image_1076 : _GEN_1138; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1140 = 12'h435 == _T_46[11:0] ? image_1077 : _GEN_1139; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1141 = 12'h436 == _T_46[11:0] ? image_1078 : _GEN_1140; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1142 = 12'h437 == _T_46[11:0] ? image_1079 : _GEN_1141; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1143 = 12'h438 == _T_46[11:0] ? image_1080 : _GEN_1142; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1144 = 12'h439 == _T_46[11:0] ? image_1081 : _GEN_1143; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1145 = 12'h43a == _T_46[11:0] ? image_1082 : _GEN_1144; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1146 = 12'h43b == _T_46[11:0] ? image_1083 : _GEN_1145; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1147 = 12'h43c == _T_46[11:0] ? image_1084 : _GEN_1146; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1148 = 12'h43d == _T_46[11:0] ? image_1085 : _GEN_1147; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1149 = 12'h43e == _T_46[11:0] ? 4'h0 : _GEN_1148; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1150 = 12'h43f == _T_46[11:0] ? 4'h0 : _GEN_1149; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1151 = 12'h440 == _T_46[11:0] ? image_1088 : _GEN_1150; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1152 = 12'h441 == _T_46[11:0] ? image_1089 : _GEN_1151; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1153 = 12'h442 == _T_46[11:0] ? image_1090 : _GEN_1152; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1154 = 12'h443 == _T_46[11:0] ? image_1091 : _GEN_1153; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1155 = 12'h444 == _T_46[11:0] ? image_1092 : _GEN_1154; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1156 = 12'h445 == _T_46[11:0] ? image_1093 : _GEN_1155; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1157 = 12'h446 == _T_46[11:0] ? image_1094 : _GEN_1156; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1158 = 12'h447 == _T_46[11:0] ? image_1095 : _GEN_1157; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1159 = 12'h448 == _T_46[11:0] ? image_1096 : _GEN_1158; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1160 = 12'h449 == _T_46[11:0] ? image_1097 : _GEN_1159; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1161 = 12'h44a == _T_46[11:0] ? image_1098 : _GEN_1160; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1162 = 12'h44b == _T_46[11:0] ? image_1099 : _GEN_1161; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1163 = 12'h44c == _T_46[11:0] ? image_1100 : _GEN_1162; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1164 = 12'h44d == _T_46[11:0] ? image_1101 : _GEN_1163; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1165 = 12'h44e == _T_46[11:0] ? image_1102 : _GEN_1164; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1166 = 12'h44f == _T_46[11:0] ? image_1103 : _GEN_1165; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1167 = 12'h450 == _T_46[11:0] ? image_1104 : _GEN_1166; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1168 = 12'h451 == _T_46[11:0] ? image_1105 : _GEN_1167; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1169 = 12'h452 == _T_46[11:0] ? image_1106 : _GEN_1168; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1170 = 12'h453 == _T_46[11:0] ? image_1107 : _GEN_1169; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1171 = 12'h454 == _T_46[11:0] ? image_1108 : _GEN_1170; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1172 = 12'h455 == _T_46[11:0] ? image_1109 : _GEN_1171; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1173 = 12'h456 == _T_46[11:0] ? image_1110 : _GEN_1172; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1174 = 12'h457 == _T_46[11:0] ? image_1111 : _GEN_1173; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1175 = 12'h458 == _T_46[11:0] ? image_1112 : _GEN_1174; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1176 = 12'h459 == _T_46[11:0] ? image_1113 : _GEN_1175; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1177 = 12'h45a == _T_46[11:0] ? image_1114 : _GEN_1176; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1178 = 12'h45b == _T_46[11:0] ? image_1115 : _GEN_1177; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1179 = 12'h45c == _T_46[11:0] ? image_1116 : _GEN_1178; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1180 = 12'h45d == _T_46[11:0] ? image_1117 : _GEN_1179; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1181 = 12'h45e == _T_46[11:0] ? image_1118 : _GEN_1180; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1182 = 12'h45f == _T_46[11:0] ? image_1119 : _GEN_1181; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1183 = 12'h460 == _T_46[11:0] ? image_1120 : _GEN_1182; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1184 = 12'h461 == _T_46[11:0] ? image_1121 : _GEN_1183; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1185 = 12'h462 == _T_46[11:0] ? image_1122 : _GEN_1184; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1186 = 12'h463 == _T_46[11:0] ? image_1123 : _GEN_1185; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1187 = 12'h464 == _T_46[11:0] ? image_1124 : _GEN_1186; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1188 = 12'h465 == _T_46[11:0] ? image_1125 : _GEN_1187; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1189 = 12'h466 == _T_46[11:0] ? image_1126 : _GEN_1188; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1190 = 12'h467 == _T_46[11:0] ? image_1127 : _GEN_1189; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1191 = 12'h468 == _T_46[11:0] ? image_1128 : _GEN_1190; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1192 = 12'h469 == _T_46[11:0] ? image_1129 : _GEN_1191; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1193 = 12'h46a == _T_46[11:0] ? image_1130 : _GEN_1192; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1194 = 12'h46b == _T_46[11:0] ? image_1131 : _GEN_1193; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1195 = 12'h46c == _T_46[11:0] ? image_1132 : _GEN_1194; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1196 = 12'h46d == _T_46[11:0] ? image_1133 : _GEN_1195; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1197 = 12'h46e == _T_46[11:0] ? image_1134 : _GEN_1196; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1198 = 12'h46f == _T_46[11:0] ? image_1135 : _GEN_1197; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1199 = 12'h470 == _T_46[11:0] ? image_1136 : _GEN_1198; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1200 = 12'h471 == _T_46[11:0] ? image_1137 : _GEN_1199; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1201 = 12'h472 == _T_46[11:0] ? image_1138 : _GEN_1200; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1202 = 12'h473 == _T_46[11:0] ? image_1139 : _GEN_1201; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1203 = 12'h474 == _T_46[11:0] ? image_1140 : _GEN_1202; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1204 = 12'h475 == _T_46[11:0] ? image_1141 : _GEN_1203; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1205 = 12'h476 == _T_46[11:0] ? image_1142 : _GEN_1204; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1206 = 12'h477 == _T_46[11:0] ? image_1143 : _GEN_1205; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1207 = 12'h478 == _T_46[11:0] ? image_1144 : _GEN_1206; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1208 = 12'h479 == _T_46[11:0] ? image_1145 : _GEN_1207; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1209 = 12'h47a == _T_46[11:0] ? image_1146 : _GEN_1208; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1210 = 12'h47b == _T_46[11:0] ? image_1147 : _GEN_1209; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1211 = 12'h47c == _T_46[11:0] ? image_1148 : _GEN_1210; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1212 = 12'h47d == _T_46[11:0] ? 4'h0 : _GEN_1211; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1213 = 12'h47e == _T_46[11:0] ? 4'h0 : _GEN_1212; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1214 = 12'h47f == _T_46[11:0] ? 4'h0 : _GEN_1213; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1215 = 12'h480 == _T_46[11:0] ? image_1152 : _GEN_1214; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1216 = 12'h481 == _T_46[11:0] ? image_1153 : _GEN_1215; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1217 = 12'h482 == _T_46[11:0] ? image_1154 : _GEN_1216; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1218 = 12'h483 == _T_46[11:0] ? image_1155 : _GEN_1217; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1219 = 12'h484 == _T_46[11:0] ? image_1156 : _GEN_1218; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1220 = 12'h485 == _T_46[11:0] ? image_1157 : _GEN_1219; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1221 = 12'h486 == _T_46[11:0] ? image_1158 : _GEN_1220; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1222 = 12'h487 == _T_46[11:0] ? image_1159 : _GEN_1221; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1223 = 12'h488 == _T_46[11:0] ? image_1160 : _GEN_1222; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1224 = 12'h489 == _T_46[11:0] ? image_1161 : _GEN_1223; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1225 = 12'h48a == _T_46[11:0] ? image_1162 : _GEN_1224; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1226 = 12'h48b == _T_46[11:0] ? image_1163 : _GEN_1225; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1227 = 12'h48c == _T_46[11:0] ? image_1164 : _GEN_1226; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1228 = 12'h48d == _T_46[11:0] ? image_1165 : _GEN_1227; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1229 = 12'h48e == _T_46[11:0] ? image_1166 : _GEN_1228; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1230 = 12'h48f == _T_46[11:0] ? image_1167 : _GEN_1229; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1231 = 12'h490 == _T_46[11:0] ? image_1168 : _GEN_1230; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1232 = 12'h491 == _T_46[11:0] ? image_1169 : _GEN_1231; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1233 = 12'h492 == _T_46[11:0] ? image_1170 : _GEN_1232; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1234 = 12'h493 == _T_46[11:0] ? image_1171 : _GEN_1233; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1235 = 12'h494 == _T_46[11:0] ? image_1172 : _GEN_1234; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1236 = 12'h495 == _T_46[11:0] ? image_1173 : _GEN_1235; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1237 = 12'h496 == _T_46[11:0] ? image_1174 : _GEN_1236; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1238 = 12'h497 == _T_46[11:0] ? image_1175 : _GEN_1237; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1239 = 12'h498 == _T_46[11:0] ? image_1176 : _GEN_1238; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1240 = 12'h499 == _T_46[11:0] ? image_1177 : _GEN_1239; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1241 = 12'h49a == _T_46[11:0] ? image_1178 : _GEN_1240; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1242 = 12'h49b == _T_46[11:0] ? image_1179 : _GEN_1241; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1243 = 12'h49c == _T_46[11:0] ? image_1180 : _GEN_1242; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1244 = 12'h49d == _T_46[11:0] ? image_1181 : _GEN_1243; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1245 = 12'h49e == _T_46[11:0] ? image_1182 : _GEN_1244; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1246 = 12'h49f == _T_46[11:0] ? image_1183 : _GEN_1245; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1247 = 12'h4a0 == _T_46[11:0] ? image_1184 : _GEN_1246; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1248 = 12'h4a1 == _T_46[11:0] ? image_1185 : _GEN_1247; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1249 = 12'h4a2 == _T_46[11:0] ? image_1186 : _GEN_1248; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1250 = 12'h4a3 == _T_46[11:0] ? image_1187 : _GEN_1249; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1251 = 12'h4a4 == _T_46[11:0] ? image_1188 : _GEN_1250; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1252 = 12'h4a5 == _T_46[11:0] ? image_1189 : _GEN_1251; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1253 = 12'h4a6 == _T_46[11:0] ? image_1190 : _GEN_1252; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1254 = 12'h4a7 == _T_46[11:0] ? image_1191 : _GEN_1253; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1255 = 12'h4a8 == _T_46[11:0] ? image_1192 : _GEN_1254; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1256 = 12'h4a9 == _T_46[11:0] ? image_1193 : _GEN_1255; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1257 = 12'h4aa == _T_46[11:0] ? image_1194 : _GEN_1256; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1258 = 12'h4ab == _T_46[11:0] ? image_1195 : _GEN_1257; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1259 = 12'h4ac == _T_46[11:0] ? image_1196 : _GEN_1258; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1260 = 12'h4ad == _T_46[11:0] ? image_1197 : _GEN_1259; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1261 = 12'h4ae == _T_46[11:0] ? image_1198 : _GEN_1260; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1262 = 12'h4af == _T_46[11:0] ? image_1199 : _GEN_1261; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1263 = 12'h4b0 == _T_46[11:0] ? image_1200 : _GEN_1262; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1264 = 12'h4b1 == _T_46[11:0] ? image_1201 : _GEN_1263; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1265 = 12'h4b2 == _T_46[11:0] ? image_1202 : _GEN_1264; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1266 = 12'h4b3 == _T_46[11:0] ? image_1203 : _GEN_1265; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1267 = 12'h4b4 == _T_46[11:0] ? image_1204 : _GEN_1266; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1268 = 12'h4b5 == _T_46[11:0] ? image_1205 : _GEN_1267; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1269 = 12'h4b6 == _T_46[11:0] ? image_1206 : _GEN_1268; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1270 = 12'h4b7 == _T_46[11:0] ? image_1207 : _GEN_1269; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1271 = 12'h4b8 == _T_46[11:0] ? image_1208 : _GEN_1270; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1272 = 12'h4b9 == _T_46[11:0] ? 4'h0 : _GEN_1271; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1273 = 12'h4ba == _T_46[11:0] ? 4'h0 : _GEN_1272; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1274 = 12'h4bb == _T_46[11:0] ? 4'h0 : _GEN_1273; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1275 = 12'h4bc == _T_46[11:0] ? 4'h0 : _GEN_1274; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1276 = 12'h4bd == _T_46[11:0] ? 4'h0 : _GEN_1275; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1277 = 12'h4be == _T_46[11:0] ? 4'h0 : _GEN_1276; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1278 = 12'h4bf == _T_46[11:0] ? 4'h0 : _GEN_1277; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1279 = 12'h4c0 == _T_46[11:0] ? image_1216 : _GEN_1278; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1280 = 12'h4c1 == _T_46[11:0] ? image_1217 : _GEN_1279; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1281 = 12'h4c2 == _T_46[11:0] ? image_1218 : _GEN_1280; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1282 = 12'h4c3 == _T_46[11:0] ? image_1219 : _GEN_1281; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1283 = 12'h4c4 == _T_46[11:0] ? image_1220 : _GEN_1282; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1284 = 12'h4c5 == _T_46[11:0] ? image_1221 : _GEN_1283; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1285 = 12'h4c6 == _T_46[11:0] ? image_1222 : _GEN_1284; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1286 = 12'h4c7 == _T_46[11:0] ? image_1223 : _GEN_1285; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1287 = 12'h4c8 == _T_46[11:0] ? image_1224 : _GEN_1286; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1288 = 12'h4c9 == _T_46[11:0] ? image_1225 : _GEN_1287; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1289 = 12'h4ca == _T_46[11:0] ? image_1226 : _GEN_1288; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1290 = 12'h4cb == _T_46[11:0] ? image_1227 : _GEN_1289; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1291 = 12'h4cc == _T_46[11:0] ? image_1228 : _GEN_1290; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1292 = 12'h4cd == _T_46[11:0] ? image_1229 : _GEN_1291; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1293 = 12'h4ce == _T_46[11:0] ? image_1230 : _GEN_1292; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1294 = 12'h4cf == _T_46[11:0] ? image_1231 : _GEN_1293; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1295 = 12'h4d0 == _T_46[11:0] ? image_1232 : _GEN_1294; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1296 = 12'h4d1 == _T_46[11:0] ? image_1233 : _GEN_1295; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1297 = 12'h4d2 == _T_46[11:0] ? image_1234 : _GEN_1296; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1298 = 12'h4d3 == _T_46[11:0] ? image_1235 : _GEN_1297; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1299 = 12'h4d4 == _T_46[11:0] ? image_1236 : _GEN_1298; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1300 = 12'h4d5 == _T_46[11:0] ? image_1237 : _GEN_1299; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1301 = 12'h4d6 == _T_46[11:0] ? image_1238 : _GEN_1300; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1302 = 12'h4d7 == _T_46[11:0] ? image_1239 : _GEN_1301; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1303 = 12'h4d8 == _T_46[11:0] ? image_1240 : _GEN_1302; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1304 = 12'h4d9 == _T_46[11:0] ? image_1241 : _GEN_1303; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1305 = 12'h4da == _T_46[11:0] ? image_1242 : _GEN_1304; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1306 = 12'h4db == _T_46[11:0] ? image_1243 : _GEN_1305; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1307 = 12'h4dc == _T_46[11:0] ? image_1244 : _GEN_1306; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1308 = 12'h4dd == _T_46[11:0] ? image_1245 : _GEN_1307; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1309 = 12'h4de == _T_46[11:0] ? image_1246 : _GEN_1308; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1310 = 12'h4df == _T_46[11:0] ? image_1247 : _GEN_1309; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1311 = 12'h4e0 == _T_46[11:0] ? image_1248 : _GEN_1310; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1312 = 12'h4e1 == _T_46[11:0] ? image_1249 : _GEN_1311; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1313 = 12'h4e2 == _T_46[11:0] ? image_1250 : _GEN_1312; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1314 = 12'h4e3 == _T_46[11:0] ? image_1251 : _GEN_1313; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1315 = 12'h4e4 == _T_46[11:0] ? image_1252 : _GEN_1314; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1316 = 12'h4e5 == _T_46[11:0] ? image_1253 : _GEN_1315; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1317 = 12'h4e6 == _T_46[11:0] ? image_1254 : _GEN_1316; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1318 = 12'h4e7 == _T_46[11:0] ? image_1255 : _GEN_1317; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1319 = 12'h4e8 == _T_46[11:0] ? image_1256 : _GEN_1318; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1320 = 12'h4e9 == _T_46[11:0] ? image_1257 : _GEN_1319; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1321 = 12'h4ea == _T_46[11:0] ? image_1258 : _GEN_1320; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1322 = 12'h4eb == _T_46[11:0] ? image_1259 : _GEN_1321; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1323 = 12'h4ec == _T_46[11:0] ? image_1260 : _GEN_1322; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1324 = 12'h4ed == _T_46[11:0] ? image_1261 : _GEN_1323; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1325 = 12'h4ee == _T_46[11:0] ? image_1262 : _GEN_1324; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1326 = 12'h4ef == _T_46[11:0] ? image_1263 : _GEN_1325; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1327 = 12'h4f0 == _T_46[11:0] ? image_1264 : _GEN_1326; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1328 = 12'h4f1 == _T_46[11:0] ? image_1265 : _GEN_1327; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1329 = 12'h4f2 == _T_46[11:0] ? image_1266 : _GEN_1328; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1330 = 12'h4f3 == _T_46[11:0] ? image_1267 : _GEN_1329; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1331 = 12'h4f4 == _T_46[11:0] ? image_1268 : _GEN_1330; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1332 = 12'h4f5 == _T_46[11:0] ? image_1269 : _GEN_1331; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1333 = 12'h4f6 == _T_46[11:0] ? image_1270 : _GEN_1332; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1334 = 12'h4f7 == _T_46[11:0] ? image_1271 : _GEN_1333; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1335 = 12'h4f8 == _T_46[11:0] ? image_1272 : _GEN_1334; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1336 = 12'h4f9 == _T_46[11:0] ? image_1273 : _GEN_1335; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1337 = 12'h4fa == _T_46[11:0] ? image_1274 : _GEN_1336; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1338 = 12'h4fb == _T_46[11:0] ? image_1275 : _GEN_1337; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1339 = 12'h4fc == _T_46[11:0] ? 4'h0 : _GEN_1338; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1340 = 12'h4fd == _T_46[11:0] ? 4'h0 : _GEN_1339; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1341 = 12'h4fe == _T_46[11:0] ? 4'h0 : _GEN_1340; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1342 = 12'h4ff == _T_46[11:0] ? 4'h0 : _GEN_1341; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1343 = 12'h500 == _T_46[11:0] ? image_1280 : _GEN_1342; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1344 = 12'h501 == _T_46[11:0] ? image_1281 : _GEN_1343; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1345 = 12'h502 == _T_46[11:0] ? image_1282 : _GEN_1344; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1346 = 12'h503 == _T_46[11:0] ? image_1283 : _GEN_1345; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1347 = 12'h504 == _T_46[11:0] ? image_1284 : _GEN_1346; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1348 = 12'h505 == _T_46[11:0] ? image_1285 : _GEN_1347; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1349 = 12'h506 == _T_46[11:0] ? image_1286 : _GEN_1348; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1350 = 12'h507 == _T_46[11:0] ? image_1287 : _GEN_1349; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1351 = 12'h508 == _T_46[11:0] ? image_1288 : _GEN_1350; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1352 = 12'h509 == _T_46[11:0] ? image_1289 : _GEN_1351; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1353 = 12'h50a == _T_46[11:0] ? image_1290 : _GEN_1352; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1354 = 12'h50b == _T_46[11:0] ? image_1291 : _GEN_1353; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1355 = 12'h50c == _T_46[11:0] ? image_1292 : _GEN_1354; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1356 = 12'h50d == _T_46[11:0] ? image_1293 : _GEN_1355; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1357 = 12'h50e == _T_46[11:0] ? image_1294 : _GEN_1356; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1358 = 12'h50f == _T_46[11:0] ? image_1295 : _GEN_1357; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1359 = 12'h510 == _T_46[11:0] ? image_1296 : _GEN_1358; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1360 = 12'h511 == _T_46[11:0] ? image_1297 : _GEN_1359; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1361 = 12'h512 == _T_46[11:0] ? image_1298 : _GEN_1360; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1362 = 12'h513 == _T_46[11:0] ? image_1299 : _GEN_1361; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1363 = 12'h514 == _T_46[11:0] ? image_1300 : _GEN_1362; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1364 = 12'h515 == _T_46[11:0] ? image_1301 : _GEN_1363; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1365 = 12'h516 == _T_46[11:0] ? image_1302 : _GEN_1364; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1366 = 12'h517 == _T_46[11:0] ? image_1303 : _GEN_1365; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1367 = 12'h518 == _T_46[11:0] ? image_1304 : _GEN_1366; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1368 = 12'h519 == _T_46[11:0] ? image_1305 : _GEN_1367; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1369 = 12'h51a == _T_46[11:0] ? image_1306 : _GEN_1368; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1370 = 12'h51b == _T_46[11:0] ? image_1307 : _GEN_1369; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1371 = 12'h51c == _T_46[11:0] ? image_1308 : _GEN_1370; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1372 = 12'h51d == _T_46[11:0] ? image_1309 : _GEN_1371; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1373 = 12'h51e == _T_46[11:0] ? image_1310 : _GEN_1372; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1374 = 12'h51f == _T_46[11:0] ? image_1311 : _GEN_1373; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1375 = 12'h520 == _T_46[11:0] ? image_1312 : _GEN_1374; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1376 = 12'h521 == _T_46[11:0] ? image_1313 : _GEN_1375; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1377 = 12'h522 == _T_46[11:0] ? image_1314 : _GEN_1376; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1378 = 12'h523 == _T_46[11:0] ? image_1315 : _GEN_1377; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1379 = 12'h524 == _T_46[11:0] ? image_1316 : _GEN_1378; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1380 = 12'h525 == _T_46[11:0] ? image_1317 : _GEN_1379; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1381 = 12'h526 == _T_46[11:0] ? image_1318 : _GEN_1380; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1382 = 12'h527 == _T_46[11:0] ? image_1319 : _GEN_1381; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1383 = 12'h528 == _T_46[11:0] ? image_1320 : _GEN_1382; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1384 = 12'h529 == _T_46[11:0] ? image_1321 : _GEN_1383; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1385 = 12'h52a == _T_46[11:0] ? image_1322 : _GEN_1384; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1386 = 12'h52b == _T_46[11:0] ? image_1323 : _GEN_1385; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1387 = 12'h52c == _T_46[11:0] ? image_1324 : _GEN_1386; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1388 = 12'h52d == _T_46[11:0] ? image_1325 : _GEN_1387; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1389 = 12'h52e == _T_46[11:0] ? image_1326 : _GEN_1388; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1390 = 12'h52f == _T_46[11:0] ? image_1327 : _GEN_1389; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1391 = 12'h530 == _T_46[11:0] ? image_1328 : _GEN_1390; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1392 = 12'h531 == _T_46[11:0] ? image_1329 : _GEN_1391; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1393 = 12'h532 == _T_46[11:0] ? image_1330 : _GEN_1392; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1394 = 12'h533 == _T_46[11:0] ? image_1331 : _GEN_1393; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1395 = 12'h534 == _T_46[11:0] ? image_1332 : _GEN_1394; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1396 = 12'h535 == _T_46[11:0] ? image_1333 : _GEN_1395; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1397 = 12'h536 == _T_46[11:0] ? image_1334 : _GEN_1396; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1398 = 12'h537 == _T_46[11:0] ? image_1335 : _GEN_1397; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1399 = 12'h538 == _T_46[11:0] ? image_1336 : _GEN_1398; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1400 = 12'h539 == _T_46[11:0] ? image_1337 : _GEN_1399; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1401 = 12'h53a == _T_46[11:0] ? image_1338 : _GEN_1400; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1402 = 12'h53b == _T_46[11:0] ? image_1339 : _GEN_1401; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1403 = 12'h53c == _T_46[11:0] ? image_1340 : _GEN_1402; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1404 = 12'h53d == _T_46[11:0] ? image_1341 : _GEN_1403; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1405 = 12'h53e == _T_46[11:0] ? 4'h0 : _GEN_1404; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1406 = 12'h53f == _T_46[11:0] ? 4'h0 : _GEN_1405; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1407 = 12'h540 == _T_46[11:0] ? image_1344 : _GEN_1406; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1408 = 12'h541 == _T_46[11:0] ? image_1345 : _GEN_1407; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1409 = 12'h542 == _T_46[11:0] ? image_1346 : _GEN_1408; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1410 = 12'h543 == _T_46[11:0] ? image_1347 : _GEN_1409; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1411 = 12'h544 == _T_46[11:0] ? image_1348 : _GEN_1410; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1412 = 12'h545 == _T_46[11:0] ? image_1349 : _GEN_1411; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1413 = 12'h546 == _T_46[11:0] ? image_1350 : _GEN_1412; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1414 = 12'h547 == _T_46[11:0] ? image_1351 : _GEN_1413; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1415 = 12'h548 == _T_46[11:0] ? image_1352 : _GEN_1414; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1416 = 12'h549 == _T_46[11:0] ? image_1353 : _GEN_1415; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1417 = 12'h54a == _T_46[11:0] ? image_1354 : _GEN_1416; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1418 = 12'h54b == _T_46[11:0] ? image_1355 : _GEN_1417; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1419 = 12'h54c == _T_46[11:0] ? image_1356 : _GEN_1418; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1420 = 12'h54d == _T_46[11:0] ? image_1357 : _GEN_1419; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1421 = 12'h54e == _T_46[11:0] ? image_1358 : _GEN_1420; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1422 = 12'h54f == _T_46[11:0] ? image_1359 : _GEN_1421; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1423 = 12'h550 == _T_46[11:0] ? image_1360 : _GEN_1422; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1424 = 12'h551 == _T_46[11:0] ? image_1361 : _GEN_1423; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1425 = 12'h552 == _T_46[11:0] ? image_1362 : _GEN_1424; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1426 = 12'h553 == _T_46[11:0] ? image_1363 : _GEN_1425; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1427 = 12'h554 == _T_46[11:0] ? image_1364 : _GEN_1426; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1428 = 12'h555 == _T_46[11:0] ? image_1365 : _GEN_1427; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1429 = 12'h556 == _T_46[11:0] ? image_1366 : _GEN_1428; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1430 = 12'h557 == _T_46[11:0] ? image_1367 : _GEN_1429; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1431 = 12'h558 == _T_46[11:0] ? image_1368 : _GEN_1430; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1432 = 12'h559 == _T_46[11:0] ? image_1369 : _GEN_1431; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1433 = 12'h55a == _T_46[11:0] ? image_1370 : _GEN_1432; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1434 = 12'h55b == _T_46[11:0] ? image_1371 : _GEN_1433; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1435 = 12'h55c == _T_46[11:0] ? image_1372 : _GEN_1434; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1436 = 12'h55d == _T_46[11:0] ? image_1373 : _GEN_1435; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1437 = 12'h55e == _T_46[11:0] ? image_1374 : _GEN_1436; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1438 = 12'h55f == _T_46[11:0] ? image_1375 : _GEN_1437; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1439 = 12'h560 == _T_46[11:0] ? image_1376 : _GEN_1438; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1440 = 12'h561 == _T_46[11:0] ? image_1377 : _GEN_1439; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1441 = 12'h562 == _T_46[11:0] ? image_1378 : _GEN_1440; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1442 = 12'h563 == _T_46[11:0] ? image_1379 : _GEN_1441; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1443 = 12'h564 == _T_46[11:0] ? image_1380 : _GEN_1442; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1444 = 12'h565 == _T_46[11:0] ? image_1381 : _GEN_1443; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1445 = 12'h566 == _T_46[11:0] ? image_1382 : _GEN_1444; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1446 = 12'h567 == _T_46[11:0] ? image_1383 : _GEN_1445; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1447 = 12'h568 == _T_46[11:0] ? image_1384 : _GEN_1446; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1448 = 12'h569 == _T_46[11:0] ? image_1385 : _GEN_1447; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1449 = 12'h56a == _T_46[11:0] ? image_1386 : _GEN_1448; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1450 = 12'h56b == _T_46[11:0] ? image_1387 : _GEN_1449; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1451 = 12'h56c == _T_46[11:0] ? image_1388 : _GEN_1450; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1452 = 12'h56d == _T_46[11:0] ? image_1389 : _GEN_1451; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1453 = 12'h56e == _T_46[11:0] ? image_1390 : _GEN_1452; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1454 = 12'h56f == _T_46[11:0] ? image_1391 : _GEN_1453; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1455 = 12'h570 == _T_46[11:0] ? image_1392 : _GEN_1454; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1456 = 12'h571 == _T_46[11:0] ? image_1393 : _GEN_1455; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1457 = 12'h572 == _T_46[11:0] ? image_1394 : _GEN_1456; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1458 = 12'h573 == _T_46[11:0] ? image_1395 : _GEN_1457; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1459 = 12'h574 == _T_46[11:0] ? image_1396 : _GEN_1458; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1460 = 12'h575 == _T_46[11:0] ? image_1397 : _GEN_1459; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1461 = 12'h576 == _T_46[11:0] ? image_1398 : _GEN_1460; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1462 = 12'h577 == _T_46[11:0] ? image_1399 : _GEN_1461; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1463 = 12'h578 == _T_46[11:0] ? image_1400 : _GEN_1462; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1464 = 12'h579 == _T_46[11:0] ? image_1401 : _GEN_1463; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1465 = 12'h57a == _T_46[11:0] ? image_1402 : _GEN_1464; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1466 = 12'h57b == _T_46[11:0] ? image_1403 : _GEN_1465; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1467 = 12'h57c == _T_46[11:0] ? image_1404 : _GEN_1466; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1468 = 12'h57d == _T_46[11:0] ? image_1405 : _GEN_1467; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1469 = 12'h57e == _T_46[11:0] ? 4'h0 : _GEN_1468; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1470 = 12'h57f == _T_46[11:0] ? 4'h0 : _GEN_1469; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1471 = 12'h580 == _T_46[11:0] ? image_1408 : _GEN_1470; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1472 = 12'h581 == _T_46[11:0] ? image_1409 : _GEN_1471; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1473 = 12'h582 == _T_46[11:0] ? image_1410 : _GEN_1472; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1474 = 12'h583 == _T_46[11:0] ? image_1411 : _GEN_1473; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1475 = 12'h584 == _T_46[11:0] ? image_1412 : _GEN_1474; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1476 = 12'h585 == _T_46[11:0] ? image_1413 : _GEN_1475; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1477 = 12'h586 == _T_46[11:0] ? image_1414 : _GEN_1476; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1478 = 12'h587 == _T_46[11:0] ? image_1415 : _GEN_1477; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1479 = 12'h588 == _T_46[11:0] ? image_1416 : _GEN_1478; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1480 = 12'h589 == _T_46[11:0] ? image_1417 : _GEN_1479; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1481 = 12'h58a == _T_46[11:0] ? image_1418 : _GEN_1480; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1482 = 12'h58b == _T_46[11:0] ? image_1419 : _GEN_1481; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1483 = 12'h58c == _T_46[11:0] ? image_1420 : _GEN_1482; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1484 = 12'h58d == _T_46[11:0] ? image_1421 : _GEN_1483; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1485 = 12'h58e == _T_46[11:0] ? image_1422 : _GEN_1484; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1486 = 12'h58f == _T_46[11:0] ? image_1423 : _GEN_1485; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1487 = 12'h590 == _T_46[11:0] ? image_1424 : _GEN_1486; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1488 = 12'h591 == _T_46[11:0] ? image_1425 : _GEN_1487; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1489 = 12'h592 == _T_46[11:0] ? image_1426 : _GEN_1488; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1490 = 12'h593 == _T_46[11:0] ? image_1427 : _GEN_1489; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1491 = 12'h594 == _T_46[11:0] ? image_1428 : _GEN_1490; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1492 = 12'h595 == _T_46[11:0] ? image_1429 : _GEN_1491; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1493 = 12'h596 == _T_46[11:0] ? image_1430 : _GEN_1492; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1494 = 12'h597 == _T_46[11:0] ? image_1431 : _GEN_1493; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1495 = 12'h598 == _T_46[11:0] ? image_1432 : _GEN_1494; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1496 = 12'h599 == _T_46[11:0] ? image_1433 : _GEN_1495; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1497 = 12'h59a == _T_46[11:0] ? image_1434 : _GEN_1496; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1498 = 12'h59b == _T_46[11:0] ? image_1435 : _GEN_1497; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1499 = 12'h59c == _T_46[11:0] ? image_1436 : _GEN_1498; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1500 = 12'h59d == _T_46[11:0] ? image_1437 : _GEN_1499; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1501 = 12'h59e == _T_46[11:0] ? image_1438 : _GEN_1500; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1502 = 12'h59f == _T_46[11:0] ? image_1439 : _GEN_1501; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1503 = 12'h5a0 == _T_46[11:0] ? image_1440 : _GEN_1502; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1504 = 12'h5a1 == _T_46[11:0] ? image_1441 : _GEN_1503; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1505 = 12'h5a2 == _T_46[11:0] ? image_1442 : _GEN_1504; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1506 = 12'h5a3 == _T_46[11:0] ? image_1443 : _GEN_1505; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1507 = 12'h5a4 == _T_46[11:0] ? image_1444 : _GEN_1506; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1508 = 12'h5a5 == _T_46[11:0] ? image_1445 : _GEN_1507; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1509 = 12'h5a6 == _T_46[11:0] ? image_1446 : _GEN_1508; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1510 = 12'h5a7 == _T_46[11:0] ? image_1447 : _GEN_1509; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1511 = 12'h5a8 == _T_46[11:0] ? image_1448 : _GEN_1510; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1512 = 12'h5a9 == _T_46[11:0] ? image_1449 : _GEN_1511; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1513 = 12'h5aa == _T_46[11:0] ? image_1450 : _GEN_1512; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1514 = 12'h5ab == _T_46[11:0] ? image_1451 : _GEN_1513; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1515 = 12'h5ac == _T_46[11:0] ? image_1452 : _GEN_1514; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1516 = 12'h5ad == _T_46[11:0] ? image_1453 : _GEN_1515; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1517 = 12'h5ae == _T_46[11:0] ? image_1454 : _GEN_1516; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1518 = 12'h5af == _T_46[11:0] ? image_1455 : _GEN_1517; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1519 = 12'h5b0 == _T_46[11:0] ? image_1456 : _GEN_1518; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1520 = 12'h5b1 == _T_46[11:0] ? image_1457 : _GEN_1519; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1521 = 12'h5b2 == _T_46[11:0] ? image_1458 : _GEN_1520; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1522 = 12'h5b3 == _T_46[11:0] ? image_1459 : _GEN_1521; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1523 = 12'h5b4 == _T_46[11:0] ? image_1460 : _GEN_1522; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1524 = 12'h5b5 == _T_46[11:0] ? image_1461 : _GEN_1523; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1525 = 12'h5b6 == _T_46[11:0] ? image_1462 : _GEN_1524; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1526 = 12'h5b7 == _T_46[11:0] ? image_1463 : _GEN_1525; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1527 = 12'h5b8 == _T_46[11:0] ? image_1464 : _GEN_1526; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1528 = 12'h5b9 == _T_46[11:0] ? image_1465 : _GEN_1527; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1529 = 12'h5ba == _T_46[11:0] ? image_1466 : _GEN_1528; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1530 = 12'h5bb == _T_46[11:0] ? image_1467 : _GEN_1529; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1531 = 12'h5bc == _T_46[11:0] ? image_1468 : _GEN_1530; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1532 = 12'h5bd == _T_46[11:0] ? image_1469 : _GEN_1531; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1533 = 12'h5be == _T_46[11:0] ? 4'h0 : _GEN_1532; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1534 = 12'h5bf == _T_46[11:0] ? 4'h0 : _GEN_1533; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1535 = 12'h5c0 == _T_46[11:0] ? image_1472 : _GEN_1534; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1536 = 12'h5c1 == _T_46[11:0] ? image_1473 : _GEN_1535; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1537 = 12'h5c2 == _T_46[11:0] ? image_1474 : _GEN_1536; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1538 = 12'h5c3 == _T_46[11:0] ? image_1475 : _GEN_1537; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1539 = 12'h5c4 == _T_46[11:0] ? image_1476 : _GEN_1538; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1540 = 12'h5c5 == _T_46[11:0] ? image_1477 : _GEN_1539; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1541 = 12'h5c6 == _T_46[11:0] ? image_1478 : _GEN_1540; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1542 = 12'h5c7 == _T_46[11:0] ? image_1479 : _GEN_1541; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1543 = 12'h5c8 == _T_46[11:0] ? image_1480 : _GEN_1542; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1544 = 12'h5c9 == _T_46[11:0] ? image_1481 : _GEN_1543; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1545 = 12'h5ca == _T_46[11:0] ? image_1482 : _GEN_1544; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1546 = 12'h5cb == _T_46[11:0] ? image_1483 : _GEN_1545; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1547 = 12'h5cc == _T_46[11:0] ? image_1484 : _GEN_1546; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1548 = 12'h5cd == _T_46[11:0] ? image_1485 : _GEN_1547; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1549 = 12'h5ce == _T_46[11:0] ? image_1486 : _GEN_1548; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1550 = 12'h5cf == _T_46[11:0] ? image_1487 : _GEN_1549; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1551 = 12'h5d0 == _T_46[11:0] ? image_1488 : _GEN_1550; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1552 = 12'h5d1 == _T_46[11:0] ? image_1489 : _GEN_1551; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1553 = 12'h5d2 == _T_46[11:0] ? image_1490 : _GEN_1552; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1554 = 12'h5d3 == _T_46[11:0] ? image_1491 : _GEN_1553; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1555 = 12'h5d4 == _T_46[11:0] ? image_1492 : _GEN_1554; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1556 = 12'h5d5 == _T_46[11:0] ? image_1493 : _GEN_1555; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1557 = 12'h5d6 == _T_46[11:0] ? image_1494 : _GEN_1556; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1558 = 12'h5d7 == _T_46[11:0] ? image_1495 : _GEN_1557; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1559 = 12'h5d8 == _T_46[11:0] ? image_1496 : _GEN_1558; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1560 = 12'h5d9 == _T_46[11:0] ? image_1497 : _GEN_1559; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1561 = 12'h5da == _T_46[11:0] ? image_1498 : _GEN_1560; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1562 = 12'h5db == _T_46[11:0] ? image_1499 : _GEN_1561; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1563 = 12'h5dc == _T_46[11:0] ? image_1500 : _GEN_1562; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1564 = 12'h5dd == _T_46[11:0] ? image_1501 : _GEN_1563; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1565 = 12'h5de == _T_46[11:0] ? image_1502 : _GEN_1564; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1566 = 12'h5df == _T_46[11:0] ? image_1503 : _GEN_1565; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1567 = 12'h5e0 == _T_46[11:0] ? image_1504 : _GEN_1566; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1568 = 12'h5e1 == _T_46[11:0] ? image_1505 : _GEN_1567; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1569 = 12'h5e2 == _T_46[11:0] ? image_1506 : _GEN_1568; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1570 = 12'h5e3 == _T_46[11:0] ? image_1507 : _GEN_1569; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1571 = 12'h5e4 == _T_46[11:0] ? image_1508 : _GEN_1570; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1572 = 12'h5e5 == _T_46[11:0] ? image_1509 : _GEN_1571; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1573 = 12'h5e6 == _T_46[11:0] ? image_1510 : _GEN_1572; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1574 = 12'h5e7 == _T_46[11:0] ? image_1511 : _GEN_1573; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1575 = 12'h5e8 == _T_46[11:0] ? image_1512 : _GEN_1574; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1576 = 12'h5e9 == _T_46[11:0] ? image_1513 : _GEN_1575; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1577 = 12'h5ea == _T_46[11:0] ? image_1514 : _GEN_1576; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1578 = 12'h5eb == _T_46[11:0] ? image_1515 : _GEN_1577; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1579 = 12'h5ec == _T_46[11:0] ? image_1516 : _GEN_1578; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1580 = 12'h5ed == _T_46[11:0] ? image_1517 : _GEN_1579; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1581 = 12'h5ee == _T_46[11:0] ? image_1518 : _GEN_1580; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1582 = 12'h5ef == _T_46[11:0] ? image_1519 : _GEN_1581; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1583 = 12'h5f0 == _T_46[11:0] ? image_1520 : _GEN_1582; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1584 = 12'h5f1 == _T_46[11:0] ? image_1521 : _GEN_1583; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1585 = 12'h5f2 == _T_46[11:0] ? image_1522 : _GEN_1584; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1586 = 12'h5f3 == _T_46[11:0] ? image_1523 : _GEN_1585; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1587 = 12'h5f4 == _T_46[11:0] ? image_1524 : _GEN_1586; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1588 = 12'h5f5 == _T_46[11:0] ? image_1525 : _GEN_1587; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1589 = 12'h5f6 == _T_46[11:0] ? image_1526 : _GEN_1588; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1590 = 12'h5f7 == _T_46[11:0] ? image_1527 : _GEN_1589; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1591 = 12'h5f8 == _T_46[11:0] ? image_1528 : _GEN_1590; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1592 = 12'h5f9 == _T_46[11:0] ? image_1529 : _GEN_1591; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1593 = 12'h5fa == _T_46[11:0] ? image_1530 : _GEN_1592; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1594 = 12'h5fb == _T_46[11:0] ? image_1531 : _GEN_1593; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1595 = 12'h5fc == _T_46[11:0] ? image_1532 : _GEN_1594; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1596 = 12'h5fd == _T_46[11:0] ? image_1533 : _GEN_1595; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1597 = 12'h5fe == _T_46[11:0] ? 4'h0 : _GEN_1596; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1598 = 12'h5ff == _T_46[11:0] ? 4'h0 : _GEN_1597; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1599 = 12'h600 == _T_46[11:0] ? image_1536 : _GEN_1598; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1600 = 12'h601 == _T_46[11:0] ? image_1537 : _GEN_1599; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1601 = 12'h602 == _T_46[11:0] ? image_1538 : _GEN_1600; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1602 = 12'h603 == _T_46[11:0] ? image_1539 : _GEN_1601; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1603 = 12'h604 == _T_46[11:0] ? image_1540 : _GEN_1602; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1604 = 12'h605 == _T_46[11:0] ? image_1541 : _GEN_1603; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1605 = 12'h606 == _T_46[11:0] ? image_1542 : _GEN_1604; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1606 = 12'h607 == _T_46[11:0] ? image_1543 : _GEN_1605; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1607 = 12'h608 == _T_46[11:0] ? image_1544 : _GEN_1606; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1608 = 12'h609 == _T_46[11:0] ? image_1545 : _GEN_1607; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1609 = 12'h60a == _T_46[11:0] ? image_1546 : _GEN_1608; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1610 = 12'h60b == _T_46[11:0] ? image_1547 : _GEN_1609; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1611 = 12'h60c == _T_46[11:0] ? image_1548 : _GEN_1610; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1612 = 12'h60d == _T_46[11:0] ? image_1549 : _GEN_1611; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1613 = 12'h60e == _T_46[11:0] ? image_1550 : _GEN_1612; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1614 = 12'h60f == _T_46[11:0] ? image_1551 : _GEN_1613; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1615 = 12'h610 == _T_46[11:0] ? image_1552 : _GEN_1614; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1616 = 12'h611 == _T_46[11:0] ? image_1553 : _GEN_1615; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1617 = 12'h612 == _T_46[11:0] ? image_1554 : _GEN_1616; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1618 = 12'h613 == _T_46[11:0] ? image_1555 : _GEN_1617; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1619 = 12'h614 == _T_46[11:0] ? image_1556 : _GEN_1618; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1620 = 12'h615 == _T_46[11:0] ? image_1557 : _GEN_1619; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1621 = 12'h616 == _T_46[11:0] ? image_1558 : _GEN_1620; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1622 = 12'h617 == _T_46[11:0] ? image_1559 : _GEN_1621; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1623 = 12'h618 == _T_46[11:0] ? image_1560 : _GEN_1622; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1624 = 12'h619 == _T_46[11:0] ? image_1561 : _GEN_1623; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1625 = 12'h61a == _T_46[11:0] ? image_1562 : _GEN_1624; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1626 = 12'h61b == _T_46[11:0] ? image_1563 : _GEN_1625; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1627 = 12'h61c == _T_46[11:0] ? image_1564 : _GEN_1626; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1628 = 12'h61d == _T_46[11:0] ? image_1565 : _GEN_1627; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1629 = 12'h61e == _T_46[11:0] ? image_1566 : _GEN_1628; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1630 = 12'h61f == _T_46[11:0] ? image_1567 : _GEN_1629; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1631 = 12'h620 == _T_46[11:0] ? image_1568 : _GEN_1630; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1632 = 12'h621 == _T_46[11:0] ? image_1569 : _GEN_1631; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1633 = 12'h622 == _T_46[11:0] ? image_1570 : _GEN_1632; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1634 = 12'h623 == _T_46[11:0] ? image_1571 : _GEN_1633; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1635 = 12'h624 == _T_46[11:0] ? image_1572 : _GEN_1634; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1636 = 12'h625 == _T_46[11:0] ? image_1573 : _GEN_1635; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1637 = 12'h626 == _T_46[11:0] ? image_1574 : _GEN_1636; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1638 = 12'h627 == _T_46[11:0] ? image_1575 : _GEN_1637; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1639 = 12'h628 == _T_46[11:0] ? image_1576 : _GEN_1638; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1640 = 12'h629 == _T_46[11:0] ? image_1577 : _GEN_1639; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1641 = 12'h62a == _T_46[11:0] ? image_1578 : _GEN_1640; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1642 = 12'h62b == _T_46[11:0] ? image_1579 : _GEN_1641; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1643 = 12'h62c == _T_46[11:0] ? image_1580 : _GEN_1642; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1644 = 12'h62d == _T_46[11:0] ? image_1581 : _GEN_1643; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1645 = 12'h62e == _T_46[11:0] ? image_1582 : _GEN_1644; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1646 = 12'h62f == _T_46[11:0] ? image_1583 : _GEN_1645; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1647 = 12'h630 == _T_46[11:0] ? image_1584 : _GEN_1646; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1648 = 12'h631 == _T_46[11:0] ? image_1585 : _GEN_1647; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1649 = 12'h632 == _T_46[11:0] ? image_1586 : _GEN_1648; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1650 = 12'h633 == _T_46[11:0] ? image_1587 : _GEN_1649; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1651 = 12'h634 == _T_46[11:0] ? image_1588 : _GEN_1650; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1652 = 12'h635 == _T_46[11:0] ? image_1589 : _GEN_1651; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1653 = 12'h636 == _T_46[11:0] ? image_1590 : _GEN_1652; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1654 = 12'h637 == _T_46[11:0] ? image_1591 : _GEN_1653; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1655 = 12'h638 == _T_46[11:0] ? image_1592 : _GEN_1654; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1656 = 12'h639 == _T_46[11:0] ? image_1593 : _GEN_1655; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1657 = 12'h63a == _T_46[11:0] ? image_1594 : _GEN_1656; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1658 = 12'h63b == _T_46[11:0] ? image_1595 : _GEN_1657; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1659 = 12'h63c == _T_46[11:0] ? image_1596 : _GEN_1658; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1660 = 12'h63d == _T_46[11:0] ? image_1597 : _GEN_1659; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1661 = 12'h63e == _T_46[11:0] ? 4'h0 : _GEN_1660; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1662 = 12'h63f == _T_46[11:0] ? 4'h0 : _GEN_1661; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1663 = 12'h640 == _T_46[11:0] ? image_1600 : _GEN_1662; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1664 = 12'h641 == _T_46[11:0] ? image_1601 : _GEN_1663; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1665 = 12'h642 == _T_46[11:0] ? image_1602 : _GEN_1664; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1666 = 12'h643 == _T_46[11:0] ? image_1603 : _GEN_1665; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1667 = 12'h644 == _T_46[11:0] ? image_1604 : _GEN_1666; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1668 = 12'h645 == _T_46[11:0] ? image_1605 : _GEN_1667; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1669 = 12'h646 == _T_46[11:0] ? image_1606 : _GEN_1668; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1670 = 12'h647 == _T_46[11:0] ? image_1607 : _GEN_1669; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1671 = 12'h648 == _T_46[11:0] ? image_1608 : _GEN_1670; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1672 = 12'h649 == _T_46[11:0] ? image_1609 : _GEN_1671; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1673 = 12'h64a == _T_46[11:0] ? image_1610 : _GEN_1672; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1674 = 12'h64b == _T_46[11:0] ? image_1611 : _GEN_1673; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1675 = 12'h64c == _T_46[11:0] ? image_1612 : _GEN_1674; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1676 = 12'h64d == _T_46[11:0] ? image_1613 : _GEN_1675; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1677 = 12'h64e == _T_46[11:0] ? image_1614 : _GEN_1676; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1678 = 12'h64f == _T_46[11:0] ? image_1615 : _GEN_1677; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1679 = 12'h650 == _T_46[11:0] ? image_1616 : _GEN_1678; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1680 = 12'h651 == _T_46[11:0] ? image_1617 : _GEN_1679; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1681 = 12'h652 == _T_46[11:0] ? image_1618 : _GEN_1680; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1682 = 12'h653 == _T_46[11:0] ? image_1619 : _GEN_1681; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1683 = 12'h654 == _T_46[11:0] ? image_1620 : _GEN_1682; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1684 = 12'h655 == _T_46[11:0] ? image_1621 : _GEN_1683; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1685 = 12'h656 == _T_46[11:0] ? image_1622 : _GEN_1684; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1686 = 12'h657 == _T_46[11:0] ? image_1623 : _GEN_1685; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1687 = 12'h658 == _T_46[11:0] ? image_1624 : _GEN_1686; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1688 = 12'h659 == _T_46[11:0] ? image_1625 : _GEN_1687; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1689 = 12'h65a == _T_46[11:0] ? image_1626 : _GEN_1688; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1690 = 12'h65b == _T_46[11:0] ? image_1627 : _GEN_1689; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1691 = 12'h65c == _T_46[11:0] ? image_1628 : _GEN_1690; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1692 = 12'h65d == _T_46[11:0] ? image_1629 : _GEN_1691; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1693 = 12'h65e == _T_46[11:0] ? image_1630 : _GEN_1692; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1694 = 12'h65f == _T_46[11:0] ? image_1631 : _GEN_1693; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1695 = 12'h660 == _T_46[11:0] ? image_1632 : _GEN_1694; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1696 = 12'h661 == _T_46[11:0] ? image_1633 : _GEN_1695; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1697 = 12'h662 == _T_46[11:0] ? image_1634 : _GEN_1696; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1698 = 12'h663 == _T_46[11:0] ? image_1635 : _GEN_1697; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1699 = 12'h664 == _T_46[11:0] ? image_1636 : _GEN_1698; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1700 = 12'h665 == _T_46[11:0] ? image_1637 : _GEN_1699; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1701 = 12'h666 == _T_46[11:0] ? image_1638 : _GEN_1700; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1702 = 12'h667 == _T_46[11:0] ? image_1639 : _GEN_1701; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1703 = 12'h668 == _T_46[11:0] ? image_1640 : _GEN_1702; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1704 = 12'h669 == _T_46[11:0] ? image_1641 : _GEN_1703; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1705 = 12'h66a == _T_46[11:0] ? image_1642 : _GEN_1704; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1706 = 12'h66b == _T_46[11:0] ? image_1643 : _GEN_1705; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1707 = 12'h66c == _T_46[11:0] ? image_1644 : _GEN_1706; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1708 = 12'h66d == _T_46[11:0] ? image_1645 : _GEN_1707; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1709 = 12'h66e == _T_46[11:0] ? image_1646 : _GEN_1708; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1710 = 12'h66f == _T_46[11:0] ? image_1647 : _GEN_1709; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1711 = 12'h670 == _T_46[11:0] ? image_1648 : _GEN_1710; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1712 = 12'h671 == _T_46[11:0] ? image_1649 : _GEN_1711; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1713 = 12'h672 == _T_46[11:0] ? image_1650 : _GEN_1712; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1714 = 12'h673 == _T_46[11:0] ? image_1651 : _GEN_1713; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1715 = 12'h674 == _T_46[11:0] ? image_1652 : _GEN_1714; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1716 = 12'h675 == _T_46[11:0] ? image_1653 : _GEN_1715; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1717 = 12'h676 == _T_46[11:0] ? image_1654 : _GEN_1716; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1718 = 12'h677 == _T_46[11:0] ? image_1655 : _GEN_1717; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1719 = 12'h678 == _T_46[11:0] ? image_1656 : _GEN_1718; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1720 = 12'h679 == _T_46[11:0] ? image_1657 : _GEN_1719; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1721 = 12'h67a == _T_46[11:0] ? image_1658 : _GEN_1720; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1722 = 12'h67b == _T_46[11:0] ? image_1659 : _GEN_1721; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1723 = 12'h67c == _T_46[11:0] ? image_1660 : _GEN_1722; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1724 = 12'h67d == _T_46[11:0] ? 4'h0 : _GEN_1723; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1725 = 12'h67e == _T_46[11:0] ? 4'h0 : _GEN_1724; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1726 = 12'h67f == _T_46[11:0] ? 4'h0 : _GEN_1725; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1727 = 12'h680 == _T_46[11:0] ? image_1664 : _GEN_1726; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1728 = 12'h681 == _T_46[11:0] ? image_1665 : _GEN_1727; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1729 = 12'h682 == _T_46[11:0] ? image_1666 : _GEN_1728; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1730 = 12'h683 == _T_46[11:0] ? image_1667 : _GEN_1729; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1731 = 12'h684 == _T_46[11:0] ? image_1668 : _GEN_1730; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1732 = 12'h685 == _T_46[11:0] ? image_1669 : _GEN_1731; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1733 = 12'h686 == _T_46[11:0] ? image_1670 : _GEN_1732; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1734 = 12'h687 == _T_46[11:0] ? image_1671 : _GEN_1733; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1735 = 12'h688 == _T_46[11:0] ? image_1672 : _GEN_1734; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1736 = 12'h689 == _T_46[11:0] ? image_1673 : _GEN_1735; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1737 = 12'h68a == _T_46[11:0] ? image_1674 : _GEN_1736; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1738 = 12'h68b == _T_46[11:0] ? image_1675 : _GEN_1737; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1739 = 12'h68c == _T_46[11:0] ? image_1676 : _GEN_1738; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1740 = 12'h68d == _T_46[11:0] ? image_1677 : _GEN_1739; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1741 = 12'h68e == _T_46[11:0] ? image_1678 : _GEN_1740; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1742 = 12'h68f == _T_46[11:0] ? image_1679 : _GEN_1741; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1743 = 12'h690 == _T_46[11:0] ? image_1680 : _GEN_1742; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1744 = 12'h691 == _T_46[11:0] ? image_1681 : _GEN_1743; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1745 = 12'h692 == _T_46[11:0] ? image_1682 : _GEN_1744; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1746 = 12'h693 == _T_46[11:0] ? image_1683 : _GEN_1745; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1747 = 12'h694 == _T_46[11:0] ? image_1684 : _GEN_1746; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1748 = 12'h695 == _T_46[11:0] ? image_1685 : _GEN_1747; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1749 = 12'h696 == _T_46[11:0] ? image_1686 : _GEN_1748; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1750 = 12'h697 == _T_46[11:0] ? image_1687 : _GEN_1749; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1751 = 12'h698 == _T_46[11:0] ? image_1688 : _GEN_1750; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1752 = 12'h699 == _T_46[11:0] ? image_1689 : _GEN_1751; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1753 = 12'h69a == _T_46[11:0] ? image_1690 : _GEN_1752; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1754 = 12'h69b == _T_46[11:0] ? image_1691 : _GEN_1753; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1755 = 12'h69c == _T_46[11:0] ? image_1692 : _GEN_1754; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1756 = 12'h69d == _T_46[11:0] ? image_1693 : _GEN_1755; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1757 = 12'h69e == _T_46[11:0] ? image_1694 : _GEN_1756; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1758 = 12'h69f == _T_46[11:0] ? image_1695 : _GEN_1757; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1759 = 12'h6a0 == _T_46[11:0] ? image_1696 : _GEN_1758; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1760 = 12'h6a1 == _T_46[11:0] ? image_1697 : _GEN_1759; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1761 = 12'h6a2 == _T_46[11:0] ? image_1698 : _GEN_1760; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1762 = 12'h6a3 == _T_46[11:0] ? image_1699 : _GEN_1761; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1763 = 12'h6a4 == _T_46[11:0] ? image_1700 : _GEN_1762; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1764 = 12'h6a5 == _T_46[11:0] ? image_1701 : _GEN_1763; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1765 = 12'h6a6 == _T_46[11:0] ? image_1702 : _GEN_1764; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1766 = 12'h6a7 == _T_46[11:0] ? image_1703 : _GEN_1765; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1767 = 12'h6a8 == _T_46[11:0] ? image_1704 : _GEN_1766; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1768 = 12'h6a9 == _T_46[11:0] ? image_1705 : _GEN_1767; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1769 = 12'h6aa == _T_46[11:0] ? image_1706 : _GEN_1768; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1770 = 12'h6ab == _T_46[11:0] ? image_1707 : _GEN_1769; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1771 = 12'h6ac == _T_46[11:0] ? image_1708 : _GEN_1770; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1772 = 12'h6ad == _T_46[11:0] ? image_1709 : _GEN_1771; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1773 = 12'h6ae == _T_46[11:0] ? image_1710 : _GEN_1772; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1774 = 12'h6af == _T_46[11:0] ? image_1711 : _GEN_1773; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1775 = 12'h6b0 == _T_46[11:0] ? image_1712 : _GEN_1774; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1776 = 12'h6b1 == _T_46[11:0] ? image_1713 : _GEN_1775; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1777 = 12'h6b2 == _T_46[11:0] ? image_1714 : _GEN_1776; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1778 = 12'h6b3 == _T_46[11:0] ? image_1715 : _GEN_1777; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1779 = 12'h6b4 == _T_46[11:0] ? image_1716 : _GEN_1778; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1780 = 12'h6b5 == _T_46[11:0] ? image_1717 : _GEN_1779; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1781 = 12'h6b6 == _T_46[11:0] ? image_1718 : _GEN_1780; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1782 = 12'h6b7 == _T_46[11:0] ? image_1719 : _GEN_1781; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1783 = 12'h6b8 == _T_46[11:0] ? image_1720 : _GEN_1782; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1784 = 12'h6b9 == _T_46[11:0] ? image_1721 : _GEN_1783; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1785 = 12'h6ba == _T_46[11:0] ? image_1722 : _GEN_1784; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1786 = 12'h6bb == _T_46[11:0] ? image_1723 : _GEN_1785; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1787 = 12'h6bc == _T_46[11:0] ? 4'h0 : _GEN_1786; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1788 = 12'h6bd == _T_46[11:0] ? 4'h0 : _GEN_1787; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1789 = 12'h6be == _T_46[11:0] ? 4'h0 : _GEN_1788; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1790 = 12'h6bf == _T_46[11:0] ? 4'h0 : _GEN_1789; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1791 = 12'h6c0 == _T_46[11:0] ? image_1728 : _GEN_1790; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1792 = 12'h6c1 == _T_46[11:0] ? image_1729 : _GEN_1791; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1793 = 12'h6c2 == _T_46[11:0] ? image_1730 : _GEN_1792; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1794 = 12'h6c3 == _T_46[11:0] ? image_1731 : _GEN_1793; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1795 = 12'h6c4 == _T_46[11:0] ? image_1732 : _GEN_1794; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1796 = 12'h6c5 == _T_46[11:0] ? image_1733 : _GEN_1795; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1797 = 12'h6c6 == _T_46[11:0] ? image_1734 : _GEN_1796; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1798 = 12'h6c7 == _T_46[11:0] ? image_1735 : _GEN_1797; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1799 = 12'h6c8 == _T_46[11:0] ? image_1736 : _GEN_1798; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1800 = 12'h6c9 == _T_46[11:0] ? image_1737 : _GEN_1799; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1801 = 12'h6ca == _T_46[11:0] ? image_1738 : _GEN_1800; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1802 = 12'h6cb == _T_46[11:0] ? image_1739 : _GEN_1801; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1803 = 12'h6cc == _T_46[11:0] ? image_1740 : _GEN_1802; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1804 = 12'h6cd == _T_46[11:0] ? image_1741 : _GEN_1803; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1805 = 12'h6ce == _T_46[11:0] ? image_1742 : _GEN_1804; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1806 = 12'h6cf == _T_46[11:0] ? image_1743 : _GEN_1805; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1807 = 12'h6d0 == _T_46[11:0] ? image_1744 : _GEN_1806; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1808 = 12'h6d1 == _T_46[11:0] ? image_1745 : _GEN_1807; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1809 = 12'h6d2 == _T_46[11:0] ? image_1746 : _GEN_1808; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1810 = 12'h6d3 == _T_46[11:0] ? image_1747 : _GEN_1809; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1811 = 12'h6d4 == _T_46[11:0] ? image_1748 : _GEN_1810; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1812 = 12'h6d5 == _T_46[11:0] ? image_1749 : _GEN_1811; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1813 = 12'h6d6 == _T_46[11:0] ? image_1750 : _GEN_1812; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1814 = 12'h6d7 == _T_46[11:0] ? image_1751 : _GEN_1813; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1815 = 12'h6d8 == _T_46[11:0] ? image_1752 : _GEN_1814; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1816 = 12'h6d9 == _T_46[11:0] ? image_1753 : _GEN_1815; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1817 = 12'h6da == _T_46[11:0] ? image_1754 : _GEN_1816; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1818 = 12'h6db == _T_46[11:0] ? image_1755 : _GEN_1817; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1819 = 12'h6dc == _T_46[11:0] ? image_1756 : _GEN_1818; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1820 = 12'h6dd == _T_46[11:0] ? image_1757 : _GEN_1819; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1821 = 12'h6de == _T_46[11:0] ? image_1758 : _GEN_1820; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1822 = 12'h6df == _T_46[11:0] ? image_1759 : _GEN_1821; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1823 = 12'h6e0 == _T_46[11:0] ? image_1760 : _GEN_1822; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1824 = 12'h6e1 == _T_46[11:0] ? image_1761 : _GEN_1823; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1825 = 12'h6e2 == _T_46[11:0] ? image_1762 : _GEN_1824; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1826 = 12'h6e3 == _T_46[11:0] ? image_1763 : _GEN_1825; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1827 = 12'h6e4 == _T_46[11:0] ? image_1764 : _GEN_1826; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1828 = 12'h6e5 == _T_46[11:0] ? image_1765 : _GEN_1827; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1829 = 12'h6e6 == _T_46[11:0] ? image_1766 : _GEN_1828; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1830 = 12'h6e7 == _T_46[11:0] ? image_1767 : _GEN_1829; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1831 = 12'h6e8 == _T_46[11:0] ? image_1768 : _GEN_1830; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1832 = 12'h6e9 == _T_46[11:0] ? image_1769 : _GEN_1831; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1833 = 12'h6ea == _T_46[11:0] ? image_1770 : _GEN_1832; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1834 = 12'h6eb == _T_46[11:0] ? image_1771 : _GEN_1833; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1835 = 12'h6ec == _T_46[11:0] ? image_1772 : _GEN_1834; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1836 = 12'h6ed == _T_46[11:0] ? image_1773 : _GEN_1835; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1837 = 12'h6ee == _T_46[11:0] ? image_1774 : _GEN_1836; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1838 = 12'h6ef == _T_46[11:0] ? image_1775 : _GEN_1837; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1839 = 12'h6f0 == _T_46[11:0] ? image_1776 : _GEN_1838; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1840 = 12'h6f1 == _T_46[11:0] ? image_1777 : _GEN_1839; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1841 = 12'h6f2 == _T_46[11:0] ? image_1778 : _GEN_1840; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1842 = 12'h6f3 == _T_46[11:0] ? image_1779 : _GEN_1841; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1843 = 12'h6f4 == _T_46[11:0] ? image_1780 : _GEN_1842; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1844 = 12'h6f5 == _T_46[11:0] ? image_1781 : _GEN_1843; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1845 = 12'h6f6 == _T_46[11:0] ? image_1782 : _GEN_1844; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1846 = 12'h6f7 == _T_46[11:0] ? image_1783 : _GEN_1845; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1847 = 12'h6f8 == _T_46[11:0] ? image_1784 : _GEN_1846; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1848 = 12'h6f9 == _T_46[11:0] ? image_1785 : _GEN_1847; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1849 = 12'h6fa == _T_46[11:0] ? image_1786 : _GEN_1848; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1850 = 12'h6fb == _T_46[11:0] ? 4'h0 : _GEN_1849; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1851 = 12'h6fc == _T_46[11:0] ? 4'h0 : _GEN_1850; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1852 = 12'h6fd == _T_46[11:0] ? 4'h0 : _GEN_1851; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1853 = 12'h6fe == _T_46[11:0] ? 4'h0 : _GEN_1852; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1854 = 12'h6ff == _T_46[11:0] ? 4'h0 : _GEN_1853; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1855 = 12'h700 == _T_46[11:0] ? 4'h0 : _GEN_1854; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1856 = 12'h701 == _T_46[11:0] ? image_1793 : _GEN_1855; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1857 = 12'h702 == _T_46[11:0] ? image_1794 : _GEN_1856; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1858 = 12'h703 == _T_46[11:0] ? image_1795 : _GEN_1857; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1859 = 12'h704 == _T_46[11:0] ? image_1796 : _GEN_1858; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1860 = 12'h705 == _T_46[11:0] ? image_1797 : _GEN_1859; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1861 = 12'h706 == _T_46[11:0] ? image_1798 : _GEN_1860; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1862 = 12'h707 == _T_46[11:0] ? image_1799 : _GEN_1861; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1863 = 12'h708 == _T_46[11:0] ? image_1800 : _GEN_1862; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1864 = 12'h709 == _T_46[11:0] ? image_1801 : _GEN_1863; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1865 = 12'h70a == _T_46[11:0] ? image_1802 : _GEN_1864; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1866 = 12'h70b == _T_46[11:0] ? image_1803 : _GEN_1865; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1867 = 12'h70c == _T_46[11:0] ? image_1804 : _GEN_1866; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1868 = 12'h70d == _T_46[11:0] ? image_1805 : _GEN_1867; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1869 = 12'h70e == _T_46[11:0] ? image_1806 : _GEN_1868; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1870 = 12'h70f == _T_46[11:0] ? image_1807 : _GEN_1869; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1871 = 12'h710 == _T_46[11:0] ? image_1808 : _GEN_1870; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1872 = 12'h711 == _T_46[11:0] ? image_1809 : _GEN_1871; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1873 = 12'h712 == _T_46[11:0] ? image_1810 : _GEN_1872; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1874 = 12'h713 == _T_46[11:0] ? image_1811 : _GEN_1873; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1875 = 12'h714 == _T_46[11:0] ? image_1812 : _GEN_1874; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1876 = 12'h715 == _T_46[11:0] ? image_1813 : _GEN_1875; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1877 = 12'h716 == _T_46[11:0] ? image_1814 : _GEN_1876; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1878 = 12'h717 == _T_46[11:0] ? image_1815 : _GEN_1877; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1879 = 12'h718 == _T_46[11:0] ? image_1816 : _GEN_1878; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1880 = 12'h719 == _T_46[11:0] ? image_1817 : _GEN_1879; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1881 = 12'h71a == _T_46[11:0] ? image_1818 : _GEN_1880; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1882 = 12'h71b == _T_46[11:0] ? image_1819 : _GEN_1881; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1883 = 12'h71c == _T_46[11:0] ? image_1820 : _GEN_1882; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1884 = 12'h71d == _T_46[11:0] ? image_1821 : _GEN_1883; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1885 = 12'h71e == _T_46[11:0] ? image_1822 : _GEN_1884; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1886 = 12'h71f == _T_46[11:0] ? image_1823 : _GEN_1885; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1887 = 12'h720 == _T_46[11:0] ? image_1824 : _GEN_1886; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1888 = 12'h721 == _T_46[11:0] ? image_1825 : _GEN_1887; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1889 = 12'h722 == _T_46[11:0] ? image_1826 : _GEN_1888; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1890 = 12'h723 == _T_46[11:0] ? image_1827 : _GEN_1889; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1891 = 12'h724 == _T_46[11:0] ? image_1828 : _GEN_1890; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1892 = 12'h725 == _T_46[11:0] ? image_1829 : _GEN_1891; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1893 = 12'h726 == _T_46[11:0] ? image_1830 : _GEN_1892; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1894 = 12'h727 == _T_46[11:0] ? image_1831 : _GEN_1893; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1895 = 12'h728 == _T_46[11:0] ? image_1832 : _GEN_1894; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1896 = 12'h729 == _T_46[11:0] ? image_1833 : _GEN_1895; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1897 = 12'h72a == _T_46[11:0] ? image_1834 : _GEN_1896; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1898 = 12'h72b == _T_46[11:0] ? image_1835 : _GEN_1897; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1899 = 12'h72c == _T_46[11:0] ? image_1836 : _GEN_1898; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1900 = 12'h72d == _T_46[11:0] ? image_1837 : _GEN_1899; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1901 = 12'h72e == _T_46[11:0] ? image_1838 : _GEN_1900; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1902 = 12'h72f == _T_46[11:0] ? image_1839 : _GEN_1901; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1903 = 12'h730 == _T_46[11:0] ? image_1840 : _GEN_1902; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1904 = 12'h731 == _T_46[11:0] ? image_1841 : _GEN_1903; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1905 = 12'h732 == _T_46[11:0] ? image_1842 : _GEN_1904; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1906 = 12'h733 == _T_46[11:0] ? image_1843 : _GEN_1905; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1907 = 12'h734 == _T_46[11:0] ? image_1844 : _GEN_1906; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1908 = 12'h735 == _T_46[11:0] ? image_1845 : _GEN_1907; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1909 = 12'h736 == _T_46[11:0] ? image_1846 : _GEN_1908; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1910 = 12'h737 == _T_46[11:0] ? image_1847 : _GEN_1909; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1911 = 12'h738 == _T_46[11:0] ? image_1848 : _GEN_1910; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1912 = 12'h739 == _T_46[11:0] ? image_1849 : _GEN_1911; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1913 = 12'h73a == _T_46[11:0] ? 4'h0 : _GEN_1912; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1914 = 12'h73b == _T_46[11:0] ? 4'h0 : _GEN_1913; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1915 = 12'h73c == _T_46[11:0] ? 4'h0 : _GEN_1914; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1916 = 12'h73d == _T_46[11:0] ? 4'h0 : _GEN_1915; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1917 = 12'h73e == _T_46[11:0] ? 4'h0 : _GEN_1916; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1918 = 12'h73f == _T_46[11:0] ? 4'h0 : _GEN_1917; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1919 = 12'h740 == _T_46[11:0] ? 4'h0 : _GEN_1918; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1920 = 12'h741 == _T_46[11:0] ? image_1857 : _GEN_1919; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1921 = 12'h742 == _T_46[11:0] ? image_1858 : _GEN_1920; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1922 = 12'h743 == _T_46[11:0] ? image_1859 : _GEN_1921; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1923 = 12'h744 == _T_46[11:0] ? image_1860 : _GEN_1922; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1924 = 12'h745 == _T_46[11:0] ? image_1861 : _GEN_1923; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1925 = 12'h746 == _T_46[11:0] ? image_1862 : _GEN_1924; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1926 = 12'h747 == _T_46[11:0] ? image_1863 : _GEN_1925; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1927 = 12'h748 == _T_46[11:0] ? image_1864 : _GEN_1926; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1928 = 12'h749 == _T_46[11:0] ? image_1865 : _GEN_1927; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1929 = 12'h74a == _T_46[11:0] ? image_1866 : _GEN_1928; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1930 = 12'h74b == _T_46[11:0] ? image_1867 : _GEN_1929; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1931 = 12'h74c == _T_46[11:0] ? image_1868 : _GEN_1930; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1932 = 12'h74d == _T_46[11:0] ? image_1869 : _GEN_1931; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1933 = 12'h74e == _T_46[11:0] ? image_1870 : _GEN_1932; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1934 = 12'h74f == _T_46[11:0] ? image_1871 : _GEN_1933; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1935 = 12'h750 == _T_46[11:0] ? image_1872 : _GEN_1934; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1936 = 12'h751 == _T_46[11:0] ? image_1873 : _GEN_1935; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1937 = 12'h752 == _T_46[11:0] ? image_1874 : _GEN_1936; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1938 = 12'h753 == _T_46[11:0] ? image_1875 : _GEN_1937; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1939 = 12'h754 == _T_46[11:0] ? image_1876 : _GEN_1938; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1940 = 12'h755 == _T_46[11:0] ? image_1877 : _GEN_1939; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1941 = 12'h756 == _T_46[11:0] ? image_1878 : _GEN_1940; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1942 = 12'h757 == _T_46[11:0] ? image_1879 : _GEN_1941; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1943 = 12'h758 == _T_46[11:0] ? image_1880 : _GEN_1942; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1944 = 12'h759 == _T_46[11:0] ? image_1881 : _GEN_1943; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1945 = 12'h75a == _T_46[11:0] ? image_1882 : _GEN_1944; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1946 = 12'h75b == _T_46[11:0] ? image_1883 : _GEN_1945; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1947 = 12'h75c == _T_46[11:0] ? image_1884 : _GEN_1946; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1948 = 12'h75d == _T_46[11:0] ? image_1885 : _GEN_1947; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1949 = 12'h75e == _T_46[11:0] ? image_1886 : _GEN_1948; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1950 = 12'h75f == _T_46[11:0] ? image_1887 : _GEN_1949; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1951 = 12'h760 == _T_46[11:0] ? image_1888 : _GEN_1950; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1952 = 12'h761 == _T_46[11:0] ? image_1889 : _GEN_1951; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1953 = 12'h762 == _T_46[11:0] ? image_1890 : _GEN_1952; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1954 = 12'h763 == _T_46[11:0] ? image_1891 : _GEN_1953; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1955 = 12'h764 == _T_46[11:0] ? image_1892 : _GEN_1954; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1956 = 12'h765 == _T_46[11:0] ? image_1893 : _GEN_1955; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1957 = 12'h766 == _T_46[11:0] ? image_1894 : _GEN_1956; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1958 = 12'h767 == _T_46[11:0] ? image_1895 : _GEN_1957; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1959 = 12'h768 == _T_46[11:0] ? image_1896 : _GEN_1958; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1960 = 12'h769 == _T_46[11:0] ? image_1897 : _GEN_1959; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1961 = 12'h76a == _T_46[11:0] ? image_1898 : _GEN_1960; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1962 = 12'h76b == _T_46[11:0] ? image_1899 : _GEN_1961; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1963 = 12'h76c == _T_46[11:0] ? image_1900 : _GEN_1962; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1964 = 12'h76d == _T_46[11:0] ? image_1901 : _GEN_1963; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1965 = 12'h76e == _T_46[11:0] ? image_1902 : _GEN_1964; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1966 = 12'h76f == _T_46[11:0] ? image_1903 : _GEN_1965; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1967 = 12'h770 == _T_46[11:0] ? image_1904 : _GEN_1966; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1968 = 12'h771 == _T_46[11:0] ? image_1905 : _GEN_1967; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1969 = 12'h772 == _T_46[11:0] ? image_1906 : _GEN_1968; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1970 = 12'h773 == _T_46[11:0] ? image_1907 : _GEN_1969; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1971 = 12'h774 == _T_46[11:0] ? image_1908 : _GEN_1970; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1972 = 12'h775 == _T_46[11:0] ? image_1909 : _GEN_1971; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1973 = 12'h776 == _T_46[11:0] ? image_1910 : _GEN_1972; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1974 = 12'h777 == _T_46[11:0] ? image_1911 : _GEN_1973; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1975 = 12'h778 == _T_46[11:0] ? image_1912 : _GEN_1974; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1976 = 12'h779 == _T_46[11:0] ? image_1913 : _GEN_1975; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1977 = 12'h77a == _T_46[11:0] ? 4'h0 : _GEN_1976; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1978 = 12'h77b == _T_46[11:0] ? 4'h0 : _GEN_1977; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1979 = 12'h77c == _T_46[11:0] ? 4'h0 : _GEN_1978; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1980 = 12'h77d == _T_46[11:0] ? 4'h0 : _GEN_1979; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1981 = 12'h77e == _T_46[11:0] ? 4'h0 : _GEN_1980; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1982 = 12'h77f == _T_46[11:0] ? 4'h0 : _GEN_1981; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1983 = 12'h780 == _T_46[11:0] ? 4'h0 : _GEN_1982; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1984 = 12'h781 == _T_46[11:0] ? image_1921 : _GEN_1983; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1985 = 12'h782 == _T_46[11:0] ? image_1922 : _GEN_1984; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1986 = 12'h783 == _T_46[11:0] ? image_1923 : _GEN_1985; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1987 = 12'h784 == _T_46[11:0] ? image_1924 : _GEN_1986; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1988 = 12'h785 == _T_46[11:0] ? image_1925 : _GEN_1987; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1989 = 12'h786 == _T_46[11:0] ? image_1926 : _GEN_1988; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1990 = 12'h787 == _T_46[11:0] ? image_1927 : _GEN_1989; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1991 = 12'h788 == _T_46[11:0] ? image_1928 : _GEN_1990; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1992 = 12'h789 == _T_46[11:0] ? image_1929 : _GEN_1991; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1993 = 12'h78a == _T_46[11:0] ? image_1930 : _GEN_1992; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1994 = 12'h78b == _T_46[11:0] ? image_1931 : _GEN_1993; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1995 = 12'h78c == _T_46[11:0] ? image_1932 : _GEN_1994; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1996 = 12'h78d == _T_46[11:0] ? image_1933 : _GEN_1995; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1997 = 12'h78e == _T_46[11:0] ? image_1934 : _GEN_1996; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1998 = 12'h78f == _T_46[11:0] ? image_1935 : _GEN_1997; // @[Filter.scala 138:46]
  wire [3:0] _GEN_1999 = 12'h790 == _T_46[11:0] ? image_1936 : _GEN_1998; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2000 = 12'h791 == _T_46[11:0] ? image_1937 : _GEN_1999; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2001 = 12'h792 == _T_46[11:0] ? image_1938 : _GEN_2000; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2002 = 12'h793 == _T_46[11:0] ? image_1939 : _GEN_2001; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2003 = 12'h794 == _T_46[11:0] ? image_1940 : _GEN_2002; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2004 = 12'h795 == _T_46[11:0] ? image_1941 : _GEN_2003; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2005 = 12'h796 == _T_46[11:0] ? image_1942 : _GEN_2004; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2006 = 12'h797 == _T_46[11:0] ? image_1943 : _GEN_2005; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2007 = 12'h798 == _T_46[11:0] ? image_1944 : _GEN_2006; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2008 = 12'h799 == _T_46[11:0] ? image_1945 : _GEN_2007; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2009 = 12'h79a == _T_46[11:0] ? image_1946 : _GEN_2008; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2010 = 12'h79b == _T_46[11:0] ? image_1947 : _GEN_2009; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2011 = 12'h79c == _T_46[11:0] ? image_1948 : _GEN_2010; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2012 = 12'h79d == _T_46[11:0] ? image_1949 : _GEN_2011; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2013 = 12'h79e == _T_46[11:0] ? image_1950 : _GEN_2012; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2014 = 12'h79f == _T_46[11:0] ? image_1951 : _GEN_2013; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2015 = 12'h7a0 == _T_46[11:0] ? image_1952 : _GEN_2014; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2016 = 12'h7a1 == _T_46[11:0] ? image_1953 : _GEN_2015; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2017 = 12'h7a2 == _T_46[11:0] ? image_1954 : _GEN_2016; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2018 = 12'h7a3 == _T_46[11:0] ? image_1955 : _GEN_2017; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2019 = 12'h7a4 == _T_46[11:0] ? image_1956 : _GEN_2018; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2020 = 12'h7a5 == _T_46[11:0] ? image_1957 : _GEN_2019; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2021 = 12'h7a6 == _T_46[11:0] ? image_1958 : _GEN_2020; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2022 = 12'h7a7 == _T_46[11:0] ? image_1959 : _GEN_2021; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2023 = 12'h7a8 == _T_46[11:0] ? image_1960 : _GEN_2022; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2024 = 12'h7a9 == _T_46[11:0] ? image_1961 : _GEN_2023; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2025 = 12'h7aa == _T_46[11:0] ? image_1962 : _GEN_2024; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2026 = 12'h7ab == _T_46[11:0] ? image_1963 : _GEN_2025; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2027 = 12'h7ac == _T_46[11:0] ? image_1964 : _GEN_2026; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2028 = 12'h7ad == _T_46[11:0] ? image_1965 : _GEN_2027; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2029 = 12'h7ae == _T_46[11:0] ? image_1966 : _GEN_2028; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2030 = 12'h7af == _T_46[11:0] ? image_1967 : _GEN_2029; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2031 = 12'h7b0 == _T_46[11:0] ? image_1968 : _GEN_2030; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2032 = 12'h7b1 == _T_46[11:0] ? image_1969 : _GEN_2031; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2033 = 12'h7b2 == _T_46[11:0] ? image_1970 : _GEN_2032; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2034 = 12'h7b3 == _T_46[11:0] ? image_1971 : _GEN_2033; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2035 = 12'h7b4 == _T_46[11:0] ? image_1972 : _GEN_2034; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2036 = 12'h7b5 == _T_46[11:0] ? image_1973 : _GEN_2035; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2037 = 12'h7b6 == _T_46[11:0] ? image_1974 : _GEN_2036; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2038 = 12'h7b7 == _T_46[11:0] ? image_1975 : _GEN_2037; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2039 = 12'h7b8 == _T_46[11:0] ? image_1976 : _GEN_2038; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2040 = 12'h7b9 == _T_46[11:0] ? image_1977 : _GEN_2039; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2041 = 12'h7ba == _T_46[11:0] ? 4'h0 : _GEN_2040; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2042 = 12'h7bb == _T_46[11:0] ? 4'h0 : _GEN_2041; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2043 = 12'h7bc == _T_46[11:0] ? 4'h0 : _GEN_2042; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2044 = 12'h7bd == _T_46[11:0] ? 4'h0 : _GEN_2043; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2045 = 12'h7be == _T_46[11:0] ? 4'h0 : _GEN_2044; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2046 = 12'h7bf == _T_46[11:0] ? 4'h0 : _GEN_2045; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2047 = 12'h7c0 == _T_46[11:0] ? 4'h0 : _GEN_2046; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2048 = 12'h7c1 == _T_46[11:0] ? image_1985 : _GEN_2047; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2049 = 12'h7c2 == _T_46[11:0] ? image_1986 : _GEN_2048; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2050 = 12'h7c3 == _T_46[11:0] ? image_1987 : _GEN_2049; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2051 = 12'h7c4 == _T_46[11:0] ? image_1988 : _GEN_2050; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2052 = 12'h7c5 == _T_46[11:0] ? image_1989 : _GEN_2051; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2053 = 12'h7c6 == _T_46[11:0] ? image_1990 : _GEN_2052; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2054 = 12'h7c7 == _T_46[11:0] ? image_1991 : _GEN_2053; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2055 = 12'h7c8 == _T_46[11:0] ? image_1992 : _GEN_2054; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2056 = 12'h7c9 == _T_46[11:0] ? image_1993 : _GEN_2055; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2057 = 12'h7ca == _T_46[11:0] ? image_1994 : _GEN_2056; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2058 = 12'h7cb == _T_46[11:0] ? image_1995 : _GEN_2057; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2059 = 12'h7cc == _T_46[11:0] ? image_1996 : _GEN_2058; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2060 = 12'h7cd == _T_46[11:0] ? image_1997 : _GEN_2059; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2061 = 12'h7ce == _T_46[11:0] ? image_1998 : _GEN_2060; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2062 = 12'h7cf == _T_46[11:0] ? image_1999 : _GEN_2061; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2063 = 12'h7d0 == _T_46[11:0] ? image_2000 : _GEN_2062; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2064 = 12'h7d1 == _T_46[11:0] ? image_2001 : _GEN_2063; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2065 = 12'h7d2 == _T_46[11:0] ? image_2002 : _GEN_2064; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2066 = 12'h7d3 == _T_46[11:0] ? image_2003 : _GEN_2065; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2067 = 12'h7d4 == _T_46[11:0] ? image_2004 : _GEN_2066; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2068 = 12'h7d5 == _T_46[11:0] ? image_2005 : _GEN_2067; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2069 = 12'h7d6 == _T_46[11:0] ? image_2006 : _GEN_2068; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2070 = 12'h7d7 == _T_46[11:0] ? image_2007 : _GEN_2069; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2071 = 12'h7d8 == _T_46[11:0] ? image_2008 : _GEN_2070; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2072 = 12'h7d9 == _T_46[11:0] ? image_2009 : _GEN_2071; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2073 = 12'h7da == _T_46[11:0] ? image_2010 : _GEN_2072; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2074 = 12'h7db == _T_46[11:0] ? image_2011 : _GEN_2073; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2075 = 12'h7dc == _T_46[11:0] ? image_2012 : _GEN_2074; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2076 = 12'h7dd == _T_46[11:0] ? image_2013 : _GEN_2075; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2077 = 12'h7de == _T_46[11:0] ? image_2014 : _GEN_2076; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2078 = 12'h7df == _T_46[11:0] ? image_2015 : _GEN_2077; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2079 = 12'h7e0 == _T_46[11:0] ? image_2016 : _GEN_2078; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2080 = 12'h7e1 == _T_46[11:0] ? image_2017 : _GEN_2079; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2081 = 12'h7e2 == _T_46[11:0] ? image_2018 : _GEN_2080; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2082 = 12'h7e3 == _T_46[11:0] ? image_2019 : _GEN_2081; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2083 = 12'h7e4 == _T_46[11:0] ? image_2020 : _GEN_2082; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2084 = 12'h7e5 == _T_46[11:0] ? image_2021 : _GEN_2083; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2085 = 12'h7e6 == _T_46[11:0] ? image_2022 : _GEN_2084; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2086 = 12'h7e7 == _T_46[11:0] ? image_2023 : _GEN_2085; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2087 = 12'h7e8 == _T_46[11:0] ? image_2024 : _GEN_2086; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2088 = 12'h7e9 == _T_46[11:0] ? image_2025 : _GEN_2087; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2089 = 12'h7ea == _T_46[11:0] ? image_2026 : _GEN_2088; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2090 = 12'h7eb == _T_46[11:0] ? image_2027 : _GEN_2089; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2091 = 12'h7ec == _T_46[11:0] ? image_2028 : _GEN_2090; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2092 = 12'h7ed == _T_46[11:0] ? image_2029 : _GEN_2091; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2093 = 12'h7ee == _T_46[11:0] ? image_2030 : _GEN_2092; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2094 = 12'h7ef == _T_46[11:0] ? image_2031 : _GEN_2093; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2095 = 12'h7f0 == _T_46[11:0] ? image_2032 : _GEN_2094; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2096 = 12'h7f1 == _T_46[11:0] ? image_2033 : _GEN_2095; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2097 = 12'h7f2 == _T_46[11:0] ? image_2034 : _GEN_2096; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2098 = 12'h7f3 == _T_46[11:0] ? image_2035 : _GEN_2097; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2099 = 12'h7f4 == _T_46[11:0] ? image_2036 : _GEN_2098; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2100 = 12'h7f5 == _T_46[11:0] ? image_2037 : _GEN_2099; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2101 = 12'h7f6 == _T_46[11:0] ? image_2038 : _GEN_2100; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2102 = 12'h7f7 == _T_46[11:0] ? image_2039 : _GEN_2101; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2103 = 12'h7f8 == _T_46[11:0] ? image_2040 : _GEN_2102; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2104 = 12'h7f9 == _T_46[11:0] ? image_2041 : _GEN_2103; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2105 = 12'h7fa == _T_46[11:0] ? 4'h0 : _GEN_2104; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2106 = 12'h7fb == _T_46[11:0] ? 4'h0 : _GEN_2105; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2107 = 12'h7fc == _T_46[11:0] ? 4'h0 : _GEN_2106; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2108 = 12'h7fd == _T_46[11:0] ? 4'h0 : _GEN_2107; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2109 = 12'h7fe == _T_46[11:0] ? 4'h0 : _GEN_2108; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2110 = 12'h7ff == _T_46[11:0] ? 4'h0 : _GEN_2109; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2111 = 12'h800 == _T_46[11:0] ? 4'h0 : _GEN_2110; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2112 = 12'h801 == _T_46[11:0] ? image_2049 : _GEN_2111; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2113 = 12'h802 == _T_46[11:0] ? image_2050 : _GEN_2112; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2114 = 12'h803 == _T_46[11:0] ? image_2051 : _GEN_2113; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2115 = 12'h804 == _T_46[11:0] ? image_2052 : _GEN_2114; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2116 = 12'h805 == _T_46[11:0] ? image_2053 : _GEN_2115; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2117 = 12'h806 == _T_46[11:0] ? image_2054 : _GEN_2116; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2118 = 12'h807 == _T_46[11:0] ? image_2055 : _GEN_2117; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2119 = 12'h808 == _T_46[11:0] ? image_2056 : _GEN_2118; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2120 = 12'h809 == _T_46[11:0] ? image_2057 : _GEN_2119; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2121 = 12'h80a == _T_46[11:0] ? image_2058 : _GEN_2120; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2122 = 12'h80b == _T_46[11:0] ? image_2059 : _GEN_2121; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2123 = 12'h80c == _T_46[11:0] ? image_2060 : _GEN_2122; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2124 = 12'h80d == _T_46[11:0] ? image_2061 : _GEN_2123; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2125 = 12'h80e == _T_46[11:0] ? image_2062 : _GEN_2124; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2126 = 12'h80f == _T_46[11:0] ? image_2063 : _GEN_2125; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2127 = 12'h810 == _T_46[11:0] ? image_2064 : _GEN_2126; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2128 = 12'h811 == _T_46[11:0] ? image_2065 : _GEN_2127; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2129 = 12'h812 == _T_46[11:0] ? image_2066 : _GEN_2128; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2130 = 12'h813 == _T_46[11:0] ? image_2067 : _GEN_2129; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2131 = 12'h814 == _T_46[11:0] ? image_2068 : _GEN_2130; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2132 = 12'h815 == _T_46[11:0] ? image_2069 : _GEN_2131; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2133 = 12'h816 == _T_46[11:0] ? image_2070 : _GEN_2132; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2134 = 12'h817 == _T_46[11:0] ? image_2071 : _GEN_2133; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2135 = 12'h818 == _T_46[11:0] ? image_2072 : _GEN_2134; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2136 = 12'h819 == _T_46[11:0] ? image_2073 : _GEN_2135; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2137 = 12'h81a == _T_46[11:0] ? image_2074 : _GEN_2136; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2138 = 12'h81b == _T_46[11:0] ? image_2075 : _GEN_2137; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2139 = 12'h81c == _T_46[11:0] ? image_2076 : _GEN_2138; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2140 = 12'h81d == _T_46[11:0] ? image_2077 : _GEN_2139; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2141 = 12'h81e == _T_46[11:0] ? image_2078 : _GEN_2140; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2142 = 12'h81f == _T_46[11:0] ? image_2079 : _GEN_2141; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2143 = 12'h820 == _T_46[11:0] ? image_2080 : _GEN_2142; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2144 = 12'h821 == _T_46[11:0] ? image_2081 : _GEN_2143; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2145 = 12'h822 == _T_46[11:0] ? image_2082 : _GEN_2144; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2146 = 12'h823 == _T_46[11:0] ? image_2083 : _GEN_2145; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2147 = 12'h824 == _T_46[11:0] ? image_2084 : _GEN_2146; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2148 = 12'h825 == _T_46[11:0] ? image_2085 : _GEN_2147; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2149 = 12'h826 == _T_46[11:0] ? image_2086 : _GEN_2148; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2150 = 12'h827 == _T_46[11:0] ? image_2087 : _GEN_2149; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2151 = 12'h828 == _T_46[11:0] ? image_2088 : _GEN_2150; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2152 = 12'h829 == _T_46[11:0] ? image_2089 : _GEN_2151; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2153 = 12'h82a == _T_46[11:0] ? image_2090 : _GEN_2152; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2154 = 12'h82b == _T_46[11:0] ? image_2091 : _GEN_2153; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2155 = 12'h82c == _T_46[11:0] ? image_2092 : _GEN_2154; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2156 = 12'h82d == _T_46[11:0] ? image_2093 : _GEN_2155; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2157 = 12'h82e == _T_46[11:0] ? image_2094 : _GEN_2156; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2158 = 12'h82f == _T_46[11:0] ? image_2095 : _GEN_2157; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2159 = 12'h830 == _T_46[11:0] ? image_2096 : _GEN_2158; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2160 = 12'h831 == _T_46[11:0] ? image_2097 : _GEN_2159; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2161 = 12'h832 == _T_46[11:0] ? image_2098 : _GEN_2160; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2162 = 12'h833 == _T_46[11:0] ? image_2099 : _GEN_2161; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2163 = 12'h834 == _T_46[11:0] ? image_2100 : _GEN_2162; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2164 = 12'h835 == _T_46[11:0] ? image_2101 : _GEN_2163; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2165 = 12'h836 == _T_46[11:0] ? image_2102 : _GEN_2164; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2166 = 12'h837 == _T_46[11:0] ? image_2103 : _GEN_2165; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2167 = 12'h838 == _T_46[11:0] ? image_2104 : _GEN_2166; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2168 = 12'h839 == _T_46[11:0] ? image_2105 : _GEN_2167; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2169 = 12'h83a == _T_46[11:0] ? image_2106 : _GEN_2168; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2170 = 12'h83b == _T_46[11:0] ? 4'h0 : _GEN_2169; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2171 = 12'h83c == _T_46[11:0] ? 4'h0 : _GEN_2170; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2172 = 12'h83d == _T_46[11:0] ? 4'h0 : _GEN_2171; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2173 = 12'h83e == _T_46[11:0] ? 4'h0 : _GEN_2172; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2174 = 12'h83f == _T_46[11:0] ? 4'h0 : _GEN_2173; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2175 = 12'h840 == _T_46[11:0] ? 4'h0 : _GEN_2174; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2176 = 12'h841 == _T_46[11:0] ? 4'h0 : _GEN_2175; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2177 = 12'h842 == _T_46[11:0] ? image_2114 : _GEN_2176; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2178 = 12'h843 == _T_46[11:0] ? image_2115 : _GEN_2177; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2179 = 12'h844 == _T_46[11:0] ? image_2116 : _GEN_2178; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2180 = 12'h845 == _T_46[11:0] ? image_2117 : _GEN_2179; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2181 = 12'h846 == _T_46[11:0] ? image_2118 : _GEN_2180; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2182 = 12'h847 == _T_46[11:0] ? image_2119 : _GEN_2181; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2183 = 12'h848 == _T_46[11:0] ? image_2120 : _GEN_2182; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2184 = 12'h849 == _T_46[11:0] ? image_2121 : _GEN_2183; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2185 = 12'h84a == _T_46[11:0] ? image_2122 : _GEN_2184; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2186 = 12'h84b == _T_46[11:0] ? image_2123 : _GEN_2185; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2187 = 12'h84c == _T_46[11:0] ? image_2124 : _GEN_2186; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2188 = 12'h84d == _T_46[11:0] ? image_2125 : _GEN_2187; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2189 = 12'h84e == _T_46[11:0] ? image_2126 : _GEN_2188; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2190 = 12'h84f == _T_46[11:0] ? image_2127 : _GEN_2189; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2191 = 12'h850 == _T_46[11:0] ? image_2128 : _GEN_2190; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2192 = 12'h851 == _T_46[11:0] ? image_2129 : _GEN_2191; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2193 = 12'h852 == _T_46[11:0] ? image_2130 : _GEN_2192; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2194 = 12'h853 == _T_46[11:0] ? image_2131 : _GEN_2193; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2195 = 12'h854 == _T_46[11:0] ? image_2132 : _GEN_2194; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2196 = 12'h855 == _T_46[11:0] ? image_2133 : _GEN_2195; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2197 = 12'h856 == _T_46[11:0] ? image_2134 : _GEN_2196; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2198 = 12'h857 == _T_46[11:0] ? image_2135 : _GEN_2197; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2199 = 12'h858 == _T_46[11:0] ? image_2136 : _GEN_2198; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2200 = 12'h859 == _T_46[11:0] ? image_2137 : _GEN_2199; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2201 = 12'h85a == _T_46[11:0] ? image_2138 : _GEN_2200; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2202 = 12'h85b == _T_46[11:0] ? image_2139 : _GEN_2201; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2203 = 12'h85c == _T_46[11:0] ? image_2140 : _GEN_2202; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2204 = 12'h85d == _T_46[11:0] ? image_2141 : _GEN_2203; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2205 = 12'h85e == _T_46[11:0] ? image_2142 : _GEN_2204; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2206 = 12'h85f == _T_46[11:0] ? image_2143 : _GEN_2205; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2207 = 12'h860 == _T_46[11:0] ? image_2144 : _GEN_2206; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2208 = 12'h861 == _T_46[11:0] ? image_2145 : _GEN_2207; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2209 = 12'h862 == _T_46[11:0] ? image_2146 : _GEN_2208; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2210 = 12'h863 == _T_46[11:0] ? image_2147 : _GEN_2209; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2211 = 12'h864 == _T_46[11:0] ? image_2148 : _GEN_2210; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2212 = 12'h865 == _T_46[11:0] ? image_2149 : _GEN_2211; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2213 = 12'h866 == _T_46[11:0] ? image_2150 : _GEN_2212; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2214 = 12'h867 == _T_46[11:0] ? image_2151 : _GEN_2213; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2215 = 12'h868 == _T_46[11:0] ? image_2152 : _GEN_2214; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2216 = 12'h869 == _T_46[11:0] ? image_2153 : _GEN_2215; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2217 = 12'h86a == _T_46[11:0] ? image_2154 : _GEN_2216; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2218 = 12'h86b == _T_46[11:0] ? image_2155 : _GEN_2217; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2219 = 12'h86c == _T_46[11:0] ? image_2156 : _GEN_2218; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2220 = 12'h86d == _T_46[11:0] ? image_2157 : _GEN_2219; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2221 = 12'h86e == _T_46[11:0] ? image_2158 : _GEN_2220; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2222 = 12'h86f == _T_46[11:0] ? image_2159 : _GEN_2221; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2223 = 12'h870 == _T_46[11:0] ? image_2160 : _GEN_2222; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2224 = 12'h871 == _T_46[11:0] ? image_2161 : _GEN_2223; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2225 = 12'h872 == _T_46[11:0] ? image_2162 : _GEN_2224; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2226 = 12'h873 == _T_46[11:0] ? image_2163 : _GEN_2225; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2227 = 12'h874 == _T_46[11:0] ? image_2164 : _GEN_2226; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2228 = 12'h875 == _T_46[11:0] ? image_2165 : _GEN_2227; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2229 = 12'h876 == _T_46[11:0] ? image_2166 : _GEN_2228; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2230 = 12'h877 == _T_46[11:0] ? image_2167 : _GEN_2229; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2231 = 12'h878 == _T_46[11:0] ? image_2168 : _GEN_2230; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2232 = 12'h879 == _T_46[11:0] ? image_2169 : _GEN_2231; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2233 = 12'h87a == _T_46[11:0] ? image_2170 : _GEN_2232; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2234 = 12'h87b == _T_46[11:0] ? 4'h0 : _GEN_2233; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2235 = 12'h87c == _T_46[11:0] ? 4'h0 : _GEN_2234; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2236 = 12'h87d == _T_46[11:0] ? 4'h0 : _GEN_2235; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2237 = 12'h87e == _T_46[11:0] ? 4'h0 : _GEN_2236; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2238 = 12'h87f == _T_46[11:0] ? 4'h0 : _GEN_2237; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2239 = 12'h880 == _T_46[11:0] ? 4'h0 : _GEN_2238; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2240 = 12'h881 == _T_46[11:0] ? image_2177 : _GEN_2239; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2241 = 12'h882 == _T_46[11:0] ? image_2178 : _GEN_2240; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2242 = 12'h883 == _T_46[11:0] ? image_2179 : _GEN_2241; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2243 = 12'h884 == _T_46[11:0] ? image_2180 : _GEN_2242; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2244 = 12'h885 == _T_46[11:0] ? image_2181 : _GEN_2243; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2245 = 12'h886 == _T_46[11:0] ? image_2182 : _GEN_2244; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2246 = 12'h887 == _T_46[11:0] ? image_2183 : _GEN_2245; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2247 = 12'h888 == _T_46[11:0] ? image_2184 : _GEN_2246; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2248 = 12'h889 == _T_46[11:0] ? image_2185 : _GEN_2247; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2249 = 12'h88a == _T_46[11:0] ? image_2186 : _GEN_2248; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2250 = 12'h88b == _T_46[11:0] ? image_2187 : _GEN_2249; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2251 = 12'h88c == _T_46[11:0] ? image_2188 : _GEN_2250; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2252 = 12'h88d == _T_46[11:0] ? image_2189 : _GEN_2251; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2253 = 12'h88e == _T_46[11:0] ? image_2190 : _GEN_2252; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2254 = 12'h88f == _T_46[11:0] ? image_2191 : _GEN_2253; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2255 = 12'h890 == _T_46[11:0] ? image_2192 : _GEN_2254; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2256 = 12'h891 == _T_46[11:0] ? image_2193 : _GEN_2255; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2257 = 12'h892 == _T_46[11:0] ? image_2194 : _GEN_2256; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2258 = 12'h893 == _T_46[11:0] ? image_2195 : _GEN_2257; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2259 = 12'h894 == _T_46[11:0] ? image_2196 : _GEN_2258; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2260 = 12'h895 == _T_46[11:0] ? image_2197 : _GEN_2259; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2261 = 12'h896 == _T_46[11:0] ? image_2198 : _GEN_2260; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2262 = 12'h897 == _T_46[11:0] ? image_2199 : _GEN_2261; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2263 = 12'h898 == _T_46[11:0] ? image_2200 : _GEN_2262; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2264 = 12'h899 == _T_46[11:0] ? image_2201 : _GEN_2263; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2265 = 12'h89a == _T_46[11:0] ? image_2202 : _GEN_2264; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2266 = 12'h89b == _T_46[11:0] ? image_2203 : _GEN_2265; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2267 = 12'h89c == _T_46[11:0] ? image_2204 : _GEN_2266; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2268 = 12'h89d == _T_46[11:0] ? image_2205 : _GEN_2267; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2269 = 12'h89e == _T_46[11:0] ? image_2206 : _GEN_2268; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2270 = 12'h89f == _T_46[11:0] ? image_2207 : _GEN_2269; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2271 = 12'h8a0 == _T_46[11:0] ? image_2208 : _GEN_2270; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2272 = 12'h8a1 == _T_46[11:0] ? image_2209 : _GEN_2271; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2273 = 12'h8a2 == _T_46[11:0] ? image_2210 : _GEN_2272; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2274 = 12'h8a3 == _T_46[11:0] ? image_2211 : _GEN_2273; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2275 = 12'h8a4 == _T_46[11:0] ? image_2212 : _GEN_2274; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2276 = 12'h8a5 == _T_46[11:0] ? image_2213 : _GEN_2275; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2277 = 12'h8a6 == _T_46[11:0] ? image_2214 : _GEN_2276; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2278 = 12'h8a7 == _T_46[11:0] ? image_2215 : _GEN_2277; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2279 = 12'h8a8 == _T_46[11:0] ? image_2216 : _GEN_2278; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2280 = 12'h8a9 == _T_46[11:0] ? image_2217 : _GEN_2279; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2281 = 12'h8aa == _T_46[11:0] ? image_2218 : _GEN_2280; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2282 = 12'h8ab == _T_46[11:0] ? image_2219 : _GEN_2281; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2283 = 12'h8ac == _T_46[11:0] ? image_2220 : _GEN_2282; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2284 = 12'h8ad == _T_46[11:0] ? image_2221 : _GEN_2283; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2285 = 12'h8ae == _T_46[11:0] ? image_2222 : _GEN_2284; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2286 = 12'h8af == _T_46[11:0] ? image_2223 : _GEN_2285; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2287 = 12'h8b0 == _T_46[11:0] ? image_2224 : _GEN_2286; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2288 = 12'h8b1 == _T_46[11:0] ? image_2225 : _GEN_2287; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2289 = 12'h8b2 == _T_46[11:0] ? image_2226 : _GEN_2288; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2290 = 12'h8b3 == _T_46[11:0] ? image_2227 : _GEN_2289; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2291 = 12'h8b4 == _T_46[11:0] ? image_2228 : _GEN_2290; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2292 = 12'h8b5 == _T_46[11:0] ? image_2229 : _GEN_2291; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2293 = 12'h8b6 == _T_46[11:0] ? image_2230 : _GEN_2292; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2294 = 12'h8b7 == _T_46[11:0] ? image_2231 : _GEN_2293; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2295 = 12'h8b8 == _T_46[11:0] ? image_2232 : _GEN_2294; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2296 = 12'h8b9 == _T_46[11:0] ? image_2233 : _GEN_2295; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2297 = 12'h8ba == _T_46[11:0] ? image_2234 : _GEN_2296; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2298 = 12'h8bb == _T_46[11:0] ? 4'h0 : _GEN_2297; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2299 = 12'h8bc == _T_46[11:0] ? 4'h0 : _GEN_2298; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2300 = 12'h8bd == _T_46[11:0] ? 4'h0 : _GEN_2299; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2301 = 12'h8be == _T_46[11:0] ? 4'h0 : _GEN_2300; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2302 = 12'h8bf == _T_46[11:0] ? 4'h0 : _GEN_2301; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2303 = 12'h8c0 == _T_46[11:0] ? 4'h0 : _GEN_2302; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2304 = 12'h8c1 == _T_46[11:0] ? 4'h0 : _GEN_2303; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2305 = 12'h8c2 == _T_46[11:0] ? 4'h0 : _GEN_2304; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2306 = 12'h8c3 == _T_46[11:0] ? image_2243 : _GEN_2305; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2307 = 12'h8c4 == _T_46[11:0] ? image_2244 : _GEN_2306; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2308 = 12'h8c5 == _T_46[11:0] ? image_2245 : _GEN_2307; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2309 = 12'h8c6 == _T_46[11:0] ? image_2246 : _GEN_2308; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2310 = 12'h8c7 == _T_46[11:0] ? image_2247 : _GEN_2309; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2311 = 12'h8c8 == _T_46[11:0] ? image_2248 : _GEN_2310; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2312 = 12'h8c9 == _T_46[11:0] ? image_2249 : _GEN_2311; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2313 = 12'h8ca == _T_46[11:0] ? image_2250 : _GEN_2312; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2314 = 12'h8cb == _T_46[11:0] ? image_2251 : _GEN_2313; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2315 = 12'h8cc == _T_46[11:0] ? image_2252 : _GEN_2314; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2316 = 12'h8cd == _T_46[11:0] ? image_2253 : _GEN_2315; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2317 = 12'h8ce == _T_46[11:0] ? image_2254 : _GEN_2316; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2318 = 12'h8cf == _T_46[11:0] ? image_2255 : _GEN_2317; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2319 = 12'h8d0 == _T_46[11:0] ? image_2256 : _GEN_2318; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2320 = 12'h8d1 == _T_46[11:0] ? image_2257 : _GEN_2319; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2321 = 12'h8d2 == _T_46[11:0] ? image_2258 : _GEN_2320; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2322 = 12'h8d3 == _T_46[11:0] ? image_2259 : _GEN_2321; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2323 = 12'h8d4 == _T_46[11:0] ? image_2260 : _GEN_2322; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2324 = 12'h8d5 == _T_46[11:0] ? image_2261 : _GEN_2323; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2325 = 12'h8d6 == _T_46[11:0] ? image_2262 : _GEN_2324; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2326 = 12'h8d7 == _T_46[11:0] ? image_2263 : _GEN_2325; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2327 = 12'h8d8 == _T_46[11:0] ? image_2264 : _GEN_2326; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2328 = 12'h8d9 == _T_46[11:0] ? image_2265 : _GEN_2327; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2329 = 12'h8da == _T_46[11:0] ? image_2266 : _GEN_2328; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2330 = 12'h8db == _T_46[11:0] ? image_2267 : _GEN_2329; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2331 = 12'h8dc == _T_46[11:0] ? image_2268 : _GEN_2330; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2332 = 12'h8dd == _T_46[11:0] ? image_2269 : _GEN_2331; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2333 = 12'h8de == _T_46[11:0] ? image_2270 : _GEN_2332; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2334 = 12'h8df == _T_46[11:0] ? image_2271 : _GEN_2333; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2335 = 12'h8e0 == _T_46[11:0] ? image_2272 : _GEN_2334; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2336 = 12'h8e1 == _T_46[11:0] ? image_2273 : _GEN_2335; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2337 = 12'h8e2 == _T_46[11:0] ? image_2274 : _GEN_2336; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2338 = 12'h8e3 == _T_46[11:0] ? image_2275 : _GEN_2337; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2339 = 12'h8e4 == _T_46[11:0] ? image_2276 : _GEN_2338; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2340 = 12'h8e5 == _T_46[11:0] ? image_2277 : _GEN_2339; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2341 = 12'h8e6 == _T_46[11:0] ? image_2278 : _GEN_2340; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2342 = 12'h8e7 == _T_46[11:0] ? image_2279 : _GEN_2341; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2343 = 12'h8e8 == _T_46[11:0] ? image_2280 : _GEN_2342; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2344 = 12'h8e9 == _T_46[11:0] ? image_2281 : _GEN_2343; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2345 = 12'h8ea == _T_46[11:0] ? image_2282 : _GEN_2344; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2346 = 12'h8eb == _T_46[11:0] ? image_2283 : _GEN_2345; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2347 = 12'h8ec == _T_46[11:0] ? image_2284 : _GEN_2346; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2348 = 12'h8ed == _T_46[11:0] ? image_2285 : _GEN_2347; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2349 = 12'h8ee == _T_46[11:0] ? image_2286 : _GEN_2348; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2350 = 12'h8ef == _T_46[11:0] ? image_2287 : _GEN_2349; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2351 = 12'h8f0 == _T_46[11:0] ? image_2288 : _GEN_2350; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2352 = 12'h8f1 == _T_46[11:0] ? image_2289 : _GEN_2351; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2353 = 12'h8f2 == _T_46[11:0] ? image_2290 : _GEN_2352; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2354 = 12'h8f3 == _T_46[11:0] ? image_2291 : _GEN_2353; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2355 = 12'h8f4 == _T_46[11:0] ? image_2292 : _GEN_2354; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2356 = 12'h8f5 == _T_46[11:0] ? image_2293 : _GEN_2355; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2357 = 12'h8f6 == _T_46[11:0] ? image_2294 : _GEN_2356; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2358 = 12'h8f7 == _T_46[11:0] ? image_2295 : _GEN_2357; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2359 = 12'h8f8 == _T_46[11:0] ? image_2296 : _GEN_2358; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2360 = 12'h8f9 == _T_46[11:0] ? image_2297 : _GEN_2359; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2361 = 12'h8fa == _T_46[11:0] ? image_2298 : _GEN_2360; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2362 = 12'h8fb == _T_46[11:0] ? 4'h0 : _GEN_2361; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2363 = 12'h8fc == _T_46[11:0] ? 4'h0 : _GEN_2362; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2364 = 12'h8fd == _T_46[11:0] ? 4'h0 : _GEN_2363; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2365 = 12'h8fe == _T_46[11:0] ? 4'h0 : _GEN_2364; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2366 = 12'h8ff == _T_46[11:0] ? 4'h0 : _GEN_2365; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2367 = 12'h900 == _T_46[11:0] ? 4'h0 : _GEN_2366; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2368 = 12'h901 == _T_46[11:0] ? 4'h0 : _GEN_2367; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2369 = 12'h902 == _T_46[11:0] ? 4'h0 : _GEN_2368; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2370 = 12'h903 == _T_46[11:0] ? image_2307 : _GEN_2369; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2371 = 12'h904 == _T_46[11:0] ? image_2308 : _GEN_2370; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2372 = 12'h905 == _T_46[11:0] ? image_2309 : _GEN_2371; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2373 = 12'h906 == _T_46[11:0] ? image_2310 : _GEN_2372; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2374 = 12'h907 == _T_46[11:0] ? image_2311 : _GEN_2373; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2375 = 12'h908 == _T_46[11:0] ? image_2312 : _GEN_2374; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2376 = 12'h909 == _T_46[11:0] ? image_2313 : _GEN_2375; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2377 = 12'h90a == _T_46[11:0] ? image_2314 : _GEN_2376; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2378 = 12'h90b == _T_46[11:0] ? image_2315 : _GEN_2377; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2379 = 12'h90c == _T_46[11:0] ? image_2316 : _GEN_2378; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2380 = 12'h90d == _T_46[11:0] ? image_2317 : _GEN_2379; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2381 = 12'h90e == _T_46[11:0] ? image_2318 : _GEN_2380; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2382 = 12'h90f == _T_46[11:0] ? image_2319 : _GEN_2381; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2383 = 12'h910 == _T_46[11:0] ? image_2320 : _GEN_2382; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2384 = 12'h911 == _T_46[11:0] ? image_2321 : _GEN_2383; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2385 = 12'h912 == _T_46[11:0] ? image_2322 : _GEN_2384; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2386 = 12'h913 == _T_46[11:0] ? image_2323 : _GEN_2385; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2387 = 12'h914 == _T_46[11:0] ? image_2324 : _GEN_2386; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2388 = 12'h915 == _T_46[11:0] ? image_2325 : _GEN_2387; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2389 = 12'h916 == _T_46[11:0] ? image_2326 : _GEN_2388; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2390 = 12'h917 == _T_46[11:0] ? image_2327 : _GEN_2389; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2391 = 12'h918 == _T_46[11:0] ? image_2328 : _GEN_2390; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2392 = 12'h919 == _T_46[11:0] ? image_2329 : _GEN_2391; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2393 = 12'h91a == _T_46[11:0] ? image_2330 : _GEN_2392; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2394 = 12'h91b == _T_46[11:0] ? image_2331 : _GEN_2393; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2395 = 12'h91c == _T_46[11:0] ? image_2332 : _GEN_2394; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2396 = 12'h91d == _T_46[11:0] ? image_2333 : _GEN_2395; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2397 = 12'h91e == _T_46[11:0] ? image_2334 : _GEN_2396; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2398 = 12'h91f == _T_46[11:0] ? image_2335 : _GEN_2397; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2399 = 12'h920 == _T_46[11:0] ? image_2336 : _GEN_2398; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2400 = 12'h921 == _T_46[11:0] ? image_2337 : _GEN_2399; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2401 = 12'h922 == _T_46[11:0] ? image_2338 : _GEN_2400; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2402 = 12'h923 == _T_46[11:0] ? image_2339 : _GEN_2401; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2403 = 12'h924 == _T_46[11:0] ? image_2340 : _GEN_2402; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2404 = 12'h925 == _T_46[11:0] ? image_2341 : _GEN_2403; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2405 = 12'h926 == _T_46[11:0] ? image_2342 : _GEN_2404; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2406 = 12'h927 == _T_46[11:0] ? image_2343 : _GEN_2405; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2407 = 12'h928 == _T_46[11:0] ? image_2344 : _GEN_2406; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2408 = 12'h929 == _T_46[11:0] ? image_2345 : _GEN_2407; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2409 = 12'h92a == _T_46[11:0] ? image_2346 : _GEN_2408; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2410 = 12'h92b == _T_46[11:0] ? image_2347 : _GEN_2409; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2411 = 12'h92c == _T_46[11:0] ? image_2348 : _GEN_2410; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2412 = 12'h92d == _T_46[11:0] ? image_2349 : _GEN_2411; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2413 = 12'h92e == _T_46[11:0] ? image_2350 : _GEN_2412; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2414 = 12'h92f == _T_46[11:0] ? image_2351 : _GEN_2413; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2415 = 12'h930 == _T_46[11:0] ? image_2352 : _GEN_2414; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2416 = 12'h931 == _T_46[11:0] ? image_2353 : _GEN_2415; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2417 = 12'h932 == _T_46[11:0] ? image_2354 : _GEN_2416; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2418 = 12'h933 == _T_46[11:0] ? image_2355 : _GEN_2417; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2419 = 12'h934 == _T_46[11:0] ? image_2356 : _GEN_2418; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2420 = 12'h935 == _T_46[11:0] ? image_2357 : _GEN_2419; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2421 = 12'h936 == _T_46[11:0] ? image_2358 : _GEN_2420; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2422 = 12'h937 == _T_46[11:0] ? image_2359 : _GEN_2421; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2423 = 12'h938 == _T_46[11:0] ? image_2360 : _GEN_2422; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2424 = 12'h939 == _T_46[11:0] ? image_2361 : _GEN_2423; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2425 = 12'h93a == _T_46[11:0] ? image_2362 : _GEN_2424; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2426 = 12'h93b == _T_46[11:0] ? 4'h0 : _GEN_2425; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2427 = 12'h93c == _T_46[11:0] ? 4'h0 : _GEN_2426; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2428 = 12'h93d == _T_46[11:0] ? 4'h0 : _GEN_2427; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2429 = 12'h93e == _T_46[11:0] ? 4'h0 : _GEN_2428; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2430 = 12'h93f == _T_46[11:0] ? 4'h0 : _GEN_2429; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2431 = 12'h940 == _T_46[11:0] ? 4'h0 : _GEN_2430; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2432 = 12'h941 == _T_46[11:0] ? 4'h0 : _GEN_2431; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2433 = 12'h942 == _T_46[11:0] ? 4'h0 : _GEN_2432; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2434 = 12'h943 == _T_46[11:0] ? 4'h0 : _GEN_2433; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2435 = 12'h944 == _T_46[11:0] ? image_2372 : _GEN_2434; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2436 = 12'h945 == _T_46[11:0] ? image_2373 : _GEN_2435; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2437 = 12'h946 == _T_46[11:0] ? image_2374 : _GEN_2436; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2438 = 12'h947 == _T_46[11:0] ? image_2375 : _GEN_2437; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2439 = 12'h948 == _T_46[11:0] ? image_2376 : _GEN_2438; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2440 = 12'h949 == _T_46[11:0] ? image_2377 : _GEN_2439; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2441 = 12'h94a == _T_46[11:0] ? image_2378 : _GEN_2440; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2442 = 12'h94b == _T_46[11:0] ? image_2379 : _GEN_2441; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2443 = 12'h94c == _T_46[11:0] ? image_2380 : _GEN_2442; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2444 = 12'h94d == _T_46[11:0] ? image_2381 : _GEN_2443; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2445 = 12'h94e == _T_46[11:0] ? image_2382 : _GEN_2444; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2446 = 12'h94f == _T_46[11:0] ? image_2383 : _GEN_2445; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2447 = 12'h950 == _T_46[11:0] ? image_2384 : _GEN_2446; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2448 = 12'h951 == _T_46[11:0] ? image_2385 : _GEN_2447; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2449 = 12'h952 == _T_46[11:0] ? image_2386 : _GEN_2448; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2450 = 12'h953 == _T_46[11:0] ? image_2387 : _GEN_2449; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2451 = 12'h954 == _T_46[11:0] ? image_2388 : _GEN_2450; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2452 = 12'h955 == _T_46[11:0] ? image_2389 : _GEN_2451; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2453 = 12'h956 == _T_46[11:0] ? image_2390 : _GEN_2452; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2454 = 12'h957 == _T_46[11:0] ? image_2391 : _GEN_2453; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2455 = 12'h958 == _T_46[11:0] ? image_2392 : _GEN_2454; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2456 = 12'h959 == _T_46[11:0] ? image_2393 : _GEN_2455; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2457 = 12'h95a == _T_46[11:0] ? image_2394 : _GEN_2456; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2458 = 12'h95b == _T_46[11:0] ? image_2395 : _GEN_2457; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2459 = 12'h95c == _T_46[11:0] ? image_2396 : _GEN_2458; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2460 = 12'h95d == _T_46[11:0] ? image_2397 : _GEN_2459; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2461 = 12'h95e == _T_46[11:0] ? image_2398 : _GEN_2460; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2462 = 12'h95f == _T_46[11:0] ? image_2399 : _GEN_2461; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2463 = 12'h960 == _T_46[11:0] ? image_2400 : _GEN_2462; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2464 = 12'h961 == _T_46[11:0] ? image_2401 : _GEN_2463; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2465 = 12'h962 == _T_46[11:0] ? image_2402 : _GEN_2464; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2466 = 12'h963 == _T_46[11:0] ? image_2403 : _GEN_2465; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2467 = 12'h964 == _T_46[11:0] ? image_2404 : _GEN_2466; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2468 = 12'h965 == _T_46[11:0] ? image_2405 : _GEN_2467; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2469 = 12'h966 == _T_46[11:0] ? image_2406 : _GEN_2468; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2470 = 12'h967 == _T_46[11:0] ? image_2407 : _GEN_2469; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2471 = 12'h968 == _T_46[11:0] ? image_2408 : _GEN_2470; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2472 = 12'h969 == _T_46[11:0] ? image_2409 : _GEN_2471; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2473 = 12'h96a == _T_46[11:0] ? image_2410 : _GEN_2472; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2474 = 12'h96b == _T_46[11:0] ? image_2411 : _GEN_2473; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2475 = 12'h96c == _T_46[11:0] ? image_2412 : _GEN_2474; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2476 = 12'h96d == _T_46[11:0] ? image_2413 : _GEN_2475; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2477 = 12'h96e == _T_46[11:0] ? image_2414 : _GEN_2476; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2478 = 12'h96f == _T_46[11:0] ? image_2415 : _GEN_2477; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2479 = 12'h970 == _T_46[11:0] ? image_2416 : _GEN_2478; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2480 = 12'h971 == _T_46[11:0] ? image_2417 : _GEN_2479; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2481 = 12'h972 == _T_46[11:0] ? image_2418 : _GEN_2480; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2482 = 12'h973 == _T_46[11:0] ? image_2419 : _GEN_2481; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2483 = 12'h974 == _T_46[11:0] ? image_2420 : _GEN_2482; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2484 = 12'h975 == _T_46[11:0] ? image_2421 : _GEN_2483; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2485 = 12'h976 == _T_46[11:0] ? image_2422 : _GEN_2484; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2486 = 12'h977 == _T_46[11:0] ? image_2423 : _GEN_2485; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2487 = 12'h978 == _T_46[11:0] ? image_2424 : _GEN_2486; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2488 = 12'h979 == _T_46[11:0] ? image_2425 : _GEN_2487; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2489 = 12'h97a == _T_46[11:0] ? image_2426 : _GEN_2488; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2490 = 12'h97b == _T_46[11:0] ? 4'h0 : _GEN_2489; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2491 = 12'h97c == _T_46[11:0] ? 4'h0 : _GEN_2490; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2492 = 12'h97d == _T_46[11:0] ? 4'h0 : _GEN_2491; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2493 = 12'h97e == _T_46[11:0] ? 4'h0 : _GEN_2492; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2494 = 12'h97f == _T_46[11:0] ? 4'h0 : _GEN_2493; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2495 = 12'h980 == _T_46[11:0] ? 4'h0 : _GEN_2494; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2496 = 12'h981 == _T_46[11:0] ? 4'h0 : _GEN_2495; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2497 = 12'h982 == _T_46[11:0] ? 4'h0 : _GEN_2496; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2498 = 12'h983 == _T_46[11:0] ? 4'h0 : _GEN_2497; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2499 = 12'h984 == _T_46[11:0] ? 4'h0 : _GEN_2498; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2500 = 12'h985 == _T_46[11:0] ? image_2437 : _GEN_2499; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2501 = 12'h986 == _T_46[11:0] ? image_2438 : _GEN_2500; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2502 = 12'h987 == _T_46[11:0] ? image_2439 : _GEN_2501; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2503 = 12'h988 == _T_46[11:0] ? image_2440 : _GEN_2502; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2504 = 12'h989 == _T_46[11:0] ? image_2441 : _GEN_2503; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2505 = 12'h98a == _T_46[11:0] ? image_2442 : _GEN_2504; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2506 = 12'h98b == _T_46[11:0] ? image_2443 : _GEN_2505; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2507 = 12'h98c == _T_46[11:0] ? image_2444 : _GEN_2506; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2508 = 12'h98d == _T_46[11:0] ? image_2445 : _GEN_2507; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2509 = 12'h98e == _T_46[11:0] ? image_2446 : _GEN_2508; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2510 = 12'h98f == _T_46[11:0] ? image_2447 : _GEN_2509; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2511 = 12'h990 == _T_46[11:0] ? image_2448 : _GEN_2510; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2512 = 12'h991 == _T_46[11:0] ? image_2449 : _GEN_2511; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2513 = 12'h992 == _T_46[11:0] ? image_2450 : _GEN_2512; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2514 = 12'h993 == _T_46[11:0] ? image_2451 : _GEN_2513; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2515 = 12'h994 == _T_46[11:0] ? image_2452 : _GEN_2514; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2516 = 12'h995 == _T_46[11:0] ? image_2453 : _GEN_2515; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2517 = 12'h996 == _T_46[11:0] ? image_2454 : _GEN_2516; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2518 = 12'h997 == _T_46[11:0] ? image_2455 : _GEN_2517; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2519 = 12'h998 == _T_46[11:0] ? image_2456 : _GEN_2518; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2520 = 12'h999 == _T_46[11:0] ? image_2457 : _GEN_2519; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2521 = 12'h99a == _T_46[11:0] ? image_2458 : _GEN_2520; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2522 = 12'h99b == _T_46[11:0] ? image_2459 : _GEN_2521; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2523 = 12'h99c == _T_46[11:0] ? image_2460 : _GEN_2522; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2524 = 12'h99d == _T_46[11:0] ? image_2461 : _GEN_2523; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2525 = 12'h99e == _T_46[11:0] ? image_2462 : _GEN_2524; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2526 = 12'h99f == _T_46[11:0] ? image_2463 : _GEN_2525; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2527 = 12'h9a0 == _T_46[11:0] ? image_2464 : _GEN_2526; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2528 = 12'h9a1 == _T_46[11:0] ? image_2465 : _GEN_2527; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2529 = 12'h9a2 == _T_46[11:0] ? image_2466 : _GEN_2528; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2530 = 12'h9a3 == _T_46[11:0] ? image_2467 : _GEN_2529; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2531 = 12'h9a4 == _T_46[11:0] ? image_2468 : _GEN_2530; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2532 = 12'h9a5 == _T_46[11:0] ? image_2469 : _GEN_2531; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2533 = 12'h9a6 == _T_46[11:0] ? image_2470 : _GEN_2532; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2534 = 12'h9a7 == _T_46[11:0] ? image_2471 : _GEN_2533; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2535 = 12'h9a8 == _T_46[11:0] ? image_2472 : _GEN_2534; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2536 = 12'h9a9 == _T_46[11:0] ? image_2473 : _GEN_2535; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2537 = 12'h9aa == _T_46[11:0] ? image_2474 : _GEN_2536; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2538 = 12'h9ab == _T_46[11:0] ? image_2475 : _GEN_2537; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2539 = 12'h9ac == _T_46[11:0] ? image_2476 : _GEN_2538; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2540 = 12'h9ad == _T_46[11:0] ? image_2477 : _GEN_2539; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2541 = 12'h9ae == _T_46[11:0] ? image_2478 : _GEN_2540; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2542 = 12'h9af == _T_46[11:0] ? image_2479 : _GEN_2541; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2543 = 12'h9b0 == _T_46[11:0] ? image_2480 : _GEN_2542; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2544 = 12'h9b1 == _T_46[11:0] ? image_2481 : _GEN_2543; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2545 = 12'h9b2 == _T_46[11:0] ? image_2482 : _GEN_2544; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2546 = 12'h9b3 == _T_46[11:0] ? image_2483 : _GEN_2545; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2547 = 12'h9b4 == _T_46[11:0] ? image_2484 : _GEN_2546; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2548 = 12'h9b5 == _T_46[11:0] ? image_2485 : _GEN_2547; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2549 = 12'h9b6 == _T_46[11:0] ? image_2486 : _GEN_2548; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2550 = 12'h9b7 == _T_46[11:0] ? image_2487 : _GEN_2549; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2551 = 12'h9b8 == _T_46[11:0] ? image_2488 : _GEN_2550; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2552 = 12'h9b9 == _T_46[11:0] ? image_2489 : _GEN_2551; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2553 = 12'h9ba == _T_46[11:0] ? image_2490 : _GEN_2552; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2554 = 12'h9bb == _T_46[11:0] ? 4'h0 : _GEN_2553; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2555 = 12'h9bc == _T_46[11:0] ? 4'h0 : _GEN_2554; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2556 = 12'h9bd == _T_46[11:0] ? 4'h0 : _GEN_2555; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2557 = 12'h9be == _T_46[11:0] ? 4'h0 : _GEN_2556; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2558 = 12'h9bf == _T_46[11:0] ? 4'h0 : _GEN_2557; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2559 = 12'h9c0 == _T_46[11:0] ? 4'h0 : _GEN_2558; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2560 = 12'h9c1 == _T_46[11:0] ? 4'h0 : _GEN_2559; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2561 = 12'h9c2 == _T_46[11:0] ? 4'h0 : _GEN_2560; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2562 = 12'h9c3 == _T_46[11:0] ? 4'h0 : _GEN_2561; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2563 = 12'h9c4 == _T_46[11:0] ? 4'h0 : _GEN_2562; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2564 = 12'h9c5 == _T_46[11:0] ? 4'h0 : _GEN_2563; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2565 = 12'h9c6 == _T_46[11:0] ? image_2502 : _GEN_2564; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2566 = 12'h9c7 == _T_46[11:0] ? image_2503 : _GEN_2565; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2567 = 12'h9c8 == _T_46[11:0] ? image_2504 : _GEN_2566; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2568 = 12'h9c9 == _T_46[11:0] ? image_2505 : _GEN_2567; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2569 = 12'h9ca == _T_46[11:0] ? image_2506 : _GEN_2568; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2570 = 12'h9cb == _T_46[11:0] ? image_2507 : _GEN_2569; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2571 = 12'h9cc == _T_46[11:0] ? image_2508 : _GEN_2570; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2572 = 12'h9cd == _T_46[11:0] ? image_2509 : _GEN_2571; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2573 = 12'h9ce == _T_46[11:0] ? image_2510 : _GEN_2572; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2574 = 12'h9cf == _T_46[11:0] ? image_2511 : _GEN_2573; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2575 = 12'h9d0 == _T_46[11:0] ? image_2512 : _GEN_2574; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2576 = 12'h9d1 == _T_46[11:0] ? image_2513 : _GEN_2575; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2577 = 12'h9d2 == _T_46[11:0] ? image_2514 : _GEN_2576; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2578 = 12'h9d3 == _T_46[11:0] ? image_2515 : _GEN_2577; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2579 = 12'h9d4 == _T_46[11:0] ? image_2516 : _GEN_2578; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2580 = 12'h9d5 == _T_46[11:0] ? image_2517 : _GEN_2579; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2581 = 12'h9d6 == _T_46[11:0] ? image_2518 : _GEN_2580; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2582 = 12'h9d7 == _T_46[11:0] ? image_2519 : _GEN_2581; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2583 = 12'h9d8 == _T_46[11:0] ? image_2520 : _GEN_2582; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2584 = 12'h9d9 == _T_46[11:0] ? image_2521 : _GEN_2583; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2585 = 12'h9da == _T_46[11:0] ? image_2522 : _GEN_2584; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2586 = 12'h9db == _T_46[11:0] ? image_2523 : _GEN_2585; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2587 = 12'h9dc == _T_46[11:0] ? image_2524 : _GEN_2586; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2588 = 12'h9dd == _T_46[11:0] ? image_2525 : _GEN_2587; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2589 = 12'h9de == _T_46[11:0] ? image_2526 : _GEN_2588; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2590 = 12'h9df == _T_46[11:0] ? image_2527 : _GEN_2589; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2591 = 12'h9e0 == _T_46[11:0] ? image_2528 : _GEN_2590; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2592 = 12'h9e1 == _T_46[11:0] ? image_2529 : _GEN_2591; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2593 = 12'h9e2 == _T_46[11:0] ? image_2530 : _GEN_2592; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2594 = 12'h9e3 == _T_46[11:0] ? image_2531 : _GEN_2593; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2595 = 12'h9e4 == _T_46[11:0] ? image_2532 : _GEN_2594; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2596 = 12'h9e5 == _T_46[11:0] ? image_2533 : _GEN_2595; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2597 = 12'h9e6 == _T_46[11:0] ? image_2534 : _GEN_2596; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2598 = 12'h9e7 == _T_46[11:0] ? image_2535 : _GEN_2597; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2599 = 12'h9e8 == _T_46[11:0] ? image_2536 : _GEN_2598; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2600 = 12'h9e9 == _T_46[11:0] ? image_2537 : _GEN_2599; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2601 = 12'h9ea == _T_46[11:0] ? image_2538 : _GEN_2600; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2602 = 12'h9eb == _T_46[11:0] ? image_2539 : _GEN_2601; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2603 = 12'h9ec == _T_46[11:0] ? image_2540 : _GEN_2602; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2604 = 12'h9ed == _T_46[11:0] ? image_2541 : _GEN_2603; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2605 = 12'h9ee == _T_46[11:0] ? image_2542 : _GEN_2604; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2606 = 12'h9ef == _T_46[11:0] ? image_2543 : _GEN_2605; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2607 = 12'h9f0 == _T_46[11:0] ? image_2544 : _GEN_2606; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2608 = 12'h9f1 == _T_46[11:0] ? image_2545 : _GEN_2607; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2609 = 12'h9f2 == _T_46[11:0] ? image_2546 : _GEN_2608; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2610 = 12'h9f3 == _T_46[11:0] ? image_2547 : _GEN_2609; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2611 = 12'h9f4 == _T_46[11:0] ? image_2548 : _GEN_2610; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2612 = 12'h9f5 == _T_46[11:0] ? image_2549 : _GEN_2611; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2613 = 12'h9f6 == _T_46[11:0] ? image_2550 : _GEN_2612; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2614 = 12'h9f7 == _T_46[11:0] ? image_2551 : _GEN_2613; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2615 = 12'h9f8 == _T_46[11:0] ? image_2552 : _GEN_2614; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2616 = 12'h9f9 == _T_46[11:0] ? image_2553 : _GEN_2615; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2617 = 12'h9fa == _T_46[11:0] ? image_2554 : _GEN_2616; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2618 = 12'h9fb == _T_46[11:0] ? 4'h0 : _GEN_2617; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2619 = 12'h9fc == _T_46[11:0] ? 4'h0 : _GEN_2618; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2620 = 12'h9fd == _T_46[11:0] ? 4'h0 : _GEN_2619; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2621 = 12'h9fe == _T_46[11:0] ? 4'h0 : _GEN_2620; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2622 = 12'h9ff == _T_46[11:0] ? 4'h0 : _GEN_2621; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2623 = 12'ha00 == _T_46[11:0] ? 4'h0 : _GEN_2622; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2624 = 12'ha01 == _T_46[11:0] ? 4'h0 : _GEN_2623; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2625 = 12'ha02 == _T_46[11:0] ? 4'h0 : _GEN_2624; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2626 = 12'ha03 == _T_46[11:0] ? 4'h0 : _GEN_2625; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2627 = 12'ha04 == _T_46[11:0] ? 4'h0 : _GEN_2626; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2628 = 12'ha05 == _T_46[11:0] ? 4'h0 : _GEN_2627; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2629 = 12'ha06 == _T_46[11:0] ? 4'h0 : _GEN_2628; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2630 = 12'ha07 == _T_46[11:0] ? image_2567 : _GEN_2629; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2631 = 12'ha08 == _T_46[11:0] ? image_2568 : _GEN_2630; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2632 = 12'ha09 == _T_46[11:0] ? image_2569 : _GEN_2631; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2633 = 12'ha0a == _T_46[11:0] ? image_2570 : _GEN_2632; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2634 = 12'ha0b == _T_46[11:0] ? image_2571 : _GEN_2633; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2635 = 12'ha0c == _T_46[11:0] ? image_2572 : _GEN_2634; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2636 = 12'ha0d == _T_46[11:0] ? image_2573 : _GEN_2635; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2637 = 12'ha0e == _T_46[11:0] ? image_2574 : _GEN_2636; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2638 = 12'ha0f == _T_46[11:0] ? image_2575 : _GEN_2637; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2639 = 12'ha10 == _T_46[11:0] ? image_2576 : _GEN_2638; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2640 = 12'ha11 == _T_46[11:0] ? image_2577 : _GEN_2639; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2641 = 12'ha12 == _T_46[11:0] ? image_2578 : _GEN_2640; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2642 = 12'ha13 == _T_46[11:0] ? image_2579 : _GEN_2641; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2643 = 12'ha14 == _T_46[11:0] ? image_2580 : _GEN_2642; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2644 = 12'ha15 == _T_46[11:0] ? image_2581 : _GEN_2643; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2645 = 12'ha16 == _T_46[11:0] ? image_2582 : _GEN_2644; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2646 = 12'ha17 == _T_46[11:0] ? image_2583 : _GEN_2645; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2647 = 12'ha18 == _T_46[11:0] ? image_2584 : _GEN_2646; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2648 = 12'ha19 == _T_46[11:0] ? image_2585 : _GEN_2647; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2649 = 12'ha1a == _T_46[11:0] ? image_2586 : _GEN_2648; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2650 = 12'ha1b == _T_46[11:0] ? image_2587 : _GEN_2649; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2651 = 12'ha1c == _T_46[11:0] ? image_2588 : _GEN_2650; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2652 = 12'ha1d == _T_46[11:0] ? image_2589 : _GEN_2651; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2653 = 12'ha1e == _T_46[11:0] ? image_2590 : _GEN_2652; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2654 = 12'ha1f == _T_46[11:0] ? image_2591 : _GEN_2653; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2655 = 12'ha20 == _T_46[11:0] ? image_2592 : _GEN_2654; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2656 = 12'ha21 == _T_46[11:0] ? image_2593 : _GEN_2655; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2657 = 12'ha22 == _T_46[11:0] ? image_2594 : _GEN_2656; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2658 = 12'ha23 == _T_46[11:0] ? image_2595 : _GEN_2657; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2659 = 12'ha24 == _T_46[11:0] ? image_2596 : _GEN_2658; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2660 = 12'ha25 == _T_46[11:0] ? image_2597 : _GEN_2659; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2661 = 12'ha26 == _T_46[11:0] ? image_2598 : _GEN_2660; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2662 = 12'ha27 == _T_46[11:0] ? image_2599 : _GEN_2661; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2663 = 12'ha28 == _T_46[11:0] ? image_2600 : _GEN_2662; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2664 = 12'ha29 == _T_46[11:0] ? image_2601 : _GEN_2663; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2665 = 12'ha2a == _T_46[11:0] ? image_2602 : _GEN_2664; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2666 = 12'ha2b == _T_46[11:0] ? image_2603 : _GEN_2665; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2667 = 12'ha2c == _T_46[11:0] ? image_2604 : _GEN_2666; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2668 = 12'ha2d == _T_46[11:0] ? image_2605 : _GEN_2667; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2669 = 12'ha2e == _T_46[11:0] ? image_2606 : _GEN_2668; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2670 = 12'ha2f == _T_46[11:0] ? image_2607 : _GEN_2669; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2671 = 12'ha30 == _T_46[11:0] ? image_2608 : _GEN_2670; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2672 = 12'ha31 == _T_46[11:0] ? image_2609 : _GEN_2671; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2673 = 12'ha32 == _T_46[11:0] ? image_2610 : _GEN_2672; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2674 = 12'ha33 == _T_46[11:0] ? image_2611 : _GEN_2673; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2675 = 12'ha34 == _T_46[11:0] ? image_2612 : _GEN_2674; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2676 = 12'ha35 == _T_46[11:0] ? image_2613 : _GEN_2675; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2677 = 12'ha36 == _T_46[11:0] ? image_2614 : _GEN_2676; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2678 = 12'ha37 == _T_46[11:0] ? image_2615 : _GEN_2677; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2679 = 12'ha38 == _T_46[11:0] ? image_2616 : _GEN_2678; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2680 = 12'ha39 == _T_46[11:0] ? image_2617 : _GEN_2679; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2681 = 12'ha3a == _T_46[11:0] ? image_2618 : _GEN_2680; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2682 = 12'ha3b == _T_46[11:0] ? 4'h0 : _GEN_2681; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2683 = 12'ha3c == _T_46[11:0] ? 4'h0 : _GEN_2682; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2684 = 12'ha3d == _T_46[11:0] ? 4'h0 : _GEN_2683; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2685 = 12'ha3e == _T_46[11:0] ? 4'h0 : _GEN_2684; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2686 = 12'ha3f == _T_46[11:0] ? 4'h0 : _GEN_2685; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2687 = 12'ha40 == _T_46[11:0] ? 4'h0 : _GEN_2686; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2688 = 12'ha41 == _T_46[11:0] ? 4'h0 : _GEN_2687; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2689 = 12'ha42 == _T_46[11:0] ? 4'h0 : _GEN_2688; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2690 = 12'ha43 == _T_46[11:0] ? 4'h0 : _GEN_2689; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2691 = 12'ha44 == _T_46[11:0] ? 4'h0 : _GEN_2690; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2692 = 12'ha45 == _T_46[11:0] ? 4'h0 : _GEN_2691; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2693 = 12'ha46 == _T_46[11:0] ? 4'h0 : _GEN_2692; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2694 = 12'ha47 == _T_46[11:0] ? 4'h0 : _GEN_2693; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2695 = 12'ha48 == _T_46[11:0] ? image_2632 : _GEN_2694; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2696 = 12'ha49 == _T_46[11:0] ? image_2633 : _GEN_2695; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2697 = 12'ha4a == _T_46[11:0] ? image_2634 : _GEN_2696; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2698 = 12'ha4b == _T_46[11:0] ? image_2635 : _GEN_2697; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2699 = 12'ha4c == _T_46[11:0] ? image_2636 : _GEN_2698; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2700 = 12'ha4d == _T_46[11:0] ? image_2637 : _GEN_2699; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2701 = 12'ha4e == _T_46[11:0] ? image_2638 : _GEN_2700; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2702 = 12'ha4f == _T_46[11:0] ? image_2639 : _GEN_2701; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2703 = 12'ha50 == _T_46[11:0] ? image_2640 : _GEN_2702; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2704 = 12'ha51 == _T_46[11:0] ? image_2641 : _GEN_2703; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2705 = 12'ha52 == _T_46[11:0] ? image_2642 : _GEN_2704; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2706 = 12'ha53 == _T_46[11:0] ? image_2643 : _GEN_2705; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2707 = 12'ha54 == _T_46[11:0] ? image_2644 : _GEN_2706; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2708 = 12'ha55 == _T_46[11:0] ? image_2645 : _GEN_2707; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2709 = 12'ha56 == _T_46[11:0] ? image_2646 : _GEN_2708; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2710 = 12'ha57 == _T_46[11:0] ? image_2647 : _GEN_2709; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2711 = 12'ha58 == _T_46[11:0] ? image_2648 : _GEN_2710; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2712 = 12'ha59 == _T_46[11:0] ? image_2649 : _GEN_2711; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2713 = 12'ha5a == _T_46[11:0] ? image_2650 : _GEN_2712; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2714 = 12'ha5b == _T_46[11:0] ? image_2651 : _GEN_2713; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2715 = 12'ha5c == _T_46[11:0] ? image_2652 : _GEN_2714; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2716 = 12'ha5d == _T_46[11:0] ? image_2653 : _GEN_2715; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2717 = 12'ha5e == _T_46[11:0] ? image_2654 : _GEN_2716; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2718 = 12'ha5f == _T_46[11:0] ? image_2655 : _GEN_2717; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2719 = 12'ha60 == _T_46[11:0] ? image_2656 : _GEN_2718; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2720 = 12'ha61 == _T_46[11:0] ? image_2657 : _GEN_2719; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2721 = 12'ha62 == _T_46[11:0] ? image_2658 : _GEN_2720; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2722 = 12'ha63 == _T_46[11:0] ? image_2659 : _GEN_2721; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2723 = 12'ha64 == _T_46[11:0] ? image_2660 : _GEN_2722; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2724 = 12'ha65 == _T_46[11:0] ? image_2661 : _GEN_2723; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2725 = 12'ha66 == _T_46[11:0] ? image_2662 : _GEN_2724; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2726 = 12'ha67 == _T_46[11:0] ? image_2663 : _GEN_2725; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2727 = 12'ha68 == _T_46[11:0] ? image_2664 : _GEN_2726; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2728 = 12'ha69 == _T_46[11:0] ? image_2665 : _GEN_2727; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2729 = 12'ha6a == _T_46[11:0] ? image_2666 : _GEN_2728; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2730 = 12'ha6b == _T_46[11:0] ? image_2667 : _GEN_2729; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2731 = 12'ha6c == _T_46[11:0] ? image_2668 : _GEN_2730; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2732 = 12'ha6d == _T_46[11:0] ? image_2669 : _GEN_2731; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2733 = 12'ha6e == _T_46[11:0] ? image_2670 : _GEN_2732; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2734 = 12'ha6f == _T_46[11:0] ? image_2671 : _GEN_2733; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2735 = 12'ha70 == _T_46[11:0] ? image_2672 : _GEN_2734; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2736 = 12'ha71 == _T_46[11:0] ? image_2673 : _GEN_2735; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2737 = 12'ha72 == _T_46[11:0] ? image_2674 : _GEN_2736; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2738 = 12'ha73 == _T_46[11:0] ? image_2675 : _GEN_2737; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2739 = 12'ha74 == _T_46[11:0] ? image_2676 : _GEN_2738; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2740 = 12'ha75 == _T_46[11:0] ? image_2677 : _GEN_2739; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2741 = 12'ha76 == _T_46[11:0] ? image_2678 : _GEN_2740; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2742 = 12'ha77 == _T_46[11:0] ? image_2679 : _GEN_2741; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2743 = 12'ha78 == _T_46[11:0] ? image_2680 : _GEN_2742; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2744 = 12'ha79 == _T_46[11:0] ? image_2681 : _GEN_2743; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2745 = 12'ha7a == _T_46[11:0] ? image_2682 : _GEN_2744; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2746 = 12'ha7b == _T_46[11:0] ? 4'h0 : _GEN_2745; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2747 = 12'ha7c == _T_46[11:0] ? 4'h0 : _GEN_2746; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2748 = 12'ha7d == _T_46[11:0] ? 4'h0 : _GEN_2747; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2749 = 12'ha7e == _T_46[11:0] ? 4'h0 : _GEN_2748; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2750 = 12'ha7f == _T_46[11:0] ? 4'h0 : _GEN_2749; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2751 = 12'ha80 == _T_46[11:0] ? 4'h0 : _GEN_2750; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2752 = 12'ha81 == _T_46[11:0] ? 4'h0 : _GEN_2751; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2753 = 12'ha82 == _T_46[11:0] ? 4'h0 : _GEN_2752; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2754 = 12'ha83 == _T_46[11:0] ? 4'h0 : _GEN_2753; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2755 = 12'ha84 == _T_46[11:0] ? 4'h0 : _GEN_2754; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2756 = 12'ha85 == _T_46[11:0] ? 4'h0 : _GEN_2755; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2757 = 12'ha86 == _T_46[11:0] ? 4'h0 : _GEN_2756; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2758 = 12'ha87 == _T_46[11:0] ? 4'h0 : _GEN_2757; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2759 = 12'ha88 == _T_46[11:0] ? 4'h0 : _GEN_2758; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2760 = 12'ha89 == _T_46[11:0] ? image_2697 : _GEN_2759; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2761 = 12'ha8a == _T_46[11:0] ? image_2698 : _GEN_2760; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2762 = 12'ha8b == _T_46[11:0] ? image_2699 : _GEN_2761; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2763 = 12'ha8c == _T_46[11:0] ? image_2700 : _GEN_2762; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2764 = 12'ha8d == _T_46[11:0] ? image_2701 : _GEN_2763; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2765 = 12'ha8e == _T_46[11:0] ? image_2702 : _GEN_2764; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2766 = 12'ha8f == _T_46[11:0] ? image_2703 : _GEN_2765; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2767 = 12'ha90 == _T_46[11:0] ? image_2704 : _GEN_2766; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2768 = 12'ha91 == _T_46[11:0] ? image_2705 : _GEN_2767; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2769 = 12'ha92 == _T_46[11:0] ? image_2706 : _GEN_2768; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2770 = 12'ha93 == _T_46[11:0] ? image_2707 : _GEN_2769; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2771 = 12'ha94 == _T_46[11:0] ? image_2708 : _GEN_2770; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2772 = 12'ha95 == _T_46[11:0] ? image_2709 : _GEN_2771; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2773 = 12'ha96 == _T_46[11:0] ? image_2710 : _GEN_2772; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2774 = 12'ha97 == _T_46[11:0] ? image_2711 : _GEN_2773; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2775 = 12'ha98 == _T_46[11:0] ? image_2712 : _GEN_2774; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2776 = 12'ha99 == _T_46[11:0] ? image_2713 : _GEN_2775; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2777 = 12'ha9a == _T_46[11:0] ? image_2714 : _GEN_2776; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2778 = 12'ha9b == _T_46[11:0] ? image_2715 : _GEN_2777; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2779 = 12'ha9c == _T_46[11:0] ? image_2716 : _GEN_2778; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2780 = 12'ha9d == _T_46[11:0] ? image_2717 : _GEN_2779; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2781 = 12'ha9e == _T_46[11:0] ? image_2718 : _GEN_2780; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2782 = 12'ha9f == _T_46[11:0] ? image_2719 : _GEN_2781; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2783 = 12'haa0 == _T_46[11:0] ? image_2720 : _GEN_2782; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2784 = 12'haa1 == _T_46[11:0] ? image_2721 : _GEN_2783; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2785 = 12'haa2 == _T_46[11:0] ? image_2722 : _GEN_2784; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2786 = 12'haa3 == _T_46[11:0] ? image_2723 : _GEN_2785; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2787 = 12'haa4 == _T_46[11:0] ? image_2724 : _GEN_2786; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2788 = 12'haa5 == _T_46[11:0] ? image_2725 : _GEN_2787; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2789 = 12'haa6 == _T_46[11:0] ? image_2726 : _GEN_2788; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2790 = 12'haa7 == _T_46[11:0] ? image_2727 : _GEN_2789; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2791 = 12'haa8 == _T_46[11:0] ? image_2728 : _GEN_2790; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2792 = 12'haa9 == _T_46[11:0] ? image_2729 : _GEN_2791; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2793 = 12'haaa == _T_46[11:0] ? image_2730 : _GEN_2792; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2794 = 12'haab == _T_46[11:0] ? image_2731 : _GEN_2793; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2795 = 12'haac == _T_46[11:0] ? image_2732 : _GEN_2794; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2796 = 12'haad == _T_46[11:0] ? image_2733 : _GEN_2795; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2797 = 12'haae == _T_46[11:0] ? image_2734 : _GEN_2796; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2798 = 12'haaf == _T_46[11:0] ? image_2735 : _GEN_2797; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2799 = 12'hab0 == _T_46[11:0] ? image_2736 : _GEN_2798; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2800 = 12'hab1 == _T_46[11:0] ? image_2737 : _GEN_2799; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2801 = 12'hab2 == _T_46[11:0] ? image_2738 : _GEN_2800; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2802 = 12'hab3 == _T_46[11:0] ? image_2739 : _GEN_2801; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2803 = 12'hab4 == _T_46[11:0] ? image_2740 : _GEN_2802; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2804 = 12'hab5 == _T_46[11:0] ? image_2741 : _GEN_2803; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2805 = 12'hab6 == _T_46[11:0] ? image_2742 : _GEN_2804; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2806 = 12'hab7 == _T_46[11:0] ? image_2743 : _GEN_2805; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2807 = 12'hab8 == _T_46[11:0] ? image_2744 : _GEN_2806; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2808 = 12'hab9 == _T_46[11:0] ? image_2745 : _GEN_2807; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2809 = 12'haba == _T_46[11:0] ? 4'h0 : _GEN_2808; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2810 = 12'habb == _T_46[11:0] ? 4'h0 : _GEN_2809; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2811 = 12'habc == _T_46[11:0] ? 4'h0 : _GEN_2810; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2812 = 12'habd == _T_46[11:0] ? 4'h0 : _GEN_2811; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2813 = 12'habe == _T_46[11:0] ? 4'h0 : _GEN_2812; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2814 = 12'habf == _T_46[11:0] ? 4'h0 : _GEN_2813; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2815 = 12'hac0 == _T_46[11:0] ? 4'h0 : _GEN_2814; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2816 = 12'hac1 == _T_46[11:0] ? 4'h0 : _GEN_2815; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2817 = 12'hac2 == _T_46[11:0] ? 4'h0 : _GEN_2816; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2818 = 12'hac3 == _T_46[11:0] ? 4'h0 : _GEN_2817; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2819 = 12'hac4 == _T_46[11:0] ? 4'h0 : _GEN_2818; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2820 = 12'hac5 == _T_46[11:0] ? 4'h0 : _GEN_2819; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2821 = 12'hac6 == _T_46[11:0] ? 4'h0 : _GEN_2820; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2822 = 12'hac7 == _T_46[11:0] ? 4'h0 : _GEN_2821; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2823 = 12'hac8 == _T_46[11:0] ? 4'h0 : _GEN_2822; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2824 = 12'hac9 == _T_46[11:0] ? 4'h0 : _GEN_2823; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2825 = 12'haca == _T_46[11:0] ? 4'h0 : _GEN_2824; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2826 = 12'hacb == _T_46[11:0] ? image_2763 : _GEN_2825; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2827 = 12'hacc == _T_46[11:0] ? image_2764 : _GEN_2826; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2828 = 12'hacd == _T_46[11:0] ? image_2765 : _GEN_2827; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2829 = 12'hace == _T_46[11:0] ? image_2766 : _GEN_2828; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2830 = 12'hacf == _T_46[11:0] ? image_2767 : _GEN_2829; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2831 = 12'had0 == _T_46[11:0] ? image_2768 : _GEN_2830; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2832 = 12'had1 == _T_46[11:0] ? image_2769 : _GEN_2831; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2833 = 12'had2 == _T_46[11:0] ? image_2770 : _GEN_2832; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2834 = 12'had3 == _T_46[11:0] ? image_2771 : _GEN_2833; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2835 = 12'had4 == _T_46[11:0] ? image_2772 : _GEN_2834; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2836 = 12'had5 == _T_46[11:0] ? image_2773 : _GEN_2835; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2837 = 12'had6 == _T_46[11:0] ? image_2774 : _GEN_2836; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2838 = 12'had7 == _T_46[11:0] ? image_2775 : _GEN_2837; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2839 = 12'had8 == _T_46[11:0] ? image_2776 : _GEN_2838; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2840 = 12'had9 == _T_46[11:0] ? image_2777 : _GEN_2839; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2841 = 12'hada == _T_46[11:0] ? image_2778 : _GEN_2840; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2842 = 12'hadb == _T_46[11:0] ? image_2779 : _GEN_2841; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2843 = 12'hadc == _T_46[11:0] ? image_2780 : _GEN_2842; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2844 = 12'hadd == _T_46[11:0] ? image_2781 : _GEN_2843; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2845 = 12'hade == _T_46[11:0] ? image_2782 : _GEN_2844; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2846 = 12'hadf == _T_46[11:0] ? image_2783 : _GEN_2845; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2847 = 12'hae0 == _T_46[11:0] ? image_2784 : _GEN_2846; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2848 = 12'hae1 == _T_46[11:0] ? image_2785 : _GEN_2847; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2849 = 12'hae2 == _T_46[11:0] ? image_2786 : _GEN_2848; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2850 = 12'hae3 == _T_46[11:0] ? image_2787 : _GEN_2849; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2851 = 12'hae4 == _T_46[11:0] ? image_2788 : _GEN_2850; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2852 = 12'hae5 == _T_46[11:0] ? image_2789 : _GEN_2851; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2853 = 12'hae6 == _T_46[11:0] ? image_2790 : _GEN_2852; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2854 = 12'hae7 == _T_46[11:0] ? image_2791 : _GEN_2853; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2855 = 12'hae8 == _T_46[11:0] ? image_2792 : _GEN_2854; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2856 = 12'hae9 == _T_46[11:0] ? image_2793 : _GEN_2855; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2857 = 12'haea == _T_46[11:0] ? image_2794 : _GEN_2856; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2858 = 12'haeb == _T_46[11:0] ? image_2795 : _GEN_2857; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2859 = 12'haec == _T_46[11:0] ? image_2796 : _GEN_2858; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2860 = 12'haed == _T_46[11:0] ? image_2797 : _GEN_2859; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2861 = 12'haee == _T_46[11:0] ? image_2798 : _GEN_2860; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2862 = 12'haef == _T_46[11:0] ? image_2799 : _GEN_2861; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2863 = 12'haf0 == _T_46[11:0] ? image_2800 : _GEN_2862; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2864 = 12'haf1 == _T_46[11:0] ? image_2801 : _GEN_2863; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2865 = 12'haf2 == _T_46[11:0] ? image_2802 : _GEN_2864; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2866 = 12'haf3 == _T_46[11:0] ? image_2803 : _GEN_2865; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2867 = 12'haf4 == _T_46[11:0] ? image_2804 : _GEN_2866; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2868 = 12'haf5 == _T_46[11:0] ? image_2805 : _GEN_2867; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2869 = 12'haf6 == _T_46[11:0] ? image_2806 : _GEN_2868; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2870 = 12'haf7 == _T_46[11:0] ? image_2807 : _GEN_2869; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2871 = 12'haf8 == _T_46[11:0] ? image_2808 : _GEN_2870; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2872 = 12'haf9 == _T_46[11:0] ? 4'h0 : _GEN_2871; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2873 = 12'hafa == _T_46[11:0] ? 4'h0 : _GEN_2872; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2874 = 12'hafb == _T_46[11:0] ? 4'h0 : _GEN_2873; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2875 = 12'hafc == _T_46[11:0] ? 4'h0 : _GEN_2874; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2876 = 12'hafd == _T_46[11:0] ? 4'h0 : _GEN_2875; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2877 = 12'hafe == _T_46[11:0] ? 4'h0 : _GEN_2876; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2878 = 12'haff == _T_46[11:0] ? 4'h0 : _GEN_2877; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2879 = 12'hb00 == _T_46[11:0] ? 4'h0 : _GEN_2878; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2880 = 12'hb01 == _T_46[11:0] ? 4'h0 : _GEN_2879; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2881 = 12'hb02 == _T_46[11:0] ? 4'h0 : _GEN_2880; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2882 = 12'hb03 == _T_46[11:0] ? 4'h0 : _GEN_2881; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2883 = 12'hb04 == _T_46[11:0] ? 4'h0 : _GEN_2882; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2884 = 12'hb05 == _T_46[11:0] ? 4'h0 : _GEN_2883; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2885 = 12'hb06 == _T_46[11:0] ? 4'h0 : _GEN_2884; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2886 = 12'hb07 == _T_46[11:0] ? 4'h0 : _GEN_2885; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2887 = 12'hb08 == _T_46[11:0] ? 4'h0 : _GEN_2886; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2888 = 12'hb09 == _T_46[11:0] ? 4'h0 : _GEN_2887; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2889 = 12'hb0a == _T_46[11:0] ? 4'h0 : _GEN_2888; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2890 = 12'hb0b == _T_46[11:0] ? 4'h0 : _GEN_2889; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2891 = 12'hb0c == _T_46[11:0] ? image_2828 : _GEN_2890; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2892 = 12'hb0d == _T_46[11:0] ? image_2829 : _GEN_2891; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2893 = 12'hb0e == _T_46[11:0] ? image_2830 : _GEN_2892; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2894 = 12'hb0f == _T_46[11:0] ? image_2831 : _GEN_2893; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2895 = 12'hb10 == _T_46[11:0] ? image_2832 : _GEN_2894; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2896 = 12'hb11 == _T_46[11:0] ? image_2833 : _GEN_2895; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2897 = 12'hb12 == _T_46[11:0] ? image_2834 : _GEN_2896; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2898 = 12'hb13 == _T_46[11:0] ? image_2835 : _GEN_2897; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2899 = 12'hb14 == _T_46[11:0] ? image_2836 : _GEN_2898; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2900 = 12'hb15 == _T_46[11:0] ? image_2837 : _GEN_2899; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2901 = 12'hb16 == _T_46[11:0] ? image_2838 : _GEN_2900; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2902 = 12'hb17 == _T_46[11:0] ? image_2839 : _GEN_2901; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2903 = 12'hb18 == _T_46[11:0] ? image_2840 : _GEN_2902; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2904 = 12'hb19 == _T_46[11:0] ? image_2841 : _GEN_2903; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2905 = 12'hb1a == _T_46[11:0] ? image_2842 : _GEN_2904; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2906 = 12'hb1b == _T_46[11:0] ? image_2843 : _GEN_2905; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2907 = 12'hb1c == _T_46[11:0] ? image_2844 : _GEN_2906; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2908 = 12'hb1d == _T_46[11:0] ? image_2845 : _GEN_2907; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2909 = 12'hb1e == _T_46[11:0] ? image_2846 : _GEN_2908; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2910 = 12'hb1f == _T_46[11:0] ? image_2847 : _GEN_2909; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2911 = 12'hb20 == _T_46[11:0] ? image_2848 : _GEN_2910; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2912 = 12'hb21 == _T_46[11:0] ? image_2849 : _GEN_2911; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2913 = 12'hb22 == _T_46[11:0] ? image_2850 : _GEN_2912; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2914 = 12'hb23 == _T_46[11:0] ? image_2851 : _GEN_2913; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2915 = 12'hb24 == _T_46[11:0] ? image_2852 : _GEN_2914; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2916 = 12'hb25 == _T_46[11:0] ? image_2853 : _GEN_2915; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2917 = 12'hb26 == _T_46[11:0] ? image_2854 : _GEN_2916; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2918 = 12'hb27 == _T_46[11:0] ? image_2855 : _GEN_2917; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2919 = 12'hb28 == _T_46[11:0] ? image_2856 : _GEN_2918; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2920 = 12'hb29 == _T_46[11:0] ? image_2857 : _GEN_2919; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2921 = 12'hb2a == _T_46[11:0] ? image_2858 : _GEN_2920; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2922 = 12'hb2b == _T_46[11:0] ? image_2859 : _GEN_2921; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2923 = 12'hb2c == _T_46[11:0] ? image_2860 : _GEN_2922; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2924 = 12'hb2d == _T_46[11:0] ? image_2861 : _GEN_2923; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2925 = 12'hb2e == _T_46[11:0] ? image_2862 : _GEN_2924; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2926 = 12'hb2f == _T_46[11:0] ? image_2863 : _GEN_2925; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2927 = 12'hb30 == _T_46[11:0] ? image_2864 : _GEN_2926; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2928 = 12'hb31 == _T_46[11:0] ? image_2865 : _GEN_2927; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2929 = 12'hb32 == _T_46[11:0] ? image_2866 : _GEN_2928; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2930 = 12'hb33 == _T_46[11:0] ? image_2867 : _GEN_2929; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2931 = 12'hb34 == _T_46[11:0] ? image_2868 : _GEN_2930; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2932 = 12'hb35 == _T_46[11:0] ? image_2869 : _GEN_2931; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2933 = 12'hb36 == _T_46[11:0] ? image_2870 : _GEN_2932; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2934 = 12'hb37 == _T_46[11:0] ? image_2871 : _GEN_2933; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2935 = 12'hb38 == _T_46[11:0] ? 4'h0 : _GEN_2934; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2936 = 12'hb39 == _T_46[11:0] ? 4'h0 : _GEN_2935; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2937 = 12'hb3a == _T_46[11:0] ? 4'h0 : _GEN_2936; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2938 = 12'hb3b == _T_46[11:0] ? 4'h0 : _GEN_2937; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2939 = 12'hb3c == _T_46[11:0] ? 4'h0 : _GEN_2938; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2940 = 12'hb3d == _T_46[11:0] ? 4'h0 : _GEN_2939; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2941 = 12'hb3e == _T_46[11:0] ? 4'h0 : _GEN_2940; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2942 = 12'hb3f == _T_46[11:0] ? 4'h0 : _GEN_2941; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2943 = 12'hb40 == _T_46[11:0] ? 4'h0 : _GEN_2942; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2944 = 12'hb41 == _T_46[11:0] ? 4'h0 : _GEN_2943; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2945 = 12'hb42 == _T_46[11:0] ? 4'h0 : _GEN_2944; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2946 = 12'hb43 == _T_46[11:0] ? 4'h0 : _GEN_2945; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2947 = 12'hb44 == _T_46[11:0] ? 4'h0 : _GEN_2946; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2948 = 12'hb45 == _T_46[11:0] ? 4'h0 : _GEN_2947; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2949 = 12'hb46 == _T_46[11:0] ? 4'h0 : _GEN_2948; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2950 = 12'hb47 == _T_46[11:0] ? 4'h0 : _GEN_2949; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2951 = 12'hb48 == _T_46[11:0] ? 4'h0 : _GEN_2950; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2952 = 12'hb49 == _T_46[11:0] ? 4'h0 : _GEN_2951; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2953 = 12'hb4a == _T_46[11:0] ? 4'h0 : _GEN_2952; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2954 = 12'hb4b == _T_46[11:0] ? 4'h0 : _GEN_2953; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2955 = 12'hb4c == _T_46[11:0] ? 4'h0 : _GEN_2954; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2956 = 12'hb4d == _T_46[11:0] ? 4'h0 : _GEN_2955; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2957 = 12'hb4e == _T_46[11:0] ? 4'h0 : _GEN_2956; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2958 = 12'hb4f == _T_46[11:0] ? image_2895 : _GEN_2957; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2959 = 12'hb50 == _T_46[11:0] ? image_2896 : _GEN_2958; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2960 = 12'hb51 == _T_46[11:0] ? image_2897 : _GEN_2959; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2961 = 12'hb52 == _T_46[11:0] ? image_2898 : _GEN_2960; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2962 = 12'hb53 == _T_46[11:0] ? image_2899 : _GEN_2961; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2963 = 12'hb54 == _T_46[11:0] ? image_2900 : _GEN_2962; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2964 = 12'hb55 == _T_46[11:0] ? image_2901 : _GEN_2963; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2965 = 12'hb56 == _T_46[11:0] ? image_2902 : _GEN_2964; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2966 = 12'hb57 == _T_46[11:0] ? image_2903 : _GEN_2965; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2967 = 12'hb58 == _T_46[11:0] ? image_2904 : _GEN_2966; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2968 = 12'hb59 == _T_46[11:0] ? image_2905 : _GEN_2967; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2969 = 12'hb5a == _T_46[11:0] ? image_2906 : _GEN_2968; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2970 = 12'hb5b == _T_46[11:0] ? image_2907 : _GEN_2969; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2971 = 12'hb5c == _T_46[11:0] ? image_2908 : _GEN_2970; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2972 = 12'hb5d == _T_46[11:0] ? image_2909 : _GEN_2971; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2973 = 12'hb5e == _T_46[11:0] ? image_2910 : _GEN_2972; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2974 = 12'hb5f == _T_46[11:0] ? image_2911 : _GEN_2973; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2975 = 12'hb60 == _T_46[11:0] ? image_2912 : _GEN_2974; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2976 = 12'hb61 == _T_46[11:0] ? image_2913 : _GEN_2975; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2977 = 12'hb62 == _T_46[11:0] ? image_2914 : _GEN_2976; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2978 = 12'hb63 == _T_46[11:0] ? image_2915 : _GEN_2977; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2979 = 12'hb64 == _T_46[11:0] ? image_2916 : _GEN_2978; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2980 = 12'hb65 == _T_46[11:0] ? image_2917 : _GEN_2979; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2981 = 12'hb66 == _T_46[11:0] ? image_2918 : _GEN_2980; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2982 = 12'hb67 == _T_46[11:0] ? image_2919 : _GEN_2981; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2983 = 12'hb68 == _T_46[11:0] ? image_2920 : _GEN_2982; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2984 = 12'hb69 == _T_46[11:0] ? image_2921 : _GEN_2983; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2985 = 12'hb6a == _T_46[11:0] ? image_2922 : _GEN_2984; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2986 = 12'hb6b == _T_46[11:0] ? image_2923 : _GEN_2985; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2987 = 12'hb6c == _T_46[11:0] ? image_2924 : _GEN_2986; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2988 = 12'hb6d == _T_46[11:0] ? image_2925 : _GEN_2987; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2989 = 12'hb6e == _T_46[11:0] ? image_2926 : _GEN_2988; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2990 = 12'hb6f == _T_46[11:0] ? image_2927 : _GEN_2989; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2991 = 12'hb70 == _T_46[11:0] ? image_2928 : _GEN_2990; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2992 = 12'hb71 == _T_46[11:0] ? image_2929 : _GEN_2991; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2993 = 12'hb72 == _T_46[11:0] ? image_2930 : _GEN_2992; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2994 = 12'hb73 == _T_46[11:0] ? image_2931 : _GEN_2993; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2995 = 12'hb74 == _T_46[11:0] ? image_2932 : _GEN_2994; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2996 = 12'hb75 == _T_46[11:0] ? image_2933 : _GEN_2995; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2997 = 12'hb76 == _T_46[11:0] ? image_2934 : _GEN_2996; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2998 = 12'hb77 == _T_46[11:0] ? 4'h0 : _GEN_2997; // @[Filter.scala 138:46]
  wire [3:0] _GEN_2999 = 12'hb78 == _T_46[11:0] ? 4'h0 : _GEN_2998; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3000 = 12'hb79 == _T_46[11:0] ? 4'h0 : _GEN_2999; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3001 = 12'hb7a == _T_46[11:0] ? 4'h0 : _GEN_3000; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3002 = 12'hb7b == _T_46[11:0] ? 4'h0 : _GEN_3001; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3003 = 12'hb7c == _T_46[11:0] ? 4'h0 : _GEN_3002; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3004 = 12'hb7d == _T_46[11:0] ? 4'h0 : _GEN_3003; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3005 = 12'hb7e == _T_46[11:0] ? 4'h0 : _GEN_3004; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3006 = 12'hb7f == _T_46[11:0] ? 4'h0 : _GEN_3005; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3007 = 12'hb80 == _T_46[11:0] ? 4'h0 : _GEN_3006; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3008 = 12'hb81 == _T_46[11:0] ? 4'h0 : _GEN_3007; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3009 = 12'hb82 == _T_46[11:0] ? 4'h0 : _GEN_3008; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3010 = 12'hb83 == _T_46[11:0] ? 4'h0 : _GEN_3009; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3011 = 12'hb84 == _T_46[11:0] ? 4'h0 : _GEN_3010; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3012 = 12'hb85 == _T_46[11:0] ? 4'h0 : _GEN_3011; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3013 = 12'hb86 == _T_46[11:0] ? 4'h0 : _GEN_3012; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3014 = 12'hb87 == _T_46[11:0] ? 4'h0 : _GEN_3013; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3015 = 12'hb88 == _T_46[11:0] ? 4'h0 : _GEN_3014; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3016 = 12'hb89 == _T_46[11:0] ? 4'h0 : _GEN_3015; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3017 = 12'hb8a == _T_46[11:0] ? 4'h0 : _GEN_3016; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3018 = 12'hb8b == _T_46[11:0] ? 4'h0 : _GEN_3017; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3019 = 12'hb8c == _T_46[11:0] ? 4'h0 : _GEN_3018; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3020 = 12'hb8d == _T_46[11:0] ? 4'h0 : _GEN_3019; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3021 = 12'hb8e == _T_46[11:0] ? 4'h0 : _GEN_3020; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3022 = 12'hb8f == _T_46[11:0] ? 4'h0 : _GEN_3021; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3023 = 12'hb90 == _T_46[11:0] ? 4'h0 : _GEN_3022; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3024 = 12'hb91 == _T_46[11:0] ? 4'h0 : _GEN_3023; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3025 = 12'hb92 == _T_46[11:0] ? 4'h0 : _GEN_3024; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3026 = 12'hb93 == _T_46[11:0] ? 4'h0 : _GEN_3025; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3027 = 12'hb94 == _T_46[11:0] ? 4'h0 : _GEN_3026; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3028 = 12'hb95 == _T_46[11:0] ? image_2965 : _GEN_3027; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3029 = 12'hb96 == _T_46[11:0] ? image_2966 : _GEN_3028; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3030 = 12'hb97 == _T_46[11:0] ? image_2967 : _GEN_3029; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3031 = 12'hb98 == _T_46[11:0] ? image_2968 : _GEN_3030; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3032 = 12'hb99 == _T_46[11:0] ? image_2969 : _GEN_3031; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3033 = 12'hb9a == _T_46[11:0] ? image_2970 : _GEN_3032; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3034 = 12'hb9b == _T_46[11:0] ? image_2971 : _GEN_3033; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3035 = 12'hb9c == _T_46[11:0] ? image_2972 : _GEN_3034; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3036 = 12'hb9d == _T_46[11:0] ? image_2973 : _GEN_3035; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3037 = 12'hb9e == _T_46[11:0] ? image_2974 : _GEN_3036; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3038 = 12'hb9f == _T_46[11:0] ? image_2975 : _GEN_3037; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3039 = 12'hba0 == _T_46[11:0] ? image_2976 : _GEN_3038; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3040 = 12'hba1 == _T_46[11:0] ? image_2977 : _GEN_3039; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3041 = 12'hba2 == _T_46[11:0] ? image_2978 : _GEN_3040; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3042 = 12'hba3 == _T_46[11:0] ? image_2979 : _GEN_3041; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3043 = 12'hba4 == _T_46[11:0] ? image_2980 : _GEN_3042; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3044 = 12'hba5 == _T_46[11:0] ? image_2981 : _GEN_3043; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3045 = 12'hba6 == _T_46[11:0] ? image_2982 : _GEN_3044; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3046 = 12'hba7 == _T_46[11:0] ? image_2983 : _GEN_3045; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3047 = 12'hba8 == _T_46[11:0] ? image_2984 : _GEN_3046; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3048 = 12'hba9 == _T_46[11:0] ? image_2985 : _GEN_3047; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3049 = 12'hbaa == _T_46[11:0] ? image_2986 : _GEN_3048; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3050 = 12'hbab == _T_46[11:0] ? image_2987 : _GEN_3049; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3051 = 12'hbac == _T_46[11:0] ? image_2988 : _GEN_3050; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3052 = 12'hbad == _T_46[11:0] ? image_2989 : _GEN_3051; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3053 = 12'hbae == _T_46[11:0] ? image_2990 : _GEN_3052; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3054 = 12'hbaf == _T_46[11:0] ? image_2991 : _GEN_3053; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3055 = 12'hbb0 == _T_46[11:0] ? image_2992 : _GEN_3054; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3056 = 12'hbb1 == _T_46[11:0] ? image_2993 : _GEN_3055; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3057 = 12'hbb2 == _T_46[11:0] ? image_2994 : _GEN_3056; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3058 = 12'hbb3 == _T_46[11:0] ? image_2995 : _GEN_3057; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3059 = 12'hbb4 == _T_46[11:0] ? image_2996 : _GEN_3058; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3060 = 12'hbb5 == _T_46[11:0] ? 4'h0 : _GEN_3059; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3061 = 12'hbb6 == _T_46[11:0] ? 4'h0 : _GEN_3060; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3062 = 12'hbb7 == _T_46[11:0] ? 4'h0 : _GEN_3061; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3063 = 12'hbb8 == _T_46[11:0] ? 4'h0 : _GEN_3062; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3064 = 12'hbb9 == _T_46[11:0] ? 4'h0 : _GEN_3063; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3065 = 12'hbba == _T_46[11:0] ? 4'h0 : _GEN_3064; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3066 = 12'hbbb == _T_46[11:0] ? 4'h0 : _GEN_3065; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3067 = 12'hbbc == _T_46[11:0] ? 4'h0 : _GEN_3066; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3068 = 12'hbbd == _T_46[11:0] ? 4'h0 : _GEN_3067; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3069 = 12'hbbe == _T_46[11:0] ? 4'h0 : _GEN_3068; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3070 = 12'hbbf == _T_46[11:0] ? 4'h0 : _GEN_3069; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3071 = 12'hbc0 == _T_46[11:0] ? 4'h0 : _GEN_3070; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3072 = 12'hbc1 == _T_46[11:0] ? 4'h0 : _GEN_3071; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3073 = 12'hbc2 == _T_46[11:0] ? 4'h0 : _GEN_3072; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3074 = 12'hbc3 == _T_46[11:0] ? 4'h0 : _GEN_3073; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3075 = 12'hbc4 == _T_46[11:0] ? 4'h0 : _GEN_3074; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3076 = 12'hbc5 == _T_46[11:0] ? 4'h0 : _GEN_3075; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3077 = 12'hbc6 == _T_46[11:0] ? 4'h0 : _GEN_3076; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3078 = 12'hbc7 == _T_46[11:0] ? 4'h0 : _GEN_3077; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3079 = 12'hbc8 == _T_46[11:0] ? 4'h0 : _GEN_3078; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3080 = 12'hbc9 == _T_46[11:0] ? 4'h0 : _GEN_3079; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3081 = 12'hbca == _T_46[11:0] ? 4'h0 : _GEN_3080; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3082 = 12'hbcb == _T_46[11:0] ? 4'h0 : _GEN_3081; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3083 = 12'hbcc == _T_46[11:0] ? 4'h0 : _GEN_3082; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3084 = 12'hbcd == _T_46[11:0] ? 4'h0 : _GEN_3083; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3085 = 12'hbce == _T_46[11:0] ? 4'h0 : _GEN_3084; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3086 = 12'hbcf == _T_46[11:0] ? 4'h0 : _GEN_3085; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3087 = 12'hbd0 == _T_46[11:0] ? 4'h0 : _GEN_3086; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3088 = 12'hbd1 == _T_46[11:0] ? 4'h0 : _GEN_3087; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3089 = 12'hbd2 == _T_46[11:0] ? 4'h0 : _GEN_3088; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3090 = 12'hbd3 == _T_46[11:0] ? 4'h0 : _GEN_3089; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3091 = 12'hbd4 == _T_46[11:0] ? 4'h0 : _GEN_3090; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3092 = 12'hbd5 == _T_46[11:0] ? 4'h0 : _GEN_3091; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3093 = 12'hbd6 == _T_46[11:0] ? 4'h0 : _GEN_3092; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3094 = 12'hbd7 == _T_46[11:0] ? 4'h0 : _GEN_3093; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3095 = 12'hbd8 == _T_46[11:0] ? 4'h0 : _GEN_3094; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3096 = 12'hbd9 == _T_46[11:0] ? 4'h0 : _GEN_3095; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3097 = 12'hbda == _T_46[11:0] ? 4'h0 : _GEN_3096; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3098 = 12'hbdb == _T_46[11:0] ? image_3035 : _GEN_3097; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3099 = 12'hbdc == _T_46[11:0] ? image_3036 : _GEN_3098; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3100 = 12'hbdd == _T_46[11:0] ? image_3037 : _GEN_3099; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3101 = 12'hbde == _T_46[11:0] ? image_3038 : _GEN_3100; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3102 = 12'hbdf == _T_46[11:0] ? image_3039 : _GEN_3101; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3103 = 12'hbe0 == _T_46[11:0] ? image_3040 : _GEN_3102; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3104 = 12'hbe1 == _T_46[11:0] ? image_3041 : _GEN_3103; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3105 = 12'hbe2 == _T_46[11:0] ? image_3042 : _GEN_3104; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3106 = 12'hbe3 == _T_46[11:0] ? image_3043 : _GEN_3105; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3107 = 12'hbe4 == _T_46[11:0] ? image_3044 : _GEN_3106; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3108 = 12'hbe5 == _T_46[11:0] ? image_3045 : _GEN_3107; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3109 = 12'hbe6 == _T_46[11:0] ? image_3046 : _GEN_3108; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3110 = 12'hbe7 == _T_46[11:0] ? image_3047 : _GEN_3109; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3111 = 12'hbe8 == _T_46[11:0] ? image_3048 : _GEN_3110; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3112 = 12'hbe9 == _T_46[11:0] ? image_3049 : _GEN_3111; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3113 = 12'hbea == _T_46[11:0] ? image_3050 : _GEN_3112; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3114 = 12'hbeb == _T_46[11:0] ? image_3051 : _GEN_3113; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3115 = 12'hbec == _T_46[11:0] ? image_3052 : _GEN_3114; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3116 = 12'hbed == _T_46[11:0] ? image_3053 : _GEN_3115; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3117 = 12'hbee == _T_46[11:0] ? image_3054 : _GEN_3116; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3118 = 12'hbef == _T_46[11:0] ? image_3055 : _GEN_3117; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3119 = 12'hbf0 == _T_46[11:0] ? image_3056 : _GEN_3118; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3120 = 12'hbf1 == _T_46[11:0] ? 4'h0 : _GEN_3119; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3121 = 12'hbf2 == _T_46[11:0] ? 4'h0 : _GEN_3120; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3122 = 12'hbf3 == _T_46[11:0] ? 4'h0 : _GEN_3121; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3123 = 12'hbf4 == _T_46[11:0] ? 4'h0 : _GEN_3122; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3124 = 12'hbf5 == _T_46[11:0] ? 4'h0 : _GEN_3123; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3125 = 12'hbf6 == _T_46[11:0] ? 4'h0 : _GEN_3124; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3126 = 12'hbf7 == _T_46[11:0] ? 4'h0 : _GEN_3125; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3127 = 12'hbf8 == _T_46[11:0] ? 4'h0 : _GEN_3126; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3128 = 12'hbf9 == _T_46[11:0] ? 4'h0 : _GEN_3127; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3129 = 12'hbfa == _T_46[11:0] ? 4'h0 : _GEN_3128; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3130 = 12'hbfb == _T_46[11:0] ? 4'h0 : _GEN_3129; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3131 = 12'hbfc == _T_46[11:0] ? 4'h0 : _GEN_3130; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3132 = 12'hbfd == _T_46[11:0] ? 4'h0 : _GEN_3131; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3133 = 12'hbfe == _T_46[11:0] ? 4'h0 : _GEN_3132; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3134 = 12'hbff == _T_46[11:0] ? 4'h0 : _GEN_3133; // @[Filter.scala 138:46]
  wire [31:0] _T_49 = pixelIndex + 32'h1; // @[Filter.scala 133:29]
  wire [31:0] _T_50 = _T_49 / 32'h40; // @[Filter.scala 133:36]
  wire [31:0] _T_52 = _T_50 + _GEN_24805; // @[Filter.scala 133:51]
  wire [31:0] _T_54 = _T_52 - 32'h1; // @[Filter.scala 133:67]
  wire [31:0] _GEN_1 = _T_49 % 32'h40; // @[Filter.scala 134:36]
  wire [6:0] _T_57 = _GEN_1[6:0]; // @[Filter.scala 134:36]
  wire [6:0] _T_59 = _T_57 + _GEN_24806; // @[Filter.scala 134:51]
  wire [6:0] _T_61 = _T_59 - 7'h1; // @[Filter.scala 134:67]
  wire  _T_63 = _T_54 >= 32'h40; // @[Filter.scala 135:27]
  wire  _T_67 = _T_61 >= 7'h30; // @[Filter.scala 135:59]
  wire  _T_68 = _T_63 | _T_67; // @[Filter.scala 135:54]
  wire [13:0] _T_69 = _T_61 * 7'h40; // @[Filter.scala 138:57]
  wire [31:0] _GEN_24810 = {{18'd0}, _T_69}; // @[Filter.scala 138:72]
  wire [31:0] _T_71 = _GEN_24810 + _T_54; // @[Filter.scala 138:72]
  wire [3:0] _GEN_3148 = 12'hc == _T_71[11:0] ? image_12 : 4'h0; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3149 = 12'hd == _T_71[11:0] ? 4'h0 : _GEN_3148; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3150 = 12'he == _T_71[11:0] ? image_14 : _GEN_3149; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3151 = 12'hf == _T_71[11:0] ? image_15 : _GEN_3150; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3152 = 12'h10 == _T_71[11:0] ? image_16 : _GEN_3151; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3153 = 12'h11 == _T_71[11:0] ? image_17 : _GEN_3152; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3154 = 12'h12 == _T_71[11:0] ? image_18 : _GEN_3153; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3155 = 12'h13 == _T_71[11:0] ? image_19 : _GEN_3154; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3156 = 12'h14 == _T_71[11:0] ? image_20 : _GEN_3155; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3157 = 12'h15 == _T_71[11:0] ? image_21 : _GEN_3156; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3158 = 12'h16 == _T_71[11:0] ? image_22 : _GEN_3157; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3159 = 12'h17 == _T_71[11:0] ? image_23 : _GEN_3158; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3160 = 12'h18 == _T_71[11:0] ? 4'h0 : _GEN_3159; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3161 = 12'h19 == _T_71[11:0] ? 4'h0 : _GEN_3160; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3162 = 12'h1a == _T_71[11:0] ? 4'h0 : _GEN_3161; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3163 = 12'h1b == _T_71[11:0] ? 4'h0 : _GEN_3162; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3164 = 12'h1c == _T_71[11:0] ? 4'h0 : _GEN_3163; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3165 = 12'h1d == _T_71[11:0] ? 4'h0 : _GEN_3164; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3166 = 12'h1e == _T_71[11:0] ? 4'h0 : _GEN_3165; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3167 = 12'h1f == _T_71[11:0] ? 4'h0 : _GEN_3166; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3168 = 12'h20 == _T_71[11:0] ? 4'h0 : _GEN_3167; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3169 = 12'h21 == _T_71[11:0] ? 4'h0 : _GEN_3168; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3170 = 12'h22 == _T_71[11:0] ? 4'h0 : _GEN_3169; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3171 = 12'h23 == _T_71[11:0] ? image_35 : _GEN_3170; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3172 = 12'h24 == _T_71[11:0] ? image_36 : _GEN_3171; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3173 = 12'h25 == _T_71[11:0] ? image_37 : _GEN_3172; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3174 = 12'h26 == _T_71[11:0] ? image_38 : _GEN_3173; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3175 = 12'h27 == _T_71[11:0] ? image_39 : _GEN_3174; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3176 = 12'h28 == _T_71[11:0] ? image_40 : _GEN_3175; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3177 = 12'h29 == _T_71[11:0] ? image_41 : _GEN_3176; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3178 = 12'h2a == _T_71[11:0] ? image_42 : _GEN_3177; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3179 = 12'h2b == _T_71[11:0] ? 4'h0 : _GEN_3178; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3180 = 12'h2c == _T_71[11:0] ? 4'h0 : _GEN_3179; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3181 = 12'h2d == _T_71[11:0] ? 4'h0 : _GEN_3180; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3182 = 12'h2e == _T_71[11:0] ? 4'h0 : _GEN_3181; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3183 = 12'h2f == _T_71[11:0] ? 4'h0 : _GEN_3182; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3184 = 12'h30 == _T_71[11:0] ? 4'h0 : _GEN_3183; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3185 = 12'h31 == _T_71[11:0] ? 4'h0 : _GEN_3184; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3186 = 12'h32 == _T_71[11:0] ? 4'h0 : _GEN_3185; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3187 = 12'h33 == _T_71[11:0] ? 4'h0 : _GEN_3186; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3188 = 12'h34 == _T_71[11:0] ? 4'h0 : _GEN_3187; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3189 = 12'h35 == _T_71[11:0] ? 4'h0 : _GEN_3188; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3190 = 12'h36 == _T_71[11:0] ? 4'h0 : _GEN_3189; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3191 = 12'h37 == _T_71[11:0] ? 4'h0 : _GEN_3190; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3192 = 12'h38 == _T_71[11:0] ? 4'h0 : _GEN_3191; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3193 = 12'h39 == _T_71[11:0] ? 4'h0 : _GEN_3192; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3194 = 12'h3a == _T_71[11:0] ? 4'h0 : _GEN_3193; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3195 = 12'h3b == _T_71[11:0] ? 4'h0 : _GEN_3194; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3196 = 12'h3c == _T_71[11:0] ? 4'h0 : _GEN_3195; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3197 = 12'h3d == _T_71[11:0] ? 4'h0 : _GEN_3196; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3198 = 12'h3e == _T_71[11:0] ? 4'h0 : _GEN_3197; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3199 = 12'h3f == _T_71[11:0] ? 4'h0 : _GEN_3198; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3200 = 12'h40 == _T_71[11:0] ? 4'h0 : _GEN_3199; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3201 = 12'h41 == _T_71[11:0] ? 4'h0 : _GEN_3200; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3202 = 12'h42 == _T_71[11:0] ? 4'h0 : _GEN_3201; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3203 = 12'h43 == _T_71[11:0] ? 4'h0 : _GEN_3202; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3204 = 12'h44 == _T_71[11:0] ? 4'h0 : _GEN_3203; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3205 = 12'h45 == _T_71[11:0] ? 4'h0 : _GEN_3204; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3206 = 12'h46 == _T_71[11:0] ? 4'h0 : _GEN_3205; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3207 = 12'h47 == _T_71[11:0] ? 4'h0 : _GEN_3206; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3208 = 12'h48 == _T_71[11:0] ? 4'h0 : _GEN_3207; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3209 = 12'h49 == _T_71[11:0] ? 4'h0 : _GEN_3208; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3210 = 12'h4a == _T_71[11:0] ? 4'h0 : _GEN_3209; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3211 = 12'h4b == _T_71[11:0] ? image_75 : _GEN_3210; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3212 = 12'h4c == _T_71[11:0] ? image_76 : _GEN_3211; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3213 = 12'h4d == _T_71[11:0] ? image_77 : _GEN_3212; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3214 = 12'h4e == _T_71[11:0] ? image_78 : _GEN_3213; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3215 = 12'h4f == _T_71[11:0] ? image_79 : _GEN_3214; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3216 = 12'h50 == _T_71[11:0] ? image_80 : _GEN_3215; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3217 = 12'h51 == _T_71[11:0] ? image_81 : _GEN_3216; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3218 = 12'h52 == _T_71[11:0] ? image_82 : _GEN_3217; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3219 = 12'h53 == _T_71[11:0] ? image_83 : _GEN_3218; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3220 = 12'h54 == _T_71[11:0] ? image_84 : _GEN_3219; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3221 = 12'h55 == _T_71[11:0] ? image_85 : _GEN_3220; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3222 = 12'h56 == _T_71[11:0] ? image_86 : _GEN_3221; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3223 = 12'h57 == _T_71[11:0] ? image_87 : _GEN_3222; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3224 = 12'h58 == _T_71[11:0] ? image_88 : _GEN_3223; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3225 = 12'h59 == _T_71[11:0] ? image_89 : _GEN_3224; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3226 = 12'h5a == _T_71[11:0] ? image_90 : _GEN_3225; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3227 = 12'h5b == _T_71[11:0] ? 4'h0 : _GEN_3226; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3228 = 12'h5c == _T_71[11:0] ? 4'h0 : _GEN_3227; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3229 = 12'h5d == _T_71[11:0] ? image_93 : _GEN_3228; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3230 = 12'h5e == _T_71[11:0] ? 4'h0 : _GEN_3229; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3231 = 12'h5f == _T_71[11:0] ? image_95 : _GEN_3230; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3232 = 12'h60 == _T_71[11:0] ? image_96 : _GEN_3231; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3233 = 12'h61 == _T_71[11:0] ? image_97 : _GEN_3232; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3234 = 12'h62 == _T_71[11:0] ? image_98 : _GEN_3233; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3235 = 12'h63 == _T_71[11:0] ? image_99 : _GEN_3234; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3236 = 12'h64 == _T_71[11:0] ? image_100 : _GEN_3235; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3237 = 12'h65 == _T_71[11:0] ? image_101 : _GEN_3236; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3238 = 12'h66 == _T_71[11:0] ? image_102 : _GEN_3237; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3239 = 12'h67 == _T_71[11:0] ? image_103 : _GEN_3238; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3240 = 12'h68 == _T_71[11:0] ? image_104 : _GEN_3239; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3241 = 12'h69 == _T_71[11:0] ? image_105 : _GEN_3240; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3242 = 12'h6a == _T_71[11:0] ? image_106 : _GEN_3241; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3243 = 12'h6b == _T_71[11:0] ? image_107 : _GEN_3242; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3244 = 12'h6c == _T_71[11:0] ? image_108 : _GEN_3243; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3245 = 12'h6d == _T_71[11:0] ? 4'h0 : _GEN_3244; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3246 = 12'h6e == _T_71[11:0] ? 4'h0 : _GEN_3245; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3247 = 12'h6f == _T_71[11:0] ? 4'h0 : _GEN_3246; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3248 = 12'h70 == _T_71[11:0] ? 4'h0 : _GEN_3247; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3249 = 12'h71 == _T_71[11:0] ? 4'h0 : _GEN_3248; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3250 = 12'h72 == _T_71[11:0] ? 4'h0 : _GEN_3249; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3251 = 12'h73 == _T_71[11:0] ? 4'h0 : _GEN_3250; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3252 = 12'h74 == _T_71[11:0] ? 4'h0 : _GEN_3251; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3253 = 12'h75 == _T_71[11:0] ? 4'h0 : _GEN_3252; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3254 = 12'h76 == _T_71[11:0] ? 4'h0 : _GEN_3253; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3255 = 12'h77 == _T_71[11:0] ? 4'h0 : _GEN_3254; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3256 = 12'h78 == _T_71[11:0] ? 4'h0 : _GEN_3255; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3257 = 12'h79 == _T_71[11:0] ? 4'h0 : _GEN_3256; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3258 = 12'h7a == _T_71[11:0] ? 4'h0 : _GEN_3257; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3259 = 12'h7b == _T_71[11:0] ? 4'h0 : _GEN_3258; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3260 = 12'h7c == _T_71[11:0] ? 4'h0 : _GEN_3259; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3261 = 12'h7d == _T_71[11:0] ? 4'h0 : _GEN_3260; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3262 = 12'h7e == _T_71[11:0] ? 4'h0 : _GEN_3261; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3263 = 12'h7f == _T_71[11:0] ? 4'h0 : _GEN_3262; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3264 = 12'h80 == _T_71[11:0] ? 4'h0 : _GEN_3263; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3265 = 12'h81 == _T_71[11:0] ? 4'h0 : _GEN_3264; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3266 = 12'h82 == _T_71[11:0] ? 4'h0 : _GEN_3265; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3267 = 12'h83 == _T_71[11:0] ? 4'h0 : _GEN_3266; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3268 = 12'h84 == _T_71[11:0] ? 4'h0 : _GEN_3267; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3269 = 12'h85 == _T_71[11:0] ? 4'h0 : _GEN_3268; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3270 = 12'h86 == _T_71[11:0] ? 4'h0 : _GEN_3269; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3271 = 12'h87 == _T_71[11:0] ? 4'h0 : _GEN_3270; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3272 = 12'h88 == _T_71[11:0] ? image_136 : _GEN_3271; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3273 = 12'h89 == _T_71[11:0] ? image_137 : _GEN_3272; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3274 = 12'h8a == _T_71[11:0] ? image_138 : _GEN_3273; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3275 = 12'h8b == _T_71[11:0] ? image_139 : _GEN_3274; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3276 = 12'h8c == _T_71[11:0] ? image_140 : _GEN_3275; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3277 = 12'h8d == _T_71[11:0] ? image_141 : _GEN_3276; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3278 = 12'h8e == _T_71[11:0] ? image_142 : _GEN_3277; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3279 = 12'h8f == _T_71[11:0] ? image_143 : _GEN_3278; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3280 = 12'h90 == _T_71[11:0] ? image_144 : _GEN_3279; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3281 = 12'h91 == _T_71[11:0] ? image_145 : _GEN_3280; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3282 = 12'h92 == _T_71[11:0] ? image_146 : _GEN_3281; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3283 = 12'h93 == _T_71[11:0] ? image_147 : _GEN_3282; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3284 = 12'h94 == _T_71[11:0] ? image_148 : _GEN_3283; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3285 = 12'h95 == _T_71[11:0] ? image_149 : _GEN_3284; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3286 = 12'h96 == _T_71[11:0] ? image_150 : _GEN_3285; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3287 = 12'h97 == _T_71[11:0] ? image_151 : _GEN_3286; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3288 = 12'h98 == _T_71[11:0] ? image_152 : _GEN_3287; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3289 = 12'h99 == _T_71[11:0] ? image_153 : _GEN_3288; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3290 = 12'h9a == _T_71[11:0] ? image_154 : _GEN_3289; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3291 = 12'h9b == _T_71[11:0] ? image_155 : _GEN_3290; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3292 = 12'h9c == _T_71[11:0] ? 4'h0 : _GEN_3291; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3293 = 12'h9d == _T_71[11:0] ? image_157 : _GEN_3292; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3294 = 12'h9e == _T_71[11:0] ? image_158 : _GEN_3293; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3295 = 12'h9f == _T_71[11:0] ? image_159 : _GEN_3294; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3296 = 12'ha0 == _T_71[11:0] ? image_160 : _GEN_3295; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3297 = 12'ha1 == _T_71[11:0] ? image_161 : _GEN_3296; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3298 = 12'ha2 == _T_71[11:0] ? image_162 : _GEN_3297; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3299 = 12'ha3 == _T_71[11:0] ? image_163 : _GEN_3298; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3300 = 12'ha4 == _T_71[11:0] ? image_164 : _GEN_3299; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3301 = 12'ha5 == _T_71[11:0] ? image_165 : _GEN_3300; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3302 = 12'ha6 == _T_71[11:0] ? image_166 : _GEN_3301; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3303 = 12'ha7 == _T_71[11:0] ? image_167 : _GEN_3302; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3304 = 12'ha8 == _T_71[11:0] ? image_168 : _GEN_3303; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3305 = 12'ha9 == _T_71[11:0] ? image_169 : _GEN_3304; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3306 = 12'haa == _T_71[11:0] ? image_170 : _GEN_3305; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3307 = 12'hab == _T_71[11:0] ? image_171 : _GEN_3306; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3308 = 12'hac == _T_71[11:0] ? image_172 : _GEN_3307; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3309 = 12'had == _T_71[11:0] ? image_173 : _GEN_3308; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3310 = 12'hae == _T_71[11:0] ? image_174 : _GEN_3309; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3311 = 12'haf == _T_71[11:0] ? image_175 : _GEN_3310; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3312 = 12'hb0 == _T_71[11:0] ? image_176 : _GEN_3311; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3313 = 12'hb1 == _T_71[11:0] ? image_177 : _GEN_3312; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3314 = 12'hb2 == _T_71[11:0] ? image_178 : _GEN_3313; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3315 = 12'hb3 == _T_71[11:0] ? image_179 : _GEN_3314; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3316 = 12'hb4 == _T_71[11:0] ? 4'h0 : _GEN_3315; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3317 = 12'hb5 == _T_71[11:0] ? 4'h0 : _GEN_3316; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3318 = 12'hb6 == _T_71[11:0] ? 4'h0 : _GEN_3317; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3319 = 12'hb7 == _T_71[11:0] ? 4'h0 : _GEN_3318; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3320 = 12'hb8 == _T_71[11:0] ? 4'h0 : _GEN_3319; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3321 = 12'hb9 == _T_71[11:0] ? 4'h0 : _GEN_3320; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3322 = 12'hba == _T_71[11:0] ? 4'h0 : _GEN_3321; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3323 = 12'hbb == _T_71[11:0] ? 4'h0 : _GEN_3322; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3324 = 12'hbc == _T_71[11:0] ? 4'h0 : _GEN_3323; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3325 = 12'hbd == _T_71[11:0] ? 4'h0 : _GEN_3324; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3326 = 12'hbe == _T_71[11:0] ? 4'h0 : _GEN_3325; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3327 = 12'hbf == _T_71[11:0] ? 4'h0 : _GEN_3326; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3328 = 12'hc0 == _T_71[11:0] ? 4'h0 : _GEN_3327; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3329 = 12'hc1 == _T_71[11:0] ? 4'h0 : _GEN_3328; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3330 = 12'hc2 == _T_71[11:0] ? 4'h0 : _GEN_3329; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3331 = 12'hc3 == _T_71[11:0] ? 4'h0 : _GEN_3330; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3332 = 12'hc4 == _T_71[11:0] ? 4'h0 : _GEN_3331; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3333 = 12'hc5 == _T_71[11:0] ? 4'h0 : _GEN_3332; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3334 = 12'hc6 == _T_71[11:0] ? 4'h0 : _GEN_3333; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3335 = 12'hc7 == _T_71[11:0] ? image_199 : _GEN_3334; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3336 = 12'hc8 == _T_71[11:0] ? image_200 : _GEN_3335; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3337 = 12'hc9 == _T_71[11:0] ? image_201 : _GEN_3336; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3338 = 12'hca == _T_71[11:0] ? image_202 : _GEN_3337; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3339 = 12'hcb == _T_71[11:0] ? image_203 : _GEN_3338; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3340 = 12'hcc == _T_71[11:0] ? image_204 : _GEN_3339; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3341 = 12'hcd == _T_71[11:0] ? image_205 : _GEN_3340; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3342 = 12'hce == _T_71[11:0] ? image_206 : _GEN_3341; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3343 = 12'hcf == _T_71[11:0] ? image_207 : _GEN_3342; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3344 = 12'hd0 == _T_71[11:0] ? image_208 : _GEN_3343; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3345 = 12'hd1 == _T_71[11:0] ? image_209 : _GEN_3344; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3346 = 12'hd2 == _T_71[11:0] ? image_210 : _GEN_3345; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3347 = 12'hd3 == _T_71[11:0] ? image_211 : _GEN_3346; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3348 = 12'hd4 == _T_71[11:0] ? image_212 : _GEN_3347; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3349 = 12'hd5 == _T_71[11:0] ? image_213 : _GEN_3348; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3350 = 12'hd6 == _T_71[11:0] ? image_214 : _GEN_3349; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3351 = 12'hd7 == _T_71[11:0] ? image_215 : _GEN_3350; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3352 = 12'hd8 == _T_71[11:0] ? image_216 : _GEN_3351; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3353 = 12'hd9 == _T_71[11:0] ? image_217 : _GEN_3352; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3354 = 12'hda == _T_71[11:0] ? image_218 : _GEN_3353; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3355 = 12'hdb == _T_71[11:0] ? image_219 : _GEN_3354; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3356 = 12'hdc == _T_71[11:0] ? image_220 : _GEN_3355; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3357 = 12'hdd == _T_71[11:0] ? image_221 : _GEN_3356; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3358 = 12'hde == _T_71[11:0] ? image_222 : _GEN_3357; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3359 = 12'hdf == _T_71[11:0] ? image_223 : _GEN_3358; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3360 = 12'he0 == _T_71[11:0] ? image_224 : _GEN_3359; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3361 = 12'he1 == _T_71[11:0] ? image_225 : _GEN_3360; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3362 = 12'he2 == _T_71[11:0] ? image_226 : _GEN_3361; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3363 = 12'he3 == _T_71[11:0] ? image_227 : _GEN_3362; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3364 = 12'he4 == _T_71[11:0] ? image_228 : _GEN_3363; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3365 = 12'he5 == _T_71[11:0] ? image_229 : _GEN_3364; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3366 = 12'he6 == _T_71[11:0] ? image_230 : _GEN_3365; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3367 = 12'he7 == _T_71[11:0] ? image_231 : _GEN_3366; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3368 = 12'he8 == _T_71[11:0] ? image_232 : _GEN_3367; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3369 = 12'he9 == _T_71[11:0] ? image_233 : _GEN_3368; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3370 = 12'hea == _T_71[11:0] ? image_234 : _GEN_3369; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3371 = 12'heb == _T_71[11:0] ? image_235 : _GEN_3370; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3372 = 12'hec == _T_71[11:0] ? image_236 : _GEN_3371; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3373 = 12'hed == _T_71[11:0] ? image_237 : _GEN_3372; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3374 = 12'hee == _T_71[11:0] ? image_238 : _GEN_3373; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3375 = 12'hef == _T_71[11:0] ? image_239 : _GEN_3374; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3376 = 12'hf0 == _T_71[11:0] ? image_240 : _GEN_3375; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3377 = 12'hf1 == _T_71[11:0] ? image_241 : _GEN_3376; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3378 = 12'hf2 == _T_71[11:0] ? image_242 : _GEN_3377; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3379 = 12'hf3 == _T_71[11:0] ? image_243 : _GEN_3378; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3380 = 12'hf4 == _T_71[11:0] ? image_244 : _GEN_3379; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3381 = 12'hf5 == _T_71[11:0] ? image_245 : _GEN_3380; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3382 = 12'hf6 == _T_71[11:0] ? image_246 : _GEN_3381; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3383 = 12'hf7 == _T_71[11:0] ? 4'h0 : _GEN_3382; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3384 = 12'hf8 == _T_71[11:0] ? 4'h0 : _GEN_3383; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3385 = 12'hf9 == _T_71[11:0] ? 4'h0 : _GEN_3384; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3386 = 12'hfa == _T_71[11:0] ? 4'h0 : _GEN_3385; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3387 = 12'hfb == _T_71[11:0] ? 4'h0 : _GEN_3386; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3388 = 12'hfc == _T_71[11:0] ? 4'h0 : _GEN_3387; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3389 = 12'hfd == _T_71[11:0] ? 4'h0 : _GEN_3388; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3390 = 12'hfe == _T_71[11:0] ? 4'h0 : _GEN_3389; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3391 = 12'hff == _T_71[11:0] ? 4'h0 : _GEN_3390; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3392 = 12'h100 == _T_71[11:0] ? 4'h0 : _GEN_3391; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3393 = 12'h101 == _T_71[11:0] ? 4'h0 : _GEN_3392; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3394 = 12'h102 == _T_71[11:0] ? 4'h0 : _GEN_3393; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3395 = 12'h103 == _T_71[11:0] ? 4'h0 : _GEN_3394; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3396 = 12'h104 == _T_71[11:0] ? 4'h0 : _GEN_3395; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3397 = 12'h105 == _T_71[11:0] ? 4'h0 : _GEN_3396; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3398 = 12'h106 == _T_71[11:0] ? image_262 : _GEN_3397; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3399 = 12'h107 == _T_71[11:0] ? image_263 : _GEN_3398; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3400 = 12'h108 == _T_71[11:0] ? image_264 : _GEN_3399; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3401 = 12'h109 == _T_71[11:0] ? image_265 : _GEN_3400; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3402 = 12'h10a == _T_71[11:0] ? image_266 : _GEN_3401; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3403 = 12'h10b == _T_71[11:0] ? image_267 : _GEN_3402; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3404 = 12'h10c == _T_71[11:0] ? image_268 : _GEN_3403; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3405 = 12'h10d == _T_71[11:0] ? image_269 : _GEN_3404; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3406 = 12'h10e == _T_71[11:0] ? image_270 : _GEN_3405; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3407 = 12'h10f == _T_71[11:0] ? image_271 : _GEN_3406; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3408 = 12'h110 == _T_71[11:0] ? image_272 : _GEN_3407; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3409 = 12'h111 == _T_71[11:0] ? image_273 : _GEN_3408; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3410 = 12'h112 == _T_71[11:0] ? image_274 : _GEN_3409; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3411 = 12'h113 == _T_71[11:0] ? image_275 : _GEN_3410; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3412 = 12'h114 == _T_71[11:0] ? image_276 : _GEN_3411; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3413 = 12'h115 == _T_71[11:0] ? image_277 : _GEN_3412; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3414 = 12'h116 == _T_71[11:0] ? image_278 : _GEN_3413; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3415 = 12'h117 == _T_71[11:0] ? image_279 : _GEN_3414; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3416 = 12'h118 == _T_71[11:0] ? image_280 : _GEN_3415; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3417 = 12'h119 == _T_71[11:0] ? image_281 : _GEN_3416; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3418 = 12'h11a == _T_71[11:0] ? image_282 : _GEN_3417; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3419 = 12'h11b == _T_71[11:0] ? image_283 : _GEN_3418; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3420 = 12'h11c == _T_71[11:0] ? image_284 : _GEN_3419; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3421 = 12'h11d == _T_71[11:0] ? image_285 : _GEN_3420; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3422 = 12'h11e == _T_71[11:0] ? image_286 : _GEN_3421; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3423 = 12'h11f == _T_71[11:0] ? image_287 : _GEN_3422; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3424 = 12'h120 == _T_71[11:0] ? image_288 : _GEN_3423; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3425 = 12'h121 == _T_71[11:0] ? image_289 : _GEN_3424; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3426 = 12'h122 == _T_71[11:0] ? image_290 : _GEN_3425; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3427 = 12'h123 == _T_71[11:0] ? image_291 : _GEN_3426; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3428 = 12'h124 == _T_71[11:0] ? image_292 : _GEN_3427; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3429 = 12'h125 == _T_71[11:0] ? image_293 : _GEN_3428; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3430 = 12'h126 == _T_71[11:0] ? image_294 : _GEN_3429; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3431 = 12'h127 == _T_71[11:0] ? image_295 : _GEN_3430; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3432 = 12'h128 == _T_71[11:0] ? image_296 : _GEN_3431; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3433 = 12'h129 == _T_71[11:0] ? image_297 : _GEN_3432; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3434 = 12'h12a == _T_71[11:0] ? image_298 : _GEN_3433; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3435 = 12'h12b == _T_71[11:0] ? image_299 : _GEN_3434; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3436 = 12'h12c == _T_71[11:0] ? image_300 : _GEN_3435; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3437 = 12'h12d == _T_71[11:0] ? image_301 : _GEN_3436; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3438 = 12'h12e == _T_71[11:0] ? image_302 : _GEN_3437; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3439 = 12'h12f == _T_71[11:0] ? image_303 : _GEN_3438; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3440 = 12'h130 == _T_71[11:0] ? image_304 : _GEN_3439; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3441 = 12'h131 == _T_71[11:0] ? image_305 : _GEN_3440; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3442 = 12'h132 == _T_71[11:0] ? image_306 : _GEN_3441; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3443 = 12'h133 == _T_71[11:0] ? image_307 : _GEN_3442; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3444 = 12'h134 == _T_71[11:0] ? image_308 : _GEN_3443; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3445 = 12'h135 == _T_71[11:0] ? image_309 : _GEN_3444; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3446 = 12'h136 == _T_71[11:0] ? image_310 : _GEN_3445; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3447 = 12'h137 == _T_71[11:0] ? image_311 : _GEN_3446; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3448 = 12'h138 == _T_71[11:0] ? image_312 : _GEN_3447; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3449 = 12'h139 == _T_71[11:0] ? image_313 : _GEN_3448; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3450 = 12'h13a == _T_71[11:0] ? image_314 : _GEN_3449; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3451 = 12'h13b == _T_71[11:0] ? image_315 : _GEN_3450; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3452 = 12'h13c == _T_71[11:0] ? 4'h0 : _GEN_3451; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3453 = 12'h13d == _T_71[11:0] ? 4'h0 : _GEN_3452; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3454 = 12'h13e == _T_71[11:0] ? 4'h0 : _GEN_3453; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3455 = 12'h13f == _T_71[11:0] ? 4'h0 : _GEN_3454; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3456 = 12'h140 == _T_71[11:0] ? 4'h0 : _GEN_3455; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3457 = 12'h141 == _T_71[11:0] ? 4'h0 : _GEN_3456; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3458 = 12'h142 == _T_71[11:0] ? 4'h0 : _GEN_3457; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3459 = 12'h143 == _T_71[11:0] ? 4'h0 : _GEN_3458; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3460 = 12'h144 == _T_71[11:0] ? 4'h0 : _GEN_3459; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3461 = 12'h145 == _T_71[11:0] ? image_325 : _GEN_3460; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3462 = 12'h146 == _T_71[11:0] ? image_326 : _GEN_3461; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3463 = 12'h147 == _T_71[11:0] ? image_327 : _GEN_3462; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3464 = 12'h148 == _T_71[11:0] ? image_328 : _GEN_3463; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3465 = 12'h149 == _T_71[11:0] ? image_329 : _GEN_3464; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3466 = 12'h14a == _T_71[11:0] ? image_330 : _GEN_3465; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3467 = 12'h14b == _T_71[11:0] ? image_331 : _GEN_3466; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3468 = 12'h14c == _T_71[11:0] ? image_332 : _GEN_3467; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3469 = 12'h14d == _T_71[11:0] ? image_333 : _GEN_3468; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3470 = 12'h14e == _T_71[11:0] ? image_334 : _GEN_3469; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3471 = 12'h14f == _T_71[11:0] ? image_335 : _GEN_3470; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3472 = 12'h150 == _T_71[11:0] ? image_336 : _GEN_3471; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3473 = 12'h151 == _T_71[11:0] ? image_337 : _GEN_3472; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3474 = 12'h152 == _T_71[11:0] ? image_338 : _GEN_3473; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3475 = 12'h153 == _T_71[11:0] ? image_339 : _GEN_3474; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3476 = 12'h154 == _T_71[11:0] ? image_340 : _GEN_3475; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3477 = 12'h155 == _T_71[11:0] ? image_341 : _GEN_3476; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3478 = 12'h156 == _T_71[11:0] ? image_342 : _GEN_3477; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3479 = 12'h157 == _T_71[11:0] ? image_343 : _GEN_3478; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3480 = 12'h158 == _T_71[11:0] ? image_344 : _GEN_3479; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3481 = 12'h159 == _T_71[11:0] ? image_345 : _GEN_3480; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3482 = 12'h15a == _T_71[11:0] ? image_346 : _GEN_3481; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3483 = 12'h15b == _T_71[11:0] ? image_347 : _GEN_3482; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3484 = 12'h15c == _T_71[11:0] ? image_348 : _GEN_3483; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3485 = 12'h15d == _T_71[11:0] ? image_349 : _GEN_3484; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3486 = 12'h15e == _T_71[11:0] ? image_350 : _GEN_3485; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3487 = 12'h15f == _T_71[11:0] ? image_351 : _GEN_3486; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3488 = 12'h160 == _T_71[11:0] ? image_352 : _GEN_3487; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3489 = 12'h161 == _T_71[11:0] ? image_353 : _GEN_3488; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3490 = 12'h162 == _T_71[11:0] ? image_354 : _GEN_3489; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3491 = 12'h163 == _T_71[11:0] ? image_355 : _GEN_3490; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3492 = 12'h164 == _T_71[11:0] ? image_356 : _GEN_3491; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3493 = 12'h165 == _T_71[11:0] ? image_357 : _GEN_3492; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3494 = 12'h166 == _T_71[11:0] ? image_358 : _GEN_3493; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3495 = 12'h167 == _T_71[11:0] ? image_359 : _GEN_3494; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3496 = 12'h168 == _T_71[11:0] ? image_360 : _GEN_3495; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3497 = 12'h169 == _T_71[11:0] ? image_361 : _GEN_3496; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3498 = 12'h16a == _T_71[11:0] ? image_362 : _GEN_3497; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3499 = 12'h16b == _T_71[11:0] ? image_363 : _GEN_3498; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3500 = 12'h16c == _T_71[11:0] ? image_364 : _GEN_3499; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3501 = 12'h16d == _T_71[11:0] ? image_365 : _GEN_3500; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3502 = 12'h16e == _T_71[11:0] ? image_366 : _GEN_3501; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3503 = 12'h16f == _T_71[11:0] ? image_367 : _GEN_3502; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3504 = 12'h170 == _T_71[11:0] ? image_368 : _GEN_3503; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3505 = 12'h171 == _T_71[11:0] ? image_369 : _GEN_3504; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3506 = 12'h172 == _T_71[11:0] ? image_370 : _GEN_3505; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3507 = 12'h173 == _T_71[11:0] ? image_371 : _GEN_3506; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3508 = 12'h174 == _T_71[11:0] ? image_372 : _GEN_3507; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3509 = 12'h175 == _T_71[11:0] ? image_373 : _GEN_3508; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3510 = 12'h176 == _T_71[11:0] ? image_374 : _GEN_3509; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3511 = 12'h177 == _T_71[11:0] ? image_375 : _GEN_3510; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3512 = 12'h178 == _T_71[11:0] ? image_376 : _GEN_3511; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3513 = 12'h179 == _T_71[11:0] ? image_377 : _GEN_3512; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3514 = 12'h17a == _T_71[11:0] ? image_378 : _GEN_3513; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3515 = 12'h17b == _T_71[11:0] ? image_379 : _GEN_3514; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3516 = 12'h17c == _T_71[11:0] ? 4'h0 : _GEN_3515; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3517 = 12'h17d == _T_71[11:0] ? 4'h0 : _GEN_3516; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3518 = 12'h17e == _T_71[11:0] ? 4'h0 : _GEN_3517; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3519 = 12'h17f == _T_71[11:0] ? 4'h0 : _GEN_3518; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3520 = 12'h180 == _T_71[11:0] ? 4'h0 : _GEN_3519; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3521 = 12'h181 == _T_71[11:0] ? 4'h0 : _GEN_3520; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3522 = 12'h182 == _T_71[11:0] ? 4'h0 : _GEN_3521; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3523 = 12'h183 == _T_71[11:0] ? 4'h0 : _GEN_3522; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3524 = 12'h184 == _T_71[11:0] ? image_388 : _GEN_3523; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3525 = 12'h185 == _T_71[11:0] ? image_389 : _GEN_3524; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3526 = 12'h186 == _T_71[11:0] ? image_390 : _GEN_3525; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3527 = 12'h187 == _T_71[11:0] ? image_391 : _GEN_3526; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3528 = 12'h188 == _T_71[11:0] ? image_392 : _GEN_3527; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3529 = 12'h189 == _T_71[11:0] ? image_393 : _GEN_3528; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3530 = 12'h18a == _T_71[11:0] ? image_394 : _GEN_3529; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3531 = 12'h18b == _T_71[11:0] ? image_395 : _GEN_3530; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3532 = 12'h18c == _T_71[11:0] ? image_396 : _GEN_3531; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3533 = 12'h18d == _T_71[11:0] ? image_397 : _GEN_3532; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3534 = 12'h18e == _T_71[11:0] ? image_398 : _GEN_3533; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3535 = 12'h18f == _T_71[11:0] ? image_399 : _GEN_3534; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3536 = 12'h190 == _T_71[11:0] ? image_400 : _GEN_3535; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3537 = 12'h191 == _T_71[11:0] ? image_401 : _GEN_3536; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3538 = 12'h192 == _T_71[11:0] ? image_402 : _GEN_3537; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3539 = 12'h193 == _T_71[11:0] ? image_403 : _GEN_3538; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3540 = 12'h194 == _T_71[11:0] ? image_404 : _GEN_3539; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3541 = 12'h195 == _T_71[11:0] ? image_405 : _GEN_3540; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3542 = 12'h196 == _T_71[11:0] ? image_406 : _GEN_3541; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3543 = 12'h197 == _T_71[11:0] ? image_407 : _GEN_3542; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3544 = 12'h198 == _T_71[11:0] ? image_408 : _GEN_3543; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3545 = 12'h199 == _T_71[11:0] ? image_409 : _GEN_3544; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3546 = 12'h19a == _T_71[11:0] ? image_410 : _GEN_3545; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3547 = 12'h19b == _T_71[11:0] ? image_411 : _GEN_3546; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3548 = 12'h19c == _T_71[11:0] ? image_412 : _GEN_3547; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3549 = 12'h19d == _T_71[11:0] ? image_413 : _GEN_3548; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3550 = 12'h19e == _T_71[11:0] ? image_414 : _GEN_3549; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3551 = 12'h19f == _T_71[11:0] ? image_415 : _GEN_3550; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3552 = 12'h1a0 == _T_71[11:0] ? image_416 : _GEN_3551; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3553 = 12'h1a1 == _T_71[11:0] ? image_417 : _GEN_3552; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3554 = 12'h1a2 == _T_71[11:0] ? image_418 : _GEN_3553; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3555 = 12'h1a3 == _T_71[11:0] ? image_419 : _GEN_3554; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3556 = 12'h1a4 == _T_71[11:0] ? image_420 : _GEN_3555; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3557 = 12'h1a5 == _T_71[11:0] ? image_421 : _GEN_3556; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3558 = 12'h1a6 == _T_71[11:0] ? image_422 : _GEN_3557; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3559 = 12'h1a7 == _T_71[11:0] ? image_423 : _GEN_3558; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3560 = 12'h1a8 == _T_71[11:0] ? image_424 : _GEN_3559; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3561 = 12'h1a9 == _T_71[11:0] ? image_425 : _GEN_3560; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3562 = 12'h1aa == _T_71[11:0] ? image_426 : _GEN_3561; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3563 = 12'h1ab == _T_71[11:0] ? image_427 : _GEN_3562; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3564 = 12'h1ac == _T_71[11:0] ? image_428 : _GEN_3563; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3565 = 12'h1ad == _T_71[11:0] ? image_429 : _GEN_3564; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3566 = 12'h1ae == _T_71[11:0] ? image_430 : _GEN_3565; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3567 = 12'h1af == _T_71[11:0] ? image_431 : _GEN_3566; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3568 = 12'h1b0 == _T_71[11:0] ? image_432 : _GEN_3567; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3569 = 12'h1b1 == _T_71[11:0] ? image_433 : _GEN_3568; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3570 = 12'h1b2 == _T_71[11:0] ? image_434 : _GEN_3569; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3571 = 12'h1b3 == _T_71[11:0] ? image_435 : _GEN_3570; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3572 = 12'h1b4 == _T_71[11:0] ? image_436 : _GEN_3571; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3573 = 12'h1b5 == _T_71[11:0] ? image_437 : _GEN_3572; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3574 = 12'h1b6 == _T_71[11:0] ? image_438 : _GEN_3573; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3575 = 12'h1b7 == _T_71[11:0] ? image_439 : _GEN_3574; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3576 = 12'h1b8 == _T_71[11:0] ? image_440 : _GEN_3575; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3577 = 12'h1b9 == _T_71[11:0] ? image_441 : _GEN_3576; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3578 = 12'h1ba == _T_71[11:0] ? image_442 : _GEN_3577; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3579 = 12'h1bb == _T_71[11:0] ? image_443 : _GEN_3578; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3580 = 12'h1bc == _T_71[11:0] ? image_444 : _GEN_3579; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3581 = 12'h1bd == _T_71[11:0] ? 4'h0 : _GEN_3580; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3582 = 12'h1be == _T_71[11:0] ? 4'h0 : _GEN_3581; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3583 = 12'h1bf == _T_71[11:0] ? 4'h0 : _GEN_3582; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3584 = 12'h1c0 == _T_71[11:0] ? 4'h0 : _GEN_3583; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3585 = 12'h1c1 == _T_71[11:0] ? 4'h0 : _GEN_3584; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3586 = 12'h1c2 == _T_71[11:0] ? 4'h0 : _GEN_3585; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3587 = 12'h1c3 == _T_71[11:0] ? image_451 : _GEN_3586; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3588 = 12'h1c4 == _T_71[11:0] ? image_452 : _GEN_3587; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3589 = 12'h1c5 == _T_71[11:0] ? image_453 : _GEN_3588; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3590 = 12'h1c6 == _T_71[11:0] ? image_454 : _GEN_3589; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3591 = 12'h1c7 == _T_71[11:0] ? image_455 : _GEN_3590; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3592 = 12'h1c8 == _T_71[11:0] ? image_456 : _GEN_3591; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3593 = 12'h1c9 == _T_71[11:0] ? image_457 : _GEN_3592; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3594 = 12'h1ca == _T_71[11:0] ? image_458 : _GEN_3593; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3595 = 12'h1cb == _T_71[11:0] ? image_459 : _GEN_3594; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3596 = 12'h1cc == _T_71[11:0] ? image_460 : _GEN_3595; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3597 = 12'h1cd == _T_71[11:0] ? image_461 : _GEN_3596; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3598 = 12'h1ce == _T_71[11:0] ? image_462 : _GEN_3597; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3599 = 12'h1cf == _T_71[11:0] ? image_463 : _GEN_3598; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3600 = 12'h1d0 == _T_71[11:0] ? image_464 : _GEN_3599; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3601 = 12'h1d1 == _T_71[11:0] ? image_465 : _GEN_3600; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3602 = 12'h1d2 == _T_71[11:0] ? image_466 : _GEN_3601; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3603 = 12'h1d3 == _T_71[11:0] ? image_467 : _GEN_3602; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3604 = 12'h1d4 == _T_71[11:0] ? image_468 : _GEN_3603; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3605 = 12'h1d5 == _T_71[11:0] ? image_469 : _GEN_3604; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3606 = 12'h1d6 == _T_71[11:0] ? image_470 : _GEN_3605; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3607 = 12'h1d7 == _T_71[11:0] ? image_471 : _GEN_3606; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3608 = 12'h1d8 == _T_71[11:0] ? image_472 : _GEN_3607; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3609 = 12'h1d9 == _T_71[11:0] ? image_473 : _GEN_3608; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3610 = 12'h1da == _T_71[11:0] ? image_474 : _GEN_3609; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3611 = 12'h1db == _T_71[11:0] ? image_475 : _GEN_3610; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3612 = 12'h1dc == _T_71[11:0] ? image_476 : _GEN_3611; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3613 = 12'h1dd == _T_71[11:0] ? image_477 : _GEN_3612; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3614 = 12'h1de == _T_71[11:0] ? image_478 : _GEN_3613; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3615 = 12'h1df == _T_71[11:0] ? image_479 : _GEN_3614; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3616 = 12'h1e0 == _T_71[11:0] ? image_480 : _GEN_3615; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3617 = 12'h1e1 == _T_71[11:0] ? image_481 : _GEN_3616; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3618 = 12'h1e2 == _T_71[11:0] ? image_482 : _GEN_3617; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3619 = 12'h1e3 == _T_71[11:0] ? image_483 : _GEN_3618; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3620 = 12'h1e4 == _T_71[11:0] ? image_484 : _GEN_3619; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3621 = 12'h1e5 == _T_71[11:0] ? image_485 : _GEN_3620; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3622 = 12'h1e6 == _T_71[11:0] ? image_486 : _GEN_3621; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3623 = 12'h1e7 == _T_71[11:0] ? image_487 : _GEN_3622; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3624 = 12'h1e8 == _T_71[11:0] ? image_488 : _GEN_3623; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3625 = 12'h1e9 == _T_71[11:0] ? image_489 : _GEN_3624; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3626 = 12'h1ea == _T_71[11:0] ? image_490 : _GEN_3625; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3627 = 12'h1eb == _T_71[11:0] ? image_491 : _GEN_3626; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3628 = 12'h1ec == _T_71[11:0] ? image_492 : _GEN_3627; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3629 = 12'h1ed == _T_71[11:0] ? image_493 : _GEN_3628; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3630 = 12'h1ee == _T_71[11:0] ? image_494 : _GEN_3629; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3631 = 12'h1ef == _T_71[11:0] ? image_495 : _GEN_3630; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3632 = 12'h1f0 == _T_71[11:0] ? image_496 : _GEN_3631; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3633 = 12'h1f1 == _T_71[11:0] ? image_497 : _GEN_3632; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3634 = 12'h1f2 == _T_71[11:0] ? image_498 : _GEN_3633; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3635 = 12'h1f3 == _T_71[11:0] ? image_499 : _GEN_3634; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3636 = 12'h1f4 == _T_71[11:0] ? image_500 : _GEN_3635; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3637 = 12'h1f5 == _T_71[11:0] ? image_501 : _GEN_3636; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3638 = 12'h1f6 == _T_71[11:0] ? image_502 : _GEN_3637; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3639 = 12'h1f7 == _T_71[11:0] ? image_503 : _GEN_3638; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3640 = 12'h1f8 == _T_71[11:0] ? image_504 : _GEN_3639; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3641 = 12'h1f9 == _T_71[11:0] ? image_505 : _GEN_3640; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3642 = 12'h1fa == _T_71[11:0] ? image_506 : _GEN_3641; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3643 = 12'h1fb == _T_71[11:0] ? image_507 : _GEN_3642; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3644 = 12'h1fc == _T_71[11:0] ? image_508 : _GEN_3643; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3645 = 12'h1fd == _T_71[11:0] ? image_509 : _GEN_3644; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3646 = 12'h1fe == _T_71[11:0] ? 4'h0 : _GEN_3645; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3647 = 12'h1ff == _T_71[11:0] ? 4'h0 : _GEN_3646; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3648 = 12'h200 == _T_71[11:0] ? 4'h0 : _GEN_3647; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3649 = 12'h201 == _T_71[11:0] ? 4'h0 : _GEN_3648; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3650 = 12'h202 == _T_71[11:0] ? 4'h0 : _GEN_3649; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3651 = 12'h203 == _T_71[11:0] ? image_515 : _GEN_3650; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3652 = 12'h204 == _T_71[11:0] ? image_516 : _GEN_3651; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3653 = 12'h205 == _T_71[11:0] ? image_517 : _GEN_3652; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3654 = 12'h206 == _T_71[11:0] ? image_518 : _GEN_3653; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3655 = 12'h207 == _T_71[11:0] ? image_519 : _GEN_3654; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3656 = 12'h208 == _T_71[11:0] ? image_520 : _GEN_3655; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3657 = 12'h209 == _T_71[11:0] ? image_521 : _GEN_3656; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3658 = 12'h20a == _T_71[11:0] ? image_522 : _GEN_3657; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3659 = 12'h20b == _T_71[11:0] ? image_523 : _GEN_3658; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3660 = 12'h20c == _T_71[11:0] ? image_524 : _GEN_3659; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3661 = 12'h20d == _T_71[11:0] ? image_525 : _GEN_3660; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3662 = 12'h20e == _T_71[11:0] ? image_526 : _GEN_3661; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3663 = 12'h20f == _T_71[11:0] ? image_527 : _GEN_3662; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3664 = 12'h210 == _T_71[11:0] ? image_528 : _GEN_3663; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3665 = 12'h211 == _T_71[11:0] ? image_529 : _GEN_3664; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3666 = 12'h212 == _T_71[11:0] ? image_530 : _GEN_3665; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3667 = 12'h213 == _T_71[11:0] ? image_531 : _GEN_3666; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3668 = 12'h214 == _T_71[11:0] ? image_532 : _GEN_3667; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3669 = 12'h215 == _T_71[11:0] ? image_533 : _GEN_3668; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3670 = 12'h216 == _T_71[11:0] ? image_534 : _GEN_3669; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3671 = 12'h217 == _T_71[11:0] ? image_535 : _GEN_3670; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3672 = 12'h218 == _T_71[11:0] ? image_536 : _GEN_3671; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3673 = 12'h219 == _T_71[11:0] ? image_537 : _GEN_3672; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3674 = 12'h21a == _T_71[11:0] ? image_538 : _GEN_3673; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3675 = 12'h21b == _T_71[11:0] ? image_539 : _GEN_3674; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3676 = 12'h21c == _T_71[11:0] ? image_540 : _GEN_3675; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3677 = 12'h21d == _T_71[11:0] ? image_541 : _GEN_3676; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3678 = 12'h21e == _T_71[11:0] ? image_542 : _GEN_3677; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3679 = 12'h21f == _T_71[11:0] ? image_543 : _GEN_3678; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3680 = 12'h220 == _T_71[11:0] ? image_544 : _GEN_3679; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3681 = 12'h221 == _T_71[11:0] ? image_545 : _GEN_3680; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3682 = 12'h222 == _T_71[11:0] ? image_546 : _GEN_3681; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3683 = 12'h223 == _T_71[11:0] ? image_547 : _GEN_3682; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3684 = 12'h224 == _T_71[11:0] ? image_548 : _GEN_3683; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3685 = 12'h225 == _T_71[11:0] ? image_549 : _GEN_3684; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3686 = 12'h226 == _T_71[11:0] ? image_550 : _GEN_3685; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3687 = 12'h227 == _T_71[11:0] ? image_551 : _GEN_3686; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3688 = 12'h228 == _T_71[11:0] ? image_552 : _GEN_3687; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3689 = 12'h229 == _T_71[11:0] ? image_553 : _GEN_3688; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3690 = 12'h22a == _T_71[11:0] ? image_554 : _GEN_3689; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3691 = 12'h22b == _T_71[11:0] ? image_555 : _GEN_3690; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3692 = 12'h22c == _T_71[11:0] ? image_556 : _GEN_3691; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3693 = 12'h22d == _T_71[11:0] ? image_557 : _GEN_3692; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3694 = 12'h22e == _T_71[11:0] ? image_558 : _GEN_3693; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3695 = 12'h22f == _T_71[11:0] ? image_559 : _GEN_3694; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3696 = 12'h230 == _T_71[11:0] ? image_560 : _GEN_3695; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3697 = 12'h231 == _T_71[11:0] ? image_561 : _GEN_3696; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3698 = 12'h232 == _T_71[11:0] ? image_562 : _GEN_3697; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3699 = 12'h233 == _T_71[11:0] ? image_563 : _GEN_3698; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3700 = 12'h234 == _T_71[11:0] ? image_564 : _GEN_3699; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3701 = 12'h235 == _T_71[11:0] ? image_565 : _GEN_3700; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3702 = 12'h236 == _T_71[11:0] ? image_566 : _GEN_3701; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3703 = 12'h237 == _T_71[11:0] ? 4'h0 : _GEN_3702; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3704 = 12'h238 == _T_71[11:0] ? 4'h0 : _GEN_3703; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3705 = 12'h239 == _T_71[11:0] ? 4'h0 : _GEN_3704; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3706 = 12'h23a == _T_71[11:0] ? 4'h0 : _GEN_3705; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3707 = 12'h23b == _T_71[11:0] ? image_571 : _GEN_3706; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3708 = 12'h23c == _T_71[11:0] ? image_572 : _GEN_3707; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3709 = 12'h23d == _T_71[11:0] ? image_573 : _GEN_3708; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3710 = 12'h23e == _T_71[11:0] ? image_574 : _GEN_3709; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3711 = 12'h23f == _T_71[11:0] ? 4'h0 : _GEN_3710; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3712 = 12'h240 == _T_71[11:0] ? 4'h0 : _GEN_3711; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3713 = 12'h241 == _T_71[11:0] ? 4'h0 : _GEN_3712; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3714 = 12'h242 == _T_71[11:0] ? image_578 : _GEN_3713; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3715 = 12'h243 == _T_71[11:0] ? image_579 : _GEN_3714; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3716 = 12'h244 == _T_71[11:0] ? image_580 : _GEN_3715; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3717 = 12'h245 == _T_71[11:0] ? image_581 : _GEN_3716; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3718 = 12'h246 == _T_71[11:0] ? image_582 : _GEN_3717; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3719 = 12'h247 == _T_71[11:0] ? image_583 : _GEN_3718; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3720 = 12'h248 == _T_71[11:0] ? image_584 : _GEN_3719; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3721 = 12'h249 == _T_71[11:0] ? image_585 : _GEN_3720; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3722 = 12'h24a == _T_71[11:0] ? image_586 : _GEN_3721; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3723 = 12'h24b == _T_71[11:0] ? image_587 : _GEN_3722; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3724 = 12'h24c == _T_71[11:0] ? image_588 : _GEN_3723; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3725 = 12'h24d == _T_71[11:0] ? image_589 : _GEN_3724; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3726 = 12'h24e == _T_71[11:0] ? image_590 : _GEN_3725; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3727 = 12'h24f == _T_71[11:0] ? image_591 : _GEN_3726; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3728 = 12'h250 == _T_71[11:0] ? image_592 : _GEN_3727; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3729 = 12'h251 == _T_71[11:0] ? image_593 : _GEN_3728; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3730 = 12'h252 == _T_71[11:0] ? image_594 : _GEN_3729; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3731 = 12'h253 == _T_71[11:0] ? image_595 : _GEN_3730; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3732 = 12'h254 == _T_71[11:0] ? image_596 : _GEN_3731; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3733 = 12'h255 == _T_71[11:0] ? image_597 : _GEN_3732; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3734 = 12'h256 == _T_71[11:0] ? image_598 : _GEN_3733; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3735 = 12'h257 == _T_71[11:0] ? image_599 : _GEN_3734; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3736 = 12'h258 == _T_71[11:0] ? image_600 : _GEN_3735; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3737 = 12'h259 == _T_71[11:0] ? image_601 : _GEN_3736; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3738 = 12'h25a == _T_71[11:0] ? image_602 : _GEN_3737; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3739 = 12'h25b == _T_71[11:0] ? image_603 : _GEN_3738; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3740 = 12'h25c == _T_71[11:0] ? image_604 : _GEN_3739; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3741 = 12'h25d == _T_71[11:0] ? image_605 : _GEN_3740; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3742 = 12'h25e == _T_71[11:0] ? image_606 : _GEN_3741; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3743 = 12'h25f == _T_71[11:0] ? image_607 : _GEN_3742; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3744 = 12'h260 == _T_71[11:0] ? 4'h0 : _GEN_3743; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3745 = 12'h261 == _T_71[11:0] ? 4'h0 : _GEN_3744; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3746 = 12'h262 == _T_71[11:0] ? 4'h0 : _GEN_3745; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3747 = 12'h263 == _T_71[11:0] ? 4'h0 : _GEN_3746; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3748 = 12'h264 == _T_71[11:0] ? 4'h0 : _GEN_3747; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3749 = 12'h265 == _T_71[11:0] ? 4'h0 : _GEN_3748; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3750 = 12'h266 == _T_71[11:0] ? image_614 : _GEN_3749; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3751 = 12'h267 == _T_71[11:0] ? image_615 : _GEN_3750; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3752 = 12'h268 == _T_71[11:0] ? image_616 : _GEN_3751; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3753 = 12'h269 == _T_71[11:0] ? image_617 : _GEN_3752; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3754 = 12'h26a == _T_71[11:0] ? image_618 : _GEN_3753; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3755 = 12'h26b == _T_71[11:0] ? image_619 : _GEN_3754; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3756 = 12'h26c == _T_71[11:0] ? image_620 : _GEN_3755; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3757 = 12'h26d == _T_71[11:0] ? image_621 : _GEN_3756; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3758 = 12'h26e == _T_71[11:0] ? image_622 : _GEN_3757; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3759 = 12'h26f == _T_71[11:0] ? image_623 : _GEN_3758; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3760 = 12'h270 == _T_71[11:0] ? image_624 : _GEN_3759; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3761 = 12'h271 == _T_71[11:0] ? image_625 : _GEN_3760; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3762 = 12'h272 == _T_71[11:0] ? image_626 : _GEN_3761; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3763 = 12'h273 == _T_71[11:0] ? image_627 : _GEN_3762; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3764 = 12'h274 == _T_71[11:0] ? image_628 : _GEN_3763; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3765 = 12'h275 == _T_71[11:0] ? 4'h0 : _GEN_3764; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3766 = 12'h276 == _T_71[11:0] ? 4'h0 : _GEN_3765; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3767 = 12'h277 == _T_71[11:0] ? 4'h0 : _GEN_3766; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3768 = 12'h278 == _T_71[11:0] ? 4'h0 : _GEN_3767; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3769 = 12'h279 == _T_71[11:0] ? 4'h0 : _GEN_3768; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3770 = 12'h27a == _T_71[11:0] ? 4'h0 : _GEN_3769; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3771 = 12'h27b == _T_71[11:0] ? 4'h0 : _GEN_3770; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3772 = 12'h27c == _T_71[11:0] ? image_636 : _GEN_3771; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3773 = 12'h27d == _T_71[11:0] ? image_637 : _GEN_3772; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3774 = 12'h27e == _T_71[11:0] ? image_638 : _GEN_3773; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3775 = 12'h27f == _T_71[11:0] ? image_639 : _GEN_3774; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3776 = 12'h280 == _T_71[11:0] ? 4'h0 : _GEN_3775; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3777 = 12'h281 == _T_71[11:0] ? 4'h0 : _GEN_3776; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3778 = 12'h282 == _T_71[11:0] ? image_642 : _GEN_3777; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3779 = 12'h283 == _T_71[11:0] ? image_643 : _GEN_3778; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3780 = 12'h284 == _T_71[11:0] ? image_644 : _GEN_3779; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3781 = 12'h285 == _T_71[11:0] ? image_645 : _GEN_3780; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3782 = 12'h286 == _T_71[11:0] ? image_646 : _GEN_3781; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3783 = 12'h287 == _T_71[11:0] ? image_647 : _GEN_3782; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3784 = 12'h288 == _T_71[11:0] ? image_648 : _GEN_3783; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3785 = 12'h289 == _T_71[11:0] ? image_649 : _GEN_3784; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3786 = 12'h28a == _T_71[11:0] ? image_650 : _GEN_3785; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3787 = 12'h28b == _T_71[11:0] ? image_651 : _GEN_3786; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3788 = 12'h28c == _T_71[11:0] ? image_652 : _GEN_3787; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3789 = 12'h28d == _T_71[11:0] ? image_653 : _GEN_3788; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3790 = 12'h28e == _T_71[11:0] ? image_654 : _GEN_3789; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3791 = 12'h28f == _T_71[11:0] ? image_655 : _GEN_3790; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3792 = 12'h290 == _T_71[11:0] ? image_656 : _GEN_3791; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3793 = 12'h291 == _T_71[11:0] ? image_657 : _GEN_3792; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3794 = 12'h292 == _T_71[11:0] ? image_658 : _GEN_3793; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3795 = 12'h293 == _T_71[11:0] ? image_659 : _GEN_3794; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3796 = 12'h294 == _T_71[11:0] ? image_660 : _GEN_3795; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3797 = 12'h295 == _T_71[11:0] ? image_661 : _GEN_3796; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3798 = 12'h296 == _T_71[11:0] ? image_662 : _GEN_3797; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3799 = 12'h297 == _T_71[11:0] ? image_663 : _GEN_3798; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3800 = 12'h298 == _T_71[11:0] ? image_664 : _GEN_3799; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3801 = 12'h299 == _T_71[11:0] ? image_665 : _GEN_3800; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3802 = 12'h29a == _T_71[11:0] ? image_666 : _GEN_3801; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3803 = 12'h29b == _T_71[11:0] ? image_667 : _GEN_3802; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3804 = 12'h29c == _T_71[11:0] ? image_668 : _GEN_3803; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3805 = 12'h29d == _T_71[11:0] ? image_669 : _GEN_3804; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3806 = 12'h29e == _T_71[11:0] ? image_670 : _GEN_3805; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3807 = 12'h29f == _T_71[11:0] ? 4'h0 : _GEN_3806; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3808 = 12'h2a0 == _T_71[11:0] ? 4'h0 : _GEN_3807; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3809 = 12'h2a1 == _T_71[11:0] ? 4'h0 : _GEN_3808; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3810 = 12'h2a2 == _T_71[11:0] ? 4'h0 : _GEN_3809; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3811 = 12'h2a3 == _T_71[11:0] ? 4'h0 : _GEN_3810; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3812 = 12'h2a4 == _T_71[11:0] ? 4'h0 : _GEN_3811; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3813 = 12'h2a5 == _T_71[11:0] ? 4'h0 : _GEN_3812; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3814 = 12'h2a6 == _T_71[11:0] ? 4'h0 : _GEN_3813; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3815 = 12'h2a7 == _T_71[11:0] ? image_679 : _GEN_3814; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3816 = 12'h2a8 == _T_71[11:0] ? image_680 : _GEN_3815; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3817 = 12'h2a9 == _T_71[11:0] ? image_681 : _GEN_3816; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3818 = 12'h2aa == _T_71[11:0] ? image_682 : _GEN_3817; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3819 = 12'h2ab == _T_71[11:0] ? image_683 : _GEN_3818; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3820 = 12'h2ac == _T_71[11:0] ? image_684 : _GEN_3819; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3821 = 12'h2ad == _T_71[11:0] ? image_685 : _GEN_3820; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3822 = 12'h2ae == _T_71[11:0] ? image_686 : _GEN_3821; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3823 = 12'h2af == _T_71[11:0] ? image_687 : _GEN_3822; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3824 = 12'h2b0 == _T_71[11:0] ? image_688 : _GEN_3823; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3825 = 12'h2b1 == _T_71[11:0] ? image_689 : _GEN_3824; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3826 = 12'h2b2 == _T_71[11:0] ? image_690 : _GEN_3825; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3827 = 12'h2b3 == _T_71[11:0] ? image_691 : _GEN_3826; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3828 = 12'h2b4 == _T_71[11:0] ? image_692 : _GEN_3827; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3829 = 12'h2b5 == _T_71[11:0] ? image_693 : _GEN_3828; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3830 = 12'h2b6 == _T_71[11:0] ? image_694 : _GEN_3829; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3831 = 12'h2b7 == _T_71[11:0] ? image_695 : _GEN_3830; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3832 = 12'h2b8 == _T_71[11:0] ? image_696 : _GEN_3831; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3833 = 12'h2b9 == _T_71[11:0] ? image_697 : _GEN_3832; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3834 = 12'h2ba == _T_71[11:0] ? image_698 : _GEN_3833; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3835 = 12'h2bb == _T_71[11:0] ? 4'h0 : _GEN_3834; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3836 = 12'h2bc == _T_71[11:0] ? 4'h0 : _GEN_3835; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3837 = 12'h2bd == _T_71[11:0] ? image_701 : _GEN_3836; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3838 = 12'h2be == _T_71[11:0] ? image_702 : _GEN_3837; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3839 = 12'h2bf == _T_71[11:0] ? image_703 : _GEN_3838; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3840 = 12'h2c0 == _T_71[11:0] ? 4'h0 : _GEN_3839; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3841 = 12'h2c1 == _T_71[11:0] ? image_705 : _GEN_3840; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3842 = 12'h2c2 == _T_71[11:0] ? image_706 : _GEN_3841; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3843 = 12'h2c3 == _T_71[11:0] ? image_707 : _GEN_3842; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3844 = 12'h2c4 == _T_71[11:0] ? image_708 : _GEN_3843; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3845 = 12'h2c5 == _T_71[11:0] ? image_709 : _GEN_3844; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3846 = 12'h2c6 == _T_71[11:0] ? image_710 : _GEN_3845; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3847 = 12'h2c7 == _T_71[11:0] ? image_711 : _GEN_3846; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3848 = 12'h2c8 == _T_71[11:0] ? image_712 : _GEN_3847; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3849 = 12'h2c9 == _T_71[11:0] ? image_713 : _GEN_3848; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3850 = 12'h2ca == _T_71[11:0] ? image_714 : _GEN_3849; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3851 = 12'h2cb == _T_71[11:0] ? image_715 : _GEN_3850; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3852 = 12'h2cc == _T_71[11:0] ? image_716 : _GEN_3851; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3853 = 12'h2cd == _T_71[11:0] ? image_717 : _GEN_3852; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3854 = 12'h2ce == _T_71[11:0] ? image_718 : _GEN_3853; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3855 = 12'h2cf == _T_71[11:0] ? image_719 : _GEN_3854; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3856 = 12'h2d0 == _T_71[11:0] ? image_720 : _GEN_3855; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3857 = 12'h2d1 == _T_71[11:0] ? image_721 : _GEN_3856; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3858 = 12'h2d2 == _T_71[11:0] ? image_722 : _GEN_3857; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3859 = 12'h2d3 == _T_71[11:0] ? image_723 : _GEN_3858; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3860 = 12'h2d4 == _T_71[11:0] ? image_724 : _GEN_3859; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3861 = 12'h2d5 == _T_71[11:0] ? image_725 : _GEN_3860; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3862 = 12'h2d6 == _T_71[11:0] ? image_726 : _GEN_3861; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3863 = 12'h2d7 == _T_71[11:0] ? image_727 : _GEN_3862; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3864 = 12'h2d8 == _T_71[11:0] ? image_728 : _GEN_3863; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3865 = 12'h2d9 == _T_71[11:0] ? image_729 : _GEN_3864; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3866 = 12'h2da == _T_71[11:0] ? image_730 : _GEN_3865; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3867 = 12'h2db == _T_71[11:0] ? image_731 : _GEN_3866; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3868 = 12'h2dc == _T_71[11:0] ? image_732 : _GEN_3867; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3869 = 12'h2dd == _T_71[11:0] ? image_733 : _GEN_3868; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3870 = 12'h2de == _T_71[11:0] ? image_734 : _GEN_3869; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3871 = 12'h2df == _T_71[11:0] ? 4'h0 : _GEN_3870; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3872 = 12'h2e0 == _T_71[11:0] ? image_736 : _GEN_3871; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3873 = 12'h2e1 == _T_71[11:0] ? image_737 : _GEN_3872; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3874 = 12'h2e2 == _T_71[11:0] ? 4'h0 : _GEN_3873; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3875 = 12'h2e3 == _T_71[11:0] ? image_739 : _GEN_3874; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3876 = 12'h2e4 == _T_71[11:0] ? image_740 : _GEN_3875; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3877 = 12'h2e5 == _T_71[11:0] ? image_741 : _GEN_3876; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3878 = 12'h2e6 == _T_71[11:0] ? 4'h0 : _GEN_3877; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3879 = 12'h2e7 == _T_71[11:0] ? 4'h0 : _GEN_3878; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3880 = 12'h2e8 == _T_71[11:0] ? image_744 : _GEN_3879; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3881 = 12'h2e9 == _T_71[11:0] ? image_745 : _GEN_3880; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3882 = 12'h2ea == _T_71[11:0] ? image_746 : _GEN_3881; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3883 = 12'h2eb == _T_71[11:0] ? image_747 : _GEN_3882; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3884 = 12'h2ec == _T_71[11:0] ? image_748 : _GEN_3883; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3885 = 12'h2ed == _T_71[11:0] ? image_749 : _GEN_3884; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3886 = 12'h2ee == _T_71[11:0] ? image_750 : _GEN_3885; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3887 = 12'h2ef == _T_71[11:0] ? image_751 : _GEN_3886; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3888 = 12'h2f0 == _T_71[11:0] ? image_752 : _GEN_3887; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3889 = 12'h2f1 == _T_71[11:0] ? image_753 : _GEN_3888; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3890 = 12'h2f2 == _T_71[11:0] ? image_754 : _GEN_3889; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3891 = 12'h2f3 == _T_71[11:0] ? image_755 : _GEN_3890; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3892 = 12'h2f4 == _T_71[11:0] ? image_756 : _GEN_3891; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3893 = 12'h2f5 == _T_71[11:0] ? 4'h0 : _GEN_3892; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3894 = 12'h2f6 == _T_71[11:0] ? image_758 : _GEN_3893; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3895 = 12'h2f7 == _T_71[11:0] ? 4'h0 : _GEN_3894; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3896 = 12'h2f8 == _T_71[11:0] ? image_760 : _GEN_3895; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3897 = 12'h2f9 == _T_71[11:0] ? image_761 : _GEN_3896; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3898 = 12'h2fa == _T_71[11:0] ? image_762 : _GEN_3897; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3899 = 12'h2fb == _T_71[11:0] ? image_763 : _GEN_3898; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3900 = 12'h2fc == _T_71[11:0] ? 4'h0 : _GEN_3899; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3901 = 12'h2fd == _T_71[11:0] ? image_765 : _GEN_3900; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3902 = 12'h2fe == _T_71[11:0] ? image_766 : _GEN_3901; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3903 = 12'h2ff == _T_71[11:0] ? image_767 : _GEN_3902; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3904 = 12'h300 == _T_71[11:0] ? image_768 : _GEN_3903; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3905 = 12'h301 == _T_71[11:0] ? image_769 : _GEN_3904; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3906 = 12'h302 == _T_71[11:0] ? image_770 : _GEN_3905; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3907 = 12'h303 == _T_71[11:0] ? image_771 : _GEN_3906; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3908 = 12'h304 == _T_71[11:0] ? image_772 : _GEN_3907; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3909 = 12'h305 == _T_71[11:0] ? image_773 : _GEN_3908; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3910 = 12'h306 == _T_71[11:0] ? image_774 : _GEN_3909; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3911 = 12'h307 == _T_71[11:0] ? image_775 : _GEN_3910; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3912 = 12'h308 == _T_71[11:0] ? image_776 : _GEN_3911; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3913 = 12'h309 == _T_71[11:0] ? image_777 : _GEN_3912; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3914 = 12'h30a == _T_71[11:0] ? image_778 : _GEN_3913; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3915 = 12'h30b == _T_71[11:0] ? image_779 : _GEN_3914; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3916 = 12'h30c == _T_71[11:0] ? image_780 : _GEN_3915; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3917 = 12'h30d == _T_71[11:0] ? image_781 : _GEN_3916; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3918 = 12'h30e == _T_71[11:0] ? image_782 : _GEN_3917; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3919 = 12'h30f == _T_71[11:0] ? image_783 : _GEN_3918; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3920 = 12'h310 == _T_71[11:0] ? image_784 : _GEN_3919; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3921 = 12'h311 == _T_71[11:0] ? image_785 : _GEN_3920; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3922 = 12'h312 == _T_71[11:0] ? image_786 : _GEN_3921; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3923 = 12'h313 == _T_71[11:0] ? image_787 : _GEN_3922; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3924 = 12'h314 == _T_71[11:0] ? image_788 : _GEN_3923; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3925 = 12'h315 == _T_71[11:0] ? image_789 : _GEN_3924; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3926 = 12'h316 == _T_71[11:0] ? image_790 : _GEN_3925; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3927 = 12'h317 == _T_71[11:0] ? image_791 : _GEN_3926; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3928 = 12'h318 == _T_71[11:0] ? image_792 : _GEN_3927; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3929 = 12'h319 == _T_71[11:0] ? image_793 : _GEN_3928; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3930 = 12'h31a == _T_71[11:0] ? image_794 : _GEN_3929; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3931 = 12'h31b == _T_71[11:0] ? image_795 : _GEN_3930; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3932 = 12'h31c == _T_71[11:0] ? image_796 : _GEN_3931; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3933 = 12'h31d == _T_71[11:0] ? image_797 : _GEN_3932; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3934 = 12'h31e == _T_71[11:0] ? 4'h0 : _GEN_3933; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3935 = 12'h31f == _T_71[11:0] ? 4'h0 : _GEN_3934; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3936 = 12'h320 == _T_71[11:0] ? image_800 : _GEN_3935; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3937 = 12'h321 == _T_71[11:0] ? image_801 : _GEN_3936; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3938 = 12'h322 == _T_71[11:0] ? image_802 : _GEN_3937; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3939 = 12'h323 == _T_71[11:0] ? image_803 : _GEN_3938; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3940 = 12'h324 == _T_71[11:0] ? image_804 : _GEN_3939; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3941 = 12'h325 == _T_71[11:0] ? image_805 : _GEN_3940; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3942 = 12'h326 == _T_71[11:0] ? image_806 : _GEN_3941; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3943 = 12'h327 == _T_71[11:0] ? 4'h0 : _GEN_3942; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3944 = 12'h328 == _T_71[11:0] ? image_808 : _GEN_3943; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3945 = 12'h329 == _T_71[11:0] ? image_809 : _GEN_3944; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3946 = 12'h32a == _T_71[11:0] ? image_810 : _GEN_3945; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3947 = 12'h32b == _T_71[11:0] ? image_811 : _GEN_3946; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3948 = 12'h32c == _T_71[11:0] ? image_812 : _GEN_3947; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3949 = 12'h32d == _T_71[11:0] ? image_813 : _GEN_3948; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3950 = 12'h32e == _T_71[11:0] ? image_814 : _GEN_3949; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3951 = 12'h32f == _T_71[11:0] ? image_815 : _GEN_3950; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3952 = 12'h330 == _T_71[11:0] ? image_816 : _GEN_3951; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3953 = 12'h331 == _T_71[11:0] ? image_817 : _GEN_3952; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3954 = 12'h332 == _T_71[11:0] ? image_818 : _GEN_3953; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3955 = 12'h333 == _T_71[11:0] ? image_819 : _GEN_3954; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3956 = 12'h334 == _T_71[11:0] ? image_820 : _GEN_3955; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3957 = 12'h335 == _T_71[11:0] ? 4'h0 : _GEN_3956; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3958 = 12'h336 == _T_71[11:0] ? image_822 : _GEN_3957; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3959 = 12'h337 == _T_71[11:0] ? image_823 : _GEN_3958; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3960 = 12'h338 == _T_71[11:0] ? image_824 : _GEN_3959; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3961 = 12'h339 == _T_71[11:0] ? image_825 : _GEN_3960; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3962 = 12'h33a == _T_71[11:0] ? image_826 : _GEN_3961; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3963 = 12'h33b == _T_71[11:0] ? 4'h0 : _GEN_3962; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3964 = 12'h33c == _T_71[11:0] ? image_828 : _GEN_3963; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3965 = 12'h33d == _T_71[11:0] ? image_829 : _GEN_3964; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3966 = 12'h33e == _T_71[11:0] ? image_830 : _GEN_3965; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3967 = 12'h33f == _T_71[11:0] ? image_831 : _GEN_3966; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3968 = 12'h340 == _T_71[11:0] ? 4'h0 : _GEN_3967; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3969 = 12'h341 == _T_71[11:0] ? image_833 : _GEN_3968; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3970 = 12'h342 == _T_71[11:0] ? image_834 : _GEN_3969; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3971 = 12'h343 == _T_71[11:0] ? image_835 : _GEN_3970; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3972 = 12'h344 == _T_71[11:0] ? image_836 : _GEN_3971; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3973 = 12'h345 == _T_71[11:0] ? image_837 : _GEN_3972; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3974 = 12'h346 == _T_71[11:0] ? image_838 : _GEN_3973; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3975 = 12'h347 == _T_71[11:0] ? image_839 : _GEN_3974; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3976 = 12'h348 == _T_71[11:0] ? image_840 : _GEN_3975; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3977 = 12'h349 == _T_71[11:0] ? image_841 : _GEN_3976; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3978 = 12'h34a == _T_71[11:0] ? image_842 : _GEN_3977; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3979 = 12'h34b == _T_71[11:0] ? image_843 : _GEN_3978; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3980 = 12'h34c == _T_71[11:0] ? image_844 : _GEN_3979; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3981 = 12'h34d == _T_71[11:0] ? image_845 : _GEN_3980; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3982 = 12'h34e == _T_71[11:0] ? image_846 : _GEN_3981; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3983 = 12'h34f == _T_71[11:0] ? image_847 : _GEN_3982; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3984 = 12'h350 == _T_71[11:0] ? image_848 : _GEN_3983; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3985 = 12'h351 == _T_71[11:0] ? image_849 : _GEN_3984; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3986 = 12'h352 == _T_71[11:0] ? image_850 : _GEN_3985; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3987 = 12'h353 == _T_71[11:0] ? image_851 : _GEN_3986; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3988 = 12'h354 == _T_71[11:0] ? image_852 : _GEN_3987; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3989 = 12'h355 == _T_71[11:0] ? image_853 : _GEN_3988; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3990 = 12'h356 == _T_71[11:0] ? image_854 : _GEN_3989; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3991 = 12'h357 == _T_71[11:0] ? image_855 : _GEN_3990; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3992 = 12'h358 == _T_71[11:0] ? image_856 : _GEN_3991; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3993 = 12'h359 == _T_71[11:0] ? image_857 : _GEN_3992; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3994 = 12'h35a == _T_71[11:0] ? image_858 : _GEN_3993; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3995 = 12'h35b == _T_71[11:0] ? image_859 : _GEN_3994; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3996 = 12'h35c == _T_71[11:0] ? image_860 : _GEN_3995; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3997 = 12'h35d == _T_71[11:0] ? image_861 : _GEN_3996; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3998 = 12'h35e == _T_71[11:0] ? image_862 : _GEN_3997; // @[Filter.scala 138:46]
  wire [3:0] _GEN_3999 = 12'h35f == _T_71[11:0] ? 4'h0 : _GEN_3998; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4000 = 12'h360 == _T_71[11:0] ? 4'h0 : _GEN_3999; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4001 = 12'h361 == _T_71[11:0] ? image_865 : _GEN_4000; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4002 = 12'h362 == _T_71[11:0] ? image_866 : _GEN_4001; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4003 = 12'h363 == _T_71[11:0] ? image_867 : _GEN_4002; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4004 = 12'h364 == _T_71[11:0] ? image_868 : _GEN_4003; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4005 = 12'h365 == _T_71[11:0] ? image_869 : _GEN_4004; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4006 = 12'h366 == _T_71[11:0] ? 4'h0 : _GEN_4005; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4007 = 12'h367 == _T_71[11:0] ? 4'h0 : _GEN_4006; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4008 = 12'h368 == _T_71[11:0] ? image_872 : _GEN_4007; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4009 = 12'h369 == _T_71[11:0] ? image_873 : _GEN_4008; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4010 = 12'h36a == _T_71[11:0] ? image_874 : _GEN_4009; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4011 = 12'h36b == _T_71[11:0] ? image_875 : _GEN_4010; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4012 = 12'h36c == _T_71[11:0] ? image_876 : _GEN_4011; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4013 = 12'h36d == _T_71[11:0] ? image_877 : _GEN_4012; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4014 = 12'h36e == _T_71[11:0] ? image_878 : _GEN_4013; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4015 = 12'h36f == _T_71[11:0] ? image_879 : _GEN_4014; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4016 = 12'h370 == _T_71[11:0] ? image_880 : _GEN_4015; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4017 = 12'h371 == _T_71[11:0] ? image_881 : _GEN_4016; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4018 = 12'h372 == _T_71[11:0] ? image_882 : _GEN_4017; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4019 = 12'h373 == _T_71[11:0] ? image_883 : _GEN_4018; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4020 = 12'h374 == _T_71[11:0] ? image_884 : _GEN_4019; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4021 = 12'h375 == _T_71[11:0] ? image_885 : _GEN_4020; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4022 = 12'h376 == _T_71[11:0] ? 4'h0 : _GEN_4021; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4023 = 12'h377 == _T_71[11:0] ? 4'h0 : _GEN_4022; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4024 = 12'h378 == _T_71[11:0] ? 4'h0 : _GEN_4023; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4025 = 12'h379 == _T_71[11:0] ? 4'h0 : _GEN_4024; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4026 = 12'h37a == _T_71[11:0] ? 4'h0 : _GEN_4025; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4027 = 12'h37b == _T_71[11:0] ? image_891 : _GEN_4026; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4028 = 12'h37c == _T_71[11:0] ? image_892 : _GEN_4027; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4029 = 12'h37d == _T_71[11:0] ? image_893 : _GEN_4028; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4030 = 12'h37e == _T_71[11:0] ? image_894 : _GEN_4029; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4031 = 12'h37f == _T_71[11:0] ? image_895 : _GEN_4030; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4032 = 12'h380 == _T_71[11:0] ? 4'h0 : _GEN_4031; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4033 = 12'h381 == _T_71[11:0] ? image_897 : _GEN_4032; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4034 = 12'h382 == _T_71[11:0] ? image_898 : _GEN_4033; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4035 = 12'h383 == _T_71[11:0] ? image_899 : _GEN_4034; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4036 = 12'h384 == _T_71[11:0] ? image_900 : _GEN_4035; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4037 = 12'h385 == _T_71[11:0] ? image_901 : _GEN_4036; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4038 = 12'h386 == _T_71[11:0] ? image_902 : _GEN_4037; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4039 = 12'h387 == _T_71[11:0] ? image_903 : _GEN_4038; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4040 = 12'h388 == _T_71[11:0] ? image_904 : _GEN_4039; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4041 = 12'h389 == _T_71[11:0] ? image_905 : _GEN_4040; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4042 = 12'h38a == _T_71[11:0] ? image_906 : _GEN_4041; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4043 = 12'h38b == _T_71[11:0] ? image_907 : _GEN_4042; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4044 = 12'h38c == _T_71[11:0] ? image_908 : _GEN_4043; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4045 = 12'h38d == _T_71[11:0] ? image_909 : _GEN_4044; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4046 = 12'h38e == _T_71[11:0] ? image_910 : _GEN_4045; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4047 = 12'h38f == _T_71[11:0] ? image_911 : _GEN_4046; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4048 = 12'h390 == _T_71[11:0] ? image_912 : _GEN_4047; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4049 = 12'h391 == _T_71[11:0] ? image_913 : _GEN_4048; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4050 = 12'h392 == _T_71[11:0] ? image_914 : _GEN_4049; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4051 = 12'h393 == _T_71[11:0] ? image_915 : _GEN_4050; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4052 = 12'h394 == _T_71[11:0] ? image_916 : _GEN_4051; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4053 = 12'h395 == _T_71[11:0] ? image_917 : _GEN_4052; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4054 = 12'h396 == _T_71[11:0] ? image_918 : _GEN_4053; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4055 = 12'h397 == _T_71[11:0] ? image_919 : _GEN_4054; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4056 = 12'h398 == _T_71[11:0] ? image_920 : _GEN_4055; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4057 = 12'h399 == _T_71[11:0] ? image_921 : _GEN_4056; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4058 = 12'h39a == _T_71[11:0] ? image_922 : _GEN_4057; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4059 = 12'h39b == _T_71[11:0] ? image_923 : _GEN_4058; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4060 = 12'h39c == _T_71[11:0] ? image_924 : _GEN_4059; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4061 = 12'h39d == _T_71[11:0] ? image_925 : _GEN_4060; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4062 = 12'h39e == _T_71[11:0] ? image_926 : _GEN_4061; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4063 = 12'h39f == _T_71[11:0] ? image_927 : _GEN_4062; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4064 = 12'h3a0 == _T_71[11:0] ? 4'h0 : _GEN_4063; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4065 = 12'h3a1 == _T_71[11:0] ? image_929 : _GEN_4064; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4066 = 12'h3a2 == _T_71[11:0] ? image_930 : _GEN_4065; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4067 = 12'h3a3 == _T_71[11:0] ? 4'h0 : _GEN_4066; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4068 = 12'h3a4 == _T_71[11:0] ? 4'h0 : _GEN_4067; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4069 = 12'h3a5 == _T_71[11:0] ? 4'h0 : _GEN_4068; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4070 = 12'h3a6 == _T_71[11:0] ? 4'h0 : _GEN_4069; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4071 = 12'h3a7 == _T_71[11:0] ? image_935 : _GEN_4070; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4072 = 12'h3a8 == _T_71[11:0] ? image_936 : _GEN_4071; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4073 = 12'h3a9 == _T_71[11:0] ? image_937 : _GEN_4072; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4074 = 12'h3aa == _T_71[11:0] ? image_938 : _GEN_4073; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4075 = 12'h3ab == _T_71[11:0] ? image_939 : _GEN_4074; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4076 = 12'h3ac == _T_71[11:0] ? image_940 : _GEN_4075; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4077 = 12'h3ad == _T_71[11:0] ? image_941 : _GEN_4076; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4078 = 12'h3ae == _T_71[11:0] ? image_942 : _GEN_4077; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4079 = 12'h3af == _T_71[11:0] ? image_943 : _GEN_4078; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4080 = 12'h3b0 == _T_71[11:0] ? image_944 : _GEN_4079; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4081 = 12'h3b1 == _T_71[11:0] ? image_945 : _GEN_4080; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4082 = 12'h3b2 == _T_71[11:0] ? image_946 : _GEN_4081; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4083 = 12'h3b3 == _T_71[11:0] ? image_947 : _GEN_4082; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4084 = 12'h3b4 == _T_71[11:0] ? image_948 : _GEN_4083; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4085 = 12'h3b5 == _T_71[11:0] ? image_949 : _GEN_4084; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4086 = 12'h3b6 == _T_71[11:0] ? image_950 : _GEN_4085; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4087 = 12'h3b7 == _T_71[11:0] ? image_951 : _GEN_4086; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4088 = 12'h3b8 == _T_71[11:0] ? image_952 : _GEN_4087; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4089 = 12'h3b9 == _T_71[11:0] ? image_953 : _GEN_4088; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4090 = 12'h3ba == _T_71[11:0] ? image_954 : _GEN_4089; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4091 = 12'h3bb == _T_71[11:0] ? image_955 : _GEN_4090; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4092 = 12'h3bc == _T_71[11:0] ? image_956 : _GEN_4091; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4093 = 12'h3bd == _T_71[11:0] ? image_957 : _GEN_4092; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4094 = 12'h3be == _T_71[11:0] ? image_958 : _GEN_4093; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4095 = 12'h3bf == _T_71[11:0] ? image_959 : _GEN_4094; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4096 = 12'h3c0 == _T_71[11:0] ? 4'h0 : _GEN_4095; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4097 = 12'h3c1 == _T_71[11:0] ? image_961 : _GEN_4096; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4098 = 12'h3c2 == _T_71[11:0] ? image_962 : _GEN_4097; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4099 = 12'h3c3 == _T_71[11:0] ? image_963 : _GEN_4098; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4100 = 12'h3c4 == _T_71[11:0] ? image_964 : _GEN_4099; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4101 = 12'h3c5 == _T_71[11:0] ? image_965 : _GEN_4100; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4102 = 12'h3c6 == _T_71[11:0] ? image_966 : _GEN_4101; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4103 = 12'h3c7 == _T_71[11:0] ? image_967 : _GEN_4102; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4104 = 12'h3c8 == _T_71[11:0] ? image_968 : _GEN_4103; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4105 = 12'h3c9 == _T_71[11:0] ? image_969 : _GEN_4104; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4106 = 12'h3ca == _T_71[11:0] ? image_970 : _GEN_4105; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4107 = 12'h3cb == _T_71[11:0] ? image_971 : _GEN_4106; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4108 = 12'h3cc == _T_71[11:0] ? image_972 : _GEN_4107; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4109 = 12'h3cd == _T_71[11:0] ? image_973 : _GEN_4108; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4110 = 12'h3ce == _T_71[11:0] ? image_974 : _GEN_4109; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4111 = 12'h3cf == _T_71[11:0] ? image_975 : _GEN_4110; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4112 = 12'h3d0 == _T_71[11:0] ? image_976 : _GEN_4111; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4113 = 12'h3d1 == _T_71[11:0] ? image_977 : _GEN_4112; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4114 = 12'h3d2 == _T_71[11:0] ? image_978 : _GEN_4113; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4115 = 12'h3d3 == _T_71[11:0] ? image_979 : _GEN_4114; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4116 = 12'h3d4 == _T_71[11:0] ? image_980 : _GEN_4115; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4117 = 12'h3d5 == _T_71[11:0] ? image_981 : _GEN_4116; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4118 = 12'h3d6 == _T_71[11:0] ? image_982 : _GEN_4117; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4119 = 12'h3d7 == _T_71[11:0] ? image_983 : _GEN_4118; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4120 = 12'h3d8 == _T_71[11:0] ? image_984 : _GEN_4119; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4121 = 12'h3d9 == _T_71[11:0] ? image_985 : _GEN_4120; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4122 = 12'h3da == _T_71[11:0] ? image_986 : _GEN_4121; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4123 = 12'h3db == _T_71[11:0] ? image_987 : _GEN_4122; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4124 = 12'h3dc == _T_71[11:0] ? image_988 : _GEN_4123; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4125 = 12'h3dd == _T_71[11:0] ? image_989 : _GEN_4124; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4126 = 12'h3de == _T_71[11:0] ? image_990 : _GEN_4125; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4127 = 12'h3df == _T_71[11:0] ? image_991 : _GEN_4126; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4128 = 12'h3e0 == _T_71[11:0] ? image_992 : _GEN_4127; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4129 = 12'h3e1 == _T_71[11:0] ? 4'h0 : _GEN_4128; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4130 = 12'h3e2 == _T_71[11:0] ? 4'h0 : _GEN_4129; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4131 = 12'h3e3 == _T_71[11:0] ? 4'h0 : _GEN_4130; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4132 = 12'h3e4 == _T_71[11:0] ? 4'h0 : _GEN_4131; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4133 = 12'h3e5 == _T_71[11:0] ? image_997 : _GEN_4132; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4134 = 12'h3e6 == _T_71[11:0] ? image_998 : _GEN_4133; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4135 = 12'h3e7 == _T_71[11:0] ? image_999 : _GEN_4134; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4136 = 12'h3e8 == _T_71[11:0] ? image_1000 : _GEN_4135; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4137 = 12'h3e9 == _T_71[11:0] ? image_1001 : _GEN_4136; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4138 = 12'h3ea == _T_71[11:0] ? image_1002 : _GEN_4137; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4139 = 12'h3eb == _T_71[11:0] ? image_1003 : _GEN_4138; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4140 = 12'h3ec == _T_71[11:0] ? image_1004 : _GEN_4139; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4141 = 12'h3ed == _T_71[11:0] ? image_1005 : _GEN_4140; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4142 = 12'h3ee == _T_71[11:0] ? image_1006 : _GEN_4141; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4143 = 12'h3ef == _T_71[11:0] ? image_1007 : _GEN_4142; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4144 = 12'h3f0 == _T_71[11:0] ? image_1008 : _GEN_4143; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4145 = 12'h3f1 == _T_71[11:0] ? image_1009 : _GEN_4144; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4146 = 12'h3f2 == _T_71[11:0] ? image_1010 : _GEN_4145; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4147 = 12'h3f3 == _T_71[11:0] ? image_1011 : _GEN_4146; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4148 = 12'h3f4 == _T_71[11:0] ? image_1012 : _GEN_4147; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4149 = 12'h3f5 == _T_71[11:0] ? image_1013 : _GEN_4148; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4150 = 12'h3f6 == _T_71[11:0] ? image_1014 : _GEN_4149; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4151 = 12'h3f7 == _T_71[11:0] ? image_1015 : _GEN_4150; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4152 = 12'h3f8 == _T_71[11:0] ? image_1016 : _GEN_4151; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4153 = 12'h3f9 == _T_71[11:0] ? image_1017 : _GEN_4152; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4154 = 12'h3fa == _T_71[11:0] ? image_1018 : _GEN_4153; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4155 = 12'h3fb == _T_71[11:0] ? image_1019 : _GEN_4154; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4156 = 12'h3fc == _T_71[11:0] ? image_1020 : _GEN_4155; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4157 = 12'h3fd == _T_71[11:0] ? 4'h0 : _GEN_4156; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4158 = 12'h3fe == _T_71[11:0] ? 4'h0 : _GEN_4157; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4159 = 12'h3ff == _T_71[11:0] ? 4'h0 : _GEN_4158; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4160 = 12'h400 == _T_71[11:0] ? image_1024 : _GEN_4159; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4161 = 12'h401 == _T_71[11:0] ? image_1025 : _GEN_4160; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4162 = 12'h402 == _T_71[11:0] ? image_1026 : _GEN_4161; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4163 = 12'h403 == _T_71[11:0] ? image_1027 : _GEN_4162; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4164 = 12'h404 == _T_71[11:0] ? image_1028 : _GEN_4163; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4165 = 12'h405 == _T_71[11:0] ? image_1029 : _GEN_4164; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4166 = 12'h406 == _T_71[11:0] ? image_1030 : _GEN_4165; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4167 = 12'h407 == _T_71[11:0] ? image_1031 : _GEN_4166; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4168 = 12'h408 == _T_71[11:0] ? image_1032 : _GEN_4167; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4169 = 12'h409 == _T_71[11:0] ? image_1033 : _GEN_4168; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4170 = 12'h40a == _T_71[11:0] ? image_1034 : _GEN_4169; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4171 = 12'h40b == _T_71[11:0] ? image_1035 : _GEN_4170; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4172 = 12'h40c == _T_71[11:0] ? image_1036 : _GEN_4171; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4173 = 12'h40d == _T_71[11:0] ? image_1037 : _GEN_4172; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4174 = 12'h40e == _T_71[11:0] ? image_1038 : _GEN_4173; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4175 = 12'h40f == _T_71[11:0] ? image_1039 : _GEN_4174; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4176 = 12'h410 == _T_71[11:0] ? image_1040 : _GEN_4175; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4177 = 12'h411 == _T_71[11:0] ? image_1041 : _GEN_4176; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4178 = 12'h412 == _T_71[11:0] ? image_1042 : _GEN_4177; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4179 = 12'h413 == _T_71[11:0] ? image_1043 : _GEN_4178; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4180 = 12'h414 == _T_71[11:0] ? image_1044 : _GEN_4179; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4181 = 12'h415 == _T_71[11:0] ? image_1045 : _GEN_4180; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4182 = 12'h416 == _T_71[11:0] ? image_1046 : _GEN_4181; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4183 = 12'h417 == _T_71[11:0] ? image_1047 : _GEN_4182; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4184 = 12'h418 == _T_71[11:0] ? image_1048 : _GEN_4183; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4185 = 12'h419 == _T_71[11:0] ? image_1049 : _GEN_4184; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4186 = 12'h41a == _T_71[11:0] ? image_1050 : _GEN_4185; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4187 = 12'h41b == _T_71[11:0] ? image_1051 : _GEN_4186; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4188 = 12'h41c == _T_71[11:0] ? image_1052 : _GEN_4187; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4189 = 12'h41d == _T_71[11:0] ? image_1053 : _GEN_4188; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4190 = 12'h41e == _T_71[11:0] ? image_1054 : _GEN_4189; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4191 = 12'h41f == _T_71[11:0] ? image_1055 : _GEN_4190; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4192 = 12'h420 == _T_71[11:0] ? image_1056 : _GEN_4191; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4193 = 12'h421 == _T_71[11:0] ? image_1057 : _GEN_4192; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4194 = 12'h422 == _T_71[11:0] ? image_1058 : _GEN_4193; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4195 = 12'h423 == _T_71[11:0] ? image_1059 : _GEN_4194; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4196 = 12'h424 == _T_71[11:0] ? image_1060 : _GEN_4195; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4197 = 12'h425 == _T_71[11:0] ? image_1061 : _GEN_4196; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4198 = 12'h426 == _T_71[11:0] ? image_1062 : _GEN_4197; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4199 = 12'h427 == _T_71[11:0] ? image_1063 : _GEN_4198; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4200 = 12'h428 == _T_71[11:0] ? image_1064 : _GEN_4199; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4201 = 12'h429 == _T_71[11:0] ? image_1065 : _GEN_4200; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4202 = 12'h42a == _T_71[11:0] ? image_1066 : _GEN_4201; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4203 = 12'h42b == _T_71[11:0] ? image_1067 : _GEN_4202; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4204 = 12'h42c == _T_71[11:0] ? image_1068 : _GEN_4203; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4205 = 12'h42d == _T_71[11:0] ? image_1069 : _GEN_4204; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4206 = 12'h42e == _T_71[11:0] ? image_1070 : _GEN_4205; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4207 = 12'h42f == _T_71[11:0] ? image_1071 : _GEN_4206; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4208 = 12'h430 == _T_71[11:0] ? image_1072 : _GEN_4207; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4209 = 12'h431 == _T_71[11:0] ? image_1073 : _GEN_4208; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4210 = 12'h432 == _T_71[11:0] ? image_1074 : _GEN_4209; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4211 = 12'h433 == _T_71[11:0] ? image_1075 : _GEN_4210; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4212 = 12'h434 == _T_71[11:0] ? image_1076 : _GEN_4211; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4213 = 12'h435 == _T_71[11:0] ? image_1077 : _GEN_4212; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4214 = 12'h436 == _T_71[11:0] ? image_1078 : _GEN_4213; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4215 = 12'h437 == _T_71[11:0] ? image_1079 : _GEN_4214; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4216 = 12'h438 == _T_71[11:0] ? image_1080 : _GEN_4215; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4217 = 12'h439 == _T_71[11:0] ? image_1081 : _GEN_4216; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4218 = 12'h43a == _T_71[11:0] ? image_1082 : _GEN_4217; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4219 = 12'h43b == _T_71[11:0] ? image_1083 : _GEN_4218; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4220 = 12'h43c == _T_71[11:0] ? image_1084 : _GEN_4219; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4221 = 12'h43d == _T_71[11:0] ? image_1085 : _GEN_4220; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4222 = 12'h43e == _T_71[11:0] ? 4'h0 : _GEN_4221; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4223 = 12'h43f == _T_71[11:0] ? 4'h0 : _GEN_4222; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4224 = 12'h440 == _T_71[11:0] ? image_1088 : _GEN_4223; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4225 = 12'h441 == _T_71[11:0] ? image_1089 : _GEN_4224; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4226 = 12'h442 == _T_71[11:0] ? image_1090 : _GEN_4225; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4227 = 12'h443 == _T_71[11:0] ? image_1091 : _GEN_4226; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4228 = 12'h444 == _T_71[11:0] ? image_1092 : _GEN_4227; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4229 = 12'h445 == _T_71[11:0] ? image_1093 : _GEN_4228; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4230 = 12'h446 == _T_71[11:0] ? image_1094 : _GEN_4229; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4231 = 12'h447 == _T_71[11:0] ? image_1095 : _GEN_4230; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4232 = 12'h448 == _T_71[11:0] ? image_1096 : _GEN_4231; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4233 = 12'h449 == _T_71[11:0] ? image_1097 : _GEN_4232; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4234 = 12'h44a == _T_71[11:0] ? image_1098 : _GEN_4233; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4235 = 12'h44b == _T_71[11:0] ? image_1099 : _GEN_4234; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4236 = 12'h44c == _T_71[11:0] ? image_1100 : _GEN_4235; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4237 = 12'h44d == _T_71[11:0] ? image_1101 : _GEN_4236; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4238 = 12'h44e == _T_71[11:0] ? image_1102 : _GEN_4237; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4239 = 12'h44f == _T_71[11:0] ? image_1103 : _GEN_4238; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4240 = 12'h450 == _T_71[11:0] ? image_1104 : _GEN_4239; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4241 = 12'h451 == _T_71[11:0] ? image_1105 : _GEN_4240; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4242 = 12'h452 == _T_71[11:0] ? image_1106 : _GEN_4241; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4243 = 12'h453 == _T_71[11:0] ? image_1107 : _GEN_4242; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4244 = 12'h454 == _T_71[11:0] ? image_1108 : _GEN_4243; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4245 = 12'h455 == _T_71[11:0] ? image_1109 : _GEN_4244; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4246 = 12'h456 == _T_71[11:0] ? image_1110 : _GEN_4245; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4247 = 12'h457 == _T_71[11:0] ? image_1111 : _GEN_4246; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4248 = 12'h458 == _T_71[11:0] ? image_1112 : _GEN_4247; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4249 = 12'h459 == _T_71[11:0] ? image_1113 : _GEN_4248; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4250 = 12'h45a == _T_71[11:0] ? image_1114 : _GEN_4249; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4251 = 12'h45b == _T_71[11:0] ? image_1115 : _GEN_4250; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4252 = 12'h45c == _T_71[11:0] ? image_1116 : _GEN_4251; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4253 = 12'h45d == _T_71[11:0] ? image_1117 : _GEN_4252; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4254 = 12'h45e == _T_71[11:0] ? image_1118 : _GEN_4253; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4255 = 12'h45f == _T_71[11:0] ? image_1119 : _GEN_4254; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4256 = 12'h460 == _T_71[11:0] ? image_1120 : _GEN_4255; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4257 = 12'h461 == _T_71[11:0] ? image_1121 : _GEN_4256; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4258 = 12'h462 == _T_71[11:0] ? image_1122 : _GEN_4257; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4259 = 12'h463 == _T_71[11:0] ? image_1123 : _GEN_4258; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4260 = 12'h464 == _T_71[11:0] ? image_1124 : _GEN_4259; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4261 = 12'h465 == _T_71[11:0] ? image_1125 : _GEN_4260; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4262 = 12'h466 == _T_71[11:0] ? image_1126 : _GEN_4261; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4263 = 12'h467 == _T_71[11:0] ? image_1127 : _GEN_4262; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4264 = 12'h468 == _T_71[11:0] ? image_1128 : _GEN_4263; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4265 = 12'h469 == _T_71[11:0] ? image_1129 : _GEN_4264; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4266 = 12'h46a == _T_71[11:0] ? image_1130 : _GEN_4265; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4267 = 12'h46b == _T_71[11:0] ? image_1131 : _GEN_4266; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4268 = 12'h46c == _T_71[11:0] ? image_1132 : _GEN_4267; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4269 = 12'h46d == _T_71[11:0] ? image_1133 : _GEN_4268; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4270 = 12'h46e == _T_71[11:0] ? image_1134 : _GEN_4269; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4271 = 12'h46f == _T_71[11:0] ? image_1135 : _GEN_4270; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4272 = 12'h470 == _T_71[11:0] ? image_1136 : _GEN_4271; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4273 = 12'h471 == _T_71[11:0] ? image_1137 : _GEN_4272; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4274 = 12'h472 == _T_71[11:0] ? image_1138 : _GEN_4273; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4275 = 12'h473 == _T_71[11:0] ? image_1139 : _GEN_4274; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4276 = 12'h474 == _T_71[11:0] ? image_1140 : _GEN_4275; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4277 = 12'h475 == _T_71[11:0] ? image_1141 : _GEN_4276; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4278 = 12'h476 == _T_71[11:0] ? image_1142 : _GEN_4277; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4279 = 12'h477 == _T_71[11:0] ? image_1143 : _GEN_4278; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4280 = 12'h478 == _T_71[11:0] ? image_1144 : _GEN_4279; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4281 = 12'h479 == _T_71[11:0] ? image_1145 : _GEN_4280; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4282 = 12'h47a == _T_71[11:0] ? image_1146 : _GEN_4281; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4283 = 12'h47b == _T_71[11:0] ? image_1147 : _GEN_4282; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4284 = 12'h47c == _T_71[11:0] ? image_1148 : _GEN_4283; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4285 = 12'h47d == _T_71[11:0] ? 4'h0 : _GEN_4284; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4286 = 12'h47e == _T_71[11:0] ? 4'h0 : _GEN_4285; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4287 = 12'h47f == _T_71[11:0] ? 4'h0 : _GEN_4286; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4288 = 12'h480 == _T_71[11:0] ? image_1152 : _GEN_4287; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4289 = 12'h481 == _T_71[11:0] ? image_1153 : _GEN_4288; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4290 = 12'h482 == _T_71[11:0] ? image_1154 : _GEN_4289; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4291 = 12'h483 == _T_71[11:0] ? image_1155 : _GEN_4290; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4292 = 12'h484 == _T_71[11:0] ? image_1156 : _GEN_4291; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4293 = 12'h485 == _T_71[11:0] ? image_1157 : _GEN_4292; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4294 = 12'h486 == _T_71[11:0] ? image_1158 : _GEN_4293; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4295 = 12'h487 == _T_71[11:0] ? image_1159 : _GEN_4294; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4296 = 12'h488 == _T_71[11:0] ? image_1160 : _GEN_4295; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4297 = 12'h489 == _T_71[11:0] ? image_1161 : _GEN_4296; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4298 = 12'h48a == _T_71[11:0] ? image_1162 : _GEN_4297; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4299 = 12'h48b == _T_71[11:0] ? image_1163 : _GEN_4298; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4300 = 12'h48c == _T_71[11:0] ? image_1164 : _GEN_4299; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4301 = 12'h48d == _T_71[11:0] ? image_1165 : _GEN_4300; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4302 = 12'h48e == _T_71[11:0] ? image_1166 : _GEN_4301; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4303 = 12'h48f == _T_71[11:0] ? image_1167 : _GEN_4302; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4304 = 12'h490 == _T_71[11:0] ? image_1168 : _GEN_4303; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4305 = 12'h491 == _T_71[11:0] ? image_1169 : _GEN_4304; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4306 = 12'h492 == _T_71[11:0] ? image_1170 : _GEN_4305; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4307 = 12'h493 == _T_71[11:0] ? image_1171 : _GEN_4306; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4308 = 12'h494 == _T_71[11:0] ? image_1172 : _GEN_4307; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4309 = 12'h495 == _T_71[11:0] ? image_1173 : _GEN_4308; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4310 = 12'h496 == _T_71[11:0] ? image_1174 : _GEN_4309; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4311 = 12'h497 == _T_71[11:0] ? image_1175 : _GEN_4310; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4312 = 12'h498 == _T_71[11:0] ? image_1176 : _GEN_4311; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4313 = 12'h499 == _T_71[11:0] ? image_1177 : _GEN_4312; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4314 = 12'h49a == _T_71[11:0] ? image_1178 : _GEN_4313; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4315 = 12'h49b == _T_71[11:0] ? image_1179 : _GEN_4314; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4316 = 12'h49c == _T_71[11:0] ? image_1180 : _GEN_4315; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4317 = 12'h49d == _T_71[11:0] ? image_1181 : _GEN_4316; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4318 = 12'h49e == _T_71[11:0] ? image_1182 : _GEN_4317; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4319 = 12'h49f == _T_71[11:0] ? image_1183 : _GEN_4318; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4320 = 12'h4a0 == _T_71[11:0] ? image_1184 : _GEN_4319; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4321 = 12'h4a1 == _T_71[11:0] ? image_1185 : _GEN_4320; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4322 = 12'h4a2 == _T_71[11:0] ? image_1186 : _GEN_4321; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4323 = 12'h4a3 == _T_71[11:0] ? image_1187 : _GEN_4322; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4324 = 12'h4a4 == _T_71[11:0] ? image_1188 : _GEN_4323; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4325 = 12'h4a5 == _T_71[11:0] ? image_1189 : _GEN_4324; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4326 = 12'h4a6 == _T_71[11:0] ? image_1190 : _GEN_4325; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4327 = 12'h4a7 == _T_71[11:0] ? image_1191 : _GEN_4326; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4328 = 12'h4a8 == _T_71[11:0] ? image_1192 : _GEN_4327; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4329 = 12'h4a9 == _T_71[11:0] ? image_1193 : _GEN_4328; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4330 = 12'h4aa == _T_71[11:0] ? image_1194 : _GEN_4329; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4331 = 12'h4ab == _T_71[11:0] ? image_1195 : _GEN_4330; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4332 = 12'h4ac == _T_71[11:0] ? image_1196 : _GEN_4331; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4333 = 12'h4ad == _T_71[11:0] ? image_1197 : _GEN_4332; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4334 = 12'h4ae == _T_71[11:0] ? image_1198 : _GEN_4333; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4335 = 12'h4af == _T_71[11:0] ? image_1199 : _GEN_4334; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4336 = 12'h4b0 == _T_71[11:0] ? image_1200 : _GEN_4335; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4337 = 12'h4b1 == _T_71[11:0] ? image_1201 : _GEN_4336; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4338 = 12'h4b2 == _T_71[11:0] ? image_1202 : _GEN_4337; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4339 = 12'h4b3 == _T_71[11:0] ? image_1203 : _GEN_4338; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4340 = 12'h4b4 == _T_71[11:0] ? image_1204 : _GEN_4339; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4341 = 12'h4b5 == _T_71[11:0] ? image_1205 : _GEN_4340; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4342 = 12'h4b6 == _T_71[11:0] ? image_1206 : _GEN_4341; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4343 = 12'h4b7 == _T_71[11:0] ? image_1207 : _GEN_4342; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4344 = 12'h4b8 == _T_71[11:0] ? image_1208 : _GEN_4343; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4345 = 12'h4b9 == _T_71[11:0] ? 4'h0 : _GEN_4344; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4346 = 12'h4ba == _T_71[11:0] ? 4'h0 : _GEN_4345; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4347 = 12'h4bb == _T_71[11:0] ? 4'h0 : _GEN_4346; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4348 = 12'h4bc == _T_71[11:0] ? 4'h0 : _GEN_4347; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4349 = 12'h4bd == _T_71[11:0] ? 4'h0 : _GEN_4348; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4350 = 12'h4be == _T_71[11:0] ? 4'h0 : _GEN_4349; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4351 = 12'h4bf == _T_71[11:0] ? 4'h0 : _GEN_4350; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4352 = 12'h4c0 == _T_71[11:0] ? image_1216 : _GEN_4351; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4353 = 12'h4c1 == _T_71[11:0] ? image_1217 : _GEN_4352; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4354 = 12'h4c2 == _T_71[11:0] ? image_1218 : _GEN_4353; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4355 = 12'h4c3 == _T_71[11:0] ? image_1219 : _GEN_4354; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4356 = 12'h4c4 == _T_71[11:0] ? image_1220 : _GEN_4355; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4357 = 12'h4c5 == _T_71[11:0] ? image_1221 : _GEN_4356; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4358 = 12'h4c6 == _T_71[11:0] ? image_1222 : _GEN_4357; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4359 = 12'h4c7 == _T_71[11:0] ? image_1223 : _GEN_4358; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4360 = 12'h4c8 == _T_71[11:0] ? image_1224 : _GEN_4359; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4361 = 12'h4c9 == _T_71[11:0] ? image_1225 : _GEN_4360; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4362 = 12'h4ca == _T_71[11:0] ? image_1226 : _GEN_4361; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4363 = 12'h4cb == _T_71[11:0] ? image_1227 : _GEN_4362; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4364 = 12'h4cc == _T_71[11:0] ? image_1228 : _GEN_4363; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4365 = 12'h4cd == _T_71[11:0] ? image_1229 : _GEN_4364; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4366 = 12'h4ce == _T_71[11:0] ? image_1230 : _GEN_4365; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4367 = 12'h4cf == _T_71[11:0] ? image_1231 : _GEN_4366; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4368 = 12'h4d0 == _T_71[11:0] ? image_1232 : _GEN_4367; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4369 = 12'h4d1 == _T_71[11:0] ? image_1233 : _GEN_4368; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4370 = 12'h4d2 == _T_71[11:0] ? image_1234 : _GEN_4369; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4371 = 12'h4d3 == _T_71[11:0] ? image_1235 : _GEN_4370; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4372 = 12'h4d4 == _T_71[11:0] ? image_1236 : _GEN_4371; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4373 = 12'h4d5 == _T_71[11:0] ? image_1237 : _GEN_4372; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4374 = 12'h4d6 == _T_71[11:0] ? image_1238 : _GEN_4373; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4375 = 12'h4d7 == _T_71[11:0] ? image_1239 : _GEN_4374; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4376 = 12'h4d8 == _T_71[11:0] ? image_1240 : _GEN_4375; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4377 = 12'h4d9 == _T_71[11:0] ? image_1241 : _GEN_4376; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4378 = 12'h4da == _T_71[11:0] ? image_1242 : _GEN_4377; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4379 = 12'h4db == _T_71[11:0] ? image_1243 : _GEN_4378; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4380 = 12'h4dc == _T_71[11:0] ? image_1244 : _GEN_4379; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4381 = 12'h4dd == _T_71[11:0] ? image_1245 : _GEN_4380; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4382 = 12'h4de == _T_71[11:0] ? image_1246 : _GEN_4381; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4383 = 12'h4df == _T_71[11:0] ? image_1247 : _GEN_4382; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4384 = 12'h4e0 == _T_71[11:0] ? image_1248 : _GEN_4383; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4385 = 12'h4e1 == _T_71[11:0] ? image_1249 : _GEN_4384; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4386 = 12'h4e2 == _T_71[11:0] ? image_1250 : _GEN_4385; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4387 = 12'h4e3 == _T_71[11:0] ? image_1251 : _GEN_4386; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4388 = 12'h4e4 == _T_71[11:0] ? image_1252 : _GEN_4387; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4389 = 12'h4e5 == _T_71[11:0] ? image_1253 : _GEN_4388; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4390 = 12'h4e6 == _T_71[11:0] ? image_1254 : _GEN_4389; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4391 = 12'h4e7 == _T_71[11:0] ? image_1255 : _GEN_4390; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4392 = 12'h4e8 == _T_71[11:0] ? image_1256 : _GEN_4391; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4393 = 12'h4e9 == _T_71[11:0] ? image_1257 : _GEN_4392; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4394 = 12'h4ea == _T_71[11:0] ? image_1258 : _GEN_4393; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4395 = 12'h4eb == _T_71[11:0] ? image_1259 : _GEN_4394; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4396 = 12'h4ec == _T_71[11:0] ? image_1260 : _GEN_4395; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4397 = 12'h4ed == _T_71[11:0] ? image_1261 : _GEN_4396; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4398 = 12'h4ee == _T_71[11:0] ? image_1262 : _GEN_4397; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4399 = 12'h4ef == _T_71[11:0] ? image_1263 : _GEN_4398; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4400 = 12'h4f0 == _T_71[11:0] ? image_1264 : _GEN_4399; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4401 = 12'h4f1 == _T_71[11:0] ? image_1265 : _GEN_4400; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4402 = 12'h4f2 == _T_71[11:0] ? image_1266 : _GEN_4401; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4403 = 12'h4f3 == _T_71[11:0] ? image_1267 : _GEN_4402; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4404 = 12'h4f4 == _T_71[11:0] ? image_1268 : _GEN_4403; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4405 = 12'h4f5 == _T_71[11:0] ? image_1269 : _GEN_4404; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4406 = 12'h4f6 == _T_71[11:0] ? image_1270 : _GEN_4405; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4407 = 12'h4f7 == _T_71[11:0] ? image_1271 : _GEN_4406; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4408 = 12'h4f8 == _T_71[11:0] ? image_1272 : _GEN_4407; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4409 = 12'h4f9 == _T_71[11:0] ? image_1273 : _GEN_4408; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4410 = 12'h4fa == _T_71[11:0] ? image_1274 : _GEN_4409; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4411 = 12'h4fb == _T_71[11:0] ? image_1275 : _GEN_4410; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4412 = 12'h4fc == _T_71[11:0] ? 4'h0 : _GEN_4411; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4413 = 12'h4fd == _T_71[11:0] ? 4'h0 : _GEN_4412; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4414 = 12'h4fe == _T_71[11:0] ? 4'h0 : _GEN_4413; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4415 = 12'h4ff == _T_71[11:0] ? 4'h0 : _GEN_4414; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4416 = 12'h500 == _T_71[11:0] ? image_1280 : _GEN_4415; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4417 = 12'h501 == _T_71[11:0] ? image_1281 : _GEN_4416; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4418 = 12'h502 == _T_71[11:0] ? image_1282 : _GEN_4417; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4419 = 12'h503 == _T_71[11:0] ? image_1283 : _GEN_4418; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4420 = 12'h504 == _T_71[11:0] ? image_1284 : _GEN_4419; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4421 = 12'h505 == _T_71[11:0] ? image_1285 : _GEN_4420; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4422 = 12'h506 == _T_71[11:0] ? image_1286 : _GEN_4421; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4423 = 12'h507 == _T_71[11:0] ? image_1287 : _GEN_4422; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4424 = 12'h508 == _T_71[11:0] ? image_1288 : _GEN_4423; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4425 = 12'h509 == _T_71[11:0] ? image_1289 : _GEN_4424; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4426 = 12'h50a == _T_71[11:0] ? image_1290 : _GEN_4425; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4427 = 12'h50b == _T_71[11:0] ? image_1291 : _GEN_4426; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4428 = 12'h50c == _T_71[11:0] ? image_1292 : _GEN_4427; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4429 = 12'h50d == _T_71[11:0] ? image_1293 : _GEN_4428; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4430 = 12'h50e == _T_71[11:0] ? image_1294 : _GEN_4429; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4431 = 12'h50f == _T_71[11:0] ? image_1295 : _GEN_4430; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4432 = 12'h510 == _T_71[11:0] ? image_1296 : _GEN_4431; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4433 = 12'h511 == _T_71[11:0] ? image_1297 : _GEN_4432; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4434 = 12'h512 == _T_71[11:0] ? image_1298 : _GEN_4433; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4435 = 12'h513 == _T_71[11:0] ? image_1299 : _GEN_4434; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4436 = 12'h514 == _T_71[11:0] ? image_1300 : _GEN_4435; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4437 = 12'h515 == _T_71[11:0] ? image_1301 : _GEN_4436; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4438 = 12'h516 == _T_71[11:0] ? image_1302 : _GEN_4437; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4439 = 12'h517 == _T_71[11:0] ? image_1303 : _GEN_4438; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4440 = 12'h518 == _T_71[11:0] ? image_1304 : _GEN_4439; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4441 = 12'h519 == _T_71[11:0] ? image_1305 : _GEN_4440; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4442 = 12'h51a == _T_71[11:0] ? image_1306 : _GEN_4441; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4443 = 12'h51b == _T_71[11:0] ? image_1307 : _GEN_4442; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4444 = 12'h51c == _T_71[11:0] ? image_1308 : _GEN_4443; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4445 = 12'h51d == _T_71[11:0] ? image_1309 : _GEN_4444; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4446 = 12'h51e == _T_71[11:0] ? image_1310 : _GEN_4445; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4447 = 12'h51f == _T_71[11:0] ? image_1311 : _GEN_4446; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4448 = 12'h520 == _T_71[11:0] ? image_1312 : _GEN_4447; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4449 = 12'h521 == _T_71[11:0] ? image_1313 : _GEN_4448; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4450 = 12'h522 == _T_71[11:0] ? image_1314 : _GEN_4449; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4451 = 12'h523 == _T_71[11:0] ? image_1315 : _GEN_4450; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4452 = 12'h524 == _T_71[11:0] ? image_1316 : _GEN_4451; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4453 = 12'h525 == _T_71[11:0] ? image_1317 : _GEN_4452; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4454 = 12'h526 == _T_71[11:0] ? image_1318 : _GEN_4453; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4455 = 12'h527 == _T_71[11:0] ? image_1319 : _GEN_4454; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4456 = 12'h528 == _T_71[11:0] ? image_1320 : _GEN_4455; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4457 = 12'h529 == _T_71[11:0] ? image_1321 : _GEN_4456; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4458 = 12'h52a == _T_71[11:0] ? image_1322 : _GEN_4457; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4459 = 12'h52b == _T_71[11:0] ? image_1323 : _GEN_4458; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4460 = 12'h52c == _T_71[11:0] ? image_1324 : _GEN_4459; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4461 = 12'h52d == _T_71[11:0] ? image_1325 : _GEN_4460; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4462 = 12'h52e == _T_71[11:0] ? image_1326 : _GEN_4461; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4463 = 12'h52f == _T_71[11:0] ? image_1327 : _GEN_4462; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4464 = 12'h530 == _T_71[11:0] ? image_1328 : _GEN_4463; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4465 = 12'h531 == _T_71[11:0] ? image_1329 : _GEN_4464; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4466 = 12'h532 == _T_71[11:0] ? image_1330 : _GEN_4465; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4467 = 12'h533 == _T_71[11:0] ? image_1331 : _GEN_4466; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4468 = 12'h534 == _T_71[11:0] ? image_1332 : _GEN_4467; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4469 = 12'h535 == _T_71[11:0] ? image_1333 : _GEN_4468; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4470 = 12'h536 == _T_71[11:0] ? image_1334 : _GEN_4469; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4471 = 12'h537 == _T_71[11:0] ? image_1335 : _GEN_4470; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4472 = 12'h538 == _T_71[11:0] ? image_1336 : _GEN_4471; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4473 = 12'h539 == _T_71[11:0] ? image_1337 : _GEN_4472; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4474 = 12'h53a == _T_71[11:0] ? image_1338 : _GEN_4473; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4475 = 12'h53b == _T_71[11:0] ? image_1339 : _GEN_4474; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4476 = 12'h53c == _T_71[11:0] ? image_1340 : _GEN_4475; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4477 = 12'h53d == _T_71[11:0] ? image_1341 : _GEN_4476; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4478 = 12'h53e == _T_71[11:0] ? 4'h0 : _GEN_4477; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4479 = 12'h53f == _T_71[11:0] ? 4'h0 : _GEN_4478; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4480 = 12'h540 == _T_71[11:0] ? image_1344 : _GEN_4479; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4481 = 12'h541 == _T_71[11:0] ? image_1345 : _GEN_4480; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4482 = 12'h542 == _T_71[11:0] ? image_1346 : _GEN_4481; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4483 = 12'h543 == _T_71[11:0] ? image_1347 : _GEN_4482; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4484 = 12'h544 == _T_71[11:0] ? image_1348 : _GEN_4483; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4485 = 12'h545 == _T_71[11:0] ? image_1349 : _GEN_4484; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4486 = 12'h546 == _T_71[11:0] ? image_1350 : _GEN_4485; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4487 = 12'h547 == _T_71[11:0] ? image_1351 : _GEN_4486; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4488 = 12'h548 == _T_71[11:0] ? image_1352 : _GEN_4487; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4489 = 12'h549 == _T_71[11:0] ? image_1353 : _GEN_4488; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4490 = 12'h54a == _T_71[11:0] ? image_1354 : _GEN_4489; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4491 = 12'h54b == _T_71[11:0] ? image_1355 : _GEN_4490; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4492 = 12'h54c == _T_71[11:0] ? image_1356 : _GEN_4491; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4493 = 12'h54d == _T_71[11:0] ? image_1357 : _GEN_4492; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4494 = 12'h54e == _T_71[11:0] ? image_1358 : _GEN_4493; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4495 = 12'h54f == _T_71[11:0] ? image_1359 : _GEN_4494; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4496 = 12'h550 == _T_71[11:0] ? image_1360 : _GEN_4495; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4497 = 12'h551 == _T_71[11:0] ? image_1361 : _GEN_4496; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4498 = 12'h552 == _T_71[11:0] ? image_1362 : _GEN_4497; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4499 = 12'h553 == _T_71[11:0] ? image_1363 : _GEN_4498; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4500 = 12'h554 == _T_71[11:0] ? image_1364 : _GEN_4499; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4501 = 12'h555 == _T_71[11:0] ? image_1365 : _GEN_4500; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4502 = 12'h556 == _T_71[11:0] ? image_1366 : _GEN_4501; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4503 = 12'h557 == _T_71[11:0] ? image_1367 : _GEN_4502; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4504 = 12'h558 == _T_71[11:0] ? image_1368 : _GEN_4503; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4505 = 12'h559 == _T_71[11:0] ? image_1369 : _GEN_4504; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4506 = 12'h55a == _T_71[11:0] ? image_1370 : _GEN_4505; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4507 = 12'h55b == _T_71[11:0] ? image_1371 : _GEN_4506; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4508 = 12'h55c == _T_71[11:0] ? image_1372 : _GEN_4507; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4509 = 12'h55d == _T_71[11:0] ? image_1373 : _GEN_4508; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4510 = 12'h55e == _T_71[11:0] ? image_1374 : _GEN_4509; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4511 = 12'h55f == _T_71[11:0] ? image_1375 : _GEN_4510; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4512 = 12'h560 == _T_71[11:0] ? image_1376 : _GEN_4511; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4513 = 12'h561 == _T_71[11:0] ? image_1377 : _GEN_4512; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4514 = 12'h562 == _T_71[11:0] ? image_1378 : _GEN_4513; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4515 = 12'h563 == _T_71[11:0] ? image_1379 : _GEN_4514; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4516 = 12'h564 == _T_71[11:0] ? image_1380 : _GEN_4515; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4517 = 12'h565 == _T_71[11:0] ? image_1381 : _GEN_4516; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4518 = 12'h566 == _T_71[11:0] ? image_1382 : _GEN_4517; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4519 = 12'h567 == _T_71[11:0] ? image_1383 : _GEN_4518; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4520 = 12'h568 == _T_71[11:0] ? image_1384 : _GEN_4519; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4521 = 12'h569 == _T_71[11:0] ? image_1385 : _GEN_4520; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4522 = 12'h56a == _T_71[11:0] ? image_1386 : _GEN_4521; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4523 = 12'h56b == _T_71[11:0] ? image_1387 : _GEN_4522; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4524 = 12'h56c == _T_71[11:0] ? image_1388 : _GEN_4523; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4525 = 12'h56d == _T_71[11:0] ? image_1389 : _GEN_4524; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4526 = 12'h56e == _T_71[11:0] ? image_1390 : _GEN_4525; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4527 = 12'h56f == _T_71[11:0] ? image_1391 : _GEN_4526; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4528 = 12'h570 == _T_71[11:0] ? image_1392 : _GEN_4527; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4529 = 12'h571 == _T_71[11:0] ? image_1393 : _GEN_4528; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4530 = 12'h572 == _T_71[11:0] ? image_1394 : _GEN_4529; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4531 = 12'h573 == _T_71[11:0] ? image_1395 : _GEN_4530; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4532 = 12'h574 == _T_71[11:0] ? image_1396 : _GEN_4531; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4533 = 12'h575 == _T_71[11:0] ? image_1397 : _GEN_4532; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4534 = 12'h576 == _T_71[11:0] ? image_1398 : _GEN_4533; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4535 = 12'h577 == _T_71[11:0] ? image_1399 : _GEN_4534; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4536 = 12'h578 == _T_71[11:0] ? image_1400 : _GEN_4535; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4537 = 12'h579 == _T_71[11:0] ? image_1401 : _GEN_4536; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4538 = 12'h57a == _T_71[11:0] ? image_1402 : _GEN_4537; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4539 = 12'h57b == _T_71[11:0] ? image_1403 : _GEN_4538; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4540 = 12'h57c == _T_71[11:0] ? image_1404 : _GEN_4539; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4541 = 12'h57d == _T_71[11:0] ? image_1405 : _GEN_4540; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4542 = 12'h57e == _T_71[11:0] ? 4'h0 : _GEN_4541; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4543 = 12'h57f == _T_71[11:0] ? 4'h0 : _GEN_4542; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4544 = 12'h580 == _T_71[11:0] ? image_1408 : _GEN_4543; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4545 = 12'h581 == _T_71[11:0] ? image_1409 : _GEN_4544; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4546 = 12'h582 == _T_71[11:0] ? image_1410 : _GEN_4545; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4547 = 12'h583 == _T_71[11:0] ? image_1411 : _GEN_4546; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4548 = 12'h584 == _T_71[11:0] ? image_1412 : _GEN_4547; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4549 = 12'h585 == _T_71[11:0] ? image_1413 : _GEN_4548; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4550 = 12'h586 == _T_71[11:0] ? image_1414 : _GEN_4549; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4551 = 12'h587 == _T_71[11:0] ? image_1415 : _GEN_4550; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4552 = 12'h588 == _T_71[11:0] ? image_1416 : _GEN_4551; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4553 = 12'h589 == _T_71[11:0] ? image_1417 : _GEN_4552; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4554 = 12'h58a == _T_71[11:0] ? image_1418 : _GEN_4553; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4555 = 12'h58b == _T_71[11:0] ? image_1419 : _GEN_4554; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4556 = 12'h58c == _T_71[11:0] ? image_1420 : _GEN_4555; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4557 = 12'h58d == _T_71[11:0] ? image_1421 : _GEN_4556; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4558 = 12'h58e == _T_71[11:0] ? image_1422 : _GEN_4557; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4559 = 12'h58f == _T_71[11:0] ? image_1423 : _GEN_4558; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4560 = 12'h590 == _T_71[11:0] ? image_1424 : _GEN_4559; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4561 = 12'h591 == _T_71[11:0] ? image_1425 : _GEN_4560; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4562 = 12'h592 == _T_71[11:0] ? image_1426 : _GEN_4561; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4563 = 12'h593 == _T_71[11:0] ? image_1427 : _GEN_4562; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4564 = 12'h594 == _T_71[11:0] ? image_1428 : _GEN_4563; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4565 = 12'h595 == _T_71[11:0] ? image_1429 : _GEN_4564; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4566 = 12'h596 == _T_71[11:0] ? image_1430 : _GEN_4565; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4567 = 12'h597 == _T_71[11:0] ? image_1431 : _GEN_4566; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4568 = 12'h598 == _T_71[11:0] ? image_1432 : _GEN_4567; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4569 = 12'h599 == _T_71[11:0] ? image_1433 : _GEN_4568; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4570 = 12'h59a == _T_71[11:0] ? image_1434 : _GEN_4569; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4571 = 12'h59b == _T_71[11:0] ? image_1435 : _GEN_4570; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4572 = 12'h59c == _T_71[11:0] ? image_1436 : _GEN_4571; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4573 = 12'h59d == _T_71[11:0] ? image_1437 : _GEN_4572; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4574 = 12'h59e == _T_71[11:0] ? image_1438 : _GEN_4573; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4575 = 12'h59f == _T_71[11:0] ? image_1439 : _GEN_4574; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4576 = 12'h5a0 == _T_71[11:0] ? image_1440 : _GEN_4575; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4577 = 12'h5a1 == _T_71[11:0] ? image_1441 : _GEN_4576; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4578 = 12'h5a2 == _T_71[11:0] ? image_1442 : _GEN_4577; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4579 = 12'h5a3 == _T_71[11:0] ? image_1443 : _GEN_4578; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4580 = 12'h5a4 == _T_71[11:0] ? image_1444 : _GEN_4579; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4581 = 12'h5a5 == _T_71[11:0] ? image_1445 : _GEN_4580; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4582 = 12'h5a6 == _T_71[11:0] ? image_1446 : _GEN_4581; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4583 = 12'h5a7 == _T_71[11:0] ? image_1447 : _GEN_4582; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4584 = 12'h5a8 == _T_71[11:0] ? image_1448 : _GEN_4583; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4585 = 12'h5a9 == _T_71[11:0] ? image_1449 : _GEN_4584; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4586 = 12'h5aa == _T_71[11:0] ? image_1450 : _GEN_4585; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4587 = 12'h5ab == _T_71[11:0] ? image_1451 : _GEN_4586; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4588 = 12'h5ac == _T_71[11:0] ? image_1452 : _GEN_4587; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4589 = 12'h5ad == _T_71[11:0] ? image_1453 : _GEN_4588; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4590 = 12'h5ae == _T_71[11:0] ? image_1454 : _GEN_4589; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4591 = 12'h5af == _T_71[11:0] ? image_1455 : _GEN_4590; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4592 = 12'h5b0 == _T_71[11:0] ? image_1456 : _GEN_4591; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4593 = 12'h5b1 == _T_71[11:0] ? image_1457 : _GEN_4592; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4594 = 12'h5b2 == _T_71[11:0] ? image_1458 : _GEN_4593; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4595 = 12'h5b3 == _T_71[11:0] ? image_1459 : _GEN_4594; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4596 = 12'h5b4 == _T_71[11:0] ? image_1460 : _GEN_4595; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4597 = 12'h5b5 == _T_71[11:0] ? image_1461 : _GEN_4596; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4598 = 12'h5b6 == _T_71[11:0] ? image_1462 : _GEN_4597; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4599 = 12'h5b7 == _T_71[11:0] ? image_1463 : _GEN_4598; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4600 = 12'h5b8 == _T_71[11:0] ? image_1464 : _GEN_4599; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4601 = 12'h5b9 == _T_71[11:0] ? image_1465 : _GEN_4600; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4602 = 12'h5ba == _T_71[11:0] ? image_1466 : _GEN_4601; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4603 = 12'h5bb == _T_71[11:0] ? image_1467 : _GEN_4602; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4604 = 12'h5bc == _T_71[11:0] ? image_1468 : _GEN_4603; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4605 = 12'h5bd == _T_71[11:0] ? image_1469 : _GEN_4604; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4606 = 12'h5be == _T_71[11:0] ? 4'h0 : _GEN_4605; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4607 = 12'h5bf == _T_71[11:0] ? 4'h0 : _GEN_4606; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4608 = 12'h5c0 == _T_71[11:0] ? image_1472 : _GEN_4607; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4609 = 12'h5c1 == _T_71[11:0] ? image_1473 : _GEN_4608; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4610 = 12'h5c2 == _T_71[11:0] ? image_1474 : _GEN_4609; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4611 = 12'h5c3 == _T_71[11:0] ? image_1475 : _GEN_4610; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4612 = 12'h5c4 == _T_71[11:0] ? image_1476 : _GEN_4611; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4613 = 12'h5c5 == _T_71[11:0] ? image_1477 : _GEN_4612; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4614 = 12'h5c6 == _T_71[11:0] ? image_1478 : _GEN_4613; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4615 = 12'h5c7 == _T_71[11:0] ? image_1479 : _GEN_4614; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4616 = 12'h5c8 == _T_71[11:0] ? image_1480 : _GEN_4615; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4617 = 12'h5c9 == _T_71[11:0] ? image_1481 : _GEN_4616; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4618 = 12'h5ca == _T_71[11:0] ? image_1482 : _GEN_4617; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4619 = 12'h5cb == _T_71[11:0] ? image_1483 : _GEN_4618; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4620 = 12'h5cc == _T_71[11:0] ? image_1484 : _GEN_4619; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4621 = 12'h5cd == _T_71[11:0] ? image_1485 : _GEN_4620; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4622 = 12'h5ce == _T_71[11:0] ? image_1486 : _GEN_4621; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4623 = 12'h5cf == _T_71[11:0] ? image_1487 : _GEN_4622; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4624 = 12'h5d0 == _T_71[11:0] ? image_1488 : _GEN_4623; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4625 = 12'h5d1 == _T_71[11:0] ? image_1489 : _GEN_4624; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4626 = 12'h5d2 == _T_71[11:0] ? image_1490 : _GEN_4625; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4627 = 12'h5d3 == _T_71[11:0] ? image_1491 : _GEN_4626; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4628 = 12'h5d4 == _T_71[11:0] ? image_1492 : _GEN_4627; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4629 = 12'h5d5 == _T_71[11:0] ? image_1493 : _GEN_4628; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4630 = 12'h5d6 == _T_71[11:0] ? image_1494 : _GEN_4629; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4631 = 12'h5d7 == _T_71[11:0] ? image_1495 : _GEN_4630; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4632 = 12'h5d8 == _T_71[11:0] ? image_1496 : _GEN_4631; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4633 = 12'h5d9 == _T_71[11:0] ? image_1497 : _GEN_4632; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4634 = 12'h5da == _T_71[11:0] ? image_1498 : _GEN_4633; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4635 = 12'h5db == _T_71[11:0] ? image_1499 : _GEN_4634; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4636 = 12'h5dc == _T_71[11:0] ? image_1500 : _GEN_4635; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4637 = 12'h5dd == _T_71[11:0] ? image_1501 : _GEN_4636; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4638 = 12'h5de == _T_71[11:0] ? image_1502 : _GEN_4637; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4639 = 12'h5df == _T_71[11:0] ? image_1503 : _GEN_4638; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4640 = 12'h5e0 == _T_71[11:0] ? image_1504 : _GEN_4639; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4641 = 12'h5e1 == _T_71[11:0] ? image_1505 : _GEN_4640; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4642 = 12'h5e2 == _T_71[11:0] ? image_1506 : _GEN_4641; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4643 = 12'h5e3 == _T_71[11:0] ? image_1507 : _GEN_4642; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4644 = 12'h5e4 == _T_71[11:0] ? image_1508 : _GEN_4643; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4645 = 12'h5e5 == _T_71[11:0] ? image_1509 : _GEN_4644; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4646 = 12'h5e6 == _T_71[11:0] ? image_1510 : _GEN_4645; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4647 = 12'h5e7 == _T_71[11:0] ? image_1511 : _GEN_4646; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4648 = 12'h5e8 == _T_71[11:0] ? image_1512 : _GEN_4647; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4649 = 12'h5e9 == _T_71[11:0] ? image_1513 : _GEN_4648; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4650 = 12'h5ea == _T_71[11:0] ? image_1514 : _GEN_4649; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4651 = 12'h5eb == _T_71[11:0] ? image_1515 : _GEN_4650; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4652 = 12'h5ec == _T_71[11:0] ? image_1516 : _GEN_4651; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4653 = 12'h5ed == _T_71[11:0] ? image_1517 : _GEN_4652; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4654 = 12'h5ee == _T_71[11:0] ? image_1518 : _GEN_4653; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4655 = 12'h5ef == _T_71[11:0] ? image_1519 : _GEN_4654; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4656 = 12'h5f0 == _T_71[11:0] ? image_1520 : _GEN_4655; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4657 = 12'h5f1 == _T_71[11:0] ? image_1521 : _GEN_4656; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4658 = 12'h5f2 == _T_71[11:0] ? image_1522 : _GEN_4657; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4659 = 12'h5f3 == _T_71[11:0] ? image_1523 : _GEN_4658; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4660 = 12'h5f4 == _T_71[11:0] ? image_1524 : _GEN_4659; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4661 = 12'h5f5 == _T_71[11:0] ? image_1525 : _GEN_4660; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4662 = 12'h5f6 == _T_71[11:0] ? image_1526 : _GEN_4661; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4663 = 12'h5f7 == _T_71[11:0] ? image_1527 : _GEN_4662; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4664 = 12'h5f8 == _T_71[11:0] ? image_1528 : _GEN_4663; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4665 = 12'h5f9 == _T_71[11:0] ? image_1529 : _GEN_4664; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4666 = 12'h5fa == _T_71[11:0] ? image_1530 : _GEN_4665; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4667 = 12'h5fb == _T_71[11:0] ? image_1531 : _GEN_4666; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4668 = 12'h5fc == _T_71[11:0] ? image_1532 : _GEN_4667; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4669 = 12'h5fd == _T_71[11:0] ? image_1533 : _GEN_4668; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4670 = 12'h5fe == _T_71[11:0] ? 4'h0 : _GEN_4669; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4671 = 12'h5ff == _T_71[11:0] ? 4'h0 : _GEN_4670; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4672 = 12'h600 == _T_71[11:0] ? image_1536 : _GEN_4671; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4673 = 12'h601 == _T_71[11:0] ? image_1537 : _GEN_4672; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4674 = 12'h602 == _T_71[11:0] ? image_1538 : _GEN_4673; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4675 = 12'h603 == _T_71[11:0] ? image_1539 : _GEN_4674; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4676 = 12'h604 == _T_71[11:0] ? image_1540 : _GEN_4675; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4677 = 12'h605 == _T_71[11:0] ? image_1541 : _GEN_4676; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4678 = 12'h606 == _T_71[11:0] ? image_1542 : _GEN_4677; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4679 = 12'h607 == _T_71[11:0] ? image_1543 : _GEN_4678; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4680 = 12'h608 == _T_71[11:0] ? image_1544 : _GEN_4679; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4681 = 12'h609 == _T_71[11:0] ? image_1545 : _GEN_4680; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4682 = 12'h60a == _T_71[11:0] ? image_1546 : _GEN_4681; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4683 = 12'h60b == _T_71[11:0] ? image_1547 : _GEN_4682; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4684 = 12'h60c == _T_71[11:0] ? image_1548 : _GEN_4683; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4685 = 12'h60d == _T_71[11:0] ? image_1549 : _GEN_4684; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4686 = 12'h60e == _T_71[11:0] ? image_1550 : _GEN_4685; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4687 = 12'h60f == _T_71[11:0] ? image_1551 : _GEN_4686; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4688 = 12'h610 == _T_71[11:0] ? image_1552 : _GEN_4687; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4689 = 12'h611 == _T_71[11:0] ? image_1553 : _GEN_4688; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4690 = 12'h612 == _T_71[11:0] ? image_1554 : _GEN_4689; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4691 = 12'h613 == _T_71[11:0] ? image_1555 : _GEN_4690; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4692 = 12'h614 == _T_71[11:0] ? image_1556 : _GEN_4691; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4693 = 12'h615 == _T_71[11:0] ? image_1557 : _GEN_4692; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4694 = 12'h616 == _T_71[11:0] ? image_1558 : _GEN_4693; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4695 = 12'h617 == _T_71[11:0] ? image_1559 : _GEN_4694; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4696 = 12'h618 == _T_71[11:0] ? image_1560 : _GEN_4695; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4697 = 12'h619 == _T_71[11:0] ? image_1561 : _GEN_4696; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4698 = 12'h61a == _T_71[11:0] ? image_1562 : _GEN_4697; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4699 = 12'h61b == _T_71[11:0] ? image_1563 : _GEN_4698; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4700 = 12'h61c == _T_71[11:0] ? image_1564 : _GEN_4699; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4701 = 12'h61d == _T_71[11:0] ? image_1565 : _GEN_4700; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4702 = 12'h61e == _T_71[11:0] ? image_1566 : _GEN_4701; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4703 = 12'h61f == _T_71[11:0] ? image_1567 : _GEN_4702; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4704 = 12'h620 == _T_71[11:0] ? image_1568 : _GEN_4703; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4705 = 12'h621 == _T_71[11:0] ? image_1569 : _GEN_4704; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4706 = 12'h622 == _T_71[11:0] ? image_1570 : _GEN_4705; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4707 = 12'h623 == _T_71[11:0] ? image_1571 : _GEN_4706; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4708 = 12'h624 == _T_71[11:0] ? image_1572 : _GEN_4707; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4709 = 12'h625 == _T_71[11:0] ? image_1573 : _GEN_4708; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4710 = 12'h626 == _T_71[11:0] ? image_1574 : _GEN_4709; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4711 = 12'h627 == _T_71[11:0] ? image_1575 : _GEN_4710; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4712 = 12'h628 == _T_71[11:0] ? image_1576 : _GEN_4711; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4713 = 12'h629 == _T_71[11:0] ? image_1577 : _GEN_4712; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4714 = 12'h62a == _T_71[11:0] ? image_1578 : _GEN_4713; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4715 = 12'h62b == _T_71[11:0] ? image_1579 : _GEN_4714; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4716 = 12'h62c == _T_71[11:0] ? image_1580 : _GEN_4715; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4717 = 12'h62d == _T_71[11:0] ? image_1581 : _GEN_4716; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4718 = 12'h62e == _T_71[11:0] ? image_1582 : _GEN_4717; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4719 = 12'h62f == _T_71[11:0] ? image_1583 : _GEN_4718; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4720 = 12'h630 == _T_71[11:0] ? image_1584 : _GEN_4719; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4721 = 12'h631 == _T_71[11:0] ? image_1585 : _GEN_4720; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4722 = 12'h632 == _T_71[11:0] ? image_1586 : _GEN_4721; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4723 = 12'h633 == _T_71[11:0] ? image_1587 : _GEN_4722; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4724 = 12'h634 == _T_71[11:0] ? image_1588 : _GEN_4723; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4725 = 12'h635 == _T_71[11:0] ? image_1589 : _GEN_4724; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4726 = 12'h636 == _T_71[11:0] ? image_1590 : _GEN_4725; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4727 = 12'h637 == _T_71[11:0] ? image_1591 : _GEN_4726; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4728 = 12'h638 == _T_71[11:0] ? image_1592 : _GEN_4727; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4729 = 12'h639 == _T_71[11:0] ? image_1593 : _GEN_4728; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4730 = 12'h63a == _T_71[11:0] ? image_1594 : _GEN_4729; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4731 = 12'h63b == _T_71[11:0] ? image_1595 : _GEN_4730; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4732 = 12'h63c == _T_71[11:0] ? image_1596 : _GEN_4731; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4733 = 12'h63d == _T_71[11:0] ? image_1597 : _GEN_4732; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4734 = 12'h63e == _T_71[11:0] ? 4'h0 : _GEN_4733; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4735 = 12'h63f == _T_71[11:0] ? 4'h0 : _GEN_4734; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4736 = 12'h640 == _T_71[11:0] ? image_1600 : _GEN_4735; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4737 = 12'h641 == _T_71[11:0] ? image_1601 : _GEN_4736; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4738 = 12'h642 == _T_71[11:0] ? image_1602 : _GEN_4737; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4739 = 12'h643 == _T_71[11:0] ? image_1603 : _GEN_4738; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4740 = 12'h644 == _T_71[11:0] ? image_1604 : _GEN_4739; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4741 = 12'h645 == _T_71[11:0] ? image_1605 : _GEN_4740; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4742 = 12'h646 == _T_71[11:0] ? image_1606 : _GEN_4741; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4743 = 12'h647 == _T_71[11:0] ? image_1607 : _GEN_4742; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4744 = 12'h648 == _T_71[11:0] ? image_1608 : _GEN_4743; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4745 = 12'h649 == _T_71[11:0] ? image_1609 : _GEN_4744; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4746 = 12'h64a == _T_71[11:0] ? image_1610 : _GEN_4745; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4747 = 12'h64b == _T_71[11:0] ? image_1611 : _GEN_4746; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4748 = 12'h64c == _T_71[11:0] ? image_1612 : _GEN_4747; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4749 = 12'h64d == _T_71[11:0] ? image_1613 : _GEN_4748; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4750 = 12'h64e == _T_71[11:0] ? image_1614 : _GEN_4749; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4751 = 12'h64f == _T_71[11:0] ? image_1615 : _GEN_4750; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4752 = 12'h650 == _T_71[11:0] ? image_1616 : _GEN_4751; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4753 = 12'h651 == _T_71[11:0] ? image_1617 : _GEN_4752; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4754 = 12'h652 == _T_71[11:0] ? image_1618 : _GEN_4753; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4755 = 12'h653 == _T_71[11:0] ? image_1619 : _GEN_4754; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4756 = 12'h654 == _T_71[11:0] ? image_1620 : _GEN_4755; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4757 = 12'h655 == _T_71[11:0] ? image_1621 : _GEN_4756; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4758 = 12'h656 == _T_71[11:0] ? image_1622 : _GEN_4757; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4759 = 12'h657 == _T_71[11:0] ? image_1623 : _GEN_4758; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4760 = 12'h658 == _T_71[11:0] ? image_1624 : _GEN_4759; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4761 = 12'h659 == _T_71[11:0] ? image_1625 : _GEN_4760; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4762 = 12'h65a == _T_71[11:0] ? image_1626 : _GEN_4761; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4763 = 12'h65b == _T_71[11:0] ? image_1627 : _GEN_4762; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4764 = 12'h65c == _T_71[11:0] ? image_1628 : _GEN_4763; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4765 = 12'h65d == _T_71[11:0] ? image_1629 : _GEN_4764; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4766 = 12'h65e == _T_71[11:0] ? image_1630 : _GEN_4765; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4767 = 12'h65f == _T_71[11:0] ? image_1631 : _GEN_4766; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4768 = 12'h660 == _T_71[11:0] ? image_1632 : _GEN_4767; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4769 = 12'h661 == _T_71[11:0] ? image_1633 : _GEN_4768; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4770 = 12'h662 == _T_71[11:0] ? image_1634 : _GEN_4769; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4771 = 12'h663 == _T_71[11:0] ? image_1635 : _GEN_4770; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4772 = 12'h664 == _T_71[11:0] ? image_1636 : _GEN_4771; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4773 = 12'h665 == _T_71[11:0] ? image_1637 : _GEN_4772; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4774 = 12'h666 == _T_71[11:0] ? image_1638 : _GEN_4773; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4775 = 12'h667 == _T_71[11:0] ? image_1639 : _GEN_4774; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4776 = 12'h668 == _T_71[11:0] ? image_1640 : _GEN_4775; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4777 = 12'h669 == _T_71[11:0] ? image_1641 : _GEN_4776; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4778 = 12'h66a == _T_71[11:0] ? image_1642 : _GEN_4777; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4779 = 12'h66b == _T_71[11:0] ? image_1643 : _GEN_4778; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4780 = 12'h66c == _T_71[11:0] ? image_1644 : _GEN_4779; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4781 = 12'h66d == _T_71[11:0] ? image_1645 : _GEN_4780; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4782 = 12'h66e == _T_71[11:0] ? image_1646 : _GEN_4781; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4783 = 12'h66f == _T_71[11:0] ? image_1647 : _GEN_4782; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4784 = 12'h670 == _T_71[11:0] ? image_1648 : _GEN_4783; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4785 = 12'h671 == _T_71[11:0] ? image_1649 : _GEN_4784; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4786 = 12'h672 == _T_71[11:0] ? image_1650 : _GEN_4785; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4787 = 12'h673 == _T_71[11:0] ? image_1651 : _GEN_4786; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4788 = 12'h674 == _T_71[11:0] ? image_1652 : _GEN_4787; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4789 = 12'h675 == _T_71[11:0] ? image_1653 : _GEN_4788; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4790 = 12'h676 == _T_71[11:0] ? image_1654 : _GEN_4789; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4791 = 12'h677 == _T_71[11:0] ? image_1655 : _GEN_4790; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4792 = 12'h678 == _T_71[11:0] ? image_1656 : _GEN_4791; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4793 = 12'h679 == _T_71[11:0] ? image_1657 : _GEN_4792; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4794 = 12'h67a == _T_71[11:0] ? image_1658 : _GEN_4793; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4795 = 12'h67b == _T_71[11:0] ? image_1659 : _GEN_4794; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4796 = 12'h67c == _T_71[11:0] ? image_1660 : _GEN_4795; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4797 = 12'h67d == _T_71[11:0] ? 4'h0 : _GEN_4796; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4798 = 12'h67e == _T_71[11:0] ? 4'h0 : _GEN_4797; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4799 = 12'h67f == _T_71[11:0] ? 4'h0 : _GEN_4798; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4800 = 12'h680 == _T_71[11:0] ? image_1664 : _GEN_4799; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4801 = 12'h681 == _T_71[11:0] ? image_1665 : _GEN_4800; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4802 = 12'h682 == _T_71[11:0] ? image_1666 : _GEN_4801; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4803 = 12'h683 == _T_71[11:0] ? image_1667 : _GEN_4802; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4804 = 12'h684 == _T_71[11:0] ? image_1668 : _GEN_4803; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4805 = 12'h685 == _T_71[11:0] ? image_1669 : _GEN_4804; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4806 = 12'h686 == _T_71[11:0] ? image_1670 : _GEN_4805; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4807 = 12'h687 == _T_71[11:0] ? image_1671 : _GEN_4806; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4808 = 12'h688 == _T_71[11:0] ? image_1672 : _GEN_4807; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4809 = 12'h689 == _T_71[11:0] ? image_1673 : _GEN_4808; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4810 = 12'h68a == _T_71[11:0] ? image_1674 : _GEN_4809; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4811 = 12'h68b == _T_71[11:0] ? image_1675 : _GEN_4810; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4812 = 12'h68c == _T_71[11:0] ? image_1676 : _GEN_4811; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4813 = 12'h68d == _T_71[11:0] ? image_1677 : _GEN_4812; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4814 = 12'h68e == _T_71[11:0] ? image_1678 : _GEN_4813; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4815 = 12'h68f == _T_71[11:0] ? image_1679 : _GEN_4814; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4816 = 12'h690 == _T_71[11:0] ? image_1680 : _GEN_4815; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4817 = 12'h691 == _T_71[11:0] ? image_1681 : _GEN_4816; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4818 = 12'h692 == _T_71[11:0] ? image_1682 : _GEN_4817; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4819 = 12'h693 == _T_71[11:0] ? image_1683 : _GEN_4818; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4820 = 12'h694 == _T_71[11:0] ? image_1684 : _GEN_4819; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4821 = 12'h695 == _T_71[11:0] ? image_1685 : _GEN_4820; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4822 = 12'h696 == _T_71[11:0] ? image_1686 : _GEN_4821; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4823 = 12'h697 == _T_71[11:0] ? image_1687 : _GEN_4822; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4824 = 12'h698 == _T_71[11:0] ? image_1688 : _GEN_4823; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4825 = 12'h699 == _T_71[11:0] ? image_1689 : _GEN_4824; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4826 = 12'h69a == _T_71[11:0] ? image_1690 : _GEN_4825; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4827 = 12'h69b == _T_71[11:0] ? image_1691 : _GEN_4826; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4828 = 12'h69c == _T_71[11:0] ? image_1692 : _GEN_4827; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4829 = 12'h69d == _T_71[11:0] ? image_1693 : _GEN_4828; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4830 = 12'h69e == _T_71[11:0] ? image_1694 : _GEN_4829; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4831 = 12'h69f == _T_71[11:0] ? image_1695 : _GEN_4830; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4832 = 12'h6a0 == _T_71[11:0] ? image_1696 : _GEN_4831; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4833 = 12'h6a1 == _T_71[11:0] ? image_1697 : _GEN_4832; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4834 = 12'h6a2 == _T_71[11:0] ? image_1698 : _GEN_4833; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4835 = 12'h6a3 == _T_71[11:0] ? image_1699 : _GEN_4834; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4836 = 12'h6a4 == _T_71[11:0] ? image_1700 : _GEN_4835; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4837 = 12'h6a5 == _T_71[11:0] ? image_1701 : _GEN_4836; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4838 = 12'h6a6 == _T_71[11:0] ? image_1702 : _GEN_4837; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4839 = 12'h6a7 == _T_71[11:0] ? image_1703 : _GEN_4838; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4840 = 12'h6a8 == _T_71[11:0] ? image_1704 : _GEN_4839; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4841 = 12'h6a9 == _T_71[11:0] ? image_1705 : _GEN_4840; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4842 = 12'h6aa == _T_71[11:0] ? image_1706 : _GEN_4841; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4843 = 12'h6ab == _T_71[11:0] ? image_1707 : _GEN_4842; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4844 = 12'h6ac == _T_71[11:0] ? image_1708 : _GEN_4843; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4845 = 12'h6ad == _T_71[11:0] ? image_1709 : _GEN_4844; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4846 = 12'h6ae == _T_71[11:0] ? image_1710 : _GEN_4845; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4847 = 12'h6af == _T_71[11:0] ? image_1711 : _GEN_4846; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4848 = 12'h6b0 == _T_71[11:0] ? image_1712 : _GEN_4847; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4849 = 12'h6b1 == _T_71[11:0] ? image_1713 : _GEN_4848; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4850 = 12'h6b2 == _T_71[11:0] ? image_1714 : _GEN_4849; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4851 = 12'h6b3 == _T_71[11:0] ? image_1715 : _GEN_4850; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4852 = 12'h6b4 == _T_71[11:0] ? image_1716 : _GEN_4851; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4853 = 12'h6b5 == _T_71[11:0] ? image_1717 : _GEN_4852; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4854 = 12'h6b6 == _T_71[11:0] ? image_1718 : _GEN_4853; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4855 = 12'h6b7 == _T_71[11:0] ? image_1719 : _GEN_4854; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4856 = 12'h6b8 == _T_71[11:0] ? image_1720 : _GEN_4855; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4857 = 12'h6b9 == _T_71[11:0] ? image_1721 : _GEN_4856; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4858 = 12'h6ba == _T_71[11:0] ? image_1722 : _GEN_4857; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4859 = 12'h6bb == _T_71[11:0] ? image_1723 : _GEN_4858; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4860 = 12'h6bc == _T_71[11:0] ? 4'h0 : _GEN_4859; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4861 = 12'h6bd == _T_71[11:0] ? 4'h0 : _GEN_4860; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4862 = 12'h6be == _T_71[11:0] ? 4'h0 : _GEN_4861; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4863 = 12'h6bf == _T_71[11:0] ? 4'h0 : _GEN_4862; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4864 = 12'h6c0 == _T_71[11:0] ? image_1728 : _GEN_4863; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4865 = 12'h6c1 == _T_71[11:0] ? image_1729 : _GEN_4864; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4866 = 12'h6c2 == _T_71[11:0] ? image_1730 : _GEN_4865; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4867 = 12'h6c3 == _T_71[11:0] ? image_1731 : _GEN_4866; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4868 = 12'h6c4 == _T_71[11:0] ? image_1732 : _GEN_4867; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4869 = 12'h6c5 == _T_71[11:0] ? image_1733 : _GEN_4868; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4870 = 12'h6c6 == _T_71[11:0] ? image_1734 : _GEN_4869; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4871 = 12'h6c7 == _T_71[11:0] ? image_1735 : _GEN_4870; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4872 = 12'h6c8 == _T_71[11:0] ? image_1736 : _GEN_4871; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4873 = 12'h6c9 == _T_71[11:0] ? image_1737 : _GEN_4872; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4874 = 12'h6ca == _T_71[11:0] ? image_1738 : _GEN_4873; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4875 = 12'h6cb == _T_71[11:0] ? image_1739 : _GEN_4874; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4876 = 12'h6cc == _T_71[11:0] ? image_1740 : _GEN_4875; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4877 = 12'h6cd == _T_71[11:0] ? image_1741 : _GEN_4876; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4878 = 12'h6ce == _T_71[11:0] ? image_1742 : _GEN_4877; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4879 = 12'h6cf == _T_71[11:0] ? image_1743 : _GEN_4878; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4880 = 12'h6d0 == _T_71[11:0] ? image_1744 : _GEN_4879; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4881 = 12'h6d1 == _T_71[11:0] ? image_1745 : _GEN_4880; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4882 = 12'h6d2 == _T_71[11:0] ? image_1746 : _GEN_4881; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4883 = 12'h6d3 == _T_71[11:0] ? image_1747 : _GEN_4882; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4884 = 12'h6d4 == _T_71[11:0] ? image_1748 : _GEN_4883; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4885 = 12'h6d5 == _T_71[11:0] ? image_1749 : _GEN_4884; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4886 = 12'h6d6 == _T_71[11:0] ? image_1750 : _GEN_4885; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4887 = 12'h6d7 == _T_71[11:0] ? image_1751 : _GEN_4886; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4888 = 12'h6d8 == _T_71[11:0] ? image_1752 : _GEN_4887; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4889 = 12'h6d9 == _T_71[11:0] ? image_1753 : _GEN_4888; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4890 = 12'h6da == _T_71[11:0] ? image_1754 : _GEN_4889; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4891 = 12'h6db == _T_71[11:0] ? image_1755 : _GEN_4890; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4892 = 12'h6dc == _T_71[11:0] ? image_1756 : _GEN_4891; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4893 = 12'h6dd == _T_71[11:0] ? image_1757 : _GEN_4892; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4894 = 12'h6de == _T_71[11:0] ? image_1758 : _GEN_4893; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4895 = 12'h6df == _T_71[11:0] ? image_1759 : _GEN_4894; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4896 = 12'h6e0 == _T_71[11:0] ? image_1760 : _GEN_4895; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4897 = 12'h6e1 == _T_71[11:0] ? image_1761 : _GEN_4896; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4898 = 12'h6e2 == _T_71[11:0] ? image_1762 : _GEN_4897; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4899 = 12'h6e3 == _T_71[11:0] ? image_1763 : _GEN_4898; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4900 = 12'h6e4 == _T_71[11:0] ? image_1764 : _GEN_4899; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4901 = 12'h6e5 == _T_71[11:0] ? image_1765 : _GEN_4900; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4902 = 12'h6e6 == _T_71[11:0] ? image_1766 : _GEN_4901; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4903 = 12'h6e7 == _T_71[11:0] ? image_1767 : _GEN_4902; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4904 = 12'h6e8 == _T_71[11:0] ? image_1768 : _GEN_4903; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4905 = 12'h6e9 == _T_71[11:0] ? image_1769 : _GEN_4904; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4906 = 12'h6ea == _T_71[11:0] ? image_1770 : _GEN_4905; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4907 = 12'h6eb == _T_71[11:0] ? image_1771 : _GEN_4906; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4908 = 12'h6ec == _T_71[11:0] ? image_1772 : _GEN_4907; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4909 = 12'h6ed == _T_71[11:0] ? image_1773 : _GEN_4908; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4910 = 12'h6ee == _T_71[11:0] ? image_1774 : _GEN_4909; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4911 = 12'h6ef == _T_71[11:0] ? image_1775 : _GEN_4910; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4912 = 12'h6f0 == _T_71[11:0] ? image_1776 : _GEN_4911; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4913 = 12'h6f1 == _T_71[11:0] ? image_1777 : _GEN_4912; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4914 = 12'h6f2 == _T_71[11:0] ? image_1778 : _GEN_4913; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4915 = 12'h6f3 == _T_71[11:0] ? image_1779 : _GEN_4914; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4916 = 12'h6f4 == _T_71[11:0] ? image_1780 : _GEN_4915; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4917 = 12'h6f5 == _T_71[11:0] ? image_1781 : _GEN_4916; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4918 = 12'h6f6 == _T_71[11:0] ? image_1782 : _GEN_4917; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4919 = 12'h6f7 == _T_71[11:0] ? image_1783 : _GEN_4918; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4920 = 12'h6f8 == _T_71[11:0] ? image_1784 : _GEN_4919; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4921 = 12'h6f9 == _T_71[11:0] ? image_1785 : _GEN_4920; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4922 = 12'h6fa == _T_71[11:0] ? image_1786 : _GEN_4921; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4923 = 12'h6fb == _T_71[11:0] ? 4'h0 : _GEN_4922; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4924 = 12'h6fc == _T_71[11:0] ? 4'h0 : _GEN_4923; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4925 = 12'h6fd == _T_71[11:0] ? 4'h0 : _GEN_4924; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4926 = 12'h6fe == _T_71[11:0] ? 4'h0 : _GEN_4925; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4927 = 12'h6ff == _T_71[11:0] ? 4'h0 : _GEN_4926; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4928 = 12'h700 == _T_71[11:0] ? 4'h0 : _GEN_4927; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4929 = 12'h701 == _T_71[11:0] ? image_1793 : _GEN_4928; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4930 = 12'h702 == _T_71[11:0] ? image_1794 : _GEN_4929; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4931 = 12'h703 == _T_71[11:0] ? image_1795 : _GEN_4930; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4932 = 12'h704 == _T_71[11:0] ? image_1796 : _GEN_4931; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4933 = 12'h705 == _T_71[11:0] ? image_1797 : _GEN_4932; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4934 = 12'h706 == _T_71[11:0] ? image_1798 : _GEN_4933; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4935 = 12'h707 == _T_71[11:0] ? image_1799 : _GEN_4934; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4936 = 12'h708 == _T_71[11:0] ? image_1800 : _GEN_4935; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4937 = 12'h709 == _T_71[11:0] ? image_1801 : _GEN_4936; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4938 = 12'h70a == _T_71[11:0] ? image_1802 : _GEN_4937; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4939 = 12'h70b == _T_71[11:0] ? image_1803 : _GEN_4938; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4940 = 12'h70c == _T_71[11:0] ? image_1804 : _GEN_4939; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4941 = 12'h70d == _T_71[11:0] ? image_1805 : _GEN_4940; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4942 = 12'h70e == _T_71[11:0] ? image_1806 : _GEN_4941; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4943 = 12'h70f == _T_71[11:0] ? image_1807 : _GEN_4942; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4944 = 12'h710 == _T_71[11:0] ? image_1808 : _GEN_4943; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4945 = 12'h711 == _T_71[11:0] ? image_1809 : _GEN_4944; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4946 = 12'h712 == _T_71[11:0] ? image_1810 : _GEN_4945; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4947 = 12'h713 == _T_71[11:0] ? image_1811 : _GEN_4946; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4948 = 12'h714 == _T_71[11:0] ? image_1812 : _GEN_4947; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4949 = 12'h715 == _T_71[11:0] ? image_1813 : _GEN_4948; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4950 = 12'h716 == _T_71[11:0] ? image_1814 : _GEN_4949; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4951 = 12'h717 == _T_71[11:0] ? image_1815 : _GEN_4950; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4952 = 12'h718 == _T_71[11:0] ? image_1816 : _GEN_4951; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4953 = 12'h719 == _T_71[11:0] ? image_1817 : _GEN_4952; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4954 = 12'h71a == _T_71[11:0] ? image_1818 : _GEN_4953; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4955 = 12'h71b == _T_71[11:0] ? image_1819 : _GEN_4954; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4956 = 12'h71c == _T_71[11:0] ? image_1820 : _GEN_4955; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4957 = 12'h71d == _T_71[11:0] ? image_1821 : _GEN_4956; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4958 = 12'h71e == _T_71[11:0] ? image_1822 : _GEN_4957; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4959 = 12'h71f == _T_71[11:0] ? image_1823 : _GEN_4958; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4960 = 12'h720 == _T_71[11:0] ? image_1824 : _GEN_4959; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4961 = 12'h721 == _T_71[11:0] ? image_1825 : _GEN_4960; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4962 = 12'h722 == _T_71[11:0] ? image_1826 : _GEN_4961; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4963 = 12'h723 == _T_71[11:0] ? image_1827 : _GEN_4962; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4964 = 12'h724 == _T_71[11:0] ? image_1828 : _GEN_4963; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4965 = 12'h725 == _T_71[11:0] ? image_1829 : _GEN_4964; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4966 = 12'h726 == _T_71[11:0] ? image_1830 : _GEN_4965; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4967 = 12'h727 == _T_71[11:0] ? image_1831 : _GEN_4966; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4968 = 12'h728 == _T_71[11:0] ? image_1832 : _GEN_4967; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4969 = 12'h729 == _T_71[11:0] ? image_1833 : _GEN_4968; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4970 = 12'h72a == _T_71[11:0] ? image_1834 : _GEN_4969; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4971 = 12'h72b == _T_71[11:0] ? image_1835 : _GEN_4970; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4972 = 12'h72c == _T_71[11:0] ? image_1836 : _GEN_4971; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4973 = 12'h72d == _T_71[11:0] ? image_1837 : _GEN_4972; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4974 = 12'h72e == _T_71[11:0] ? image_1838 : _GEN_4973; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4975 = 12'h72f == _T_71[11:0] ? image_1839 : _GEN_4974; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4976 = 12'h730 == _T_71[11:0] ? image_1840 : _GEN_4975; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4977 = 12'h731 == _T_71[11:0] ? image_1841 : _GEN_4976; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4978 = 12'h732 == _T_71[11:0] ? image_1842 : _GEN_4977; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4979 = 12'h733 == _T_71[11:0] ? image_1843 : _GEN_4978; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4980 = 12'h734 == _T_71[11:0] ? image_1844 : _GEN_4979; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4981 = 12'h735 == _T_71[11:0] ? image_1845 : _GEN_4980; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4982 = 12'h736 == _T_71[11:0] ? image_1846 : _GEN_4981; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4983 = 12'h737 == _T_71[11:0] ? image_1847 : _GEN_4982; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4984 = 12'h738 == _T_71[11:0] ? image_1848 : _GEN_4983; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4985 = 12'h739 == _T_71[11:0] ? image_1849 : _GEN_4984; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4986 = 12'h73a == _T_71[11:0] ? 4'h0 : _GEN_4985; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4987 = 12'h73b == _T_71[11:0] ? 4'h0 : _GEN_4986; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4988 = 12'h73c == _T_71[11:0] ? 4'h0 : _GEN_4987; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4989 = 12'h73d == _T_71[11:0] ? 4'h0 : _GEN_4988; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4990 = 12'h73e == _T_71[11:0] ? 4'h0 : _GEN_4989; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4991 = 12'h73f == _T_71[11:0] ? 4'h0 : _GEN_4990; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4992 = 12'h740 == _T_71[11:0] ? 4'h0 : _GEN_4991; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4993 = 12'h741 == _T_71[11:0] ? image_1857 : _GEN_4992; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4994 = 12'h742 == _T_71[11:0] ? image_1858 : _GEN_4993; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4995 = 12'h743 == _T_71[11:0] ? image_1859 : _GEN_4994; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4996 = 12'h744 == _T_71[11:0] ? image_1860 : _GEN_4995; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4997 = 12'h745 == _T_71[11:0] ? image_1861 : _GEN_4996; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4998 = 12'h746 == _T_71[11:0] ? image_1862 : _GEN_4997; // @[Filter.scala 138:46]
  wire [3:0] _GEN_4999 = 12'h747 == _T_71[11:0] ? image_1863 : _GEN_4998; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5000 = 12'h748 == _T_71[11:0] ? image_1864 : _GEN_4999; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5001 = 12'h749 == _T_71[11:0] ? image_1865 : _GEN_5000; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5002 = 12'h74a == _T_71[11:0] ? image_1866 : _GEN_5001; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5003 = 12'h74b == _T_71[11:0] ? image_1867 : _GEN_5002; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5004 = 12'h74c == _T_71[11:0] ? image_1868 : _GEN_5003; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5005 = 12'h74d == _T_71[11:0] ? image_1869 : _GEN_5004; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5006 = 12'h74e == _T_71[11:0] ? image_1870 : _GEN_5005; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5007 = 12'h74f == _T_71[11:0] ? image_1871 : _GEN_5006; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5008 = 12'h750 == _T_71[11:0] ? image_1872 : _GEN_5007; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5009 = 12'h751 == _T_71[11:0] ? image_1873 : _GEN_5008; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5010 = 12'h752 == _T_71[11:0] ? image_1874 : _GEN_5009; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5011 = 12'h753 == _T_71[11:0] ? image_1875 : _GEN_5010; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5012 = 12'h754 == _T_71[11:0] ? image_1876 : _GEN_5011; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5013 = 12'h755 == _T_71[11:0] ? image_1877 : _GEN_5012; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5014 = 12'h756 == _T_71[11:0] ? image_1878 : _GEN_5013; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5015 = 12'h757 == _T_71[11:0] ? image_1879 : _GEN_5014; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5016 = 12'h758 == _T_71[11:0] ? image_1880 : _GEN_5015; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5017 = 12'h759 == _T_71[11:0] ? image_1881 : _GEN_5016; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5018 = 12'h75a == _T_71[11:0] ? image_1882 : _GEN_5017; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5019 = 12'h75b == _T_71[11:0] ? image_1883 : _GEN_5018; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5020 = 12'h75c == _T_71[11:0] ? image_1884 : _GEN_5019; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5021 = 12'h75d == _T_71[11:0] ? image_1885 : _GEN_5020; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5022 = 12'h75e == _T_71[11:0] ? image_1886 : _GEN_5021; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5023 = 12'h75f == _T_71[11:0] ? image_1887 : _GEN_5022; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5024 = 12'h760 == _T_71[11:0] ? image_1888 : _GEN_5023; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5025 = 12'h761 == _T_71[11:0] ? image_1889 : _GEN_5024; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5026 = 12'h762 == _T_71[11:0] ? image_1890 : _GEN_5025; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5027 = 12'h763 == _T_71[11:0] ? image_1891 : _GEN_5026; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5028 = 12'h764 == _T_71[11:0] ? image_1892 : _GEN_5027; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5029 = 12'h765 == _T_71[11:0] ? image_1893 : _GEN_5028; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5030 = 12'h766 == _T_71[11:0] ? image_1894 : _GEN_5029; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5031 = 12'h767 == _T_71[11:0] ? image_1895 : _GEN_5030; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5032 = 12'h768 == _T_71[11:0] ? image_1896 : _GEN_5031; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5033 = 12'h769 == _T_71[11:0] ? image_1897 : _GEN_5032; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5034 = 12'h76a == _T_71[11:0] ? image_1898 : _GEN_5033; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5035 = 12'h76b == _T_71[11:0] ? image_1899 : _GEN_5034; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5036 = 12'h76c == _T_71[11:0] ? image_1900 : _GEN_5035; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5037 = 12'h76d == _T_71[11:0] ? image_1901 : _GEN_5036; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5038 = 12'h76e == _T_71[11:0] ? image_1902 : _GEN_5037; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5039 = 12'h76f == _T_71[11:0] ? image_1903 : _GEN_5038; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5040 = 12'h770 == _T_71[11:0] ? image_1904 : _GEN_5039; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5041 = 12'h771 == _T_71[11:0] ? image_1905 : _GEN_5040; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5042 = 12'h772 == _T_71[11:0] ? image_1906 : _GEN_5041; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5043 = 12'h773 == _T_71[11:0] ? image_1907 : _GEN_5042; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5044 = 12'h774 == _T_71[11:0] ? image_1908 : _GEN_5043; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5045 = 12'h775 == _T_71[11:0] ? image_1909 : _GEN_5044; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5046 = 12'h776 == _T_71[11:0] ? image_1910 : _GEN_5045; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5047 = 12'h777 == _T_71[11:0] ? image_1911 : _GEN_5046; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5048 = 12'h778 == _T_71[11:0] ? image_1912 : _GEN_5047; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5049 = 12'h779 == _T_71[11:0] ? image_1913 : _GEN_5048; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5050 = 12'h77a == _T_71[11:0] ? 4'h0 : _GEN_5049; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5051 = 12'h77b == _T_71[11:0] ? 4'h0 : _GEN_5050; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5052 = 12'h77c == _T_71[11:0] ? 4'h0 : _GEN_5051; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5053 = 12'h77d == _T_71[11:0] ? 4'h0 : _GEN_5052; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5054 = 12'h77e == _T_71[11:0] ? 4'h0 : _GEN_5053; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5055 = 12'h77f == _T_71[11:0] ? 4'h0 : _GEN_5054; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5056 = 12'h780 == _T_71[11:0] ? 4'h0 : _GEN_5055; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5057 = 12'h781 == _T_71[11:0] ? image_1921 : _GEN_5056; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5058 = 12'h782 == _T_71[11:0] ? image_1922 : _GEN_5057; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5059 = 12'h783 == _T_71[11:0] ? image_1923 : _GEN_5058; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5060 = 12'h784 == _T_71[11:0] ? image_1924 : _GEN_5059; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5061 = 12'h785 == _T_71[11:0] ? image_1925 : _GEN_5060; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5062 = 12'h786 == _T_71[11:0] ? image_1926 : _GEN_5061; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5063 = 12'h787 == _T_71[11:0] ? image_1927 : _GEN_5062; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5064 = 12'h788 == _T_71[11:0] ? image_1928 : _GEN_5063; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5065 = 12'h789 == _T_71[11:0] ? image_1929 : _GEN_5064; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5066 = 12'h78a == _T_71[11:0] ? image_1930 : _GEN_5065; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5067 = 12'h78b == _T_71[11:0] ? image_1931 : _GEN_5066; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5068 = 12'h78c == _T_71[11:0] ? image_1932 : _GEN_5067; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5069 = 12'h78d == _T_71[11:0] ? image_1933 : _GEN_5068; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5070 = 12'h78e == _T_71[11:0] ? image_1934 : _GEN_5069; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5071 = 12'h78f == _T_71[11:0] ? image_1935 : _GEN_5070; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5072 = 12'h790 == _T_71[11:0] ? image_1936 : _GEN_5071; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5073 = 12'h791 == _T_71[11:0] ? image_1937 : _GEN_5072; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5074 = 12'h792 == _T_71[11:0] ? image_1938 : _GEN_5073; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5075 = 12'h793 == _T_71[11:0] ? image_1939 : _GEN_5074; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5076 = 12'h794 == _T_71[11:0] ? image_1940 : _GEN_5075; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5077 = 12'h795 == _T_71[11:0] ? image_1941 : _GEN_5076; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5078 = 12'h796 == _T_71[11:0] ? image_1942 : _GEN_5077; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5079 = 12'h797 == _T_71[11:0] ? image_1943 : _GEN_5078; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5080 = 12'h798 == _T_71[11:0] ? image_1944 : _GEN_5079; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5081 = 12'h799 == _T_71[11:0] ? image_1945 : _GEN_5080; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5082 = 12'h79a == _T_71[11:0] ? image_1946 : _GEN_5081; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5083 = 12'h79b == _T_71[11:0] ? image_1947 : _GEN_5082; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5084 = 12'h79c == _T_71[11:0] ? image_1948 : _GEN_5083; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5085 = 12'h79d == _T_71[11:0] ? image_1949 : _GEN_5084; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5086 = 12'h79e == _T_71[11:0] ? image_1950 : _GEN_5085; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5087 = 12'h79f == _T_71[11:0] ? image_1951 : _GEN_5086; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5088 = 12'h7a0 == _T_71[11:0] ? image_1952 : _GEN_5087; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5089 = 12'h7a1 == _T_71[11:0] ? image_1953 : _GEN_5088; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5090 = 12'h7a2 == _T_71[11:0] ? image_1954 : _GEN_5089; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5091 = 12'h7a3 == _T_71[11:0] ? image_1955 : _GEN_5090; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5092 = 12'h7a4 == _T_71[11:0] ? image_1956 : _GEN_5091; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5093 = 12'h7a5 == _T_71[11:0] ? image_1957 : _GEN_5092; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5094 = 12'h7a6 == _T_71[11:0] ? image_1958 : _GEN_5093; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5095 = 12'h7a7 == _T_71[11:0] ? image_1959 : _GEN_5094; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5096 = 12'h7a8 == _T_71[11:0] ? image_1960 : _GEN_5095; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5097 = 12'h7a9 == _T_71[11:0] ? image_1961 : _GEN_5096; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5098 = 12'h7aa == _T_71[11:0] ? image_1962 : _GEN_5097; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5099 = 12'h7ab == _T_71[11:0] ? image_1963 : _GEN_5098; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5100 = 12'h7ac == _T_71[11:0] ? image_1964 : _GEN_5099; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5101 = 12'h7ad == _T_71[11:0] ? image_1965 : _GEN_5100; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5102 = 12'h7ae == _T_71[11:0] ? image_1966 : _GEN_5101; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5103 = 12'h7af == _T_71[11:0] ? image_1967 : _GEN_5102; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5104 = 12'h7b0 == _T_71[11:0] ? image_1968 : _GEN_5103; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5105 = 12'h7b1 == _T_71[11:0] ? image_1969 : _GEN_5104; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5106 = 12'h7b2 == _T_71[11:0] ? image_1970 : _GEN_5105; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5107 = 12'h7b3 == _T_71[11:0] ? image_1971 : _GEN_5106; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5108 = 12'h7b4 == _T_71[11:0] ? image_1972 : _GEN_5107; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5109 = 12'h7b5 == _T_71[11:0] ? image_1973 : _GEN_5108; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5110 = 12'h7b6 == _T_71[11:0] ? image_1974 : _GEN_5109; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5111 = 12'h7b7 == _T_71[11:0] ? image_1975 : _GEN_5110; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5112 = 12'h7b8 == _T_71[11:0] ? image_1976 : _GEN_5111; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5113 = 12'h7b9 == _T_71[11:0] ? image_1977 : _GEN_5112; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5114 = 12'h7ba == _T_71[11:0] ? 4'h0 : _GEN_5113; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5115 = 12'h7bb == _T_71[11:0] ? 4'h0 : _GEN_5114; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5116 = 12'h7bc == _T_71[11:0] ? 4'h0 : _GEN_5115; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5117 = 12'h7bd == _T_71[11:0] ? 4'h0 : _GEN_5116; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5118 = 12'h7be == _T_71[11:0] ? 4'h0 : _GEN_5117; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5119 = 12'h7bf == _T_71[11:0] ? 4'h0 : _GEN_5118; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5120 = 12'h7c0 == _T_71[11:0] ? 4'h0 : _GEN_5119; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5121 = 12'h7c1 == _T_71[11:0] ? image_1985 : _GEN_5120; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5122 = 12'h7c2 == _T_71[11:0] ? image_1986 : _GEN_5121; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5123 = 12'h7c3 == _T_71[11:0] ? image_1987 : _GEN_5122; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5124 = 12'h7c4 == _T_71[11:0] ? image_1988 : _GEN_5123; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5125 = 12'h7c5 == _T_71[11:0] ? image_1989 : _GEN_5124; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5126 = 12'h7c6 == _T_71[11:0] ? image_1990 : _GEN_5125; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5127 = 12'h7c7 == _T_71[11:0] ? image_1991 : _GEN_5126; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5128 = 12'h7c8 == _T_71[11:0] ? image_1992 : _GEN_5127; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5129 = 12'h7c9 == _T_71[11:0] ? image_1993 : _GEN_5128; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5130 = 12'h7ca == _T_71[11:0] ? image_1994 : _GEN_5129; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5131 = 12'h7cb == _T_71[11:0] ? image_1995 : _GEN_5130; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5132 = 12'h7cc == _T_71[11:0] ? image_1996 : _GEN_5131; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5133 = 12'h7cd == _T_71[11:0] ? image_1997 : _GEN_5132; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5134 = 12'h7ce == _T_71[11:0] ? image_1998 : _GEN_5133; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5135 = 12'h7cf == _T_71[11:0] ? image_1999 : _GEN_5134; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5136 = 12'h7d0 == _T_71[11:0] ? image_2000 : _GEN_5135; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5137 = 12'h7d1 == _T_71[11:0] ? image_2001 : _GEN_5136; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5138 = 12'h7d2 == _T_71[11:0] ? image_2002 : _GEN_5137; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5139 = 12'h7d3 == _T_71[11:0] ? image_2003 : _GEN_5138; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5140 = 12'h7d4 == _T_71[11:0] ? image_2004 : _GEN_5139; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5141 = 12'h7d5 == _T_71[11:0] ? image_2005 : _GEN_5140; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5142 = 12'h7d6 == _T_71[11:0] ? image_2006 : _GEN_5141; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5143 = 12'h7d7 == _T_71[11:0] ? image_2007 : _GEN_5142; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5144 = 12'h7d8 == _T_71[11:0] ? image_2008 : _GEN_5143; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5145 = 12'h7d9 == _T_71[11:0] ? image_2009 : _GEN_5144; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5146 = 12'h7da == _T_71[11:0] ? image_2010 : _GEN_5145; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5147 = 12'h7db == _T_71[11:0] ? image_2011 : _GEN_5146; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5148 = 12'h7dc == _T_71[11:0] ? image_2012 : _GEN_5147; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5149 = 12'h7dd == _T_71[11:0] ? image_2013 : _GEN_5148; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5150 = 12'h7de == _T_71[11:0] ? image_2014 : _GEN_5149; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5151 = 12'h7df == _T_71[11:0] ? image_2015 : _GEN_5150; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5152 = 12'h7e0 == _T_71[11:0] ? image_2016 : _GEN_5151; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5153 = 12'h7e1 == _T_71[11:0] ? image_2017 : _GEN_5152; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5154 = 12'h7e2 == _T_71[11:0] ? image_2018 : _GEN_5153; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5155 = 12'h7e3 == _T_71[11:0] ? image_2019 : _GEN_5154; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5156 = 12'h7e4 == _T_71[11:0] ? image_2020 : _GEN_5155; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5157 = 12'h7e5 == _T_71[11:0] ? image_2021 : _GEN_5156; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5158 = 12'h7e6 == _T_71[11:0] ? image_2022 : _GEN_5157; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5159 = 12'h7e7 == _T_71[11:0] ? image_2023 : _GEN_5158; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5160 = 12'h7e8 == _T_71[11:0] ? image_2024 : _GEN_5159; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5161 = 12'h7e9 == _T_71[11:0] ? image_2025 : _GEN_5160; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5162 = 12'h7ea == _T_71[11:0] ? image_2026 : _GEN_5161; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5163 = 12'h7eb == _T_71[11:0] ? image_2027 : _GEN_5162; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5164 = 12'h7ec == _T_71[11:0] ? image_2028 : _GEN_5163; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5165 = 12'h7ed == _T_71[11:0] ? image_2029 : _GEN_5164; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5166 = 12'h7ee == _T_71[11:0] ? image_2030 : _GEN_5165; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5167 = 12'h7ef == _T_71[11:0] ? image_2031 : _GEN_5166; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5168 = 12'h7f0 == _T_71[11:0] ? image_2032 : _GEN_5167; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5169 = 12'h7f1 == _T_71[11:0] ? image_2033 : _GEN_5168; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5170 = 12'h7f2 == _T_71[11:0] ? image_2034 : _GEN_5169; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5171 = 12'h7f3 == _T_71[11:0] ? image_2035 : _GEN_5170; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5172 = 12'h7f4 == _T_71[11:0] ? image_2036 : _GEN_5171; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5173 = 12'h7f5 == _T_71[11:0] ? image_2037 : _GEN_5172; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5174 = 12'h7f6 == _T_71[11:0] ? image_2038 : _GEN_5173; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5175 = 12'h7f7 == _T_71[11:0] ? image_2039 : _GEN_5174; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5176 = 12'h7f8 == _T_71[11:0] ? image_2040 : _GEN_5175; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5177 = 12'h7f9 == _T_71[11:0] ? image_2041 : _GEN_5176; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5178 = 12'h7fa == _T_71[11:0] ? 4'h0 : _GEN_5177; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5179 = 12'h7fb == _T_71[11:0] ? 4'h0 : _GEN_5178; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5180 = 12'h7fc == _T_71[11:0] ? 4'h0 : _GEN_5179; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5181 = 12'h7fd == _T_71[11:0] ? 4'h0 : _GEN_5180; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5182 = 12'h7fe == _T_71[11:0] ? 4'h0 : _GEN_5181; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5183 = 12'h7ff == _T_71[11:0] ? 4'h0 : _GEN_5182; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5184 = 12'h800 == _T_71[11:0] ? 4'h0 : _GEN_5183; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5185 = 12'h801 == _T_71[11:0] ? image_2049 : _GEN_5184; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5186 = 12'h802 == _T_71[11:0] ? image_2050 : _GEN_5185; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5187 = 12'h803 == _T_71[11:0] ? image_2051 : _GEN_5186; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5188 = 12'h804 == _T_71[11:0] ? image_2052 : _GEN_5187; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5189 = 12'h805 == _T_71[11:0] ? image_2053 : _GEN_5188; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5190 = 12'h806 == _T_71[11:0] ? image_2054 : _GEN_5189; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5191 = 12'h807 == _T_71[11:0] ? image_2055 : _GEN_5190; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5192 = 12'h808 == _T_71[11:0] ? image_2056 : _GEN_5191; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5193 = 12'h809 == _T_71[11:0] ? image_2057 : _GEN_5192; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5194 = 12'h80a == _T_71[11:0] ? image_2058 : _GEN_5193; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5195 = 12'h80b == _T_71[11:0] ? image_2059 : _GEN_5194; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5196 = 12'h80c == _T_71[11:0] ? image_2060 : _GEN_5195; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5197 = 12'h80d == _T_71[11:0] ? image_2061 : _GEN_5196; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5198 = 12'h80e == _T_71[11:0] ? image_2062 : _GEN_5197; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5199 = 12'h80f == _T_71[11:0] ? image_2063 : _GEN_5198; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5200 = 12'h810 == _T_71[11:0] ? image_2064 : _GEN_5199; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5201 = 12'h811 == _T_71[11:0] ? image_2065 : _GEN_5200; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5202 = 12'h812 == _T_71[11:0] ? image_2066 : _GEN_5201; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5203 = 12'h813 == _T_71[11:0] ? image_2067 : _GEN_5202; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5204 = 12'h814 == _T_71[11:0] ? image_2068 : _GEN_5203; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5205 = 12'h815 == _T_71[11:0] ? image_2069 : _GEN_5204; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5206 = 12'h816 == _T_71[11:0] ? image_2070 : _GEN_5205; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5207 = 12'h817 == _T_71[11:0] ? image_2071 : _GEN_5206; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5208 = 12'h818 == _T_71[11:0] ? image_2072 : _GEN_5207; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5209 = 12'h819 == _T_71[11:0] ? image_2073 : _GEN_5208; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5210 = 12'h81a == _T_71[11:0] ? image_2074 : _GEN_5209; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5211 = 12'h81b == _T_71[11:0] ? image_2075 : _GEN_5210; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5212 = 12'h81c == _T_71[11:0] ? image_2076 : _GEN_5211; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5213 = 12'h81d == _T_71[11:0] ? image_2077 : _GEN_5212; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5214 = 12'h81e == _T_71[11:0] ? image_2078 : _GEN_5213; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5215 = 12'h81f == _T_71[11:0] ? image_2079 : _GEN_5214; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5216 = 12'h820 == _T_71[11:0] ? image_2080 : _GEN_5215; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5217 = 12'h821 == _T_71[11:0] ? image_2081 : _GEN_5216; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5218 = 12'h822 == _T_71[11:0] ? image_2082 : _GEN_5217; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5219 = 12'h823 == _T_71[11:0] ? image_2083 : _GEN_5218; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5220 = 12'h824 == _T_71[11:0] ? image_2084 : _GEN_5219; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5221 = 12'h825 == _T_71[11:0] ? image_2085 : _GEN_5220; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5222 = 12'h826 == _T_71[11:0] ? image_2086 : _GEN_5221; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5223 = 12'h827 == _T_71[11:0] ? image_2087 : _GEN_5222; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5224 = 12'h828 == _T_71[11:0] ? image_2088 : _GEN_5223; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5225 = 12'h829 == _T_71[11:0] ? image_2089 : _GEN_5224; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5226 = 12'h82a == _T_71[11:0] ? image_2090 : _GEN_5225; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5227 = 12'h82b == _T_71[11:0] ? image_2091 : _GEN_5226; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5228 = 12'h82c == _T_71[11:0] ? image_2092 : _GEN_5227; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5229 = 12'h82d == _T_71[11:0] ? image_2093 : _GEN_5228; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5230 = 12'h82e == _T_71[11:0] ? image_2094 : _GEN_5229; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5231 = 12'h82f == _T_71[11:0] ? image_2095 : _GEN_5230; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5232 = 12'h830 == _T_71[11:0] ? image_2096 : _GEN_5231; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5233 = 12'h831 == _T_71[11:0] ? image_2097 : _GEN_5232; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5234 = 12'h832 == _T_71[11:0] ? image_2098 : _GEN_5233; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5235 = 12'h833 == _T_71[11:0] ? image_2099 : _GEN_5234; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5236 = 12'h834 == _T_71[11:0] ? image_2100 : _GEN_5235; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5237 = 12'h835 == _T_71[11:0] ? image_2101 : _GEN_5236; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5238 = 12'h836 == _T_71[11:0] ? image_2102 : _GEN_5237; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5239 = 12'h837 == _T_71[11:0] ? image_2103 : _GEN_5238; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5240 = 12'h838 == _T_71[11:0] ? image_2104 : _GEN_5239; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5241 = 12'h839 == _T_71[11:0] ? image_2105 : _GEN_5240; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5242 = 12'h83a == _T_71[11:0] ? image_2106 : _GEN_5241; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5243 = 12'h83b == _T_71[11:0] ? 4'h0 : _GEN_5242; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5244 = 12'h83c == _T_71[11:0] ? 4'h0 : _GEN_5243; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5245 = 12'h83d == _T_71[11:0] ? 4'h0 : _GEN_5244; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5246 = 12'h83e == _T_71[11:0] ? 4'h0 : _GEN_5245; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5247 = 12'h83f == _T_71[11:0] ? 4'h0 : _GEN_5246; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5248 = 12'h840 == _T_71[11:0] ? 4'h0 : _GEN_5247; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5249 = 12'h841 == _T_71[11:0] ? 4'h0 : _GEN_5248; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5250 = 12'h842 == _T_71[11:0] ? image_2114 : _GEN_5249; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5251 = 12'h843 == _T_71[11:0] ? image_2115 : _GEN_5250; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5252 = 12'h844 == _T_71[11:0] ? image_2116 : _GEN_5251; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5253 = 12'h845 == _T_71[11:0] ? image_2117 : _GEN_5252; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5254 = 12'h846 == _T_71[11:0] ? image_2118 : _GEN_5253; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5255 = 12'h847 == _T_71[11:0] ? image_2119 : _GEN_5254; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5256 = 12'h848 == _T_71[11:0] ? image_2120 : _GEN_5255; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5257 = 12'h849 == _T_71[11:0] ? image_2121 : _GEN_5256; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5258 = 12'h84a == _T_71[11:0] ? image_2122 : _GEN_5257; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5259 = 12'h84b == _T_71[11:0] ? image_2123 : _GEN_5258; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5260 = 12'h84c == _T_71[11:0] ? image_2124 : _GEN_5259; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5261 = 12'h84d == _T_71[11:0] ? image_2125 : _GEN_5260; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5262 = 12'h84e == _T_71[11:0] ? image_2126 : _GEN_5261; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5263 = 12'h84f == _T_71[11:0] ? image_2127 : _GEN_5262; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5264 = 12'h850 == _T_71[11:0] ? image_2128 : _GEN_5263; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5265 = 12'h851 == _T_71[11:0] ? image_2129 : _GEN_5264; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5266 = 12'h852 == _T_71[11:0] ? image_2130 : _GEN_5265; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5267 = 12'h853 == _T_71[11:0] ? image_2131 : _GEN_5266; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5268 = 12'h854 == _T_71[11:0] ? image_2132 : _GEN_5267; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5269 = 12'h855 == _T_71[11:0] ? image_2133 : _GEN_5268; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5270 = 12'h856 == _T_71[11:0] ? image_2134 : _GEN_5269; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5271 = 12'h857 == _T_71[11:0] ? image_2135 : _GEN_5270; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5272 = 12'h858 == _T_71[11:0] ? image_2136 : _GEN_5271; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5273 = 12'h859 == _T_71[11:0] ? image_2137 : _GEN_5272; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5274 = 12'h85a == _T_71[11:0] ? image_2138 : _GEN_5273; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5275 = 12'h85b == _T_71[11:0] ? image_2139 : _GEN_5274; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5276 = 12'h85c == _T_71[11:0] ? image_2140 : _GEN_5275; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5277 = 12'h85d == _T_71[11:0] ? image_2141 : _GEN_5276; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5278 = 12'h85e == _T_71[11:0] ? image_2142 : _GEN_5277; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5279 = 12'h85f == _T_71[11:0] ? image_2143 : _GEN_5278; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5280 = 12'h860 == _T_71[11:0] ? image_2144 : _GEN_5279; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5281 = 12'h861 == _T_71[11:0] ? image_2145 : _GEN_5280; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5282 = 12'h862 == _T_71[11:0] ? image_2146 : _GEN_5281; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5283 = 12'h863 == _T_71[11:0] ? image_2147 : _GEN_5282; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5284 = 12'h864 == _T_71[11:0] ? image_2148 : _GEN_5283; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5285 = 12'h865 == _T_71[11:0] ? image_2149 : _GEN_5284; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5286 = 12'h866 == _T_71[11:0] ? image_2150 : _GEN_5285; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5287 = 12'h867 == _T_71[11:0] ? image_2151 : _GEN_5286; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5288 = 12'h868 == _T_71[11:0] ? image_2152 : _GEN_5287; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5289 = 12'h869 == _T_71[11:0] ? image_2153 : _GEN_5288; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5290 = 12'h86a == _T_71[11:0] ? image_2154 : _GEN_5289; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5291 = 12'h86b == _T_71[11:0] ? image_2155 : _GEN_5290; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5292 = 12'h86c == _T_71[11:0] ? image_2156 : _GEN_5291; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5293 = 12'h86d == _T_71[11:0] ? image_2157 : _GEN_5292; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5294 = 12'h86e == _T_71[11:0] ? image_2158 : _GEN_5293; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5295 = 12'h86f == _T_71[11:0] ? image_2159 : _GEN_5294; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5296 = 12'h870 == _T_71[11:0] ? image_2160 : _GEN_5295; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5297 = 12'h871 == _T_71[11:0] ? image_2161 : _GEN_5296; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5298 = 12'h872 == _T_71[11:0] ? image_2162 : _GEN_5297; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5299 = 12'h873 == _T_71[11:0] ? image_2163 : _GEN_5298; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5300 = 12'h874 == _T_71[11:0] ? image_2164 : _GEN_5299; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5301 = 12'h875 == _T_71[11:0] ? image_2165 : _GEN_5300; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5302 = 12'h876 == _T_71[11:0] ? image_2166 : _GEN_5301; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5303 = 12'h877 == _T_71[11:0] ? image_2167 : _GEN_5302; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5304 = 12'h878 == _T_71[11:0] ? image_2168 : _GEN_5303; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5305 = 12'h879 == _T_71[11:0] ? image_2169 : _GEN_5304; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5306 = 12'h87a == _T_71[11:0] ? image_2170 : _GEN_5305; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5307 = 12'h87b == _T_71[11:0] ? 4'h0 : _GEN_5306; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5308 = 12'h87c == _T_71[11:0] ? 4'h0 : _GEN_5307; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5309 = 12'h87d == _T_71[11:0] ? 4'h0 : _GEN_5308; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5310 = 12'h87e == _T_71[11:0] ? 4'h0 : _GEN_5309; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5311 = 12'h87f == _T_71[11:0] ? 4'h0 : _GEN_5310; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5312 = 12'h880 == _T_71[11:0] ? 4'h0 : _GEN_5311; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5313 = 12'h881 == _T_71[11:0] ? image_2177 : _GEN_5312; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5314 = 12'h882 == _T_71[11:0] ? image_2178 : _GEN_5313; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5315 = 12'h883 == _T_71[11:0] ? image_2179 : _GEN_5314; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5316 = 12'h884 == _T_71[11:0] ? image_2180 : _GEN_5315; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5317 = 12'h885 == _T_71[11:0] ? image_2181 : _GEN_5316; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5318 = 12'h886 == _T_71[11:0] ? image_2182 : _GEN_5317; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5319 = 12'h887 == _T_71[11:0] ? image_2183 : _GEN_5318; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5320 = 12'h888 == _T_71[11:0] ? image_2184 : _GEN_5319; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5321 = 12'h889 == _T_71[11:0] ? image_2185 : _GEN_5320; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5322 = 12'h88a == _T_71[11:0] ? image_2186 : _GEN_5321; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5323 = 12'h88b == _T_71[11:0] ? image_2187 : _GEN_5322; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5324 = 12'h88c == _T_71[11:0] ? image_2188 : _GEN_5323; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5325 = 12'h88d == _T_71[11:0] ? image_2189 : _GEN_5324; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5326 = 12'h88e == _T_71[11:0] ? image_2190 : _GEN_5325; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5327 = 12'h88f == _T_71[11:0] ? image_2191 : _GEN_5326; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5328 = 12'h890 == _T_71[11:0] ? image_2192 : _GEN_5327; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5329 = 12'h891 == _T_71[11:0] ? image_2193 : _GEN_5328; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5330 = 12'h892 == _T_71[11:0] ? image_2194 : _GEN_5329; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5331 = 12'h893 == _T_71[11:0] ? image_2195 : _GEN_5330; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5332 = 12'h894 == _T_71[11:0] ? image_2196 : _GEN_5331; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5333 = 12'h895 == _T_71[11:0] ? image_2197 : _GEN_5332; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5334 = 12'h896 == _T_71[11:0] ? image_2198 : _GEN_5333; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5335 = 12'h897 == _T_71[11:0] ? image_2199 : _GEN_5334; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5336 = 12'h898 == _T_71[11:0] ? image_2200 : _GEN_5335; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5337 = 12'h899 == _T_71[11:0] ? image_2201 : _GEN_5336; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5338 = 12'h89a == _T_71[11:0] ? image_2202 : _GEN_5337; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5339 = 12'h89b == _T_71[11:0] ? image_2203 : _GEN_5338; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5340 = 12'h89c == _T_71[11:0] ? image_2204 : _GEN_5339; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5341 = 12'h89d == _T_71[11:0] ? image_2205 : _GEN_5340; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5342 = 12'h89e == _T_71[11:0] ? image_2206 : _GEN_5341; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5343 = 12'h89f == _T_71[11:0] ? image_2207 : _GEN_5342; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5344 = 12'h8a0 == _T_71[11:0] ? image_2208 : _GEN_5343; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5345 = 12'h8a1 == _T_71[11:0] ? image_2209 : _GEN_5344; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5346 = 12'h8a2 == _T_71[11:0] ? image_2210 : _GEN_5345; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5347 = 12'h8a3 == _T_71[11:0] ? image_2211 : _GEN_5346; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5348 = 12'h8a4 == _T_71[11:0] ? image_2212 : _GEN_5347; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5349 = 12'h8a5 == _T_71[11:0] ? image_2213 : _GEN_5348; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5350 = 12'h8a6 == _T_71[11:0] ? image_2214 : _GEN_5349; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5351 = 12'h8a7 == _T_71[11:0] ? image_2215 : _GEN_5350; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5352 = 12'h8a8 == _T_71[11:0] ? image_2216 : _GEN_5351; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5353 = 12'h8a9 == _T_71[11:0] ? image_2217 : _GEN_5352; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5354 = 12'h8aa == _T_71[11:0] ? image_2218 : _GEN_5353; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5355 = 12'h8ab == _T_71[11:0] ? image_2219 : _GEN_5354; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5356 = 12'h8ac == _T_71[11:0] ? image_2220 : _GEN_5355; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5357 = 12'h8ad == _T_71[11:0] ? image_2221 : _GEN_5356; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5358 = 12'h8ae == _T_71[11:0] ? image_2222 : _GEN_5357; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5359 = 12'h8af == _T_71[11:0] ? image_2223 : _GEN_5358; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5360 = 12'h8b0 == _T_71[11:0] ? image_2224 : _GEN_5359; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5361 = 12'h8b1 == _T_71[11:0] ? image_2225 : _GEN_5360; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5362 = 12'h8b2 == _T_71[11:0] ? image_2226 : _GEN_5361; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5363 = 12'h8b3 == _T_71[11:0] ? image_2227 : _GEN_5362; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5364 = 12'h8b4 == _T_71[11:0] ? image_2228 : _GEN_5363; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5365 = 12'h8b5 == _T_71[11:0] ? image_2229 : _GEN_5364; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5366 = 12'h8b6 == _T_71[11:0] ? image_2230 : _GEN_5365; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5367 = 12'h8b7 == _T_71[11:0] ? image_2231 : _GEN_5366; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5368 = 12'h8b8 == _T_71[11:0] ? image_2232 : _GEN_5367; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5369 = 12'h8b9 == _T_71[11:0] ? image_2233 : _GEN_5368; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5370 = 12'h8ba == _T_71[11:0] ? image_2234 : _GEN_5369; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5371 = 12'h8bb == _T_71[11:0] ? 4'h0 : _GEN_5370; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5372 = 12'h8bc == _T_71[11:0] ? 4'h0 : _GEN_5371; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5373 = 12'h8bd == _T_71[11:0] ? 4'h0 : _GEN_5372; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5374 = 12'h8be == _T_71[11:0] ? 4'h0 : _GEN_5373; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5375 = 12'h8bf == _T_71[11:0] ? 4'h0 : _GEN_5374; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5376 = 12'h8c0 == _T_71[11:0] ? 4'h0 : _GEN_5375; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5377 = 12'h8c1 == _T_71[11:0] ? 4'h0 : _GEN_5376; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5378 = 12'h8c2 == _T_71[11:0] ? 4'h0 : _GEN_5377; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5379 = 12'h8c3 == _T_71[11:0] ? image_2243 : _GEN_5378; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5380 = 12'h8c4 == _T_71[11:0] ? image_2244 : _GEN_5379; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5381 = 12'h8c5 == _T_71[11:0] ? image_2245 : _GEN_5380; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5382 = 12'h8c6 == _T_71[11:0] ? image_2246 : _GEN_5381; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5383 = 12'h8c7 == _T_71[11:0] ? image_2247 : _GEN_5382; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5384 = 12'h8c8 == _T_71[11:0] ? image_2248 : _GEN_5383; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5385 = 12'h8c9 == _T_71[11:0] ? image_2249 : _GEN_5384; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5386 = 12'h8ca == _T_71[11:0] ? image_2250 : _GEN_5385; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5387 = 12'h8cb == _T_71[11:0] ? image_2251 : _GEN_5386; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5388 = 12'h8cc == _T_71[11:0] ? image_2252 : _GEN_5387; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5389 = 12'h8cd == _T_71[11:0] ? image_2253 : _GEN_5388; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5390 = 12'h8ce == _T_71[11:0] ? image_2254 : _GEN_5389; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5391 = 12'h8cf == _T_71[11:0] ? image_2255 : _GEN_5390; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5392 = 12'h8d0 == _T_71[11:0] ? image_2256 : _GEN_5391; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5393 = 12'h8d1 == _T_71[11:0] ? image_2257 : _GEN_5392; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5394 = 12'h8d2 == _T_71[11:0] ? image_2258 : _GEN_5393; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5395 = 12'h8d3 == _T_71[11:0] ? image_2259 : _GEN_5394; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5396 = 12'h8d4 == _T_71[11:0] ? image_2260 : _GEN_5395; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5397 = 12'h8d5 == _T_71[11:0] ? image_2261 : _GEN_5396; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5398 = 12'h8d6 == _T_71[11:0] ? image_2262 : _GEN_5397; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5399 = 12'h8d7 == _T_71[11:0] ? image_2263 : _GEN_5398; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5400 = 12'h8d8 == _T_71[11:0] ? image_2264 : _GEN_5399; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5401 = 12'h8d9 == _T_71[11:0] ? image_2265 : _GEN_5400; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5402 = 12'h8da == _T_71[11:0] ? image_2266 : _GEN_5401; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5403 = 12'h8db == _T_71[11:0] ? image_2267 : _GEN_5402; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5404 = 12'h8dc == _T_71[11:0] ? image_2268 : _GEN_5403; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5405 = 12'h8dd == _T_71[11:0] ? image_2269 : _GEN_5404; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5406 = 12'h8de == _T_71[11:0] ? image_2270 : _GEN_5405; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5407 = 12'h8df == _T_71[11:0] ? image_2271 : _GEN_5406; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5408 = 12'h8e0 == _T_71[11:0] ? image_2272 : _GEN_5407; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5409 = 12'h8e1 == _T_71[11:0] ? image_2273 : _GEN_5408; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5410 = 12'h8e2 == _T_71[11:0] ? image_2274 : _GEN_5409; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5411 = 12'h8e3 == _T_71[11:0] ? image_2275 : _GEN_5410; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5412 = 12'h8e4 == _T_71[11:0] ? image_2276 : _GEN_5411; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5413 = 12'h8e5 == _T_71[11:0] ? image_2277 : _GEN_5412; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5414 = 12'h8e6 == _T_71[11:0] ? image_2278 : _GEN_5413; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5415 = 12'h8e7 == _T_71[11:0] ? image_2279 : _GEN_5414; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5416 = 12'h8e8 == _T_71[11:0] ? image_2280 : _GEN_5415; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5417 = 12'h8e9 == _T_71[11:0] ? image_2281 : _GEN_5416; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5418 = 12'h8ea == _T_71[11:0] ? image_2282 : _GEN_5417; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5419 = 12'h8eb == _T_71[11:0] ? image_2283 : _GEN_5418; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5420 = 12'h8ec == _T_71[11:0] ? image_2284 : _GEN_5419; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5421 = 12'h8ed == _T_71[11:0] ? image_2285 : _GEN_5420; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5422 = 12'h8ee == _T_71[11:0] ? image_2286 : _GEN_5421; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5423 = 12'h8ef == _T_71[11:0] ? image_2287 : _GEN_5422; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5424 = 12'h8f0 == _T_71[11:0] ? image_2288 : _GEN_5423; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5425 = 12'h8f1 == _T_71[11:0] ? image_2289 : _GEN_5424; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5426 = 12'h8f2 == _T_71[11:0] ? image_2290 : _GEN_5425; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5427 = 12'h8f3 == _T_71[11:0] ? image_2291 : _GEN_5426; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5428 = 12'h8f4 == _T_71[11:0] ? image_2292 : _GEN_5427; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5429 = 12'h8f5 == _T_71[11:0] ? image_2293 : _GEN_5428; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5430 = 12'h8f6 == _T_71[11:0] ? image_2294 : _GEN_5429; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5431 = 12'h8f7 == _T_71[11:0] ? image_2295 : _GEN_5430; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5432 = 12'h8f8 == _T_71[11:0] ? image_2296 : _GEN_5431; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5433 = 12'h8f9 == _T_71[11:0] ? image_2297 : _GEN_5432; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5434 = 12'h8fa == _T_71[11:0] ? image_2298 : _GEN_5433; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5435 = 12'h8fb == _T_71[11:0] ? 4'h0 : _GEN_5434; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5436 = 12'h8fc == _T_71[11:0] ? 4'h0 : _GEN_5435; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5437 = 12'h8fd == _T_71[11:0] ? 4'h0 : _GEN_5436; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5438 = 12'h8fe == _T_71[11:0] ? 4'h0 : _GEN_5437; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5439 = 12'h8ff == _T_71[11:0] ? 4'h0 : _GEN_5438; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5440 = 12'h900 == _T_71[11:0] ? 4'h0 : _GEN_5439; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5441 = 12'h901 == _T_71[11:0] ? 4'h0 : _GEN_5440; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5442 = 12'h902 == _T_71[11:0] ? 4'h0 : _GEN_5441; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5443 = 12'h903 == _T_71[11:0] ? image_2307 : _GEN_5442; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5444 = 12'h904 == _T_71[11:0] ? image_2308 : _GEN_5443; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5445 = 12'h905 == _T_71[11:0] ? image_2309 : _GEN_5444; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5446 = 12'h906 == _T_71[11:0] ? image_2310 : _GEN_5445; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5447 = 12'h907 == _T_71[11:0] ? image_2311 : _GEN_5446; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5448 = 12'h908 == _T_71[11:0] ? image_2312 : _GEN_5447; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5449 = 12'h909 == _T_71[11:0] ? image_2313 : _GEN_5448; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5450 = 12'h90a == _T_71[11:0] ? image_2314 : _GEN_5449; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5451 = 12'h90b == _T_71[11:0] ? image_2315 : _GEN_5450; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5452 = 12'h90c == _T_71[11:0] ? image_2316 : _GEN_5451; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5453 = 12'h90d == _T_71[11:0] ? image_2317 : _GEN_5452; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5454 = 12'h90e == _T_71[11:0] ? image_2318 : _GEN_5453; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5455 = 12'h90f == _T_71[11:0] ? image_2319 : _GEN_5454; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5456 = 12'h910 == _T_71[11:0] ? image_2320 : _GEN_5455; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5457 = 12'h911 == _T_71[11:0] ? image_2321 : _GEN_5456; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5458 = 12'h912 == _T_71[11:0] ? image_2322 : _GEN_5457; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5459 = 12'h913 == _T_71[11:0] ? image_2323 : _GEN_5458; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5460 = 12'h914 == _T_71[11:0] ? image_2324 : _GEN_5459; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5461 = 12'h915 == _T_71[11:0] ? image_2325 : _GEN_5460; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5462 = 12'h916 == _T_71[11:0] ? image_2326 : _GEN_5461; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5463 = 12'h917 == _T_71[11:0] ? image_2327 : _GEN_5462; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5464 = 12'h918 == _T_71[11:0] ? image_2328 : _GEN_5463; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5465 = 12'h919 == _T_71[11:0] ? image_2329 : _GEN_5464; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5466 = 12'h91a == _T_71[11:0] ? image_2330 : _GEN_5465; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5467 = 12'h91b == _T_71[11:0] ? image_2331 : _GEN_5466; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5468 = 12'h91c == _T_71[11:0] ? image_2332 : _GEN_5467; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5469 = 12'h91d == _T_71[11:0] ? image_2333 : _GEN_5468; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5470 = 12'h91e == _T_71[11:0] ? image_2334 : _GEN_5469; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5471 = 12'h91f == _T_71[11:0] ? image_2335 : _GEN_5470; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5472 = 12'h920 == _T_71[11:0] ? image_2336 : _GEN_5471; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5473 = 12'h921 == _T_71[11:0] ? image_2337 : _GEN_5472; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5474 = 12'h922 == _T_71[11:0] ? image_2338 : _GEN_5473; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5475 = 12'h923 == _T_71[11:0] ? image_2339 : _GEN_5474; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5476 = 12'h924 == _T_71[11:0] ? image_2340 : _GEN_5475; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5477 = 12'h925 == _T_71[11:0] ? image_2341 : _GEN_5476; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5478 = 12'h926 == _T_71[11:0] ? image_2342 : _GEN_5477; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5479 = 12'h927 == _T_71[11:0] ? image_2343 : _GEN_5478; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5480 = 12'h928 == _T_71[11:0] ? image_2344 : _GEN_5479; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5481 = 12'h929 == _T_71[11:0] ? image_2345 : _GEN_5480; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5482 = 12'h92a == _T_71[11:0] ? image_2346 : _GEN_5481; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5483 = 12'h92b == _T_71[11:0] ? image_2347 : _GEN_5482; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5484 = 12'h92c == _T_71[11:0] ? image_2348 : _GEN_5483; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5485 = 12'h92d == _T_71[11:0] ? image_2349 : _GEN_5484; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5486 = 12'h92e == _T_71[11:0] ? image_2350 : _GEN_5485; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5487 = 12'h92f == _T_71[11:0] ? image_2351 : _GEN_5486; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5488 = 12'h930 == _T_71[11:0] ? image_2352 : _GEN_5487; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5489 = 12'h931 == _T_71[11:0] ? image_2353 : _GEN_5488; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5490 = 12'h932 == _T_71[11:0] ? image_2354 : _GEN_5489; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5491 = 12'h933 == _T_71[11:0] ? image_2355 : _GEN_5490; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5492 = 12'h934 == _T_71[11:0] ? image_2356 : _GEN_5491; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5493 = 12'h935 == _T_71[11:0] ? image_2357 : _GEN_5492; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5494 = 12'h936 == _T_71[11:0] ? image_2358 : _GEN_5493; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5495 = 12'h937 == _T_71[11:0] ? image_2359 : _GEN_5494; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5496 = 12'h938 == _T_71[11:0] ? image_2360 : _GEN_5495; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5497 = 12'h939 == _T_71[11:0] ? image_2361 : _GEN_5496; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5498 = 12'h93a == _T_71[11:0] ? image_2362 : _GEN_5497; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5499 = 12'h93b == _T_71[11:0] ? 4'h0 : _GEN_5498; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5500 = 12'h93c == _T_71[11:0] ? 4'h0 : _GEN_5499; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5501 = 12'h93d == _T_71[11:0] ? 4'h0 : _GEN_5500; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5502 = 12'h93e == _T_71[11:0] ? 4'h0 : _GEN_5501; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5503 = 12'h93f == _T_71[11:0] ? 4'h0 : _GEN_5502; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5504 = 12'h940 == _T_71[11:0] ? 4'h0 : _GEN_5503; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5505 = 12'h941 == _T_71[11:0] ? 4'h0 : _GEN_5504; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5506 = 12'h942 == _T_71[11:0] ? 4'h0 : _GEN_5505; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5507 = 12'h943 == _T_71[11:0] ? 4'h0 : _GEN_5506; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5508 = 12'h944 == _T_71[11:0] ? image_2372 : _GEN_5507; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5509 = 12'h945 == _T_71[11:0] ? image_2373 : _GEN_5508; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5510 = 12'h946 == _T_71[11:0] ? image_2374 : _GEN_5509; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5511 = 12'h947 == _T_71[11:0] ? image_2375 : _GEN_5510; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5512 = 12'h948 == _T_71[11:0] ? image_2376 : _GEN_5511; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5513 = 12'h949 == _T_71[11:0] ? image_2377 : _GEN_5512; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5514 = 12'h94a == _T_71[11:0] ? image_2378 : _GEN_5513; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5515 = 12'h94b == _T_71[11:0] ? image_2379 : _GEN_5514; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5516 = 12'h94c == _T_71[11:0] ? image_2380 : _GEN_5515; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5517 = 12'h94d == _T_71[11:0] ? image_2381 : _GEN_5516; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5518 = 12'h94e == _T_71[11:0] ? image_2382 : _GEN_5517; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5519 = 12'h94f == _T_71[11:0] ? image_2383 : _GEN_5518; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5520 = 12'h950 == _T_71[11:0] ? image_2384 : _GEN_5519; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5521 = 12'h951 == _T_71[11:0] ? image_2385 : _GEN_5520; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5522 = 12'h952 == _T_71[11:0] ? image_2386 : _GEN_5521; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5523 = 12'h953 == _T_71[11:0] ? image_2387 : _GEN_5522; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5524 = 12'h954 == _T_71[11:0] ? image_2388 : _GEN_5523; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5525 = 12'h955 == _T_71[11:0] ? image_2389 : _GEN_5524; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5526 = 12'h956 == _T_71[11:0] ? image_2390 : _GEN_5525; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5527 = 12'h957 == _T_71[11:0] ? image_2391 : _GEN_5526; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5528 = 12'h958 == _T_71[11:0] ? image_2392 : _GEN_5527; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5529 = 12'h959 == _T_71[11:0] ? image_2393 : _GEN_5528; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5530 = 12'h95a == _T_71[11:0] ? image_2394 : _GEN_5529; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5531 = 12'h95b == _T_71[11:0] ? image_2395 : _GEN_5530; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5532 = 12'h95c == _T_71[11:0] ? image_2396 : _GEN_5531; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5533 = 12'h95d == _T_71[11:0] ? image_2397 : _GEN_5532; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5534 = 12'h95e == _T_71[11:0] ? image_2398 : _GEN_5533; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5535 = 12'h95f == _T_71[11:0] ? image_2399 : _GEN_5534; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5536 = 12'h960 == _T_71[11:0] ? image_2400 : _GEN_5535; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5537 = 12'h961 == _T_71[11:0] ? image_2401 : _GEN_5536; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5538 = 12'h962 == _T_71[11:0] ? image_2402 : _GEN_5537; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5539 = 12'h963 == _T_71[11:0] ? image_2403 : _GEN_5538; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5540 = 12'h964 == _T_71[11:0] ? image_2404 : _GEN_5539; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5541 = 12'h965 == _T_71[11:0] ? image_2405 : _GEN_5540; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5542 = 12'h966 == _T_71[11:0] ? image_2406 : _GEN_5541; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5543 = 12'h967 == _T_71[11:0] ? image_2407 : _GEN_5542; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5544 = 12'h968 == _T_71[11:0] ? image_2408 : _GEN_5543; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5545 = 12'h969 == _T_71[11:0] ? image_2409 : _GEN_5544; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5546 = 12'h96a == _T_71[11:0] ? image_2410 : _GEN_5545; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5547 = 12'h96b == _T_71[11:0] ? image_2411 : _GEN_5546; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5548 = 12'h96c == _T_71[11:0] ? image_2412 : _GEN_5547; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5549 = 12'h96d == _T_71[11:0] ? image_2413 : _GEN_5548; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5550 = 12'h96e == _T_71[11:0] ? image_2414 : _GEN_5549; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5551 = 12'h96f == _T_71[11:0] ? image_2415 : _GEN_5550; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5552 = 12'h970 == _T_71[11:0] ? image_2416 : _GEN_5551; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5553 = 12'h971 == _T_71[11:0] ? image_2417 : _GEN_5552; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5554 = 12'h972 == _T_71[11:0] ? image_2418 : _GEN_5553; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5555 = 12'h973 == _T_71[11:0] ? image_2419 : _GEN_5554; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5556 = 12'h974 == _T_71[11:0] ? image_2420 : _GEN_5555; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5557 = 12'h975 == _T_71[11:0] ? image_2421 : _GEN_5556; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5558 = 12'h976 == _T_71[11:0] ? image_2422 : _GEN_5557; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5559 = 12'h977 == _T_71[11:0] ? image_2423 : _GEN_5558; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5560 = 12'h978 == _T_71[11:0] ? image_2424 : _GEN_5559; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5561 = 12'h979 == _T_71[11:0] ? image_2425 : _GEN_5560; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5562 = 12'h97a == _T_71[11:0] ? image_2426 : _GEN_5561; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5563 = 12'h97b == _T_71[11:0] ? 4'h0 : _GEN_5562; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5564 = 12'h97c == _T_71[11:0] ? 4'h0 : _GEN_5563; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5565 = 12'h97d == _T_71[11:0] ? 4'h0 : _GEN_5564; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5566 = 12'h97e == _T_71[11:0] ? 4'h0 : _GEN_5565; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5567 = 12'h97f == _T_71[11:0] ? 4'h0 : _GEN_5566; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5568 = 12'h980 == _T_71[11:0] ? 4'h0 : _GEN_5567; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5569 = 12'h981 == _T_71[11:0] ? 4'h0 : _GEN_5568; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5570 = 12'h982 == _T_71[11:0] ? 4'h0 : _GEN_5569; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5571 = 12'h983 == _T_71[11:0] ? 4'h0 : _GEN_5570; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5572 = 12'h984 == _T_71[11:0] ? 4'h0 : _GEN_5571; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5573 = 12'h985 == _T_71[11:0] ? image_2437 : _GEN_5572; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5574 = 12'h986 == _T_71[11:0] ? image_2438 : _GEN_5573; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5575 = 12'h987 == _T_71[11:0] ? image_2439 : _GEN_5574; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5576 = 12'h988 == _T_71[11:0] ? image_2440 : _GEN_5575; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5577 = 12'h989 == _T_71[11:0] ? image_2441 : _GEN_5576; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5578 = 12'h98a == _T_71[11:0] ? image_2442 : _GEN_5577; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5579 = 12'h98b == _T_71[11:0] ? image_2443 : _GEN_5578; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5580 = 12'h98c == _T_71[11:0] ? image_2444 : _GEN_5579; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5581 = 12'h98d == _T_71[11:0] ? image_2445 : _GEN_5580; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5582 = 12'h98e == _T_71[11:0] ? image_2446 : _GEN_5581; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5583 = 12'h98f == _T_71[11:0] ? image_2447 : _GEN_5582; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5584 = 12'h990 == _T_71[11:0] ? image_2448 : _GEN_5583; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5585 = 12'h991 == _T_71[11:0] ? image_2449 : _GEN_5584; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5586 = 12'h992 == _T_71[11:0] ? image_2450 : _GEN_5585; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5587 = 12'h993 == _T_71[11:0] ? image_2451 : _GEN_5586; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5588 = 12'h994 == _T_71[11:0] ? image_2452 : _GEN_5587; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5589 = 12'h995 == _T_71[11:0] ? image_2453 : _GEN_5588; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5590 = 12'h996 == _T_71[11:0] ? image_2454 : _GEN_5589; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5591 = 12'h997 == _T_71[11:0] ? image_2455 : _GEN_5590; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5592 = 12'h998 == _T_71[11:0] ? image_2456 : _GEN_5591; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5593 = 12'h999 == _T_71[11:0] ? image_2457 : _GEN_5592; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5594 = 12'h99a == _T_71[11:0] ? image_2458 : _GEN_5593; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5595 = 12'h99b == _T_71[11:0] ? image_2459 : _GEN_5594; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5596 = 12'h99c == _T_71[11:0] ? image_2460 : _GEN_5595; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5597 = 12'h99d == _T_71[11:0] ? image_2461 : _GEN_5596; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5598 = 12'h99e == _T_71[11:0] ? image_2462 : _GEN_5597; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5599 = 12'h99f == _T_71[11:0] ? image_2463 : _GEN_5598; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5600 = 12'h9a0 == _T_71[11:0] ? image_2464 : _GEN_5599; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5601 = 12'h9a1 == _T_71[11:0] ? image_2465 : _GEN_5600; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5602 = 12'h9a2 == _T_71[11:0] ? image_2466 : _GEN_5601; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5603 = 12'h9a3 == _T_71[11:0] ? image_2467 : _GEN_5602; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5604 = 12'h9a4 == _T_71[11:0] ? image_2468 : _GEN_5603; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5605 = 12'h9a5 == _T_71[11:0] ? image_2469 : _GEN_5604; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5606 = 12'h9a6 == _T_71[11:0] ? image_2470 : _GEN_5605; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5607 = 12'h9a7 == _T_71[11:0] ? image_2471 : _GEN_5606; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5608 = 12'h9a8 == _T_71[11:0] ? image_2472 : _GEN_5607; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5609 = 12'h9a9 == _T_71[11:0] ? image_2473 : _GEN_5608; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5610 = 12'h9aa == _T_71[11:0] ? image_2474 : _GEN_5609; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5611 = 12'h9ab == _T_71[11:0] ? image_2475 : _GEN_5610; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5612 = 12'h9ac == _T_71[11:0] ? image_2476 : _GEN_5611; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5613 = 12'h9ad == _T_71[11:0] ? image_2477 : _GEN_5612; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5614 = 12'h9ae == _T_71[11:0] ? image_2478 : _GEN_5613; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5615 = 12'h9af == _T_71[11:0] ? image_2479 : _GEN_5614; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5616 = 12'h9b0 == _T_71[11:0] ? image_2480 : _GEN_5615; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5617 = 12'h9b1 == _T_71[11:0] ? image_2481 : _GEN_5616; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5618 = 12'h9b2 == _T_71[11:0] ? image_2482 : _GEN_5617; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5619 = 12'h9b3 == _T_71[11:0] ? image_2483 : _GEN_5618; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5620 = 12'h9b4 == _T_71[11:0] ? image_2484 : _GEN_5619; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5621 = 12'h9b5 == _T_71[11:0] ? image_2485 : _GEN_5620; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5622 = 12'h9b6 == _T_71[11:0] ? image_2486 : _GEN_5621; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5623 = 12'h9b7 == _T_71[11:0] ? image_2487 : _GEN_5622; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5624 = 12'h9b8 == _T_71[11:0] ? image_2488 : _GEN_5623; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5625 = 12'h9b9 == _T_71[11:0] ? image_2489 : _GEN_5624; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5626 = 12'h9ba == _T_71[11:0] ? image_2490 : _GEN_5625; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5627 = 12'h9bb == _T_71[11:0] ? 4'h0 : _GEN_5626; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5628 = 12'h9bc == _T_71[11:0] ? 4'h0 : _GEN_5627; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5629 = 12'h9bd == _T_71[11:0] ? 4'h0 : _GEN_5628; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5630 = 12'h9be == _T_71[11:0] ? 4'h0 : _GEN_5629; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5631 = 12'h9bf == _T_71[11:0] ? 4'h0 : _GEN_5630; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5632 = 12'h9c0 == _T_71[11:0] ? 4'h0 : _GEN_5631; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5633 = 12'h9c1 == _T_71[11:0] ? 4'h0 : _GEN_5632; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5634 = 12'h9c2 == _T_71[11:0] ? 4'h0 : _GEN_5633; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5635 = 12'h9c3 == _T_71[11:0] ? 4'h0 : _GEN_5634; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5636 = 12'h9c4 == _T_71[11:0] ? 4'h0 : _GEN_5635; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5637 = 12'h9c5 == _T_71[11:0] ? 4'h0 : _GEN_5636; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5638 = 12'h9c6 == _T_71[11:0] ? image_2502 : _GEN_5637; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5639 = 12'h9c7 == _T_71[11:0] ? image_2503 : _GEN_5638; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5640 = 12'h9c8 == _T_71[11:0] ? image_2504 : _GEN_5639; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5641 = 12'h9c9 == _T_71[11:0] ? image_2505 : _GEN_5640; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5642 = 12'h9ca == _T_71[11:0] ? image_2506 : _GEN_5641; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5643 = 12'h9cb == _T_71[11:0] ? image_2507 : _GEN_5642; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5644 = 12'h9cc == _T_71[11:0] ? image_2508 : _GEN_5643; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5645 = 12'h9cd == _T_71[11:0] ? image_2509 : _GEN_5644; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5646 = 12'h9ce == _T_71[11:0] ? image_2510 : _GEN_5645; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5647 = 12'h9cf == _T_71[11:0] ? image_2511 : _GEN_5646; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5648 = 12'h9d0 == _T_71[11:0] ? image_2512 : _GEN_5647; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5649 = 12'h9d1 == _T_71[11:0] ? image_2513 : _GEN_5648; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5650 = 12'h9d2 == _T_71[11:0] ? image_2514 : _GEN_5649; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5651 = 12'h9d3 == _T_71[11:0] ? image_2515 : _GEN_5650; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5652 = 12'h9d4 == _T_71[11:0] ? image_2516 : _GEN_5651; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5653 = 12'h9d5 == _T_71[11:0] ? image_2517 : _GEN_5652; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5654 = 12'h9d6 == _T_71[11:0] ? image_2518 : _GEN_5653; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5655 = 12'h9d7 == _T_71[11:0] ? image_2519 : _GEN_5654; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5656 = 12'h9d8 == _T_71[11:0] ? image_2520 : _GEN_5655; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5657 = 12'h9d9 == _T_71[11:0] ? image_2521 : _GEN_5656; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5658 = 12'h9da == _T_71[11:0] ? image_2522 : _GEN_5657; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5659 = 12'h9db == _T_71[11:0] ? image_2523 : _GEN_5658; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5660 = 12'h9dc == _T_71[11:0] ? image_2524 : _GEN_5659; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5661 = 12'h9dd == _T_71[11:0] ? image_2525 : _GEN_5660; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5662 = 12'h9de == _T_71[11:0] ? image_2526 : _GEN_5661; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5663 = 12'h9df == _T_71[11:0] ? image_2527 : _GEN_5662; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5664 = 12'h9e0 == _T_71[11:0] ? image_2528 : _GEN_5663; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5665 = 12'h9e1 == _T_71[11:0] ? image_2529 : _GEN_5664; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5666 = 12'h9e2 == _T_71[11:0] ? image_2530 : _GEN_5665; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5667 = 12'h9e3 == _T_71[11:0] ? image_2531 : _GEN_5666; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5668 = 12'h9e4 == _T_71[11:0] ? image_2532 : _GEN_5667; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5669 = 12'h9e5 == _T_71[11:0] ? image_2533 : _GEN_5668; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5670 = 12'h9e6 == _T_71[11:0] ? image_2534 : _GEN_5669; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5671 = 12'h9e7 == _T_71[11:0] ? image_2535 : _GEN_5670; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5672 = 12'h9e8 == _T_71[11:0] ? image_2536 : _GEN_5671; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5673 = 12'h9e9 == _T_71[11:0] ? image_2537 : _GEN_5672; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5674 = 12'h9ea == _T_71[11:0] ? image_2538 : _GEN_5673; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5675 = 12'h9eb == _T_71[11:0] ? image_2539 : _GEN_5674; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5676 = 12'h9ec == _T_71[11:0] ? image_2540 : _GEN_5675; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5677 = 12'h9ed == _T_71[11:0] ? image_2541 : _GEN_5676; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5678 = 12'h9ee == _T_71[11:0] ? image_2542 : _GEN_5677; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5679 = 12'h9ef == _T_71[11:0] ? image_2543 : _GEN_5678; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5680 = 12'h9f0 == _T_71[11:0] ? image_2544 : _GEN_5679; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5681 = 12'h9f1 == _T_71[11:0] ? image_2545 : _GEN_5680; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5682 = 12'h9f2 == _T_71[11:0] ? image_2546 : _GEN_5681; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5683 = 12'h9f3 == _T_71[11:0] ? image_2547 : _GEN_5682; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5684 = 12'h9f4 == _T_71[11:0] ? image_2548 : _GEN_5683; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5685 = 12'h9f5 == _T_71[11:0] ? image_2549 : _GEN_5684; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5686 = 12'h9f6 == _T_71[11:0] ? image_2550 : _GEN_5685; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5687 = 12'h9f7 == _T_71[11:0] ? image_2551 : _GEN_5686; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5688 = 12'h9f8 == _T_71[11:0] ? image_2552 : _GEN_5687; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5689 = 12'h9f9 == _T_71[11:0] ? image_2553 : _GEN_5688; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5690 = 12'h9fa == _T_71[11:0] ? image_2554 : _GEN_5689; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5691 = 12'h9fb == _T_71[11:0] ? 4'h0 : _GEN_5690; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5692 = 12'h9fc == _T_71[11:0] ? 4'h0 : _GEN_5691; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5693 = 12'h9fd == _T_71[11:0] ? 4'h0 : _GEN_5692; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5694 = 12'h9fe == _T_71[11:0] ? 4'h0 : _GEN_5693; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5695 = 12'h9ff == _T_71[11:0] ? 4'h0 : _GEN_5694; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5696 = 12'ha00 == _T_71[11:0] ? 4'h0 : _GEN_5695; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5697 = 12'ha01 == _T_71[11:0] ? 4'h0 : _GEN_5696; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5698 = 12'ha02 == _T_71[11:0] ? 4'h0 : _GEN_5697; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5699 = 12'ha03 == _T_71[11:0] ? 4'h0 : _GEN_5698; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5700 = 12'ha04 == _T_71[11:0] ? 4'h0 : _GEN_5699; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5701 = 12'ha05 == _T_71[11:0] ? 4'h0 : _GEN_5700; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5702 = 12'ha06 == _T_71[11:0] ? 4'h0 : _GEN_5701; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5703 = 12'ha07 == _T_71[11:0] ? image_2567 : _GEN_5702; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5704 = 12'ha08 == _T_71[11:0] ? image_2568 : _GEN_5703; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5705 = 12'ha09 == _T_71[11:0] ? image_2569 : _GEN_5704; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5706 = 12'ha0a == _T_71[11:0] ? image_2570 : _GEN_5705; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5707 = 12'ha0b == _T_71[11:0] ? image_2571 : _GEN_5706; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5708 = 12'ha0c == _T_71[11:0] ? image_2572 : _GEN_5707; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5709 = 12'ha0d == _T_71[11:0] ? image_2573 : _GEN_5708; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5710 = 12'ha0e == _T_71[11:0] ? image_2574 : _GEN_5709; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5711 = 12'ha0f == _T_71[11:0] ? image_2575 : _GEN_5710; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5712 = 12'ha10 == _T_71[11:0] ? image_2576 : _GEN_5711; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5713 = 12'ha11 == _T_71[11:0] ? image_2577 : _GEN_5712; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5714 = 12'ha12 == _T_71[11:0] ? image_2578 : _GEN_5713; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5715 = 12'ha13 == _T_71[11:0] ? image_2579 : _GEN_5714; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5716 = 12'ha14 == _T_71[11:0] ? image_2580 : _GEN_5715; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5717 = 12'ha15 == _T_71[11:0] ? image_2581 : _GEN_5716; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5718 = 12'ha16 == _T_71[11:0] ? image_2582 : _GEN_5717; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5719 = 12'ha17 == _T_71[11:0] ? image_2583 : _GEN_5718; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5720 = 12'ha18 == _T_71[11:0] ? image_2584 : _GEN_5719; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5721 = 12'ha19 == _T_71[11:0] ? image_2585 : _GEN_5720; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5722 = 12'ha1a == _T_71[11:0] ? image_2586 : _GEN_5721; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5723 = 12'ha1b == _T_71[11:0] ? image_2587 : _GEN_5722; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5724 = 12'ha1c == _T_71[11:0] ? image_2588 : _GEN_5723; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5725 = 12'ha1d == _T_71[11:0] ? image_2589 : _GEN_5724; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5726 = 12'ha1e == _T_71[11:0] ? image_2590 : _GEN_5725; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5727 = 12'ha1f == _T_71[11:0] ? image_2591 : _GEN_5726; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5728 = 12'ha20 == _T_71[11:0] ? image_2592 : _GEN_5727; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5729 = 12'ha21 == _T_71[11:0] ? image_2593 : _GEN_5728; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5730 = 12'ha22 == _T_71[11:0] ? image_2594 : _GEN_5729; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5731 = 12'ha23 == _T_71[11:0] ? image_2595 : _GEN_5730; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5732 = 12'ha24 == _T_71[11:0] ? image_2596 : _GEN_5731; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5733 = 12'ha25 == _T_71[11:0] ? image_2597 : _GEN_5732; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5734 = 12'ha26 == _T_71[11:0] ? image_2598 : _GEN_5733; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5735 = 12'ha27 == _T_71[11:0] ? image_2599 : _GEN_5734; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5736 = 12'ha28 == _T_71[11:0] ? image_2600 : _GEN_5735; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5737 = 12'ha29 == _T_71[11:0] ? image_2601 : _GEN_5736; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5738 = 12'ha2a == _T_71[11:0] ? image_2602 : _GEN_5737; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5739 = 12'ha2b == _T_71[11:0] ? image_2603 : _GEN_5738; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5740 = 12'ha2c == _T_71[11:0] ? image_2604 : _GEN_5739; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5741 = 12'ha2d == _T_71[11:0] ? image_2605 : _GEN_5740; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5742 = 12'ha2e == _T_71[11:0] ? image_2606 : _GEN_5741; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5743 = 12'ha2f == _T_71[11:0] ? image_2607 : _GEN_5742; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5744 = 12'ha30 == _T_71[11:0] ? image_2608 : _GEN_5743; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5745 = 12'ha31 == _T_71[11:0] ? image_2609 : _GEN_5744; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5746 = 12'ha32 == _T_71[11:0] ? image_2610 : _GEN_5745; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5747 = 12'ha33 == _T_71[11:0] ? image_2611 : _GEN_5746; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5748 = 12'ha34 == _T_71[11:0] ? image_2612 : _GEN_5747; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5749 = 12'ha35 == _T_71[11:0] ? image_2613 : _GEN_5748; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5750 = 12'ha36 == _T_71[11:0] ? image_2614 : _GEN_5749; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5751 = 12'ha37 == _T_71[11:0] ? image_2615 : _GEN_5750; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5752 = 12'ha38 == _T_71[11:0] ? image_2616 : _GEN_5751; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5753 = 12'ha39 == _T_71[11:0] ? image_2617 : _GEN_5752; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5754 = 12'ha3a == _T_71[11:0] ? image_2618 : _GEN_5753; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5755 = 12'ha3b == _T_71[11:0] ? 4'h0 : _GEN_5754; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5756 = 12'ha3c == _T_71[11:0] ? 4'h0 : _GEN_5755; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5757 = 12'ha3d == _T_71[11:0] ? 4'h0 : _GEN_5756; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5758 = 12'ha3e == _T_71[11:0] ? 4'h0 : _GEN_5757; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5759 = 12'ha3f == _T_71[11:0] ? 4'h0 : _GEN_5758; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5760 = 12'ha40 == _T_71[11:0] ? 4'h0 : _GEN_5759; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5761 = 12'ha41 == _T_71[11:0] ? 4'h0 : _GEN_5760; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5762 = 12'ha42 == _T_71[11:0] ? 4'h0 : _GEN_5761; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5763 = 12'ha43 == _T_71[11:0] ? 4'h0 : _GEN_5762; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5764 = 12'ha44 == _T_71[11:0] ? 4'h0 : _GEN_5763; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5765 = 12'ha45 == _T_71[11:0] ? 4'h0 : _GEN_5764; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5766 = 12'ha46 == _T_71[11:0] ? 4'h0 : _GEN_5765; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5767 = 12'ha47 == _T_71[11:0] ? 4'h0 : _GEN_5766; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5768 = 12'ha48 == _T_71[11:0] ? image_2632 : _GEN_5767; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5769 = 12'ha49 == _T_71[11:0] ? image_2633 : _GEN_5768; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5770 = 12'ha4a == _T_71[11:0] ? image_2634 : _GEN_5769; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5771 = 12'ha4b == _T_71[11:0] ? image_2635 : _GEN_5770; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5772 = 12'ha4c == _T_71[11:0] ? image_2636 : _GEN_5771; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5773 = 12'ha4d == _T_71[11:0] ? image_2637 : _GEN_5772; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5774 = 12'ha4e == _T_71[11:0] ? image_2638 : _GEN_5773; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5775 = 12'ha4f == _T_71[11:0] ? image_2639 : _GEN_5774; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5776 = 12'ha50 == _T_71[11:0] ? image_2640 : _GEN_5775; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5777 = 12'ha51 == _T_71[11:0] ? image_2641 : _GEN_5776; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5778 = 12'ha52 == _T_71[11:0] ? image_2642 : _GEN_5777; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5779 = 12'ha53 == _T_71[11:0] ? image_2643 : _GEN_5778; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5780 = 12'ha54 == _T_71[11:0] ? image_2644 : _GEN_5779; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5781 = 12'ha55 == _T_71[11:0] ? image_2645 : _GEN_5780; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5782 = 12'ha56 == _T_71[11:0] ? image_2646 : _GEN_5781; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5783 = 12'ha57 == _T_71[11:0] ? image_2647 : _GEN_5782; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5784 = 12'ha58 == _T_71[11:0] ? image_2648 : _GEN_5783; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5785 = 12'ha59 == _T_71[11:0] ? image_2649 : _GEN_5784; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5786 = 12'ha5a == _T_71[11:0] ? image_2650 : _GEN_5785; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5787 = 12'ha5b == _T_71[11:0] ? image_2651 : _GEN_5786; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5788 = 12'ha5c == _T_71[11:0] ? image_2652 : _GEN_5787; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5789 = 12'ha5d == _T_71[11:0] ? image_2653 : _GEN_5788; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5790 = 12'ha5e == _T_71[11:0] ? image_2654 : _GEN_5789; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5791 = 12'ha5f == _T_71[11:0] ? image_2655 : _GEN_5790; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5792 = 12'ha60 == _T_71[11:0] ? image_2656 : _GEN_5791; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5793 = 12'ha61 == _T_71[11:0] ? image_2657 : _GEN_5792; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5794 = 12'ha62 == _T_71[11:0] ? image_2658 : _GEN_5793; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5795 = 12'ha63 == _T_71[11:0] ? image_2659 : _GEN_5794; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5796 = 12'ha64 == _T_71[11:0] ? image_2660 : _GEN_5795; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5797 = 12'ha65 == _T_71[11:0] ? image_2661 : _GEN_5796; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5798 = 12'ha66 == _T_71[11:0] ? image_2662 : _GEN_5797; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5799 = 12'ha67 == _T_71[11:0] ? image_2663 : _GEN_5798; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5800 = 12'ha68 == _T_71[11:0] ? image_2664 : _GEN_5799; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5801 = 12'ha69 == _T_71[11:0] ? image_2665 : _GEN_5800; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5802 = 12'ha6a == _T_71[11:0] ? image_2666 : _GEN_5801; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5803 = 12'ha6b == _T_71[11:0] ? image_2667 : _GEN_5802; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5804 = 12'ha6c == _T_71[11:0] ? image_2668 : _GEN_5803; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5805 = 12'ha6d == _T_71[11:0] ? image_2669 : _GEN_5804; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5806 = 12'ha6e == _T_71[11:0] ? image_2670 : _GEN_5805; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5807 = 12'ha6f == _T_71[11:0] ? image_2671 : _GEN_5806; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5808 = 12'ha70 == _T_71[11:0] ? image_2672 : _GEN_5807; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5809 = 12'ha71 == _T_71[11:0] ? image_2673 : _GEN_5808; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5810 = 12'ha72 == _T_71[11:0] ? image_2674 : _GEN_5809; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5811 = 12'ha73 == _T_71[11:0] ? image_2675 : _GEN_5810; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5812 = 12'ha74 == _T_71[11:0] ? image_2676 : _GEN_5811; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5813 = 12'ha75 == _T_71[11:0] ? image_2677 : _GEN_5812; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5814 = 12'ha76 == _T_71[11:0] ? image_2678 : _GEN_5813; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5815 = 12'ha77 == _T_71[11:0] ? image_2679 : _GEN_5814; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5816 = 12'ha78 == _T_71[11:0] ? image_2680 : _GEN_5815; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5817 = 12'ha79 == _T_71[11:0] ? image_2681 : _GEN_5816; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5818 = 12'ha7a == _T_71[11:0] ? image_2682 : _GEN_5817; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5819 = 12'ha7b == _T_71[11:0] ? 4'h0 : _GEN_5818; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5820 = 12'ha7c == _T_71[11:0] ? 4'h0 : _GEN_5819; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5821 = 12'ha7d == _T_71[11:0] ? 4'h0 : _GEN_5820; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5822 = 12'ha7e == _T_71[11:0] ? 4'h0 : _GEN_5821; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5823 = 12'ha7f == _T_71[11:0] ? 4'h0 : _GEN_5822; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5824 = 12'ha80 == _T_71[11:0] ? 4'h0 : _GEN_5823; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5825 = 12'ha81 == _T_71[11:0] ? 4'h0 : _GEN_5824; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5826 = 12'ha82 == _T_71[11:0] ? 4'h0 : _GEN_5825; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5827 = 12'ha83 == _T_71[11:0] ? 4'h0 : _GEN_5826; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5828 = 12'ha84 == _T_71[11:0] ? 4'h0 : _GEN_5827; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5829 = 12'ha85 == _T_71[11:0] ? 4'h0 : _GEN_5828; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5830 = 12'ha86 == _T_71[11:0] ? 4'h0 : _GEN_5829; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5831 = 12'ha87 == _T_71[11:0] ? 4'h0 : _GEN_5830; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5832 = 12'ha88 == _T_71[11:0] ? 4'h0 : _GEN_5831; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5833 = 12'ha89 == _T_71[11:0] ? image_2697 : _GEN_5832; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5834 = 12'ha8a == _T_71[11:0] ? image_2698 : _GEN_5833; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5835 = 12'ha8b == _T_71[11:0] ? image_2699 : _GEN_5834; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5836 = 12'ha8c == _T_71[11:0] ? image_2700 : _GEN_5835; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5837 = 12'ha8d == _T_71[11:0] ? image_2701 : _GEN_5836; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5838 = 12'ha8e == _T_71[11:0] ? image_2702 : _GEN_5837; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5839 = 12'ha8f == _T_71[11:0] ? image_2703 : _GEN_5838; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5840 = 12'ha90 == _T_71[11:0] ? image_2704 : _GEN_5839; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5841 = 12'ha91 == _T_71[11:0] ? image_2705 : _GEN_5840; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5842 = 12'ha92 == _T_71[11:0] ? image_2706 : _GEN_5841; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5843 = 12'ha93 == _T_71[11:0] ? image_2707 : _GEN_5842; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5844 = 12'ha94 == _T_71[11:0] ? image_2708 : _GEN_5843; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5845 = 12'ha95 == _T_71[11:0] ? image_2709 : _GEN_5844; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5846 = 12'ha96 == _T_71[11:0] ? image_2710 : _GEN_5845; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5847 = 12'ha97 == _T_71[11:0] ? image_2711 : _GEN_5846; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5848 = 12'ha98 == _T_71[11:0] ? image_2712 : _GEN_5847; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5849 = 12'ha99 == _T_71[11:0] ? image_2713 : _GEN_5848; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5850 = 12'ha9a == _T_71[11:0] ? image_2714 : _GEN_5849; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5851 = 12'ha9b == _T_71[11:0] ? image_2715 : _GEN_5850; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5852 = 12'ha9c == _T_71[11:0] ? image_2716 : _GEN_5851; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5853 = 12'ha9d == _T_71[11:0] ? image_2717 : _GEN_5852; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5854 = 12'ha9e == _T_71[11:0] ? image_2718 : _GEN_5853; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5855 = 12'ha9f == _T_71[11:0] ? image_2719 : _GEN_5854; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5856 = 12'haa0 == _T_71[11:0] ? image_2720 : _GEN_5855; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5857 = 12'haa1 == _T_71[11:0] ? image_2721 : _GEN_5856; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5858 = 12'haa2 == _T_71[11:0] ? image_2722 : _GEN_5857; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5859 = 12'haa3 == _T_71[11:0] ? image_2723 : _GEN_5858; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5860 = 12'haa4 == _T_71[11:0] ? image_2724 : _GEN_5859; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5861 = 12'haa5 == _T_71[11:0] ? image_2725 : _GEN_5860; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5862 = 12'haa6 == _T_71[11:0] ? image_2726 : _GEN_5861; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5863 = 12'haa7 == _T_71[11:0] ? image_2727 : _GEN_5862; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5864 = 12'haa8 == _T_71[11:0] ? image_2728 : _GEN_5863; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5865 = 12'haa9 == _T_71[11:0] ? image_2729 : _GEN_5864; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5866 = 12'haaa == _T_71[11:0] ? image_2730 : _GEN_5865; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5867 = 12'haab == _T_71[11:0] ? image_2731 : _GEN_5866; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5868 = 12'haac == _T_71[11:0] ? image_2732 : _GEN_5867; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5869 = 12'haad == _T_71[11:0] ? image_2733 : _GEN_5868; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5870 = 12'haae == _T_71[11:0] ? image_2734 : _GEN_5869; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5871 = 12'haaf == _T_71[11:0] ? image_2735 : _GEN_5870; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5872 = 12'hab0 == _T_71[11:0] ? image_2736 : _GEN_5871; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5873 = 12'hab1 == _T_71[11:0] ? image_2737 : _GEN_5872; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5874 = 12'hab2 == _T_71[11:0] ? image_2738 : _GEN_5873; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5875 = 12'hab3 == _T_71[11:0] ? image_2739 : _GEN_5874; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5876 = 12'hab4 == _T_71[11:0] ? image_2740 : _GEN_5875; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5877 = 12'hab5 == _T_71[11:0] ? image_2741 : _GEN_5876; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5878 = 12'hab6 == _T_71[11:0] ? image_2742 : _GEN_5877; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5879 = 12'hab7 == _T_71[11:0] ? image_2743 : _GEN_5878; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5880 = 12'hab8 == _T_71[11:0] ? image_2744 : _GEN_5879; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5881 = 12'hab9 == _T_71[11:0] ? image_2745 : _GEN_5880; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5882 = 12'haba == _T_71[11:0] ? 4'h0 : _GEN_5881; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5883 = 12'habb == _T_71[11:0] ? 4'h0 : _GEN_5882; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5884 = 12'habc == _T_71[11:0] ? 4'h0 : _GEN_5883; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5885 = 12'habd == _T_71[11:0] ? 4'h0 : _GEN_5884; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5886 = 12'habe == _T_71[11:0] ? 4'h0 : _GEN_5885; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5887 = 12'habf == _T_71[11:0] ? 4'h0 : _GEN_5886; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5888 = 12'hac0 == _T_71[11:0] ? 4'h0 : _GEN_5887; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5889 = 12'hac1 == _T_71[11:0] ? 4'h0 : _GEN_5888; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5890 = 12'hac2 == _T_71[11:0] ? 4'h0 : _GEN_5889; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5891 = 12'hac3 == _T_71[11:0] ? 4'h0 : _GEN_5890; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5892 = 12'hac4 == _T_71[11:0] ? 4'h0 : _GEN_5891; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5893 = 12'hac5 == _T_71[11:0] ? 4'h0 : _GEN_5892; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5894 = 12'hac6 == _T_71[11:0] ? 4'h0 : _GEN_5893; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5895 = 12'hac7 == _T_71[11:0] ? 4'h0 : _GEN_5894; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5896 = 12'hac8 == _T_71[11:0] ? 4'h0 : _GEN_5895; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5897 = 12'hac9 == _T_71[11:0] ? 4'h0 : _GEN_5896; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5898 = 12'haca == _T_71[11:0] ? 4'h0 : _GEN_5897; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5899 = 12'hacb == _T_71[11:0] ? image_2763 : _GEN_5898; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5900 = 12'hacc == _T_71[11:0] ? image_2764 : _GEN_5899; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5901 = 12'hacd == _T_71[11:0] ? image_2765 : _GEN_5900; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5902 = 12'hace == _T_71[11:0] ? image_2766 : _GEN_5901; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5903 = 12'hacf == _T_71[11:0] ? image_2767 : _GEN_5902; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5904 = 12'had0 == _T_71[11:0] ? image_2768 : _GEN_5903; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5905 = 12'had1 == _T_71[11:0] ? image_2769 : _GEN_5904; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5906 = 12'had2 == _T_71[11:0] ? image_2770 : _GEN_5905; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5907 = 12'had3 == _T_71[11:0] ? image_2771 : _GEN_5906; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5908 = 12'had4 == _T_71[11:0] ? image_2772 : _GEN_5907; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5909 = 12'had5 == _T_71[11:0] ? image_2773 : _GEN_5908; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5910 = 12'had6 == _T_71[11:0] ? image_2774 : _GEN_5909; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5911 = 12'had7 == _T_71[11:0] ? image_2775 : _GEN_5910; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5912 = 12'had8 == _T_71[11:0] ? image_2776 : _GEN_5911; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5913 = 12'had9 == _T_71[11:0] ? image_2777 : _GEN_5912; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5914 = 12'hada == _T_71[11:0] ? image_2778 : _GEN_5913; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5915 = 12'hadb == _T_71[11:0] ? image_2779 : _GEN_5914; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5916 = 12'hadc == _T_71[11:0] ? image_2780 : _GEN_5915; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5917 = 12'hadd == _T_71[11:0] ? image_2781 : _GEN_5916; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5918 = 12'hade == _T_71[11:0] ? image_2782 : _GEN_5917; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5919 = 12'hadf == _T_71[11:0] ? image_2783 : _GEN_5918; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5920 = 12'hae0 == _T_71[11:0] ? image_2784 : _GEN_5919; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5921 = 12'hae1 == _T_71[11:0] ? image_2785 : _GEN_5920; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5922 = 12'hae2 == _T_71[11:0] ? image_2786 : _GEN_5921; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5923 = 12'hae3 == _T_71[11:0] ? image_2787 : _GEN_5922; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5924 = 12'hae4 == _T_71[11:0] ? image_2788 : _GEN_5923; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5925 = 12'hae5 == _T_71[11:0] ? image_2789 : _GEN_5924; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5926 = 12'hae6 == _T_71[11:0] ? image_2790 : _GEN_5925; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5927 = 12'hae7 == _T_71[11:0] ? image_2791 : _GEN_5926; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5928 = 12'hae8 == _T_71[11:0] ? image_2792 : _GEN_5927; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5929 = 12'hae9 == _T_71[11:0] ? image_2793 : _GEN_5928; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5930 = 12'haea == _T_71[11:0] ? image_2794 : _GEN_5929; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5931 = 12'haeb == _T_71[11:0] ? image_2795 : _GEN_5930; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5932 = 12'haec == _T_71[11:0] ? image_2796 : _GEN_5931; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5933 = 12'haed == _T_71[11:0] ? image_2797 : _GEN_5932; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5934 = 12'haee == _T_71[11:0] ? image_2798 : _GEN_5933; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5935 = 12'haef == _T_71[11:0] ? image_2799 : _GEN_5934; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5936 = 12'haf0 == _T_71[11:0] ? image_2800 : _GEN_5935; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5937 = 12'haf1 == _T_71[11:0] ? image_2801 : _GEN_5936; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5938 = 12'haf2 == _T_71[11:0] ? image_2802 : _GEN_5937; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5939 = 12'haf3 == _T_71[11:0] ? image_2803 : _GEN_5938; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5940 = 12'haf4 == _T_71[11:0] ? image_2804 : _GEN_5939; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5941 = 12'haf5 == _T_71[11:0] ? image_2805 : _GEN_5940; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5942 = 12'haf6 == _T_71[11:0] ? image_2806 : _GEN_5941; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5943 = 12'haf7 == _T_71[11:0] ? image_2807 : _GEN_5942; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5944 = 12'haf8 == _T_71[11:0] ? image_2808 : _GEN_5943; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5945 = 12'haf9 == _T_71[11:0] ? 4'h0 : _GEN_5944; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5946 = 12'hafa == _T_71[11:0] ? 4'h0 : _GEN_5945; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5947 = 12'hafb == _T_71[11:0] ? 4'h0 : _GEN_5946; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5948 = 12'hafc == _T_71[11:0] ? 4'h0 : _GEN_5947; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5949 = 12'hafd == _T_71[11:0] ? 4'h0 : _GEN_5948; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5950 = 12'hafe == _T_71[11:0] ? 4'h0 : _GEN_5949; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5951 = 12'haff == _T_71[11:0] ? 4'h0 : _GEN_5950; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5952 = 12'hb00 == _T_71[11:0] ? 4'h0 : _GEN_5951; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5953 = 12'hb01 == _T_71[11:0] ? 4'h0 : _GEN_5952; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5954 = 12'hb02 == _T_71[11:0] ? 4'h0 : _GEN_5953; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5955 = 12'hb03 == _T_71[11:0] ? 4'h0 : _GEN_5954; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5956 = 12'hb04 == _T_71[11:0] ? 4'h0 : _GEN_5955; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5957 = 12'hb05 == _T_71[11:0] ? 4'h0 : _GEN_5956; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5958 = 12'hb06 == _T_71[11:0] ? 4'h0 : _GEN_5957; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5959 = 12'hb07 == _T_71[11:0] ? 4'h0 : _GEN_5958; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5960 = 12'hb08 == _T_71[11:0] ? 4'h0 : _GEN_5959; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5961 = 12'hb09 == _T_71[11:0] ? 4'h0 : _GEN_5960; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5962 = 12'hb0a == _T_71[11:0] ? 4'h0 : _GEN_5961; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5963 = 12'hb0b == _T_71[11:0] ? 4'h0 : _GEN_5962; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5964 = 12'hb0c == _T_71[11:0] ? image_2828 : _GEN_5963; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5965 = 12'hb0d == _T_71[11:0] ? image_2829 : _GEN_5964; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5966 = 12'hb0e == _T_71[11:0] ? image_2830 : _GEN_5965; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5967 = 12'hb0f == _T_71[11:0] ? image_2831 : _GEN_5966; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5968 = 12'hb10 == _T_71[11:0] ? image_2832 : _GEN_5967; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5969 = 12'hb11 == _T_71[11:0] ? image_2833 : _GEN_5968; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5970 = 12'hb12 == _T_71[11:0] ? image_2834 : _GEN_5969; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5971 = 12'hb13 == _T_71[11:0] ? image_2835 : _GEN_5970; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5972 = 12'hb14 == _T_71[11:0] ? image_2836 : _GEN_5971; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5973 = 12'hb15 == _T_71[11:0] ? image_2837 : _GEN_5972; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5974 = 12'hb16 == _T_71[11:0] ? image_2838 : _GEN_5973; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5975 = 12'hb17 == _T_71[11:0] ? image_2839 : _GEN_5974; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5976 = 12'hb18 == _T_71[11:0] ? image_2840 : _GEN_5975; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5977 = 12'hb19 == _T_71[11:0] ? image_2841 : _GEN_5976; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5978 = 12'hb1a == _T_71[11:0] ? image_2842 : _GEN_5977; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5979 = 12'hb1b == _T_71[11:0] ? image_2843 : _GEN_5978; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5980 = 12'hb1c == _T_71[11:0] ? image_2844 : _GEN_5979; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5981 = 12'hb1d == _T_71[11:0] ? image_2845 : _GEN_5980; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5982 = 12'hb1e == _T_71[11:0] ? image_2846 : _GEN_5981; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5983 = 12'hb1f == _T_71[11:0] ? image_2847 : _GEN_5982; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5984 = 12'hb20 == _T_71[11:0] ? image_2848 : _GEN_5983; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5985 = 12'hb21 == _T_71[11:0] ? image_2849 : _GEN_5984; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5986 = 12'hb22 == _T_71[11:0] ? image_2850 : _GEN_5985; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5987 = 12'hb23 == _T_71[11:0] ? image_2851 : _GEN_5986; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5988 = 12'hb24 == _T_71[11:0] ? image_2852 : _GEN_5987; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5989 = 12'hb25 == _T_71[11:0] ? image_2853 : _GEN_5988; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5990 = 12'hb26 == _T_71[11:0] ? image_2854 : _GEN_5989; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5991 = 12'hb27 == _T_71[11:0] ? image_2855 : _GEN_5990; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5992 = 12'hb28 == _T_71[11:0] ? image_2856 : _GEN_5991; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5993 = 12'hb29 == _T_71[11:0] ? image_2857 : _GEN_5992; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5994 = 12'hb2a == _T_71[11:0] ? image_2858 : _GEN_5993; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5995 = 12'hb2b == _T_71[11:0] ? image_2859 : _GEN_5994; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5996 = 12'hb2c == _T_71[11:0] ? image_2860 : _GEN_5995; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5997 = 12'hb2d == _T_71[11:0] ? image_2861 : _GEN_5996; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5998 = 12'hb2e == _T_71[11:0] ? image_2862 : _GEN_5997; // @[Filter.scala 138:46]
  wire [3:0] _GEN_5999 = 12'hb2f == _T_71[11:0] ? image_2863 : _GEN_5998; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6000 = 12'hb30 == _T_71[11:0] ? image_2864 : _GEN_5999; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6001 = 12'hb31 == _T_71[11:0] ? image_2865 : _GEN_6000; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6002 = 12'hb32 == _T_71[11:0] ? image_2866 : _GEN_6001; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6003 = 12'hb33 == _T_71[11:0] ? image_2867 : _GEN_6002; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6004 = 12'hb34 == _T_71[11:0] ? image_2868 : _GEN_6003; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6005 = 12'hb35 == _T_71[11:0] ? image_2869 : _GEN_6004; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6006 = 12'hb36 == _T_71[11:0] ? image_2870 : _GEN_6005; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6007 = 12'hb37 == _T_71[11:0] ? image_2871 : _GEN_6006; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6008 = 12'hb38 == _T_71[11:0] ? 4'h0 : _GEN_6007; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6009 = 12'hb39 == _T_71[11:0] ? 4'h0 : _GEN_6008; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6010 = 12'hb3a == _T_71[11:0] ? 4'h0 : _GEN_6009; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6011 = 12'hb3b == _T_71[11:0] ? 4'h0 : _GEN_6010; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6012 = 12'hb3c == _T_71[11:0] ? 4'h0 : _GEN_6011; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6013 = 12'hb3d == _T_71[11:0] ? 4'h0 : _GEN_6012; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6014 = 12'hb3e == _T_71[11:0] ? 4'h0 : _GEN_6013; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6015 = 12'hb3f == _T_71[11:0] ? 4'h0 : _GEN_6014; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6016 = 12'hb40 == _T_71[11:0] ? 4'h0 : _GEN_6015; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6017 = 12'hb41 == _T_71[11:0] ? 4'h0 : _GEN_6016; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6018 = 12'hb42 == _T_71[11:0] ? 4'h0 : _GEN_6017; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6019 = 12'hb43 == _T_71[11:0] ? 4'h0 : _GEN_6018; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6020 = 12'hb44 == _T_71[11:0] ? 4'h0 : _GEN_6019; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6021 = 12'hb45 == _T_71[11:0] ? 4'h0 : _GEN_6020; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6022 = 12'hb46 == _T_71[11:0] ? 4'h0 : _GEN_6021; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6023 = 12'hb47 == _T_71[11:0] ? 4'h0 : _GEN_6022; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6024 = 12'hb48 == _T_71[11:0] ? 4'h0 : _GEN_6023; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6025 = 12'hb49 == _T_71[11:0] ? 4'h0 : _GEN_6024; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6026 = 12'hb4a == _T_71[11:0] ? 4'h0 : _GEN_6025; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6027 = 12'hb4b == _T_71[11:0] ? 4'h0 : _GEN_6026; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6028 = 12'hb4c == _T_71[11:0] ? 4'h0 : _GEN_6027; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6029 = 12'hb4d == _T_71[11:0] ? 4'h0 : _GEN_6028; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6030 = 12'hb4e == _T_71[11:0] ? 4'h0 : _GEN_6029; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6031 = 12'hb4f == _T_71[11:0] ? image_2895 : _GEN_6030; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6032 = 12'hb50 == _T_71[11:0] ? image_2896 : _GEN_6031; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6033 = 12'hb51 == _T_71[11:0] ? image_2897 : _GEN_6032; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6034 = 12'hb52 == _T_71[11:0] ? image_2898 : _GEN_6033; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6035 = 12'hb53 == _T_71[11:0] ? image_2899 : _GEN_6034; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6036 = 12'hb54 == _T_71[11:0] ? image_2900 : _GEN_6035; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6037 = 12'hb55 == _T_71[11:0] ? image_2901 : _GEN_6036; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6038 = 12'hb56 == _T_71[11:0] ? image_2902 : _GEN_6037; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6039 = 12'hb57 == _T_71[11:0] ? image_2903 : _GEN_6038; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6040 = 12'hb58 == _T_71[11:0] ? image_2904 : _GEN_6039; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6041 = 12'hb59 == _T_71[11:0] ? image_2905 : _GEN_6040; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6042 = 12'hb5a == _T_71[11:0] ? image_2906 : _GEN_6041; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6043 = 12'hb5b == _T_71[11:0] ? image_2907 : _GEN_6042; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6044 = 12'hb5c == _T_71[11:0] ? image_2908 : _GEN_6043; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6045 = 12'hb5d == _T_71[11:0] ? image_2909 : _GEN_6044; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6046 = 12'hb5e == _T_71[11:0] ? image_2910 : _GEN_6045; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6047 = 12'hb5f == _T_71[11:0] ? image_2911 : _GEN_6046; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6048 = 12'hb60 == _T_71[11:0] ? image_2912 : _GEN_6047; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6049 = 12'hb61 == _T_71[11:0] ? image_2913 : _GEN_6048; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6050 = 12'hb62 == _T_71[11:0] ? image_2914 : _GEN_6049; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6051 = 12'hb63 == _T_71[11:0] ? image_2915 : _GEN_6050; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6052 = 12'hb64 == _T_71[11:0] ? image_2916 : _GEN_6051; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6053 = 12'hb65 == _T_71[11:0] ? image_2917 : _GEN_6052; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6054 = 12'hb66 == _T_71[11:0] ? image_2918 : _GEN_6053; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6055 = 12'hb67 == _T_71[11:0] ? image_2919 : _GEN_6054; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6056 = 12'hb68 == _T_71[11:0] ? image_2920 : _GEN_6055; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6057 = 12'hb69 == _T_71[11:0] ? image_2921 : _GEN_6056; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6058 = 12'hb6a == _T_71[11:0] ? image_2922 : _GEN_6057; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6059 = 12'hb6b == _T_71[11:0] ? image_2923 : _GEN_6058; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6060 = 12'hb6c == _T_71[11:0] ? image_2924 : _GEN_6059; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6061 = 12'hb6d == _T_71[11:0] ? image_2925 : _GEN_6060; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6062 = 12'hb6e == _T_71[11:0] ? image_2926 : _GEN_6061; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6063 = 12'hb6f == _T_71[11:0] ? image_2927 : _GEN_6062; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6064 = 12'hb70 == _T_71[11:0] ? image_2928 : _GEN_6063; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6065 = 12'hb71 == _T_71[11:0] ? image_2929 : _GEN_6064; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6066 = 12'hb72 == _T_71[11:0] ? image_2930 : _GEN_6065; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6067 = 12'hb73 == _T_71[11:0] ? image_2931 : _GEN_6066; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6068 = 12'hb74 == _T_71[11:0] ? image_2932 : _GEN_6067; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6069 = 12'hb75 == _T_71[11:0] ? image_2933 : _GEN_6068; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6070 = 12'hb76 == _T_71[11:0] ? image_2934 : _GEN_6069; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6071 = 12'hb77 == _T_71[11:0] ? 4'h0 : _GEN_6070; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6072 = 12'hb78 == _T_71[11:0] ? 4'h0 : _GEN_6071; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6073 = 12'hb79 == _T_71[11:0] ? 4'h0 : _GEN_6072; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6074 = 12'hb7a == _T_71[11:0] ? 4'h0 : _GEN_6073; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6075 = 12'hb7b == _T_71[11:0] ? 4'h0 : _GEN_6074; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6076 = 12'hb7c == _T_71[11:0] ? 4'h0 : _GEN_6075; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6077 = 12'hb7d == _T_71[11:0] ? 4'h0 : _GEN_6076; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6078 = 12'hb7e == _T_71[11:0] ? 4'h0 : _GEN_6077; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6079 = 12'hb7f == _T_71[11:0] ? 4'h0 : _GEN_6078; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6080 = 12'hb80 == _T_71[11:0] ? 4'h0 : _GEN_6079; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6081 = 12'hb81 == _T_71[11:0] ? 4'h0 : _GEN_6080; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6082 = 12'hb82 == _T_71[11:0] ? 4'h0 : _GEN_6081; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6083 = 12'hb83 == _T_71[11:0] ? 4'h0 : _GEN_6082; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6084 = 12'hb84 == _T_71[11:0] ? 4'h0 : _GEN_6083; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6085 = 12'hb85 == _T_71[11:0] ? 4'h0 : _GEN_6084; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6086 = 12'hb86 == _T_71[11:0] ? 4'h0 : _GEN_6085; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6087 = 12'hb87 == _T_71[11:0] ? 4'h0 : _GEN_6086; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6088 = 12'hb88 == _T_71[11:0] ? 4'h0 : _GEN_6087; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6089 = 12'hb89 == _T_71[11:0] ? 4'h0 : _GEN_6088; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6090 = 12'hb8a == _T_71[11:0] ? 4'h0 : _GEN_6089; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6091 = 12'hb8b == _T_71[11:0] ? 4'h0 : _GEN_6090; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6092 = 12'hb8c == _T_71[11:0] ? 4'h0 : _GEN_6091; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6093 = 12'hb8d == _T_71[11:0] ? 4'h0 : _GEN_6092; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6094 = 12'hb8e == _T_71[11:0] ? 4'h0 : _GEN_6093; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6095 = 12'hb8f == _T_71[11:0] ? 4'h0 : _GEN_6094; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6096 = 12'hb90 == _T_71[11:0] ? 4'h0 : _GEN_6095; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6097 = 12'hb91 == _T_71[11:0] ? 4'h0 : _GEN_6096; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6098 = 12'hb92 == _T_71[11:0] ? 4'h0 : _GEN_6097; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6099 = 12'hb93 == _T_71[11:0] ? 4'h0 : _GEN_6098; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6100 = 12'hb94 == _T_71[11:0] ? 4'h0 : _GEN_6099; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6101 = 12'hb95 == _T_71[11:0] ? image_2965 : _GEN_6100; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6102 = 12'hb96 == _T_71[11:0] ? image_2966 : _GEN_6101; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6103 = 12'hb97 == _T_71[11:0] ? image_2967 : _GEN_6102; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6104 = 12'hb98 == _T_71[11:0] ? image_2968 : _GEN_6103; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6105 = 12'hb99 == _T_71[11:0] ? image_2969 : _GEN_6104; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6106 = 12'hb9a == _T_71[11:0] ? image_2970 : _GEN_6105; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6107 = 12'hb9b == _T_71[11:0] ? image_2971 : _GEN_6106; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6108 = 12'hb9c == _T_71[11:0] ? image_2972 : _GEN_6107; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6109 = 12'hb9d == _T_71[11:0] ? image_2973 : _GEN_6108; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6110 = 12'hb9e == _T_71[11:0] ? image_2974 : _GEN_6109; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6111 = 12'hb9f == _T_71[11:0] ? image_2975 : _GEN_6110; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6112 = 12'hba0 == _T_71[11:0] ? image_2976 : _GEN_6111; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6113 = 12'hba1 == _T_71[11:0] ? image_2977 : _GEN_6112; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6114 = 12'hba2 == _T_71[11:0] ? image_2978 : _GEN_6113; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6115 = 12'hba3 == _T_71[11:0] ? image_2979 : _GEN_6114; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6116 = 12'hba4 == _T_71[11:0] ? image_2980 : _GEN_6115; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6117 = 12'hba5 == _T_71[11:0] ? image_2981 : _GEN_6116; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6118 = 12'hba6 == _T_71[11:0] ? image_2982 : _GEN_6117; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6119 = 12'hba7 == _T_71[11:0] ? image_2983 : _GEN_6118; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6120 = 12'hba8 == _T_71[11:0] ? image_2984 : _GEN_6119; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6121 = 12'hba9 == _T_71[11:0] ? image_2985 : _GEN_6120; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6122 = 12'hbaa == _T_71[11:0] ? image_2986 : _GEN_6121; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6123 = 12'hbab == _T_71[11:0] ? image_2987 : _GEN_6122; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6124 = 12'hbac == _T_71[11:0] ? image_2988 : _GEN_6123; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6125 = 12'hbad == _T_71[11:0] ? image_2989 : _GEN_6124; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6126 = 12'hbae == _T_71[11:0] ? image_2990 : _GEN_6125; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6127 = 12'hbaf == _T_71[11:0] ? image_2991 : _GEN_6126; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6128 = 12'hbb0 == _T_71[11:0] ? image_2992 : _GEN_6127; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6129 = 12'hbb1 == _T_71[11:0] ? image_2993 : _GEN_6128; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6130 = 12'hbb2 == _T_71[11:0] ? image_2994 : _GEN_6129; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6131 = 12'hbb3 == _T_71[11:0] ? image_2995 : _GEN_6130; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6132 = 12'hbb4 == _T_71[11:0] ? image_2996 : _GEN_6131; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6133 = 12'hbb5 == _T_71[11:0] ? 4'h0 : _GEN_6132; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6134 = 12'hbb6 == _T_71[11:0] ? 4'h0 : _GEN_6133; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6135 = 12'hbb7 == _T_71[11:0] ? 4'h0 : _GEN_6134; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6136 = 12'hbb8 == _T_71[11:0] ? 4'h0 : _GEN_6135; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6137 = 12'hbb9 == _T_71[11:0] ? 4'h0 : _GEN_6136; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6138 = 12'hbba == _T_71[11:0] ? 4'h0 : _GEN_6137; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6139 = 12'hbbb == _T_71[11:0] ? 4'h0 : _GEN_6138; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6140 = 12'hbbc == _T_71[11:0] ? 4'h0 : _GEN_6139; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6141 = 12'hbbd == _T_71[11:0] ? 4'h0 : _GEN_6140; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6142 = 12'hbbe == _T_71[11:0] ? 4'h0 : _GEN_6141; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6143 = 12'hbbf == _T_71[11:0] ? 4'h0 : _GEN_6142; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6144 = 12'hbc0 == _T_71[11:0] ? 4'h0 : _GEN_6143; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6145 = 12'hbc1 == _T_71[11:0] ? 4'h0 : _GEN_6144; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6146 = 12'hbc2 == _T_71[11:0] ? 4'h0 : _GEN_6145; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6147 = 12'hbc3 == _T_71[11:0] ? 4'h0 : _GEN_6146; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6148 = 12'hbc4 == _T_71[11:0] ? 4'h0 : _GEN_6147; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6149 = 12'hbc5 == _T_71[11:0] ? 4'h0 : _GEN_6148; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6150 = 12'hbc6 == _T_71[11:0] ? 4'h0 : _GEN_6149; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6151 = 12'hbc7 == _T_71[11:0] ? 4'h0 : _GEN_6150; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6152 = 12'hbc8 == _T_71[11:0] ? 4'h0 : _GEN_6151; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6153 = 12'hbc9 == _T_71[11:0] ? 4'h0 : _GEN_6152; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6154 = 12'hbca == _T_71[11:0] ? 4'h0 : _GEN_6153; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6155 = 12'hbcb == _T_71[11:0] ? 4'h0 : _GEN_6154; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6156 = 12'hbcc == _T_71[11:0] ? 4'h0 : _GEN_6155; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6157 = 12'hbcd == _T_71[11:0] ? 4'h0 : _GEN_6156; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6158 = 12'hbce == _T_71[11:0] ? 4'h0 : _GEN_6157; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6159 = 12'hbcf == _T_71[11:0] ? 4'h0 : _GEN_6158; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6160 = 12'hbd0 == _T_71[11:0] ? 4'h0 : _GEN_6159; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6161 = 12'hbd1 == _T_71[11:0] ? 4'h0 : _GEN_6160; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6162 = 12'hbd2 == _T_71[11:0] ? 4'h0 : _GEN_6161; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6163 = 12'hbd3 == _T_71[11:0] ? 4'h0 : _GEN_6162; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6164 = 12'hbd4 == _T_71[11:0] ? 4'h0 : _GEN_6163; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6165 = 12'hbd5 == _T_71[11:0] ? 4'h0 : _GEN_6164; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6166 = 12'hbd6 == _T_71[11:0] ? 4'h0 : _GEN_6165; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6167 = 12'hbd7 == _T_71[11:0] ? 4'h0 : _GEN_6166; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6168 = 12'hbd8 == _T_71[11:0] ? 4'h0 : _GEN_6167; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6169 = 12'hbd9 == _T_71[11:0] ? 4'h0 : _GEN_6168; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6170 = 12'hbda == _T_71[11:0] ? 4'h0 : _GEN_6169; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6171 = 12'hbdb == _T_71[11:0] ? image_3035 : _GEN_6170; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6172 = 12'hbdc == _T_71[11:0] ? image_3036 : _GEN_6171; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6173 = 12'hbdd == _T_71[11:0] ? image_3037 : _GEN_6172; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6174 = 12'hbde == _T_71[11:0] ? image_3038 : _GEN_6173; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6175 = 12'hbdf == _T_71[11:0] ? image_3039 : _GEN_6174; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6176 = 12'hbe0 == _T_71[11:0] ? image_3040 : _GEN_6175; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6177 = 12'hbe1 == _T_71[11:0] ? image_3041 : _GEN_6176; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6178 = 12'hbe2 == _T_71[11:0] ? image_3042 : _GEN_6177; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6179 = 12'hbe3 == _T_71[11:0] ? image_3043 : _GEN_6178; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6180 = 12'hbe4 == _T_71[11:0] ? image_3044 : _GEN_6179; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6181 = 12'hbe5 == _T_71[11:0] ? image_3045 : _GEN_6180; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6182 = 12'hbe6 == _T_71[11:0] ? image_3046 : _GEN_6181; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6183 = 12'hbe7 == _T_71[11:0] ? image_3047 : _GEN_6182; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6184 = 12'hbe8 == _T_71[11:0] ? image_3048 : _GEN_6183; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6185 = 12'hbe9 == _T_71[11:0] ? image_3049 : _GEN_6184; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6186 = 12'hbea == _T_71[11:0] ? image_3050 : _GEN_6185; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6187 = 12'hbeb == _T_71[11:0] ? image_3051 : _GEN_6186; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6188 = 12'hbec == _T_71[11:0] ? image_3052 : _GEN_6187; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6189 = 12'hbed == _T_71[11:0] ? image_3053 : _GEN_6188; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6190 = 12'hbee == _T_71[11:0] ? image_3054 : _GEN_6189; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6191 = 12'hbef == _T_71[11:0] ? image_3055 : _GEN_6190; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6192 = 12'hbf0 == _T_71[11:0] ? image_3056 : _GEN_6191; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6193 = 12'hbf1 == _T_71[11:0] ? 4'h0 : _GEN_6192; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6194 = 12'hbf2 == _T_71[11:0] ? 4'h0 : _GEN_6193; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6195 = 12'hbf3 == _T_71[11:0] ? 4'h0 : _GEN_6194; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6196 = 12'hbf4 == _T_71[11:0] ? 4'h0 : _GEN_6195; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6197 = 12'hbf5 == _T_71[11:0] ? 4'h0 : _GEN_6196; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6198 = 12'hbf6 == _T_71[11:0] ? 4'h0 : _GEN_6197; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6199 = 12'hbf7 == _T_71[11:0] ? 4'h0 : _GEN_6198; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6200 = 12'hbf8 == _T_71[11:0] ? 4'h0 : _GEN_6199; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6201 = 12'hbf9 == _T_71[11:0] ? 4'h0 : _GEN_6200; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6202 = 12'hbfa == _T_71[11:0] ? 4'h0 : _GEN_6201; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6203 = 12'hbfb == _T_71[11:0] ? 4'h0 : _GEN_6202; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6204 = 12'hbfc == _T_71[11:0] ? 4'h0 : _GEN_6203; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6205 = 12'hbfd == _T_71[11:0] ? 4'h0 : _GEN_6204; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6206 = 12'hbfe == _T_71[11:0] ? 4'h0 : _GEN_6205; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6207 = 12'hbff == _T_71[11:0] ? 4'h0 : _GEN_6206; // @[Filter.scala 138:46]
  wire [31:0] _T_74 = pixelIndex + 32'h2; // @[Filter.scala 133:29]
  wire [31:0] _T_75 = _T_74 / 32'h40; // @[Filter.scala 133:36]
  wire [31:0] _T_77 = _T_75 + _GEN_24805; // @[Filter.scala 133:51]
  wire [31:0] _T_79 = _T_77 - 32'h1; // @[Filter.scala 133:67]
  wire [31:0] _GEN_2 = _T_74 % 32'h40; // @[Filter.scala 134:36]
  wire [6:0] _T_82 = _GEN_2[6:0]; // @[Filter.scala 134:36]
  wire [6:0] _T_84 = _T_82 + _GEN_24806; // @[Filter.scala 134:51]
  wire [6:0] _T_86 = _T_84 - 7'h1; // @[Filter.scala 134:67]
  wire  _T_88 = _T_79 >= 32'h40; // @[Filter.scala 135:27]
  wire  _T_92 = _T_86 >= 7'h30; // @[Filter.scala 135:59]
  wire  _T_93 = _T_88 | _T_92; // @[Filter.scala 135:54]
  wire [13:0] _T_94 = _T_86 * 7'h40; // @[Filter.scala 138:57]
  wire [31:0] _GEN_24813 = {{18'd0}, _T_94}; // @[Filter.scala 138:72]
  wire [31:0] _T_96 = _GEN_24813 + _T_79; // @[Filter.scala 138:72]
  wire [3:0] _GEN_6221 = 12'hc == _T_96[11:0] ? image_12 : 4'h0; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6222 = 12'hd == _T_96[11:0] ? 4'h0 : _GEN_6221; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6223 = 12'he == _T_96[11:0] ? image_14 : _GEN_6222; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6224 = 12'hf == _T_96[11:0] ? image_15 : _GEN_6223; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6225 = 12'h10 == _T_96[11:0] ? image_16 : _GEN_6224; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6226 = 12'h11 == _T_96[11:0] ? image_17 : _GEN_6225; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6227 = 12'h12 == _T_96[11:0] ? image_18 : _GEN_6226; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6228 = 12'h13 == _T_96[11:0] ? image_19 : _GEN_6227; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6229 = 12'h14 == _T_96[11:0] ? image_20 : _GEN_6228; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6230 = 12'h15 == _T_96[11:0] ? image_21 : _GEN_6229; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6231 = 12'h16 == _T_96[11:0] ? image_22 : _GEN_6230; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6232 = 12'h17 == _T_96[11:0] ? image_23 : _GEN_6231; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6233 = 12'h18 == _T_96[11:0] ? 4'h0 : _GEN_6232; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6234 = 12'h19 == _T_96[11:0] ? 4'h0 : _GEN_6233; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6235 = 12'h1a == _T_96[11:0] ? 4'h0 : _GEN_6234; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6236 = 12'h1b == _T_96[11:0] ? 4'h0 : _GEN_6235; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6237 = 12'h1c == _T_96[11:0] ? 4'h0 : _GEN_6236; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6238 = 12'h1d == _T_96[11:0] ? 4'h0 : _GEN_6237; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6239 = 12'h1e == _T_96[11:0] ? 4'h0 : _GEN_6238; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6240 = 12'h1f == _T_96[11:0] ? 4'h0 : _GEN_6239; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6241 = 12'h20 == _T_96[11:0] ? 4'h0 : _GEN_6240; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6242 = 12'h21 == _T_96[11:0] ? 4'h0 : _GEN_6241; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6243 = 12'h22 == _T_96[11:0] ? 4'h0 : _GEN_6242; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6244 = 12'h23 == _T_96[11:0] ? image_35 : _GEN_6243; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6245 = 12'h24 == _T_96[11:0] ? image_36 : _GEN_6244; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6246 = 12'h25 == _T_96[11:0] ? image_37 : _GEN_6245; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6247 = 12'h26 == _T_96[11:0] ? image_38 : _GEN_6246; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6248 = 12'h27 == _T_96[11:0] ? image_39 : _GEN_6247; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6249 = 12'h28 == _T_96[11:0] ? image_40 : _GEN_6248; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6250 = 12'h29 == _T_96[11:0] ? image_41 : _GEN_6249; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6251 = 12'h2a == _T_96[11:0] ? image_42 : _GEN_6250; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6252 = 12'h2b == _T_96[11:0] ? 4'h0 : _GEN_6251; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6253 = 12'h2c == _T_96[11:0] ? 4'h0 : _GEN_6252; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6254 = 12'h2d == _T_96[11:0] ? 4'h0 : _GEN_6253; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6255 = 12'h2e == _T_96[11:0] ? 4'h0 : _GEN_6254; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6256 = 12'h2f == _T_96[11:0] ? 4'h0 : _GEN_6255; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6257 = 12'h30 == _T_96[11:0] ? 4'h0 : _GEN_6256; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6258 = 12'h31 == _T_96[11:0] ? 4'h0 : _GEN_6257; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6259 = 12'h32 == _T_96[11:0] ? 4'h0 : _GEN_6258; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6260 = 12'h33 == _T_96[11:0] ? 4'h0 : _GEN_6259; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6261 = 12'h34 == _T_96[11:0] ? 4'h0 : _GEN_6260; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6262 = 12'h35 == _T_96[11:0] ? 4'h0 : _GEN_6261; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6263 = 12'h36 == _T_96[11:0] ? 4'h0 : _GEN_6262; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6264 = 12'h37 == _T_96[11:0] ? 4'h0 : _GEN_6263; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6265 = 12'h38 == _T_96[11:0] ? 4'h0 : _GEN_6264; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6266 = 12'h39 == _T_96[11:0] ? 4'h0 : _GEN_6265; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6267 = 12'h3a == _T_96[11:0] ? 4'h0 : _GEN_6266; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6268 = 12'h3b == _T_96[11:0] ? 4'h0 : _GEN_6267; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6269 = 12'h3c == _T_96[11:0] ? 4'h0 : _GEN_6268; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6270 = 12'h3d == _T_96[11:0] ? 4'h0 : _GEN_6269; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6271 = 12'h3e == _T_96[11:0] ? 4'h0 : _GEN_6270; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6272 = 12'h3f == _T_96[11:0] ? 4'h0 : _GEN_6271; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6273 = 12'h40 == _T_96[11:0] ? 4'h0 : _GEN_6272; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6274 = 12'h41 == _T_96[11:0] ? 4'h0 : _GEN_6273; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6275 = 12'h42 == _T_96[11:0] ? 4'h0 : _GEN_6274; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6276 = 12'h43 == _T_96[11:0] ? 4'h0 : _GEN_6275; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6277 = 12'h44 == _T_96[11:0] ? 4'h0 : _GEN_6276; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6278 = 12'h45 == _T_96[11:0] ? 4'h0 : _GEN_6277; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6279 = 12'h46 == _T_96[11:0] ? 4'h0 : _GEN_6278; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6280 = 12'h47 == _T_96[11:0] ? 4'h0 : _GEN_6279; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6281 = 12'h48 == _T_96[11:0] ? 4'h0 : _GEN_6280; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6282 = 12'h49 == _T_96[11:0] ? 4'h0 : _GEN_6281; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6283 = 12'h4a == _T_96[11:0] ? 4'h0 : _GEN_6282; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6284 = 12'h4b == _T_96[11:0] ? image_75 : _GEN_6283; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6285 = 12'h4c == _T_96[11:0] ? image_76 : _GEN_6284; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6286 = 12'h4d == _T_96[11:0] ? image_77 : _GEN_6285; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6287 = 12'h4e == _T_96[11:0] ? image_78 : _GEN_6286; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6288 = 12'h4f == _T_96[11:0] ? image_79 : _GEN_6287; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6289 = 12'h50 == _T_96[11:0] ? image_80 : _GEN_6288; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6290 = 12'h51 == _T_96[11:0] ? image_81 : _GEN_6289; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6291 = 12'h52 == _T_96[11:0] ? image_82 : _GEN_6290; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6292 = 12'h53 == _T_96[11:0] ? image_83 : _GEN_6291; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6293 = 12'h54 == _T_96[11:0] ? image_84 : _GEN_6292; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6294 = 12'h55 == _T_96[11:0] ? image_85 : _GEN_6293; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6295 = 12'h56 == _T_96[11:0] ? image_86 : _GEN_6294; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6296 = 12'h57 == _T_96[11:0] ? image_87 : _GEN_6295; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6297 = 12'h58 == _T_96[11:0] ? image_88 : _GEN_6296; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6298 = 12'h59 == _T_96[11:0] ? image_89 : _GEN_6297; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6299 = 12'h5a == _T_96[11:0] ? image_90 : _GEN_6298; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6300 = 12'h5b == _T_96[11:0] ? 4'h0 : _GEN_6299; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6301 = 12'h5c == _T_96[11:0] ? 4'h0 : _GEN_6300; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6302 = 12'h5d == _T_96[11:0] ? image_93 : _GEN_6301; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6303 = 12'h5e == _T_96[11:0] ? 4'h0 : _GEN_6302; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6304 = 12'h5f == _T_96[11:0] ? image_95 : _GEN_6303; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6305 = 12'h60 == _T_96[11:0] ? image_96 : _GEN_6304; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6306 = 12'h61 == _T_96[11:0] ? image_97 : _GEN_6305; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6307 = 12'h62 == _T_96[11:0] ? image_98 : _GEN_6306; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6308 = 12'h63 == _T_96[11:0] ? image_99 : _GEN_6307; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6309 = 12'h64 == _T_96[11:0] ? image_100 : _GEN_6308; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6310 = 12'h65 == _T_96[11:0] ? image_101 : _GEN_6309; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6311 = 12'h66 == _T_96[11:0] ? image_102 : _GEN_6310; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6312 = 12'h67 == _T_96[11:0] ? image_103 : _GEN_6311; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6313 = 12'h68 == _T_96[11:0] ? image_104 : _GEN_6312; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6314 = 12'h69 == _T_96[11:0] ? image_105 : _GEN_6313; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6315 = 12'h6a == _T_96[11:0] ? image_106 : _GEN_6314; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6316 = 12'h6b == _T_96[11:0] ? image_107 : _GEN_6315; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6317 = 12'h6c == _T_96[11:0] ? image_108 : _GEN_6316; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6318 = 12'h6d == _T_96[11:0] ? 4'h0 : _GEN_6317; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6319 = 12'h6e == _T_96[11:0] ? 4'h0 : _GEN_6318; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6320 = 12'h6f == _T_96[11:0] ? 4'h0 : _GEN_6319; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6321 = 12'h70 == _T_96[11:0] ? 4'h0 : _GEN_6320; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6322 = 12'h71 == _T_96[11:0] ? 4'h0 : _GEN_6321; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6323 = 12'h72 == _T_96[11:0] ? 4'h0 : _GEN_6322; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6324 = 12'h73 == _T_96[11:0] ? 4'h0 : _GEN_6323; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6325 = 12'h74 == _T_96[11:0] ? 4'h0 : _GEN_6324; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6326 = 12'h75 == _T_96[11:0] ? 4'h0 : _GEN_6325; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6327 = 12'h76 == _T_96[11:0] ? 4'h0 : _GEN_6326; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6328 = 12'h77 == _T_96[11:0] ? 4'h0 : _GEN_6327; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6329 = 12'h78 == _T_96[11:0] ? 4'h0 : _GEN_6328; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6330 = 12'h79 == _T_96[11:0] ? 4'h0 : _GEN_6329; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6331 = 12'h7a == _T_96[11:0] ? 4'h0 : _GEN_6330; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6332 = 12'h7b == _T_96[11:0] ? 4'h0 : _GEN_6331; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6333 = 12'h7c == _T_96[11:0] ? 4'h0 : _GEN_6332; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6334 = 12'h7d == _T_96[11:0] ? 4'h0 : _GEN_6333; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6335 = 12'h7e == _T_96[11:0] ? 4'h0 : _GEN_6334; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6336 = 12'h7f == _T_96[11:0] ? 4'h0 : _GEN_6335; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6337 = 12'h80 == _T_96[11:0] ? 4'h0 : _GEN_6336; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6338 = 12'h81 == _T_96[11:0] ? 4'h0 : _GEN_6337; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6339 = 12'h82 == _T_96[11:0] ? 4'h0 : _GEN_6338; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6340 = 12'h83 == _T_96[11:0] ? 4'h0 : _GEN_6339; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6341 = 12'h84 == _T_96[11:0] ? 4'h0 : _GEN_6340; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6342 = 12'h85 == _T_96[11:0] ? 4'h0 : _GEN_6341; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6343 = 12'h86 == _T_96[11:0] ? 4'h0 : _GEN_6342; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6344 = 12'h87 == _T_96[11:0] ? 4'h0 : _GEN_6343; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6345 = 12'h88 == _T_96[11:0] ? image_136 : _GEN_6344; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6346 = 12'h89 == _T_96[11:0] ? image_137 : _GEN_6345; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6347 = 12'h8a == _T_96[11:0] ? image_138 : _GEN_6346; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6348 = 12'h8b == _T_96[11:0] ? image_139 : _GEN_6347; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6349 = 12'h8c == _T_96[11:0] ? image_140 : _GEN_6348; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6350 = 12'h8d == _T_96[11:0] ? image_141 : _GEN_6349; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6351 = 12'h8e == _T_96[11:0] ? image_142 : _GEN_6350; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6352 = 12'h8f == _T_96[11:0] ? image_143 : _GEN_6351; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6353 = 12'h90 == _T_96[11:0] ? image_144 : _GEN_6352; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6354 = 12'h91 == _T_96[11:0] ? image_145 : _GEN_6353; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6355 = 12'h92 == _T_96[11:0] ? image_146 : _GEN_6354; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6356 = 12'h93 == _T_96[11:0] ? image_147 : _GEN_6355; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6357 = 12'h94 == _T_96[11:0] ? image_148 : _GEN_6356; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6358 = 12'h95 == _T_96[11:0] ? image_149 : _GEN_6357; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6359 = 12'h96 == _T_96[11:0] ? image_150 : _GEN_6358; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6360 = 12'h97 == _T_96[11:0] ? image_151 : _GEN_6359; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6361 = 12'h98 == _T_96[11:0] ? image_152 : _GEN_6360; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6362 = 12'h99 == _T_96[11:0] ? image_153 : _GEN_6361; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6363 = 12'h9a == _T_96[11:0] ? image_154 : _GEN_6362; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6364 = 12'h9b == _T_96[11:0] ? image_155 : _GEN_6363; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6365 = 12'h9c == _T_96[11:0] ? 4'h0 : _GEN_6364; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6366 = 12'h9d == _T_96[11:0] ? image_157 : _GEN_6365; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6367 = 12'h9e == _T_96[11:0] ? image_158 : _GEN_6366; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6368 = 12'h9f == _T_96[11:0] ? image_159 : _GEN_6367; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6369 = 12'ha0 == _T_96[11:0] ? image_160 : _GEN_6368; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6370 = 12'ha1 == _T_96[11:0] ? image_161 : _GEN_6369; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6371 = 12'ha2 == _T_96[11:0] ? image_162 : _GEN_6370; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6372 = 12'ha3 == _T_96[11:0] ? image_163 : _GEN_6371; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6373 = 12'ha4 == _T_96[11:0] ? image_164 : _GEN_6372; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6374 = 12'ha5 == _T_96[11:0] ? image_165 : _GEN_6373; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6375 = 12'ha6 == _T_96[11:0] ? image_166 : _GEN_6374; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6376 = 12'ha7 == _T_96[11:0] ? image_167 : _GEN_6375; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6377 = 12'ha8 == _T_96[11:0] ? image_168 : _GEN_6376; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6378 = 12'ha9 == _T_96[11:0] ? image_169 : _GEN_6377; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6379 = 12'haa == _T_96[11:0] ? image_170 : _GEN_6378; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6380 = 12'hab == _T_96[11:0] ? image_171 : _GEN_6379; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6381 = 12'hac == _T_96[11:0] ? image_172 : _GEN_6380; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6382 = 12'had == _T_96[11:0] ? image_173 : _GEN_6381; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6383 = 12'hae == _T_96[11:0] ? image_174 : _GEN_6382; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6384 = 12'haf == _T_96[11:0] ? image_175 : _GEN_6383; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6385 = 12'hb0 == _T_96[11:0] ? image_176 : _GEN_6384; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6386 = 12'hb1 == _T_96[11:0] ? image_177 : _GEN_6385; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6387 = 12'hb2 == _T_96[11:0] ? image_178 : _GEN_6386; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6388 = 12'hb3 == _T_96[11:0] ? image_179 : _GEN_6387; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6389 = 12'hb4 == _T_96[11:0] ? 4'h0 : _GEN_6388; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6390 = 12'hb5 == _T_96[11:0] ? 4'h0 : _GEN_6389; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6391 = 12'hb6 == _T_96[11:0] ? 4'h0 : _GEN_6390; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6392 = 12'hb7 == _T_96[11:0] ? 4'h0 : _GEN_6391; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6393 = 12'hb8 == _T_96[11:0] ? 4'h0 : _GEN_6392; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6394 = 12'hb9 == _T_96[11:0] ? 4'h0 : _GEN_6393; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6395 = 12'hba == _T_96[11:0] ? 4'h0 : _GEN_6394; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6396 = 12'hbb == _T_96[11:0] ? 4'h0 : _GEN_6395; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6397 = 12'hbc == _T_96[11:0] ? 4'h0 : _GEN_6396; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6398 = 12'hbd == _T_96[11:0] ? 4'h0 : _GEN_6397; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6399 = 12'hbe == _T_96[11:0] ? 4'h0 : _GEN_6398; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6400 = 12'hbf == _T_96[11:0] ? 4'h0 : _GEN_6399; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6401 = 12'hc0 == _T_96[11:0] ? 4'h0 : _GEN_6400; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6402 = 12'hc1 == _T_96[11:0] ? 4'h0 : _GEN_6401; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6403 = 12'hc2 == _T_96[11:0] ? 4'h0 : _GEN_6402; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6404 = 12'hc3 == _T_96[11:0] ? 4'h0 : _GEN_6403; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6405 = 12'hc4 == _T_96[11:0] ? 4'h0 : _GEN_6404; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6406 = 12'hc5 == _T_96[11:0] ? 4'h0 : _GEN_6405; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6407 = 12'hc6 == _T_96[11:0] ? 4'h0 : _GEN_6406; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6408 = 12'hc7 == _T_96[11:0] ? image_199 : _GEN_6407; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6409 = 12'hc8 == _T_96[11:0] ? image_200 : _GEN_6408; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6410 = 12'hc9 == _T_96[11:0] ? image_201 : _GEN_6409; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6411 = 12'hca == _T_96[11:0] ? image_202 : _GEN_6410; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6412 = 12'hcb == _T_96[11:0] ? image_203 : _GEN_6411; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6413 = 12'hcc == _T_96[11:0] ? image_204 : _GEN_6412; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6414 = 12'hcd == _T_96[11:0] ? image_205 : _GEN_6413; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6415 = 12'hce == _T_96[11:0] ? image_206 : _GEN_6414; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6416 = 12'hcf == _T_96[11:0] ? image_207 : _GEN_6415; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6417 = 12'hd0 == _T_96[11:0] ? image_208 : _GEN_6416; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6418 = 12'hd1 == _T_96[11:0] ? image_209 : _GEN_6417; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6419 = 12'hd2 == _T_96[11:0] ? image_210 : _GEN_6418; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6420 = 12'hd3 == _T_96[11:0] ? image_211 : _GEN_6419; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6421 = 12'hd4 == _T_96[11:0] ? image_212 : _GEN_6420; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6422 = 12'hd5 == _T_96[11:0] ? image_213 : _GEN_6421; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6423 = 12'hd6 == _T_96[11:0] ? image_214 : _GEN_6422; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6424 = 12'hd7 == _T_96[11:0] ? image_215 : _GEN_6423; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6425 = 12'hd8 == _T_96[11:0] ? image_216 : _GEN_6424; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6426 = 12'hd9 == _T_96[11:0] ? image_217 : _GEN_6425; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6427 = 12'hda == _T_96[11:0] ? image_218 : _GEN_6426; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6428 = 12'hdb == _T_96[11:0] ? image_219 : _GEN_6427; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6429 = 12'hdc == _T_96[11:0] ? image_220 : _GEN_6428; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6430 = 12'hdd == _T_96[11:0] ? image_221 : _GEN_6429; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6431 = 12'hde == _T_96[11:0] ? image_222 : _GEN_6430; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6432 = 12'hdf == _T_96[11:0] ? image_223 : _GEN_6431; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6433 = 12'he0 == _T_96[11:0] ? image_224 : _GEN_6432; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6434 = 12'he1 == _T_96[11:0] ? image_225 : _GEN_6433; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6435 = 12'he2 == _T_96[11:0] ? image_226 : _GEN_6434; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6436 = 12'he3 == _T_96[11:0] ? image_227 : _GEN_6435; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6437 = 12'he4 == _T_96[11:0] ? image_228 : _GEN_6436; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6438 = 12'he5 == _T_96[11:0] ? image_229 : _GEN_6437; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6439 = 12'he6 == _T_96[11:0] ? image_230 : _GEN_6438; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6440 = 12'he7 == _T_96[11:0] ? image_231 : _GEN_6439; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6441 = 12'he8 == _T_96[11:0] ? image_232 : _GEN_6440; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6442 = 12'he9 == _T_96[11:0] ? image_233 : _GEN_6441; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6443 = 12'hea == _T_96[11:0] ? image_234 : _GEN_6442; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6444 = 12'heb == _T_96[11:0] ? image_235 : _GEN_6443; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6445 = 12'hec == _T_96[11:0] ? image_236 : _GEN_6444; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6446 = 12'hed == _T_96[11:0] ? image_237 : _GEN_6445; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6447 = 12'hee == _T_96[11:0] ? image_238 : _GEN_6446; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6448 = 12'hef == _T_96[11:0] ? image_239 : _GEN_6447; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6449 = 12'hf0 == _T_96[11:0] ? image_240 : _GEN_6448; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6450 = 12'hf1 == _T_96[11:0] ? image_241 : _GEN_6449; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6451 = 12'hf2 == _T_96[11:0] ? image_242 : _GEN_6450; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6452 = 12'hf3 == _T_96[11:0] ? image_243 : _GEN_6451; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6453 = 12'hf4 == _T_96[11:0] ? image_244 : _GEN_6452; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6454 = 12'hf5 == _T_96[11:0] ? image_245 : _GEN_6453; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6455 = 12'hf6 == _T_96[11:0] ? image_246 : _GEN_6454; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6456 = 12'hf7 == _T_96[11:0] ? 4'h0 : _GEN_6455; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6457 = 12'hf8 == _T_96[11:0] ? 4'h0 : _GEN_6456; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6458 = 12'hf9 == _T_96[11:0] ? 4'h0 : _GEN_6457; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6459 = 12'hfa == _T_96[11:0] ? 4'h0 : _GEN_6458; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6460 = 12'hfb == _T_96[11:0] ? 4'h0 : _GEN_6459; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6461 = 12'hfc == _T_96[11:0] ? 4'h0 : _GEN_6460; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6462 = 12'hfd == _T_96[11:0] ? 4'h0 : _GEN_6461; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6463 = 12'hfe == _T_96[11:0] ? 4'h0 : _GEN_6462; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6464 = 12'hff == _T_96[11:0] ? 4'h0 : _GEN_6463; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6465 = 12'h100 == _T_96[11:0] ? 4'h0 : _GEN_6464; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6466 = 12'h101 == _T_96[11:0] ? 4'h0 : _GEN_6465; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6467 = 12'h102 == _T_96[11:0] ? 4'h0 : _GEN_6466; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6468 = 12'h103 == _T_96[11:0] ? 4'h0 : _GEN_6467; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6469 = 12'h104 == _T_96[11:0] ? 4'h0 : _GEN_6468; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6470 = 12'h105 == _T_96[11:0] ? 4'h0 : _GEN_6469; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6471 = 12'h106 == _T_96[11:0] ? image_262 : _GEN_6470; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6472 = 12'h107 == _T_96[11:0] ? image_263 : _GEN_6471; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6473 = 12'h108 == _T_96[11:0] ? image_264 : _GEN_6472; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6474 = 12'h109 == _T_96[11:0] ? image_265 : _GEN_6473; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6475 = 12'h10a == _T_96[11:0] ? image_266 : _GEN_6474; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6476 = 12'h10b == _T_96[11:0] ? image_267 : _GEN_6475; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6477 = 12'h10c == _T_96[11:0] ? image_268 : _GEN_6476; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6478 = 12'h10d == _T_96[11:0] ? image_269 : _GEN_6477; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6479 = 12'h10e == _T_96[11:0] ? image_270 : _GEN_6478; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6480 = 12'h10f == _T_96[11:0] ? image_271 : _GEN_6479; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6481 = 12'h110 == _T_96[11:0] ? image_272 : _GEN_6480; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6482 = 12'h111 == _T_96[11:0] ? image_273 : _GEN_6481; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6483 = 12'h112 == _T_96[11:0] ? image_274 : _GEN_6482; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6484 = 12'h113 == _T_96[11:0] ? image_275 : _GEN_6483; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6485 = 12'h114 == _T_96[11:0] ? image_276 : _GEN_6484; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6486 = 12'h115 == _T_96[11:0] ? image_277 : _GEN_6485; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6487 = 12'h116 == _T_96[11:0] ? image_278 : _GEN_6486; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6488 = 12'h117 == _T_96[11:0] ? image_279 : _GEN_6487; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6489 = 12'h118 == _T_96[11:0] ? image_280 : _GEN_6488; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6490 = 12'h119 == _T_96[11:0] ? image_281 : _GEN_6489; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6491 = 12'h11a == _T_96[11:0] ? image_282 : _GEN_6490; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6492 = 12'h11b == _T_96[11:0] ? image_283 : _GEN_6491; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6493 = 12'h11c == _T_96[11:0] ? image_284 : _GEN_6492; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6494 = 12'h11d == _T_96[11:0] ? image_285 : _GEN_6493; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6495 = 12'h11e == _T_96[11:0] ? image_286 : _GEN_6494; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6496 = 12'h11f == _T_96[11:0] ? image_287 : _GEN_6495; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6497 = 12'h120 == _T_96[11:0] ? image_288 : _GEN_6496; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6498 = 12'h121 == _T_96[11:0] ? image_289 : _GEN_6497; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6499 = 12'h122 == _T_96[11:0] ? image_290 : _GEN_6498; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6500 = 12'h123 == _T_96[11:0] ? image_291 : _GEN_6499; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6501 = 12'h124 == _T_96[11:0] ? image_292 : _GEN_6500; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6502 = 12'h125 == _T_96[11:0] ? image_293 : _GEN_6501; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6503 = 12'h126 == _T_96[11:0] ? image_294 : _GEN_6502; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6504 = 12'h127 == _T_96[11:0] ? image_295 : _GEN_6503; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6505 = 12'h128 == _T_96[11:0] ? image_296 : _GEN_6504; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6506 = 12'h129 == _T_96[11:0] ? image_297 : _GEN_6505; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6507 = 12'h12a == _T_96[11:0] ? image_298 : _GEN_6506; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6508 = 12'h12b == _T_96[11:0] ? image_299 : _GEN_6507; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6509 = 12'h12c == _T_96[11:0] ? image_300 : _GEN_6508; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6510 = 12'h12d == _T_96[11:0] ? image_301 : _GEN_6509; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6511 = 12'h12e == _T_96[11:0] ? image_302 : _GEN_6510; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6512 = 12'h12f == _T_96[11:0] ? image_303 : _GEN_6511; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6513 = 12'h130 == _T_96[11:0] ? image_304 : _GEN_6512; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6514 = 12'h131 == _T_96[11:0] ? image_305 : _GEN_6513; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6515 = 12'h132 == _T_96[11:0] ? image_306 : _GEN_6514; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6516 = 12'h133 == _T_96[11:0] ? image_307 : _GEN_6515; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6517 = 12'h134 == _T_96[11:0] ? image_308 : _GEN_6516; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6518 = 12'h135 == _T_96[11:0] ? image_309 : _GEN_6517; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6519 = 12'h136 == _T_96[11:0] ? image_310 : _GEN_6518; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6520 = 12'h137 == _T_96[11:0] ? image_311 : _GEN_6519; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6521 = 12'h138 == _T_96[11:0] ? image_312 : _GEN_6520; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6522 = 12'h139 == _T_96[11:0] ? image_313 : _GEN_6521; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6523 = 12'h13a == _T_96[11:0] ? image_314 : _GEN_6522; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6524 = 12'h13b == _T_96[11:0] ? image_315 : _GEN_6523; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6525 = 12'h13c == _T_96[11:0] ? 4'h0 : _GEN_6524; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6526 = 12'h13d == _T_96[11:0] ? 4'h0 : _GEN_6525; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6527 = 12'h13e == _T_96[11:0] ? 4'h0 : _GEN_6526; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6528 = 12'h13f == _T_96[11:0] ? 4'h0 : _GEN_6527; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6529 = 12'h140 == _T_96[11:0] ? 4'h0 : _GEN_6528; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6530 = 12'h141 == _T_96[11:0] ? 4'h0 : _GEN_6529; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6531 = 12'h142 == _T_96[11:0] ? 4'h0 : _GEN_6530; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6532 = 12'h143 == _T_96[11:0] ? 4'h0 : _GEN_6531; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6533 = 12'h144 == _T_96[11:0] ? 4'h0 : _GEN_6532; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6534 = 12'h145 == _T_96[11:0] ? image_325 : _GEN_6533; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6535 = 12'h146 == _T_96[11:0] ? image_326 : _GEN_6534; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6536 = 12'h147 == _T_96[11:0] ? image_327 : _GEN_6535; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6537 = 12'h148 == _T_96[11:0] ? image_328 : _GEN_6536; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6538 = 12'h149 == _T_96[11:0] ? image_329 : _GEN_6537; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6539 = 12'h14a == _T_96[11:0] ? image_330 : _GEN_6538; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6540 = 12'h14b == _T_96[11:0] ? image_331 : _GEN_6539; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6541 = 12'h14c == _T_96[11:0] ? image_332 : _GEN_6540; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6542 = 12'h14d == _T_96[11:0] ? image_333 : _GEN_6541; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6543 = 12'h14e == _T_96[11:0] ? image_334 : _GEN_6542; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6544 = 12'h14f == _T_96[11:0] ? image_335 : _GEN_6543; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6545 = 12'h150 == _T_96[11:0] ? image_336 : _GEN_6544; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6546 = 12'h151 == _T_96[11:0] ? image_337 : _GEN_6545; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6547 = 12'h152 == _T_96[11:0] ? image_338 : _GEN_6546; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6548 = 12'h153 == _T_96[11:0] ? image_339 : _GEN_6547; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6549 = 12'h154 == _T_96[11:0] ? image_340 : _GEN_6548; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6550 = 12'h155 == _T_96[11:0] ? image_341 : _GEN_6549; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6551 = 12'h156 == _T_96[11:0] ? image_342 : _GEN_6550; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6552 = 12'h157 == _T_96[11:0] ? image_343 : _GEN_6551; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6553 = 12'h158 == _T_96[11:0] ? image_344 : _GEN_6552; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6554 = 12'h159 == _T_96[11:0] ? image_345 : _GEN_6553; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6555 = 12'h15a == _T_96[11:0] ? image_346 : _GEN_6554; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6556 = 12'h15b == _T_96[11:0] ? image_347 : _GEN_6555; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6557 = 12'h15c == _T_96[11:0] ? image_348 : _GEN_6556; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6558 = 12'h15d == _T_96[11:0] ? image_349 : _GEN_6557; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6559 = 12'h15e == _T_96[11:0] ? image_350 : _GEN_6558; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6560 = 12'h15f == _T_96[11:0] ? image_351 : _GEN_6559; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6561 = 12'h160 == _T_96[11:0] ? image_352 : _GEN_6560; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6562 = 12'h161 == _T_96[11:0] ? image_353 : _GEN_6561; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6563 = 12'h162 == _T_96[11:0] ? image_354 : _GEN_6562; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6564 = 12'h163 == _T_96[11:0] ? image_355 : _GEN_6563; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6565 = 12'h164 == _T_96[11:0] ? image_356 : _GEN_6564; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6566 = 12'h165 == _T_96[11:0] ? image_357 : _GEN_6565; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6567 = 12'h166 == _T_96[11:0] ? image_358 : _GEN_6566; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6568 = 12'h167 == _T_96[11:0] ? image_359 : _GEN_6567; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6569 = 12'h168 == _T_96[11:0] ? image_360 : _GEN_6568; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6570 = 12'h169 == _T_96[11:0] ? image_361 : _GEN_6569; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6571 = 12'h16a == _T_96[11:0] ? image_362 : _GEN_6570; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6572 = 12'h16b == _T_96[11:0] ? image_363 : _GEN_6571; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6573 = 12'h16c == _T_96[11:0] ? image_364 : _GEN_6572; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6574 = 12'h16d == _T_96[11:0] ? image_365 : _GEN_6573; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6575 = 12'h16e == _T_96[11:0] ? image_366 : _GEN_6574; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6576 = 12'h16f == _T_96[11:0] ? image_367 : _GEN_6575; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6577 = 12'h170 == _T_96[11:0] ? image_368 : _GEN_6576; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6578 = 12'h171 == _T_96[11:0] ? image_369 : _GEN_6577; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6579 = 12'h172 == _T_96[11:0] ? image_370 : _GEN_6578; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6580 = 12'h173 == _T_96[11:0] ? image_371 : _GEN_6579; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6581 = 12'h174 == _T_96[11:0] ? image_372 : _GEN_6580; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6582 = 12'h175 == _T_96[11:0] ? image_373 : _GEN_6581; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6583 = 12'h176 == _T_96[11:0] ? image_374 : _GEN_6582; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6584 = 12'h177 == _T_96[11:0] ? image_375 : _GEN_6583; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6585 = 12'h178 == _T_96[11:0] ? image_376 : _GEN_6584; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6586 = 12'h179 == _T_96[11:0] ? image_377 : _GEN_6585; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6587 = 12'h17a == _T_96[11:0] ? image_378 : _GEN_6586; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6588 = 12'h17b == _T_96[11:0] ? image_379 : _GEN_6587; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6589 = 12'h17c == _T_96[11:0] ? 4'h0 : _GEN_6588; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6590 = 12'h17d == _T_96[11:0] ? 4'h0 : _GEN_6589; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6591 = 12'h17e == _T_96[11:0] ? 4'h0 : _GEN_6590; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6592 = 12'h17f == _T_96[11:0] ? 4'h0 : _GEN_6591; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6593 = 12'h180 == _T_96[11:0] ? 4'h0 : _GEN_6592; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6594 = 12'h181 == _T_96[11:0] ? 4'h0 : _GEN_6593; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6595 = 12'h182 == _T_96[11:0] ? 4'h0 : _GEN_6594; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6596 = 12'h183 == _T_96[11:0] ? 4'h0 : _GEN_6595; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6597 = 12'h184 == _T_96[11:0] ? image_388 : _GEN_6596; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6598 = 12'h185 == _T_96[11:0] ? image_389 : _GEN_6597; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6599 = 12'h186 == _T_96[11:0] ? image_390 : _GEN_6598; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6600 = 12'h187 == _T_96[11:0] ? image_391 : _GEN_6599; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6601 = 12'h188 == _T_96[11:0] ? image_392 : _GEN_6600; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6602 = 12'h189 == _T_96[11:0] ? image_393 : _GEN_6601; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6603 = 12'h18a == _T_96[11:0] ? image_394 : _GEN_6602; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6604 = 12'h18b == _T_96[11:0] ? image_395 : _GEN_6603; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6605 = 12'h18c == _T_96[11:0] ? image_396 : _GEN_6604; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6606 = 12'h18d == _T_96[11:0] ? image_397 : _GEN_6605; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6607 = 12'h18e == _T_96[11:0] ? image_398 : _GEN_6606; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6608 = 12'h18f == _T_96[11:0] ? image_399 : _GEN_6607; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6609 = 12'h190 == _T_96[11:0] ? image_400 : _GEN_6608; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6610 = 12'h191 == _T_96[11:0] ? image_401 : _GEN_6609; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6611 = 12'h192 == _T_96[11:0] ? image_402 : _GEN_6610; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6612 = 12'h193 == _T_96[11:0] ? image_403 : _GEN_6611; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6613 = 12'h194 == _T_96[11:0] ? image_404 : _GEN_6612; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6614 = 12'h195 == _T_96[11:0] ? image_405 : _GEN_6613; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6615 = 12'h196 == _T_96[11:0] ? image_406 : _GEN_6614; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6616 = 12'h197 == _T_96[11:0] ? image_407 : _GEN_6615; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6617 = 12'h198 == _T_96[11:0] ? image_408 : _GEN_6616; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6618 = 12'h199 == _T_96[11:0] ? image_409 : _GEN_6617; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6619 = 12'h19a == _T_96[11:0] ? image_410 : _GEN_6618; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6620 = 12'h19b == _T_96[11:0] ? image_411 : _GEN_6619; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6621 = 12'h19c == _T_96[11:0] ? image_412 : _GEN_6620; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6622 = 12'h19d == _T_96[11:0] ? image_413 : _GEN_6621; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6623 = 12'h19e == _T_96[11:0] ? image_414 : _GEN_6622; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6624 = 12'h19f == _T_96[11:0] ? image_415 : _GEN_6623; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6625 = 12'h1a0 == _T_96[11:0] ? image_416 : _GEN_6624; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6626 = 12'h1a1 == _T_96[11:0] ? image_417 : _GEN_6625; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6627 = 12'h1a2 == _T_96[11:0] ? image_418 : _GEN_6626; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6628 = 12'h1a3 == _T_96[11:0] ? image_419 : _GEN_6627; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6629 = 12'h1a4 == _T_96[11:0] ? image_420 : _GEN_6628; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6630 = 12'h1a5 == _T_96[11:0] ? image_421 : _GEN_6629; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6631 = 12'h1a6 == _T_96[11:0] ? image_422 : _GEN_6630; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6632 = 12'h1a7 == _T_96[11:0] ? image_423 : _GEN_6631; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6633 = 12'h1a8 == _T_96[11:0] ? image_424 : _GEN_6632; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6634 = 12'h1a9 == _T_96[11:0] ? image_425 : _GEN_6633; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6635 = 12'h1aa == _T_96[11:0] ? image_426 : _GEN_6634; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6636 = 12'h1ab == _T_96[11:0] ? image_427 : _GEN_6635; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6637 = 12'h1ac == _T_96[11:0] ? image_428 : _GEN_6636; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6638 = 12'h1ad == _T_96[11:0] ? image_429 : _GEN_6637; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6639 = 12'h1ae == _T_96[11:0] ? image_430 : _GEN_6638; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6640 = 12'h1af == _T_96[11:0] ? image_431 : _GEN_6639; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6641 = 12'h1b0 == _T_96[11:0] ? image_432 : _GEN_6640; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6642 = 12'h1b1 == _T_96[11:0] ? image_433 : _GEN_6641; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6643 = 12'h1b2 == _T_96[11:0] ? image_434 : _GEN_6642; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6644 = 12'h1b3 == _T_96[11:0] ? image_435 : _GEN_6643; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6645 = 12'h1b4 == _T_96[11:0] ? image_436 : _GEN_6644; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6646 = 12'h1b5 == _T_96[11:0] ? image_437 : _GEN_6645; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6647 = 12'h1b6 == _T_96[11:0] ? image_438 : _GEN_6646; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6648 = 12'h1b7 == _T_96[11:0] ? image_439 : _GEN_6647; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6649 = 12'h1b8 == _T_96[11:0] ? image_440 : _GEN_6648; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6650 = 12'h1b9 == _T_96[11:0] ? image_441 : _GEN_6649; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6651 = 12'h1ba == _T_96[11:0] ? image_442 : _GEN_6650; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6652 = 12'h1bb == _T_96[11:0] ? image_443 : _GEN_6651; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6653 = 12'h1bc == _T_96[11:0] ? image_444 : _GEN_6652; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6654 = 12'h1bd == _T_96[11:0] ? 4'h0 : _GEN_6653; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6655 = 12'h1be == _T_96[11:0] ? 4'h0 : _GEN_6654; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6656 = 12'h1bf == _T_96[11:0] ? 4'h0 : _GEN_6655; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6657 = 12'h1c0 == _T_96[11:0] ? 4'h0 : _GEN_6656; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6658 = 12'h1c1 == _T_96[11:0] ? 4'h0 : _GEN_6657; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6659 = 12'h1c2 == _T_96[11:0] ? 4'h0 : _GEN_6658; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6660 = 12'h1c3 == _T_96[11:0] ? image_451 : _GEN_6659; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6661 = 12'h1c4 == _T_96[11:0] ? image_452 : _GEN_6660; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6662 = 12'h1c5 == _T_96[11:0] ? image_453 : _GEN_6661; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6663 = 12'h1c6 == _T_96[11:0] ? image_454 : _GEN_6662; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6664 = 12'h1c7 == _T_96[11:0] ? image_455 : _GEN_6663; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6665 = 12'h1c8 == _T_96[11:0] ? image_456 : _GEN_6664; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6666 = 12'h1c9 == _T_96[11:0] ? image_457 : _GEN_6665; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6667 = 12'h1ca == _T_96[11:0] ? image_458 : _GEN_6666; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6668 = 12'h1cb == _T_96[11:0] ? image_459 : _GEN_6667; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6669 = 12'h1cc == _T_96[11:0] ? image_460 : _GEN_6668; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6670 = 12'h1cd == _T_96[11:0] ? image_461 : _GEN_6669; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6671 = 12'h1ce == _T_96[11:0] ? image_462 : _GEN_6670; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6672 = 12'h1cf == _T_96[11:0] ? image_463 : _GEN_6671; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6673 = 12'h1d0 == _T_96[11:0] ? image_464 : _GEN_6672; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6674 = 12'h1d1 == _T_96[11:0] ? image_465 : _GEN_6673; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6675 = 12'h1d2 == _T_96[11:0] ? image_466 : _GEN_6674; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6676 = 12'h1d3 == _T_96[11:0] ? image_467 : _GEN_6675; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6677 = 12'h1d4 == _T_96[11:0] ? image_468 : _GEN_6676; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6678 = 12'h1d5 == _T_96[11:0] ? image_469 : _GEN_6677; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6679 = 12'h1d6 == _T_96[11:0] ? image_470 : _GEN_6678; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6680 = 12'h1d7 == _T_96[11:0] ? image_471 : _GEN_6679; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6681 = 12'h1d8 == _T_96[11:0] ? image_472 : _GEN_6680; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6682 = 12'h1d9 == _T_96[11:0] ? image_473 : _GEN_6681; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6683 = 12'h1da == _T_96[11:0] ? image_474 : _GEN_6682; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6684 = 12'h1db == _T_96[11:0] ? image_475 : _GEN_6683; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6685 = 12'h1dc == _T_96[11:0] ? image_476 : _GEN_6684; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6686 = 12'h1dd == _T_96[11:0] ? image_477 : _GEN_6685; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6687 = 12'h1de == _T_96[11:0] ? image_478 : _GEN_6686; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6688 = 12'h1df == _T_96[11:0] ? image_479 : _GEN_6687; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6689 = 12'h1e0 == _T_96[11:0] ? image_480 : _GEN_6688; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6690 = 12'h1e1 == _T_96[11:0] ? image_481 : _GEN_6689; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6691 = 12'h1e2 == _T_96[11:0] ? image_482 : _GEN_6690; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6692 = 12'h1e3 == _T_96[11:0] ? image_483 : _GEN_6691; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6693 = 12'h1e4 == _T_96[11:0] ? image_484 : _GEN_6692; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6694 = 12'h1e5 == _T_96[11:0] ? image_485 : _GEN_6693; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6695 = 12'h1e6 == _T_96[11:0] ? image_486 : _GEN_6694; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6696 = 12'h1e7 == _T_96[11:0] ? image_487 : _GEN_6695; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6697 = 12'h1e8 == _T_96[11:0] ? image_488 : _GEN_6696; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6698 = 12'h1e9 == _T_96[11:0] ? image_489 : _GEN_6697; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6699 = 12'h1ea == _T_96[11:0] ? image_490 : _GEN_6698; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6700 = 12'h1eb == _T_96[11:0] ? image_491 : _GEN_6699; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6701 = 12'h1ec == _T_96[11:0] ? image_492 : _GEN_6700; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6702 = 12'h1ed == _T_96[11:0] ? image_493 : _GEN_6701; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6703 = 12'h1ee == _T_96[11:0] ? image_494 : _GEN_6702; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6704 = 12'h1ef == _T_96[11:0] ? image_495 : _GEN_6703; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6705 = 12'h1f0 == _T_96[11:0] ? image_496 : _GEN_6704; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6706 = 12'h1f1 == _T_96[11:0] ? image_497 : _GEN_6705; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6707 = 12'h1f2 == _T_96[11:0] ? image_498 : _GEN_6706; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6708 = 12'h1f3 == _T_96[11:0] ? image_499 : _GEN_6707; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6709 = 12'h1f4 == _T_96[11:0] ? image_500 : _GEN_6708; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6710 = 12'h1f5 == _T_96[11:0] ? image_501 : _GEN_6709; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6711 = 12'h1f6 == _T_96[11:0] ? image_502 : _GEN_6710; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6712 = 12'h1f7 == _T_96[11:0] ? image_503 : _GEN_6711; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6713 = 12'h1f8 == _T_96[11:0] ? image_504 : _GEN_6712; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6714 = 12'h1f9 == _T_96[11:0] ? image_505 : _GEN_6713; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6715 = 12'h1fa == _T_96[11:0] ? image_506 : _GEN_6714; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6716 = 12'h1fb == _T_96[11:0] ? image_507 : _GEN_6715; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6717 = 12'h1fc == _T_96[11:0] ? image_508 : _GEN_6716; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6718 = 12'h1fd == _T_96[11:0] ? image_509 : _GEN_6717; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6719 = 12'h1fe == _T_96[11:0] ? 4'h0 : _GEN_6718; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6720 = 12'h1ff == _T_96[11:0] ? 4'h0 : _GEN_6719; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6721 = 12'h200 == _T_96[11:0] ? 4'h0 : _GEN_6720; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6722 = 12'h201 == _T_96[11:0] ? 4'h0 : _GEN_6721; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6723 = 12'h202 == _T_96[11:0] ? 4'h0 : _GEN_6722; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6724 = 12'h203 == _T_96[11:0] ? image_515 : _GEN_6723; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6725 = 12'h204 == _T_96[11:0] ? image_516 : _GEN_6724; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6726 = 12'h205 == _T_96[11:0] ? image_517 : _GEN_6725; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6727 = 12'h206 == _T_96[11:0] ? image_518 : _GEN_6726; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6728 = 12'h207 == _T_96[11:0] ? image_519 : _GEN_6727; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6729 = 12'h208 == _T_96[11:0] ? image_520 : _GEN_6728; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6730 = 12'h209 == _T_96[11:0] ? image_521 : _GEN_6729; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6731 = 12'h20a == _T_96[11:0] ? image_522 : _GEN_6730; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6732 = 12'h20b == _T_96[11:0] ? image_523 : _GEN_6731; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6733 = 12'h20c == _T_96[11:0] ? image_524 : _GEN_6732; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6734 = 12'h20d == _T_96[11:0] ? image_525 : _GEN_6733; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6735 = 12'h20e == _T_96[11:0] ? image_526 : _GEN_6734; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6736 = 12'h20f == _T_96[11:0] ? image_527 : _GEN_6735; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6737 = 12'h210 == _T_96[11:0] ? image_528 : _GEN_6736; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6738 = 12'h211 == _T_96[11:0] ? image_529 : _GEN_6737; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6739 = 12'h212 == _T_96[11:0] ? image_530 : _GEN_6738; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6740 = 12'h213 == _T_96[11:0] ? image_531 : _GEN_6739; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6741 = 12'h214 == _T_96[11:0] ? image_532 : _GEN_6740; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6742 = 12'h215 == _T_96[11:0] ? image_533 : _GEN_6741; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6743 = 12'h216 == _T_96[11:0] ? image_534 : _GEN_6742; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6744 = 12'h217 == _T_96[11:0] ? image_535 : _GEN_6743; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6745 = 12'h218 == _T_96[11:0] ? image_536 : _GEN_6744; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6746 = 12'h219 == _T_96[11:0] ? image_537 : _GEN_6745; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6747 = 12'h21a == _T_96[11:0] ? image_538 : _GEN_6746; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6748 = 12'h21b == _T_96[11:0] ? image_539 : _GEN_6747; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6749 = 12'h21c == _T_96[11:0] ? image_540 : _GEN_6748; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6750 = 12'h21d == _T_96[11:0] ? image_541 : _GEN_6749; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6751 = 12'h21e == _T_96[11:0] ? image_542 : _GEN_6750; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6752 = 12'h21f == _T_96[11:0] ? image_543 : _GEN_6751; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6753 = 12'h220 == _T_96[11:0] ? image_544 : _GEN_6752; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6754 = 12'h221 == _T_96[11:0] ? image_545 : _GEN_6753; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6755 = 12'h222 == _T_96[11:0] ? image_546 : _GEN_6754; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6756 = 12'h223 == _T_96[11:0] ? image_547 : _GEN_6755; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6757 = 12'h224 == _T_96[11:0] ? image_548 : _GEN_6756; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6758 = 12'h225 == _T_96[11:0] ? image_549 : _GEN_6757; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6759 = 12'h226 == _T_96[11:0] ? image_550 : _GEN_6758; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6760 = 12'h227 == _T_96[11:0] ? image_551 : _GEN_6759; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6761 = 12'h228 == _T_96[11:0] ? image_552 : _GEN_6760; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6762 = 12'h229 == _T_96[11:0] ? image_553 : _GEN_6761; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6763 = 12'h22a == _T_96[11:0] ? image_554 : _GEN_6762; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6764 = 12'h22b == _T_96[11:0] ? image_555 : _GEN_6763; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6765 = 12'h22c == _T_96[11:0] ? image_556 : _GEN_6764; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6766 = 12'h22d == _T_96[11:0] ? image_557 : _GEN_6765; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6767 = 12'h22e == _T_96[11:0] ? image_558 : _GEN_6766; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6768 = 12'h22f == _T_96[11:0] ? image_559 : _GEN_6767; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6769 = 12'h230 == _T_96[11:0] ? image_560 : _GEN_6768; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6770 = 12'h231 == _T_96[11:0] ? image_561 : _GEN_6769; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6771 = 12'h232 == _T_96[11:0] ? image_562 : _GEN_6770; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6772 = 12'h233 == _T_96[11:0] ? image_563 : _GEN_6771; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6773 = 12'h234 == _T_96[11:0] ? image_564 : _GEN_6772; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6774 = 12'h235 == _T_96[11:0] ? image_565 : _GEN_6773; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6775 = 12'h236 == _T_96[11:0] ? image_566 : _GEN_6774; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6776 = 12'h237 == _T_96[11:0] ? 4'h0 : _GEN_6775; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6777 = 12'h238 == _T_96[11:0] ? 4'h0 : _GEN_6776; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6778 = 12'h239 == _T_96[11:0] ? 4'h0 : _GEN_6777; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6779 = 12'h23a == _T_96[11:0] ? 4'h0 : _GEN_6778; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6780 = 12'h23b == _T_96[11:0] ? image_571 : _GEN_6779; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6781 = 12'h23c == _T_96[11:0] ? image_572 : _GEN_6780; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6782 = 12'h23d == _T_96[11:0] ? image_573 : _GEN_6781; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6783 = 12'h23e == _T_96[11:0] ? image_574 : _GEN_6782; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6784 = 12'h23f == _T_96[11:0] ? 4'h0 : _GEN_6783; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6785 = 12'h240 == _T_96[11:0] ? 4'h0 : _GEN_6784; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6786 = 12'h241 == _T_96[11:0] ? 4'h0 : _GEN_6785; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6787 = 12'h242 == _T_96[11:0] ? image_578 : _GEN_6786; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6788 = 12'h243 == _T_96[11:0] ? image_579 : _GEN_6787; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6789 = 12'h244 == _T_96[11:0] ? image_580 : _GEN_6788; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6790 = 12'h245 == _T_96[11:0] ? image_581 : _GEN_6789; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6791 = 12'h246 == _T_96[11:0] ? image_582 : _GEN_6790; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6792 = 12'h247 == _T_96[11:0] ? image_583 : _GEN_6791; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6793 = 12'h248 == _T_96[11:0] ? image_584 : _GEN_6792; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6794 = 12'h249 == _T_96[11:0] ? image_585 : _GEN_6793; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6795 = 12'h24a == _T_96[11:0] ? image_586 : _GEN_6794; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6796 = 12'h24b == _T_96[11:0] ? image_587 : _GEN_6795; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6797 = 12'h24c == _T_96[11:0] ? image_588 : _GEN_6796; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6798 = 12'h24d == _T_96[11:0] ? image_589 : _GEN_6797; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6799 = 12'h24e == _T_96[11:0] ? image_590 : _GEN_6798; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6800 = 12'h24f == _T_96[11:0] ? image_591 : _GEN_6799; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6801 = 12'h250 == _T_96[11:0] ? image_592 : _GEN_6800; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6802 = 12'h251 == _T_96[11:0] ? image_593 : _GEN_6801; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6803 = 12'h252 == _T_96[11:0] ? image_594 : _GEN_6802; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6804 = 12'h253 == _T_96[11:0] ? image_595 : _GEN_6803; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6805 = 12'h254 == _T_96[11:0] ? image_596 : _GEN_6804; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6806 = 12'h255 == _T_96[11:0] ? image_597 : _GEN_6805; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6807 = 12'h256 == _T_96[11:0] ? image_598 : _GEN_6806; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6808 = 12'h257 == _T_96[11:0] ? image_599 : _GEN_6807; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6809 = 12'h258 == _T_96[11:0] ? image_600 : _GEN_6808; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6810 = 12'h259 == _T_96[11:0] ? image_601 : _GEN_6809; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6811 = 12'h25a == _T_96[11:0] ? image_602 : _GEN_6810; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6812 = 12'h25b == _T_96[11:0] ? image_603 : _GEN_6811; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6813 = 12'h25c == _T_96[11:0] ? image_604 : _GEN_6812; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6814 = 12'h25d == _T_96[11:0] ? image_605 : _GEN_6813; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6815 = 12'h25e == _T_96[11:0] ? image_606 : _GEN_6814; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6816 = 12'h25f == _T_96[11:0] ? image_607 : _GEN_6815; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6817 = 12'h260 == _T_96[11:0] ? 4'h0 : _GEN_6816; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6818 = 12'h261 == _T_96[11:0] ? 4'h0 : _GEN_6817; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6819 = 12'h262 == _T_96[11:0] ? 4'h0 : _GEN_6818; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6820 = 12'h263 == _T_96[11:0] ? 4'h0 : _GEN_6819; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6821 = 12'h264 == _T_96[11:0] ? 4'h0 : _GEN_6820; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6822 = 12'h265 == _T_96[11:0] ? 4'h0 : _GEN_6821; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6823 = 12'h266 == _T_96[11:0] ? image_614 : _GEN_6822; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6824 = 12'h267 == _T_96[11:0] ? image_615 : _GEN_6823; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6825 = 12'h268 == _T_96[11:0] ? image_616 : _GEN_6824; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6826 = 12'h269 == _T_96[11:0] ? image_617 : _GEN_6825; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6827 = 12'h26a == _T_96[11:0] ? image_618 : _GEN_6826; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6828 = 12'h26b == _T_96[11:0] ? image_619 : _GEN_6827; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6829 = 12'h26c == _T_96[11:0] ? image_620 : _GEN_6828; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6830 = 12'h26d == _T_96[11:0] ? image_621 : _GEN_6829; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6831 = 12'h26e == _T_96[11:0] ? image_622 : _GEN_6830; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6832 = 12'h26f == _T_96[11:0] ? image_623 : _GEN_6831; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6833 = 12'h270 == _T_96[11:0] ? image_624 : _GEN_6832; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6834 = 12'h271 == _T_96[11:0] ? image_625 : _GEN_6833; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6835 = 12'h272 == _T_96[11:0] ? image_626 : _GEN_6834; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6836 = 12'h273 == _T_96[11:0] ? image_627 : _GEN_6835; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6837 = 12'h274 == _T_96[11:0] ? image_628 : _GEN_6836; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6838 = 12'h275 == _T_96[11:0] ? 4'h0 : _GEN_6837; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6839 = 12'h276 == _T_96[11:0] ? 4'h0 : _GEN_6838; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6840 = 12'h277 == _T_96[11:0] ? 4'h0 : _GEN_6839; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6841 = 12'h278 == _T_96[11:0] ? 4'h0 : _GEN_6840; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6842 = 12'h279 == _T_96[11:0] ? 4'h0 : _GEN_6841; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6843 = 12'h27a == _T_96[11:0] ? 4'h0 : _GEN_6842; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6844 = 12'h27b == _T_96[11:0] ? 4'h0 : _GEN_6843; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6845 = 12'h27c == _T_96[11:0] ? image_636 : _GEN_6844; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6846 = 12'h27d == _T_96[11:0] ? image_637 : _GEN_6845; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6847 = 12'h27e == _T_96[11:0] ? image_638 : _GEN_6846; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6848 = 12'h27f == _T_96[11:0] ? image_639 : _GEN_6847; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6849 = 12'h280 == _T_96[11:0] ? 4'h0 : _GEN_6848; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6850 = 12'h281 == _T_96[11:0] ? 4'h0 : _GEN_6849; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6851 = 12'h282 == _T_96[11:0] ? image_642 : _GEN_6850; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6852 = 12'h283 == _T_96[11:0] ? image_643 : _GEN_6851; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6853 = 12'h284 == _T_96[11:0] ? image_644 : _GEN_6852; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6854 = 12'h285 == _T_96[11:0] ? image_645 : _GEN_6853; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6855 = 12'h286 == _T_96[11:0] ? image_646 : _GEN_6854; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6856 = 12'h287 == _T_96[11:0] ? image_647 : _GEN_6855; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6857 = 12'h288 == _T_96[11:0] ? image_648 : _GEN_6856; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6858 = 12'h289 == _T_96[11:0] ? image_649 : _GEN_6857; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6859 = 12'h28a == _T_96[11:0] ? image_650 : _GEN_6858; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6860 = 12'h28b == _T_96[11:0] ? image_651 : _GEN_6859; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6861 = 12'h28c == _T_96[11:0] ? image_652 : _GEN_6860; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6862 = 12'h28d == _T_96[11:0] ? image_653 : _GEN_6861; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6863 = 12'h28e == _T_96[11:0] ? image_654 : _GEN_6862; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6864 = 12'h28f == _T_96[11:0] ? image_655 : _GEN_6863; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6865 = 12'h290 == _T_96[11:0] ? image_656 : _GEN_6864; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6866 = 12'h291 == _T_96[11:0] ? image_657 : _GEN_6865; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6867 = 12'h292 == _T_96[11:0] ? image_658 : _GEN_6866; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6868 = 12'h293 == _T_96[11:0] ? image_659 : _GEN_6867; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6869 = 12'h294 == _T_96[11:0] ? image_660 : _GEN_6868; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6870 = 12'h295 == _T_96[11:0] ? image_661 : _GEN_6869; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6871 = 12'h296 == _T_96[11:0] ? image_662 : _GEN_6870; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6872 = 12'h297 == _T_96[11:0] ? image_663 : _GEN_6871; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6873 = 12'h298 == _T_96[11:0] ? image_664 : _GEN_6872; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6874 = 12'h299 == _T_96[11:0] ? image_665 : _GEN_6873; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6875 = 12'h29a == _T_96[11:0] ? image_666 : _GEN_6874; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6876 = 12'h29b == _T_96[11:0] ? image_667 : _GEN_6875; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6877 = 12'h29c == _T_96[11:0] ? image_668 : _GEN_6876; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6878 = 12'h29d == _T_96[11:0] ? image_669 : _GEN_6877; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6879 = 12'h29e == _T_96[11:0] ? image_670 : _GEN_6878; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6880 = 12'h29f == _T_96[11:0] ? 4'h0 : _GEN_6879; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6881 = 12'h2a0 == _T_96[11:0] ? 4'h0 : _GEN_6880; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6882 = 12'h2a1 == _T_96[11:0] ? 4'h0 : _GEN_6881; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6883 = 12'h2a2 == _T_96[11:0] ? 4'h0 : _GEN_6882; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6884 = 12'h2a3 == _T_96[11:0] ? 4'h0 : _GEN_6883; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6885 = 12'h2a4 == _T_96[11:0] ? 4'h0 : _GEN_6884; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6886 = 12'h2a5 == _T_96[11:0] ? 4'h0 : _GEN_6885; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6887 = 12'h2a6 == _T_96[11:0] ? 4'h0 : _GEN_6886; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6888 = 12'h2a7 == _T_96[11:0] ? image_679 : _GEN_6887; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6889 = 12'h2a8 == _T_96[11:0] ? image_680 : _GEN_6888; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6890 = 12'h2a9 == _T_96[11:0] ? image_681 : _GEN_6889; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6891 = 12'h2aa == _T_96[11:0] ? image_682 : _GEN_6890; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6892 = 12'h2ab == _T_96[11:0] ? image_683 : _GEN_6891; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6893 = 12'h2ac == _T_96[11:0] ? image_684 : _GEN_6892; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6894 = 12'h2ad == _T_96[11:0] ? image_685 : _GEN_6893; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6895 = 12'h2ae == _T_96[11:0] ? image_686 : _GEN_6894; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6896 = 12'h2af == _T_96[11:0] ? image_687 : _GEN_6895; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6897 = 12'h2b0 == _T_96[11:0] ? image_688 : _GEN_6896; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6898 = 12'h2b1 == _T_96[11:0] ? image_689 : _GEN_6897; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6899 = 12'h2b2 == _T_96[11:0] ? image_690 : _GEN_6898; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6900 = 12'h2b3 == _T_96[11:0] ? image_691 : _GEN_6899; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6901 = 12'h2b4 == _T_96[11:0] ? image_692 : _GEN_6900; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6902 = 12'h2b5 == _T_96[11:0] ? image_693 : _GEN_6901; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6903 = 12'h2b6 == _T_96[11:0] ? image_694 : _GEN_6902; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6904 = 12'h2b7 == _T_96[11:0] ? image_695 : _GEN_6903; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6905 = 12'h2b8 == _T_96[11:0] ? image_696 : _GEN_6904; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6906 = 12'h2b9 == _T_96[11:0] ? image_697 : _GEN_6905; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6907 = 12'h2ba == _T_96[11:0] ? image_698 : _GEN_6906; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6908 = 12'h2bb == _T_96[11:0] ? 4'h0 : _GEN_6907; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6909 = 12'h2bc == _T_96[11:0] ? 4'h0 : _GEN_6908; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6910 = 12'h2bd == _T_96[11:0] ? image_701 : _GEN_6909; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6911 = 12'h2be == _T_96[11:0] ? image_702 : _GEN_6910; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6912 = 12'h2bf == _T_96[11:0] ? image_703 : _GEN_6911; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6913 = 12'h2c0 == _T_96[11:0] ? 4'h0 : _GEN_6912; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6914 = 12'h2c1 == _T_96[11:0] ? image_705 : _GEN_6913; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6915 = 12'h2c2 == _T_96[11:0] ? image_706 : _GEN_6914; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6916 = 12'h2c3 == _T_96[11:0] ? image_707 : _GEN_6915; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6917 = 12'h2c4 == _T_96[11:0] ? image_708 : _GEN_6916; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6918 = 12'h2c5 == _T_96[11:0] ? image_709 : _GEN_6917; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6919 = 12'h2c6 == _T_96[11:0] ? image_710 : _GEN_6918; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6920 = 12'h2c7 == _T_96[11:0] ? image_711 : _GEN_6919; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6921 = 12'h2c8 == _T_96[11:0] ? image_712 : _GEN_6920; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6922 = 12'h2c9 == _T_96[11:0] ? image_713 : _GEN_6921; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6923 = 12'h2ca == _T_96[11:0] ? image_714 : _GEN_6922; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6924 = 12'h2cb == _T_96[11:0] ? image_715 : _GEN_6923; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6925 = 12'h2cc == _T_96[11:0] ? image_716 : _GEN_6924; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6926 = 12'h2cd == _T_96[11:0] ? image_717 : _GEN_6925; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6927 = 12'h2ce == _T_96[11:0] ? image_718 : _GEN_6926; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6928 = 12'h2cf == _T_96[11:0] ? image_719 : _GEN_6927; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6929 = 12'h2d0 == _T_96[11:0] ? image_720 : _GEN_6928; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6930 = 12'h2d1 == _T_96[11:0] ? image_721 : _GEN_6929; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6931 = 12'h2d2 == _T_96[11:0] ? image_722 : _GEN_6930; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6932 = 12'h2d3 == _T_96[11:0] ? image_723 : _GEN_6931; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6933 = 12'h2d4 == _T_96[11:0] ? image_724 : _GEN_6932; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6934 = 12'h2d5 == _T_96[11:0] ? image_725 : _GEN_6933; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6935 = 12'h2d6 == _T_96[11:0] ? image_726 : _GEN_6934; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6936 = 12'h2d7 == _T_96[11:0] ? image_727 : _GEN_6935; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6937 = 12'h2d8 == _T_96[11:0] ? image_728 : _GEN_6936; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6938 = 12'h2d9 == _T_96[11:0] ? image_729 : _GEN_6937; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6939 = 12'h2da == _T_96[11:0] ? image_730 : _GEN_6938; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6940 = 12'h2db == _T_96[11:0] ? image_731 : _GEN_6939; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6941 = 12'h2dc == _T_96[11:0] ? image_732 : _GEN_6940; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6942 = 12'h2dd == _T_96[11:0] ? image_733 : _GEN_6941; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6943 = 12'h2de == _T_96[11:0] ? image_734 : _GEN_6942; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6944 = 12'h2df == _T_96[11:0] ? 4'h0 : _GEN_6943; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6945 = 12'h2e0 == _T_96[11:0] ? image_736 : _GEN_6944; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6946 = 12'h2e1 == _T_96[11:0] ? image_737 : _GEN_6945; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6947 = 12'h2e2 == _T_96[11:0] ? 4'h0 : _GEN_6946; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6948 = 12'h2e3 == _T_96[11:0] ? image_739 : _GEN_6947; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6949 = 12'h2e4 == _T_96[11:0] ? image_740 : _GEN_6948; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6950 = 12'h2e5 == _T_96[11:0] ? image_741 : _GEN_6949; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6951 = 12'h2e6 == _T_96[11:0] ? 4'h0 : _GEN_6950; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6952 = 12'h2e7 == _T_96[11:0] ? 4'h0 : _GEN_6951; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6953 = 12'h2e8 == _T_96[11:0] ? image_744 : _GEN_6952; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6954 = 12'h2e9 == _T_96[11:0] ? image_745 : _GEN_6953; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6955 = 12'h2ea == _T_96[11:0] ? image_746 : _GEN_6954; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6956 = 12'h2eb == _T_96[11:0] ? image_747 : _GEN_6955; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6957 = 12'h2ec == _T_96[11:0] ? image_748 : _GEN_6956; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6958 = 12'h2ed == _T_96[11:0] ? image_749 : _GEN_6957; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6959 = 12'h2ee == _T_96[11:0] ? image_750 : _GEN_6958; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6960 = 12'h2ef == _T_96[11:0] ? image_751 : _GEN_6959; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6961 = 12'h2f0 == _T_96[11:0] ? image_752 : _GEN_6960; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6962 = 12'h2f1 == _T_96[11:0] ? image_753 : _GEN_6961; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6963 = 12'h2f2 == _T_96[11:0] ? image_754 : _GEN_6962; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6964 = 12'h2f3 == _T_96[11:0] ? image_755 : _GEN_6963; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6965 = 12'h2f4 == _T_96[11:0] ? image_756 : _GEN_6964; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6966 = 12'h2f5 == _T_96[11:0] ? 4'h0 : _GEN_6965; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6967 = 12'h2f6 == _T_96[11:0] ? image_758 : _GEN_6966; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6968 = 12'h2f7 == _T_96[11:0] ? 4'h0 : _GEN_6967; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6969 = 12'h2f8 == _T_96[11:0] ? image_760 : _GEN_6968; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6970 = 12'h2f9 == _T_96[11:0] ? image_761 : _GEN_6969; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6971 = 12'h2fa == _T_96[11:0] ? image_762 : _GEN_6970; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6972 = 12'h2fb == _T_96[11:0] ? image_763 : _GEN_6971; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6973 = 12'h2fc == _T_96[11:0] ? 4'h0 : _GEN_6972; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6974 = 12'h2fd == _T_96[11:0] ? image_765 : _GEN_6973; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6975 = 12'h2fe == _T_96[11:0] ? image_766 : _GEN_6974; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6976 = 12'h2ff == _T_96[11:0] ? image_767 : _GEN_6975; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6977 = 12'h300 == _T_96[11:0] ? image_768 : _GEN_6976; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6978 = 12'h301 == _T_96[11:0] ? image_769 : _GEN_6977; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6979 = 12'h302 == _T_96[11:0] ? image_770 : _GEN_6978; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6980 = 12'h303 == _T_96[11:0] ? image_771 : _GEN_6979; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6981 = 12'h304 == _T_96[11:0] ? image_772 : _GEN_6980; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6982 = 12'h305 == _T_96[11:0] ? image_773 : _GEN_6981; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6983 = 12'h306 == _T_96[11:0] ? image_774 : _GEN_6982; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6984 = 12'h307 == _T_96[11:0] ? image_775 : _GEN_6983; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6985 = 12'h308 == _T_96[11:0] ? image_776 : _GEN_6984; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6986 = 12'h309 == _T_96[11:0] ? image_777 : _GEN_6985; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6987 = 12'h30a == _T_96[11:0] ? image_778 : _GEN_6986; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6988 = 12'h30b == _T_96[11:0] ? image_779 : _GEN_6987; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6989 = 12'h30c == _T_96[11:0] ? image_780 : _GEN_6988; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6990 = 12'h30d == _T_96[11:0] ? image_781 : _GEN_6989; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6991 = 12'h30e == _T_96[11:0] ? image_782 : _GEN_6990; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6992 = 12'h30f == _T_96[11:0] ? image_783 : _GEN_6991; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6993 = 12'h310 == _T_96[11:0] ? image_784 : _GEN_6992; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6994 = 12'h311 == _T_96[11:0] ? image_785 : _GEN_6993; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6995 = 12'h312 == _T_96[11:0] ? image_786 : _GEN_6994; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6996 = 12'h313 == _T_96[11:0] ? image_787 : _GEN_6995; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6997 = 12'h314 == _T_96[11:0] ? image_788 : _GEN_6996; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6998 = 12'h315 == _T_96[11:0] ? image_789 : _GEN_6997; // @[Filter.scala 138:46]
  wire [3:0] _GEN_6999 = 12'h316 == _T_96[11:0] ? image_790 : _GEN_6998; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7000 = 12'h317 == _T_96[11:0] ? image_791 : _GEN_6999; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7001 = 12'h318 == _T_96[11:0] ? image_792 : _GEN_7000; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7002 = 12'h319 == _T_96[11:0] ? image_793 : _GEN_7001; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7003 = 12'h31a == _T_96[11:0] ? image_794 : _GEN_7002; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7004 = 12'h31b == _T_96[11:0] ? image_795 : _GEN_7003; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7005 = 12'h31c == _T_96[11:0] ? image_796 : _GEN_7004; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7006 = 12'h31d == _T_96[11:0] ? image_797 : _GEN_7005; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7007 = 12'h31e == _T_96[11:0] ? 4'h0 : _GEN_7006; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7008 = 12'h31f == _T_96[11:0] ? 4'h0 : _GEN_7007; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7009 = 12'h320 == _T_96[11:0] ? image_800 : _GEN_7008; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7010 = 12'h321 == _T_96[11:0] ? image_801 : _GEN_7009; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7011 = 12'h322 == _T_96[11:0] ? image_802 : _GEN_7010; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7012 = 12'h323 == _T_96[11:0] ? image_803 : _GEN_7011; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7013 = 12'h324 == _T_96[11:0] ? image_804 : _GEN_7012; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7014 = 12'h325 == _T_96[11:0] ? image_805 : _GEN_7013; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7015 = 12'h326 == _T_96[11:0] ? image_806 : _GEN_7014; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7016 = 12'h327 == _T_96[11:0] ? 4'h0 : _GEN_7015; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7017 = 12'h328 == _T_96[11:0] ? image_808 : _GEN_7016; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7018 = 12'h329 == _T_96[11:0] ? image_809 : _GEN_7017; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7019 = 12'h32a == _T_96[11:0] ? image_810 : _GEN_7018; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7020 = 12'h32b == _T_96[11:0] ? image_811 : _GEN_7019; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7021 = 12'h32c == _T_96[11:0] ? image_812 : _GEN_7020; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7022 = 12'h32d == _T_96[11:0] ? image_813 : _GEN_7021; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7023 = 12'h32e == _T_96[11:0] ? image_814 : _GEN_7022; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7024 = 12'h32f == _T_96[11:0] ? image_815 : _GEN_7023; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7025 = 12'h330 == _T_96[11:0] ? image_816 : _GEN_7024; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7026 = 12'h331 == _T_96[11:0] ? image_817 : _GEN_7025; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7027 = 12'h332 == _T_96[11:0] ? image_818 : _GEN_7026; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7028 = 12'h333 == _T_96[11:0] ? image_819 : _GEN_7027; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7029 = 12'h334 == _T_96[11:0] ? image_820 : _GEN_7028; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7030 = 12'h335 == _T_96[11:0] ? 4'h0 : _GEN_7029; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7031 = 12'h336 == _T_96[11:0] ? image_822 : _GEN_7030; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7032 = 12'h337 == _T_96[11:0] ? image_823 : _GEN_7031; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7033 = 12'h338 == _T_96[11:0] ? image_824 : _GEN_7032; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7034 = 12'h339 == _T_96[11:0] ? image_825 : _GEN_7033; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7035 = 12'h33a == _T_96[11:0] ? image_826 : _GEN_7034; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7036 = 12'h33b == _T_96[11:0] ? 4'h0 : _GEN_7035; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7037 = 12'h33c == _T_96[11:0] ? image_828 : _GEN_7036; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7038 = 12'h33d == _T_96[11:0] ? image_829 : _GEN_7037; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7039 = 12'h33e == _T_96[11:0] ? image_830 : _GEN_7038; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7040 = 12'h33f == _T_96[11:0] ? image_831 : _GEN_7039; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7041 = 12'h340 == _T_96[11:0] ? 4'h0 : _GEN_7040; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7042 = 12'h341 == _T_96[11:0] ? image_833 : _GEN_7041; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7043 = 12'h342 == _T_96[11:0] ? image_834 : _GEN_7042; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7044 = 12'h343 == _T_96[11:0] ? image_835 : _GEN_7043; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7045 = 12'h344 == _T_96[11:0] ? image_836 : _GEN_7044; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7046 = 12'h345 == _T_96[11:0] ? image_837 : _GEN_7045; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7047 = 12'h346 == _T_96[11:0] ? image_838 : _GEN_7046; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7048 = 12'h347 == _T_96[11:0] ? image_839 : _GEN_7047; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7049 = 12'h348 == _T_96[11:0] ? image_840 : _GEN_7048; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7050 = 12'h349 == _T_96[11:0] ? image_841 : _GEN_7049; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7051 = 12'h34a == _T_96[11:0] ? image_842 : _GEN_7050; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7052 = 12'h34b == _T_96[11:0] ? image_843 : _GEN_7051; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7053 = 12'h34c == _T_96[11:0] ? image_844 : _GEN_7052; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7054 = 12'h34d == _T_96[11:0] ? image_845 : _GEN_7053; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7055 = 12'h34e == _T_96[11:0] ? image_846 : _GEN_7054; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7056 = 12'h34f == _T_96[11:0] ? image_847 : _GEN_7055; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7057 = 12'h350 == _T_96[11:0] ? image_848 : _GEN_7056; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7058 = 12'h351 == _T_96[11:0] ? image_849 : _GEN_7057; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7059 = 12'h352 == _T_96[11:0] ? image_850 : _GEN_7058; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7060 = 12'h353 == _T_96[11:0] ? image_851 : _GEN_7059; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7061 = 12'h354 == _T_96[11:0] ? image_852 : _GEN_7060; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7062 = 12'h355 == _T_96[11:0] ? image_853 : _GEN_7061; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7063 = 12'h356 == _T_96[11:0] ? image_854 : _GEN_7062; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7064 = 12'h357 == _T_96[11:0] ? image_855 : _GEN_7063; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7065 = 12'h358 == _T_96[11:0] ? image_856 : _GEN_7064; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7066 = 12'h359 == _T_96[11:0] ? image_857 : _GEN_7065; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7067 = 12'h35a == _T_96[11:0] ? image_858 : _GEN_7066; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7068 = 12'h35b == _T_96[11:0] ? image_859 : _GEN_7067; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7069 = 12'h35c == _T_96[11:0] ? image_860 : _GEN_7068; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7070 = 12'h35d == _T_96[11:0] ? image_861 : _GEN_7069; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7071 = 12'h35e == _T_96[11:0] ? image_862 : _GEN_7070; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7072 = 12'h35f == _T_96[11:0] ? 4'h0 : _GEN_7071; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7073 = 12'h360 == _T_96[11:0] ? 4'h0 : _GEN_7072; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7074 = 12'h361 == _T_96[11:0] ? image_865 : _GEN_7073; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7075 = 12'h362 == _T_96[11:0] ? image_866 : _GEN_7074; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7076 = 12'h363 == _T_96[11:0] ? image_867 : _GEN_7075; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7077 = 12'h364 == _T_96[11:0] ? image_868 : _GEN_7076; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7078 = 12'h365 == _T_96[11:0] ? image_869 : _GEN_7077; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7079 = 12'h366 == _T_96[11:0] ? 4'h0 : _GEN_7078; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7080 = 12'h367 == _T_96[11:0] ? 4'h0 : _GEN_7079; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7081 = 12'h368 == _T_96[11:0] ? image_872 : _GEN_7080; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7082 = 12'h369 == _T_96[11:0] ? image_873 : _GEN_7081; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7083 = 12'h36a == _T_96[11:0] ? image_874 : _GEN_7082; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7084 = 12'h36b == _T_96[11:0] ? image_875 : _GEN_7083; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7085 = 12'h36c == _T_96[11:0] ? image_876 : _GEN_7084; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7086 = 12'h36d == _T_96[11:0] ? image_877 : _GEN_7085; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7087 = 12'h36e == _T_96[11:0] ? image_878 : _GEN_7086; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7088 = 12'h36f == _T_96[11:0] ? image_879 : _GEN_7087; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7089 = 12'h370 == _T_96[11:0] ? image_880 : _GEN_7088; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7090 = 12'h371 == _T_96[11:0] ? image_881 : _GEN_7089; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7091 = 12'h372 == _T_96[11:0] ? image_882 : _GEN_7090; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7092 = 12'h373 == _T_96[11:0] ? image_883 : _GEN_7091; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7093 = 12'h374 == _T_96[11:0] ? image_884 : _GEN_7092; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7094 = 12'h375 == _T_96[11:0] ? image_885 : _GEN_7093; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7095 = 12'h376 == _T_96[11:0] ? 4'h0 : _GEN_7094; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7096 = 12'h377 == _T_96[11:0] ? 4'h0 : _GEN_7095; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7097 = 12'h378 == _T_96[11:0] ? 4'h0 : _GEN_7096; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7098 = 12'h379 == _T_96[11:0] ? 4'h0 : _GEN_7097; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7099 = 12'h37a == _T_96[11:0] ? 4'h0 : _GEN_7098; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7100 = 12'h37b == _T_96[11:0] ? image_891 : _GEN_7099; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7101 = 12'h37c == _T_96[11:0] ? image_892 : _GEN_7100; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7102 = 12'h37d == _T_96[11:0] ? image_893 : _GEN_7101; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7103 = 12'h37e == _T_96[11:0] ? image_894 : _GEN_7102; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7104 = 12'h37f == _T_96[11:0] ? image_895 : _GEN_7103; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7105 = 12'h380 == _T_96[11:0] ? 4'h0 : _GEN_7104; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7106 = 12'h381 == _T_96[11:0] ? image_897 : _GEN_7105; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7107 = 12'h382 == _T_96[11:0] ? image_898 : _GEN_7106; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7108 = 12'h383 == _T_96[11:0] ? image_899 : _GEN_7107; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7109 = 12'h384 == _T_96[11:0] ? image_900 : _GEN_7108; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7110 = 12'h385 == _T_96[11:0] ? image_901 : _GEN_7109; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7111 = 12'h386 == _T_96[11:0] ? image_902 : _GEN_7110; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7112 = 12'h387 == _T_96[11:0] ? image_903 : _GEN_7111; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7113 = 12'h388 == _T_96[11:0] ? image_904 : _GEN_7112; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7114 = 12'h389 == _T_96[11:0] ? image_905 : _GEN_7113; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7115 = 12'h38a == _T_96[11:0] ? image_906 : _GEN_7114; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7116 = 12'h38b == _T_96[11:0] ? image_907 : _GEN_7115; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7117 = 12'h38c == _T_96[11:0] ? image_908 : _GEN_7116; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7118 = 12'h38d == _T_96[11:0] ? image_909 : _GEN_7117; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7119 = 12'h38e == _T_96[11:0] ? image_910 : _GEN_7118; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7120 = 12'h38f == _T_96[11:0] ? image_911 : _GEN_7119; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7121 = 12'h390 == _T_96[11:0] ? image_912 : _GEN_7120; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7122 = 12'h391 == _T_96[11:0] ? image_913 : _GEN_7121; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7123 = 12'h392 == _T_96[11:0] ? image_914 : _GEN_7122; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7124 = 12'h393 == _T_96[11:0] ? image_915 : _GEN_7123; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7125 = 12'h394 == _T_96[11:0] ? image_916 : _GEN_7124; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7126 = 12'h395 == _T_96[11:0] ? image_917 : _GEN_7125; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7127 = 12'h396 == _T_96[11:0] ? image_918 : _GEN_7126; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7128 = 12'h397 == _T_96[11:0] ? image_919 : _GEN_7127; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7129 = 12'h398 == _T_96[11:0] ? image_920 : _GEN_7128; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7130 = 12'h399 == _T_96[11:0] ? image_921 : _GEN_7129; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7131 = 12'h39a == _T_96[11:0] ? image_922 : _GEN_7130; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7132 = 12'h39b == _T_96[11:0] ? image_923 : _GEN_7131; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7133 = 12'h39c == _T_96[11:0] ? image_924 : _GEN_7132; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7134 = 12'h39d == _T_96[11:0] ? image_925 : _GEN_7133; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7135 = 12'h39e == _T_96[11:0] ? image_926 : _GEN_7134; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7136 = 12'h39f == _T_96[11:0] ? image_927 : _GEN_7135; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7137 = 12'h3a0 == _T_96[11:0] ? 4'h0 : _GEN_7136; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7138 = 12'h3a1 == _T_96[11:0] ? image_929 : _GEN_7137; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7139 = 12'h3a2 == _T_96[11:0] ? image_930 : _GEN_7138; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7140 = 12'h3a3 == _T_96[11:0] ? 4'h0 : _GEN_7139; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7141 = 12'h3a4 == _T_96[11:0] ? 4'h0 : _GEN_7140; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7142 = 12'h3a5 == _T_96[11:0] ? 4'h0 : _GEN_7141; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7143 = 12'h3a6 == _T_96[11:0] ? 4'h0 : _GEN_7142; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7144 = 12'h3a7 == _T_96[11:0] ? image_935 : _GEN_7143; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7145 = 12'h3a8 == _T_96[11:0] ? image_936 : _GEN_7144; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7146 = 12'h3a9 == _T_96[11:0] ? image_937 : _GEN_7145; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7147 = 12'h3aa == _T_96[11:0] ? image_938 : _GEN_7146; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7148 = 12'h3ab == _T_96[11:0] ? image_939 : _GEN_7147; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7149 = 12'h3ac == _T_96[11:0] ? image_940 : _GEN_7148; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7150 = 12'h3ad == _T_96[11:0] ? image_941 : _GEN_7149; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7151 = 12'h3ae == _T_96[11:0] ? image_942 : _GEN_7150; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7152 = 12'h3af == _T_96[11:0] ? image_943 : _GEN_7151; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7153 = 12'h3b0 == _T_96[11:0] ? image_944 : _GEN_7152; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7154 = 12'h3b1 == _T_96[11:0] ? image_945 : _GEN_7153; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7155 = 12'h3b2 == _T_96[11:0] ? image_946 : _GEN_7154; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7156 = 12'h3b3 == _T_96[11:0] ? image_947 : _GEN_7155; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7157 = 12'h3b4 == _T_96[11:0] ? image_948 : _GEN_7156; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7158 = 12'h3b5 == _T_96[11:0] ? image_949 : _GEN_7157; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7159 = 12'h3b6 == _T_96[11:0] ? image_950 : _GEN_7158; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7160 = 12'h3b7 == _T_96[11:0] ? image_951 : _GEN_7159; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7161 = 12'h3b8 == _T_96[11:0] ? image_952 : _GEN_7160; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7162 = 12'h3b9 == _T_96[11:0] ? image_953 : _GEN_7161; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7163 = 12'h3ba == _T_96[11:0] ? image_954 : _GEN_7162; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7164 = 12'h3bb == _T_96[11:0] ? image_955 : _GEN_7163; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7165 = 12'h3bc == _T_96[11:0] ? image_956 : _GEN_7164; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7166 = 12'h3bd == _T_96[11:0] ? image_957 : _GEN_7165; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7167 = 12'h3be == _T_96[11:0] ? image_958 : _GEN_7166; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7168 = 12'h3bf == _T_96[11:0] ? image_959 : _GEN_7167; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7169 = 12'h3c0 == _T_96[11:0] ? 4'h0 : _GEN_7168; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7170 = 12'h3c1 == _T_96[11:0] ? image_961 : _GEN_7169; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7171 = 12'h3c2 == _T_96[11:0] ? image_962 : _GEN_7170; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7172 = 12'h3c3 == _T_96[11:0] ? image_963 : _GEN_7171; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7173 = 12'h3c4 == _T_96[11:0] ? image_964 : _GEN_7172; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7174 = 12'h3c5 == _T_96[11:0] ? image_965 : _GEN_7173; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7175 = 12'h3c6 == _T_96[11:0] ? image_966 : _GEN_7174; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7176 = 12'h3c7 == _T_96[11:0] ? image_967 : _GEN_7175; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7177 = 12'h3c8 == _T_96[11:0] ? image_968 : _GEN_7176; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7178 = 12'h3c9 == _T_96[11:0] ? image_969 : _GEN_7177; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7179 = 12'h3ca == _T_96[11:0] ? image_970 : _GEN_7178; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7180 = 12'h3cb == _T_96[11:0] ? image_971 : _GEN_7179; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7181 = 12'h3cc == _T_96[11:0] ? image_972 : _GEN_7180; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7182 = 12'h3cd == _T_96[11:0] ? image_973 : _GEN_7181; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7183 = 12'h3ce == _T_96[11:0] ? image_974 : _GEN_7182; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7184 = 12'h3cf == _T_96[11:0] ? image_975 : _GEN_7183; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7185 = 12'h3d0 == _T_96[11:0] ? image_976 : _GEN_7184; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7186 = 12'h3d1 == _T_96[11:0] ? image_977 : _GEN_7185; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7187 = 12'h3d2 == _T_96[11:0] ? image_978 : _GEN_7186; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7188 = 12'h3d3 == _T_96[11:0] ? image_979 : _GEN_7187; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7189 = 12'h3d4 == _T_96[11:0] ? image_980 : _GEN_7188; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7190 = 12'h3d5 == _T_96[11:0] ? image_981 : _GEN_7189; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7191 = 12'h3d6 == _T_96[11:0] ? image_982 : _GEN_7190; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7192 = 12'h3d7 == _T_96[11:0] ? image_983 : _GEN_7191; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7193 = 12'h3d8 == _T_96[11:0] ? image_984 : _GEN_7192; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7194 = 12'h3d9 == _T_96[11:0] ? image_985 : _GEN_7193; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7195 = 12'h3da == _T_96[11:0] ? image_986 : _GEN_7194; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7196 = 12'h3db == _T_96[11:0] ? image_987 : _GEN_7195; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7197 = 12'h3dc == _T_96[11:0] ? image_988 : _GEN_7196; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7198 = 12'h3dd == _T_96[11:0] ? image_989 : _GEN_7197; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7199 = 12'h3de == _T_96[11:0] ? image_990 : _GEN_7198; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7200 = 12'h3df == _T_96[11:0] ? image_991 : _GEN_7199; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7201 = 12'h3e0 == _T_96[11:0] ? image_992 : _GEN_7200; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7202 = 12'h3e1 == _T_96[11:0] ? 4'h0 : _GEN_7201; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7203 = 12'h3e2 == _T_96[11:0] ? 4'h0 : _GEN_7202; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7204 = 12'h3e3 == _T_96[11:0] ? 4'h0 : _GEN_7203; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7205 = 12'h3e4 == _T_96[11:0] ? 4'h0 : _GEN_7204; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7206 = 12'h3e5 == _T_96[11:0] ? image_997 : _GEN_7205; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7207 = 12'h3e6 == _T_96[11:0] ? image_998 : _GEN_7206; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7208 = 12'h3e7 == _T_96[11:0] ? image_999 : _GEN_7207; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7209 = 12'h3e8 == _T_96[11:0] ? image_1000 : _GEN_7208; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7210 = 12'h3e9 == _T_96[11:0] ? image_1001 : _GEN_7209; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7211 = 12'h3ea == _T_96[11:0] ? image_1002 : _GEN_7210; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7212 = 12'h3eb == _T_96[11:0] ? image_1003 : _GEN_7211; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7213 = 12'h3ec == _T_96[11:0] ? image_1004 : _GEN_7212; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7214 = 12'h3ed == _T_96[11:0] ? image_1005 : _GEN_7213; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7215 = 12'h3ee == _T_96[11:0] ? image_1006 : _GEN_7214; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7216 = 12'h3ef == _T_96[11:0] ? image_1007 : _GEN_7215; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7217 = 12'h3f0 == _T_96[11:0] ? image_1008 : _GEN_7216; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7218 = 12'h3f1 == _T_96[11:0] ? image_1009 : _GEN_7217; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7219 = 12'h3f2 == _T_96[11:0] ? image_1010 : _GEN_7218; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7220 = 12'h3f3 == _T_96[11:0] ? image_1011 : _GEN_7219; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7221 = 12'h3f4 == _T_96[11:0] ? image_1012 : _GEN_7220; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7222 = 12'h3f5 == _T_96[11:0] ? image_1013 : _GEN_7221; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7223 = 12'h3f6 == _T_96[11:0] ? image_1014 : _GEN_7222; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7224 = 12'h3f7 == _T_96[11:0] ? image_1015 : _GEN_7223; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7225 = 12'h3f8 == _T_96[11:0] ? image_1016 : _GEN_7224; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7226 = 12'h3f9 == _T_96[11:0] ? image_1017 : _GEN_7225; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7227 = 12'h3fa == _T_96[11:0] ? image_1018 : _GEN_7226; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7228 = 12'h3fb == _T_96[11:0] ? image_1019 : _GEN_7227; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7229 = 12'h3fc == _T_96[11:0] ? image_1020 : _GEN_7228; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7230 = 12'h3fd == _T_96[11:0] ? 4'h0 : _GEN_7229; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7231 = 12'h3fe == _T_96[11:0] ? 4'h0 : _GEN_7230; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7232 = 12'h3ff == _T_96[11:0] ? 4'h0 : _GEN_7231; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7233 = 12'h400 == _T_96[11:0] ? image_1024 : _GEN_7232; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7234 = 12'h401 == _T_96[11:0] ? image_1025 : _GEN_7233; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7235 = 12'h402 == _T_96[11:0] ? image_1026 : _GEN_7234; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7236 = 12'h403 == _T_96[11:0] ? image_1027 : _GEN_7235; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7237 = 12'h404 == _T_96[11:0] ? image_1028 : _GEN_7236; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7238 = 12'h405 == _T_96[11:0] ? image_1029 : _GEN_7237; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7239 = 12'h406 == _T_96[11:0] ? image_1030 : _GEN_7238; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7240 = 12'h407 == _T_96[11:0] ? image_1031 : _GEN_7239; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7241 = 12'h408 == _T_96[11:0] ? image_1032 : _GEN_7240; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7242 = 12'h409 == _T_96[11:0] ? image_1033 : _GEN_7241; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7243 = 12'h40a == _T_96[11:0] ? image_1034 : _GEN_7242; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7244 = 12'h40b == _T_96[11:0] ? image_1035 : _GEN_7243; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7245 = 12'h40c == _T_96[11:0] ? image_1036 : _GEN_7244; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7246 = 12'h40d == _T_96[11:0] ? image_1037 : _GEN_7245; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7247 = 12'h40e == _T_96[11:0] ? image_1038 : _GEN_7246; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7248 = 12'h40f == _T_96[11:0] ? image_1039 : _GEN_7247; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7249 = 12'h410 == _T_96[11:0] ? image_1040 : _GEN_7248; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7250 = 12'h411 == _T_96[11:0] ? image_1041 : _GEN_7249; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7251 = 12'h412 == _T_96[11:0] ? image_1042 : _GEN_7250; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7252 = 12'h413 == _T_96[11:0] ? image_1043 : _GEN_7251; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7253 = 12'h414 == _T_96[11:0] ? image_1044 : _GEN_7252; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7254 = 12'h415 == _T_96[11:0] ? image_1045 : _GEN_7253; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7255 = 12'h416 == _T_96[11:0] ? image_1046 : _GEN_7254; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7256 = 12'h417 == _T_96[11:0] ? image_1047 : _GEN_7255; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7257 = 12'h418 == _T_96[11:0] ? image_1048 : _GEN_7256; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7258 = 12'h419 == _T_96[11:0] ? image_1049 : _GEN_7257; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7259 = 12'h41a == _T_96[11:0] ? image_1050 : _GEN_7258; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7260 = 12'h41b == _T_96[11:0] ? image_1051 : _GEN_7259; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7261 = 12'h41c == _T_96[11:0] ? image_1052 : _GEN_7260; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7262 = 12'h41d == _T_96[11:0] ? image_1053 : _GEN_7261; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7263 = 12'h41e == _T_96[11:0] ? image_1054 : _GEN_7262; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7264 = 12'h41f == _T_96[11:0] ? image_1055 : _GEN_7263; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7265 = 12'h420 == _T_96[11:0] ? image_1056 : _GEN_7264; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7266 = 12'h421 == _T_96[11:0] ? image_1057 : _GEN_7265; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7267 = 12'h422 == _T_96[11:0] ? image_1058 : _GEN_7266; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7268 = 12'h423 == _T_96[11:0] ? image_1059 : _GEN_7267; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7269 = 12'h424 == _T_96[11:0] ? image_1060 : _GEN_7268; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7270 = 12'h425 == _T_96[11:0] ? image_1061 : _GEN_7269; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7271 = 12'h426 == _T_96[11:0] ? image_1062 : _GEN_7270; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7272 = 12'h427 == _T_96[11:0] ? image_1063 : _GEN_7271; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7273 = 12'h428 == _T_96[11:0] ? image_1064 : _GEN_7272; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7274 = 12'h429 == _T_96[11:0] ? image_1065 : _GEN_7273; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7275 = 12'h42a == _T_96[11:0] ? image_1066 : _GEN_7274; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7276 = 12'h42b == _T_96[11:0] ? image_1067 : _GEN_7275; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7277 = 12'h42c == _T_96[11:0] ? image_1068 : _GEN_7276; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7278 = 12'h42d == _T_96[11:0] ? image_1069 : _GEN_7277; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7279 = 12'h42e == _T_96[11:0] ? image_1070 : _GEN_7278; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7280 = 12'h42f == _T_96[11:0] ? image_1071 : _GEN_7279; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7281 = 12'h430 == _T_96[11:0] ? image_1072 : _GEN_7280; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7282 = 12'h431 == _T_96[11:0] ? image_1073 : _GEN_7281; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7283 = 12'h432 == _T_96[11:0] ? image_1074 : _GEN_7282; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7284 = 12'h433 == _T_96[11:0] ? image_1075 : _GEN_7283; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7285 = 12'h434 == _T_96[11:0] ? image_1076 : _GEN_7284; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7286 = 12'h435 == _T_96[11:0] ? image_1077 : _GEN_7285; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7287 = 12'h436 == _T_96[11:0] ? image_1078 : _GEN_7286; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7288 = 12'h437 == _T_96[11:0] ? image_1079 : _GEN_7287; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7289 = 12'h438 == _T_96[11:0] ? image_1080 : _GEN_7288; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7290 = 12'h439 == _T_96[11:0] ? image_1081 : _GEN_7289; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7291 = 12'h43a == _T_96[11:0] ? image_1082 : _GEN_7290; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7292 = 12'h43b == _T_96[11:0] ? image_1083 : _GEN_7291; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7293 = 12'h43c == _T_96[11:0] ? image_1084 : _GEN_7292; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7294 = 12'h43d == _T_96[11:0] ? image_1085 : _GEN_7293; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7295 = 12'h43e == _T_96[11:0] ? 4'h0 : _GEN_7294; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7296 = 12'h43f == _T_96[11:0] ? 4'h0 : _GEN_7295; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7297 = 12'h440 == _T_96[11:0] ? image_1088 : _GEN_7296; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7298 = 12'h441 == _T_96[11:0] ? image_1089 : _GEN_7297; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7299 = 12'h442 == _T_96[11:0] ? image_1090 : _GEN_7298; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7300 = 12'h443 == _T_96[11:0] ? image_1091 : _GEN_7299; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7301 = 12'h444 == _T_96[11:0] ? image_1092 : _GEN_7300; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7302 = 12'h445 == _T_96[11:0] ? image_1093 : _GEN_7301; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7303 = 12'h446 == _T_96[11:0] ? image_1094 : _GEN_7302; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7304 = 12'h447 == _T_96[11:0] ? image_1095 : _GEN_7303; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7305 = 12'h448 == _T_96[11:0] ? image_1096 : _GEN_7304; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7306 = 12'h449 == _T_96[11:0] ? image_1097 : _GEN_7305; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7307 = 12'h44a == _T_96[11:0] ? image_1098 : _GEN_7306; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7308 = 12'h44b == _T_96[11:0] ? image_1099 : _GEN_7307; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7309 = 12'h44c == _T_96[11:0] ? image_1100 : _GEN_7308; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7310 = 12'h44d == _T_96[11:0] ? image_1101 : _GEN_7309; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7311 = 12'h44e == _T_96[11:0] ? image_1102 : _GEN_7310; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7312 = 12'h44f == _T_96[11:0] ? image_1103 : _GEN_7311; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7313 = 12'h450 == _T_96[11:0] ? image_1104 : _GEN_7312; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7314 = 12'h451 == _T_96[11:0] ? image_1105 : _GEN_7313; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7315 = 12'h452 == _T_96[11:0] ? image_1106 : _GEN_7314; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7316 = 12'h453 == _T_96[11:0] ? image_1107 : _GEN_7315; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7317 = 12'h454 == _T_96[11:0] ? image_1108 : _GEN_7316; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7318 = 12'h455 == _T_96[11:0] ? image_1109 : _GEN_7317; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7319 = 12'h456 == _T_96[11:0] ? image_1110 : _GEN_7318; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7320 = 12'h457 == _T_96[11:0] ? image_1111 : _GEN_7319; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7321 = 12'h458 == _T_96[11:0] ? image_1112 : _GEN_7320; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7322 = 12'h459 == _T_96[11:0] ? image_1113 : _GEN_7321; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7323 = 12'h45a == _T_96[11:0] ? image_1114 : _GEN_7322; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7324 = 12'h45b == _T_96[11:0] ? image_1115 : _GEN_7323; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7325 = 12'h45c == _T_96[11:0] ? image_1116 : _GEN_7324; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7326 = 12'h45d == _T_96[11:0] ? image_1117 : _GEN_7325; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7327 = 12'h45e == _T_96[11:0] ? image_1118 : _GEN_7326; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7328 = 12'h45f == _T_96[11:0] ? image_1119 : _GEN_7327; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7329 = 12'h460 == _T_96[11:0] ? image_1120 : _GEN_7328; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7330 = 12'h461 == _T_96[11:0] ? image_1121 : _GEN_7329; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7331 = 12'h462 == _T_96[11:0] ? image_1122 : _GEN_7330; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7332 = 12'h463 == _T_96[11:0] ? image_1123 : _GEN_7331; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7333 = 12'h464 == _T_96[11:0] ? image_1124 : _GEN_7332; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7334 = 12'h465 == _T_96[11:0] ? image_1125 : _GEN_7333; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7335 = 12'h466 == _T_96[11:0] ? image_1126 : _GEN_7334; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7336 = 12'h467 == _T_96[11:0] ? image_1127 : _GEN_7335; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7337 = 12'h468 == _T_96[11:0] ? image_1128 : _GEN_7336; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7338 = 12'h469 == _T_96[11:0] ? image_1129 : _GEN_7337; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7339 = 12'h46a == _T_96[11:0] ? image_1130 : _GEN_7338; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7340 = 12'h46b == _T_96[11:0] ? image_1131 : _GEN_7339; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7341 = 12'h46c == _T_96[11:0] ? image_1132 : _GEN_7340; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7342 = 12'h46d == _T_96[11:0] ? image_1133 : _GEN_7341; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7343 = 12'h46e == _T_96[11:0] ? image_1134 : _GEN_7342; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7344 = 12'h46f == _T_96[11:0] ? image_1135 : _GEN_7343; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7345 = 12'h470 == _T_96[11:0] ? image_1136 : _GEN_7344; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7346 = 12'h471 == _T_96[11:0] ? image_1137 : _GEN_7345; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7347 = 12'h472 == _T_96[11:0] ? image_1138 : _GEN_7346; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7348 = 12'h473 == _T_96[11:0] ? image_1139 : _GEN_7347; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7349 = 12'h474 == _T_96[11:0] ? image_1140 : _GEN_7348; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7350 = 12'h475 == _T_96[11:0] ? image_1141 : _GEN_7349; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7351 = 12'h476 == _T_96[11:0] ? image_1142 : _GEN_7350; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7352 = 12'h477 == _T_96[11:0] ? image_1143 : _GEN_7351; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7353 = 12'h478 == _T_96[11:0] ? image_1144 : _GEN_7352; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7354 = 12'h479 == _T_96[11:0] ? image_1145 : _GEN_7353; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7355 = 12'h47a == _T_96[11:0] ? image_1146 : _GEN_7354; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7356 = 12'h47b == _T_96[11:0] ? image_1147 : _GEN_7355; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7357 = 12'h47c == _T_96[11:0] ? image_1148 : _GEN_7356; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7358 = 12'h47d == _T_96[11:0] ? 4'h0 : _GEN_7357; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7359 = 12'h47e == _T_96[11:0] ? 4'h0 : _GEN_7358; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7360 = 12'h47f == _T_96[11:0] ? 4'h0 : _GEN_7359; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7361 = 12'h480 == _T_96[11:0] ? image_1152 : _GEN_7360; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7362 = 12'h481 == _T_96[11:0] ? image_1153 : _GEN_7361; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7363 = 12'h482 == _T_96[11:0] ? image_1154 : _GEN_7362; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7364 = 12'h483 == _T_96[11:0] ? image_1155 : _GEN_7363; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7365 = 12'h484 == _T_96[11:0] ? image_1156 : _GEN_7364; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7366 = 12'h485 == _T_96[11:0] ? image_1157 : _GEN_7365; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7367 = 12'h486 == _T_96[11:0] ? image_1158 : _GEN_7366; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7368 = 12'h487 == _T_96[11:0] ? image_1159 : _GEN_7367; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7369 = 12'h488 == _T_96[11:0] ? image_1160 : _GEN_7368; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7370 = 12'h489 == _T_96[11:0] ? image_1161 : _GEN_7369; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7371 = 12'h48a == _T_96[11:0] ? image_1162 : _GEN_7370; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7372 = 12'h48b == _T_96[11:0] ? image_1163 : _GEN_7371; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7373 = 12'h48c == _T_96[11:0] ? image_1164 : _GEN_7372; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7374 = 12'h48d == _T_96[11:0] ? image_1165 : _GEN_7373; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7375 = 12'h48e == _T_96[11:0] ? image_1166 : _GEN_7374; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7376 = 12'h48f == _T_96[11:0] ? image_1167 : _GEN_7375; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7377 = 12'h490 == _T_96[11:0] ? image_1168 : _GEN_7376; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7378 = 12'h491 == _T_96[11:0] ? image_1169 : _GEN_7377; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7379 = 12'h492 == _T_96[11:0] ? image_1170 : _GEN_7378; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7380 = 12'h493 == _T_96[11:0] ? image_1171 : _GEN_7379; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7381 = 12'h494 == _T_96[11:0] ? image_1172 : _GEN_7380; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7382 = 12'h495 == _T_96[11:0] ? image_1173 : _GEN_7381; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7383 = 12'h496 == _T_96[11:0] ? image_1174 : _GEN_7382; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7384 = 12'h497 == _T_96[11:0] ? image_1175 : _GEN_7383; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7385 = 12'h498 == _T_96[11:0] ? image_1176 : _GEN_7384; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7386 = 12'h499 == _T_96[11:0] ? image_1177 : _GEN_7385; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7387 = 12'h49a == _T_96[11:0] ? image_1178 : _GEN_7386; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7388 = 12'h49b == _T_96[11:0] ? image_1179 : _GEN_7387; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7389 = 12'h49c == _T_96[11:0] ? image_1180 : _GEN_7388; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7390 = 12'h49d == _T_96[11:0] ? image_1181 : _GEN_7389; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7391 = 12'h49e == _T_96[11:0] ? image_1182 : _GEN_7390; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7392 = 12'h49f == _T_96[11:0] ? image_1183 : _GEN_7391; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7393 = 12'h4a0 == _T_96[11:0] ? image_1184 : _GEN_7392; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7394 = 12'h4a1 == _T_96[11:0] ? image_1185 : _GEN_7393; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7395 = 12'h4a2 == _T_96[11:0] ? image_1186 : _GEN_7394; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7396 = 12'h4a3 == _T_96[11:0] ? image_1187 : _GEN_7395; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7397 = 12'h4a4 == _T_96[11:0] ? image_1188 : _GEN_7396; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7398 = 12'h4a5 == _T_96[11:0] ? image_1189 : _GEN_7397; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7399 = 12'h4a6 == _T_96[11:0] ? image_1190 : _GEN_7398; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7400 = 12'h4a7 == _T_96[11:0] ? image_1191 : _GEN_7399; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7401 = 12'h4a8 == _T_96[11:0] ? image_1192 : _GEN_7400; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7402 = 12'h4a9 == _T_96[11:0] ? image_1193 : _GEN_7401; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7403 = 12'h4aa == _T_96[11:0] ? image_1194 : _GEN_7402; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7404 = 12'h4ab == _T_96[11:0] ? image_1195 : _GEN_7403; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7405 = 12'h4ac == _T_96[11:0] ? image_1196 : _GEN_7404; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7406 = 12'h4ad == _T_96[11:0] ? image_1197 : _GEN_7405; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7407 = 12'h4ae == _T_96[11:0] ? image_1198 : _GEN_7406; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7408 = 12'h4af == _T_96[11:0] ? image_1199 : _GEN_7407; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7409 = 12'h4b0 == _T_96[11:0] ? image_1200 : _GEN_7408; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7410 = 12'h4b1 == _T_96[11:0] ? image_1201 : _GEN_7409; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7411 = 12'h4b2 == _T_96[11:0] ? image_1202 : _GEN_7410; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7412 = 12'h4b3 == _T_96[11:0] ? image_1203 : _GEN_7411; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7413 = 12'h4b4 == _T_96[11:0] ? image_1204 : _GEN_7412; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7414 = 12'h4b5 == _T_96[11:0] ? image_1205 : _GEN_7413; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7415 = 12'h4b6 == _T_96[11:0] ? image_1206 : _GEN_7414; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7416 = 12'h4b7 == _T_96[11:0] ? image_1207 : _GEN_7415; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7417 = 12'h4b8 == _T_96[11:0] ? image_1208 : _GEN_7416; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7418 = 12'h4b9 == _T_96[11:0] ? 4'h0 : _GEN_7417; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7419 = 12'h4ba == _T_96[11:0] ? 4'h0 : _GEN_7418; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7420 = 12'h4bb == _T_96[11:0] ? 4'h0 : _GEN_7419; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7421 = 12'h4bc == _T_96[11:0] ? 4'h0 : _GEN_7420; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7422 = 12'h4bd == _T_96[11:0] ? 4'h0 : _GEN_7421; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7423 = 12'h4be == _T_96[11:0] ? 4'h0 : _GEN_7422; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7424 = 12'h4bf == _T_96[11:0] ? 4'h0 : _GEN_7423; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7425 = 12'h4c0 == _T_96[11:0] ? image_1216 : _GEN_7424; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7426 = 12'h4c1 == _T_96[11:0] ? image_1217 : _GEN_7425; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7427 = 12'h4c2 == _T_96[11:0] ? image_1218 : _GEN_7426; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7428 = 12'h4c3 == _T_96[11:0] ? image_1219 : _GEN_7427; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7429 = 12'h4c4 == _T_96[11:0] ? image_1220 : _GEN_7428; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7430 = 12'h4c5 == _T_96[11:0] ? image_1221 : _GEN_7429; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7431 = 12'h4c6 == _T_96[11:0] ? image_1222 : _GEN_7430; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7432 = 12'h4c7 == _T_96[11:0] ? image_1223 : _GEN_7431; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7433 = 12'h4c8 == _T_96[11:0] ? image_1224 : _GEN_7432; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7434 = 12'h4c9 == _T_96[11:0] ? image_1225 : _GEN_7433; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7435 = 12'h4ca == _T_96[11:0] ? image_1226 : _GEN_7434; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7436 = 12'h4cb == _T_96[11:0] ? image_1227 : _GEN_7435; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7437 = 12'h4cc == _T_96[11:0] ? image_1228 : _GEN_7436; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7438 = 12'h4cd == _T_96[11:0] ? image_1229 : _GEN_7437; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7439 = 12'h4ce == _T_96[11:0] ? image_1230 : _GEN_7438; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7440 = 12'h4cf == _T_96[11:0] ? image_1231 : _GEN_7439; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7441 = 12'h4d0 == _T_96[11:0] ? image_1232 : _GEN_7440; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7442 = 12'h4d1 == _T_96[11:0] ? image_1233 : _GEN_7441; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7443 = 12'h4d2 == _T_96[11:0] ? image_1234 : _GEN_7442; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7444 = 12'h4d3 == _T_96[11:0] ? image_1235 : _GEN_7443; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7445 = 12'h4d4 == _T_96[11:0] ? image_1236 : _GEN_7444; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7446 = 12'h4d5 == _T_96[11:0] ? image_1237 : _GEN_7445; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7447 = 12'h4d6 == _T_96[11:0] ? image_1238 : _GEN_7446; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7448 = 12'h4d7 == _T_96[11:0] ? image_1239 : _GEN_7447; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7449 = 12'h4d8 == _T_96[11:0] ? image_1240 : _GEN_7448; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7450 = 12'h4d9 == _T_96[11:0] ? image_1241 : _GEN_7449; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7451 = 12'h4da == _T_96[11:0] ? image_1242 : _GEN_7450; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7452 = 12'h4db == _T_96[11:0] ? image_1243 : _GEN_7451; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7453 = 12'h4dc == _T_96[11:0] ? image_1244 : _GEN_7452; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7454 = 12'h4dd == _T_96[11:0] ? image_1245 : _GEN_7453; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7455 = 12'h4de == _T_96[11:0] ? image_1246 : _GEN_7454; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7456 = 12'h4df == _T_96[11:0] ? image_1247 : _GEN_7455; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7457 = 12'h4e0 == _T_96[11:0] ? image_1248 : _GEN_7456; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7458 = 12'h4e1 == _T_96[11:0] ? image_1249 : _GEN_7457; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7459 = 12'h4e2 == _T_96[11:0] ? image_1250 : _GEN_7458; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7460 = 12'h4e3 == _T_96[11:0] ? image_1251 : _GEN_7459; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7461 = 12'h4e4 == _T_96[11:0] ? image_1252 : _GEN_7460; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7462 = 12'h4e5 == _T_96[11:0] ? image_1253 : _GEN_7461; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7463 = 12'h4e6 == _T_96[11:0] ? image_1254 : _GEN_7462; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7464 = 12'h4e7 == _T_96[11:0] ? image_1255 : _GEN_7463; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7465 = 12'h4e8 == _T_96[11:0] ? image_1256 : _GEN_7464; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7466 = 12'h4e9 == _T_96[11:0] ? image_1257 : _GEN_7465; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7467 = 12'h4ea == _T_96[11:0] ? image_1258 : _GEN_7466; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7468 = 12'h4eb == _T_96[11:0] ? image_1259 : _GEN_7467; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7469 = 12'h4ec == _T_96[11:0] ? image_1260 : _GEN_7468; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7470 = 12'h4ed == _T_96[11:0] ? image_1261 : _GEN_7469; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7471 = 12'h4ee == _T_96[11:0] ? image_1262 : _GEN_7470; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7472 = 12'h4ef == _T_96[11:0] ? image_1263 : _GEN_7471; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7473 = 12'h4f0 == _T_96[11:0] ? image_1264 : _GEN_7472; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7474 = 12'h4f1 == _T_96[11:0] ? image_1265 : _GEN_7473; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7475 = 12'h4f2 == _T_96[11:0] ? image_1266 : _GEN_7474; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7476 = 12'h4f3 == _T_96[11:0] ? image_1267 : _GEN_7475; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7477 = 12'h4f4 == _T_96[11:0] ? image_1268 : _GEN_7476; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7478 = 12'h4f5 == _T_96[11:0] ? image_1269 : _GEN_7477; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7479 = 12'h4f6 == _T_96[11:0] ? image_1270 : _GEN_7478; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7480 = 12'h4f7 == _T_96[11:0] ? image_1271 : _GEN_7479; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7481 = 12'h4f8 == _T_96[11:0] ? image_1272 : _GEN_7480; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7482 = 12'h4f9 == _T_96[11:0] ? image_1273 : _GEN_7481; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7483 = 12'h4fa == _T_96[11:0] ? image_1274 : _GEN_7482; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7484 = 12'h4fb == _T_96[11:0] ? image_1275 : _GEN_7483; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7485 = 12'h4fc == _T_96[11:0] ? 4'h0 : _GEN_7484; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7486 = 12'h4fd == _T_96[11:0] ? 4'h0 : _GEN_7485; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7487 = 12'h4fe == _T_96[11:0] ? 4'h0 : _GEN_7486; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7488 = 12'h4ff == _T_96[11:0] ? 4'h0 : _GEN_7487; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7489 = 12'h500 == _T_96[11:0] ? image_1280 : _GEN_7488; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7490 = 12'h501 == _T_96[11:0] ? image_1281 : _GEN_7489; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7491 = 12'h502 == _T_96[11:0] ? image_1282 : _GEN_7490; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7492 = 12'h503 == _T_96[11:0] ? image_1283 : _GEN_7491; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7493 = 12'h504 == _T_96[11:0] ? image_1284 : _GEN_7492; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7494 = 12'h505 == _T_96[11:0] ? image_1285 : _GEN_7493; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7495 = 12'h506 == _T_96[11:0] ? image_1286 : _GEN_7494; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7496 = 12'h507 == _T_96[11:0] ? image_1287 : _GEN_7495; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7497 = 12'h508 == _T_96[11:0] ? image_1288 : _GEN_7496; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7498 = 12'h509 == _T_96[11:0] ? image_1289 : _GEN_7497; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7499 = 12'h50a == _T_96[11:0] ? image_1290 : _GEN_7498; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7500 = 12'h50b == _T_96[11:0] ? image_1291 : _GEN_7499; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7501 = 12'h50c == _T_96[11:0] ? image_1292 : _GEN_7500; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7502 = 12'h50d == _T_96[11:0] ? image_1293 : _GEN_7501; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7503 = 12'h50e == _T_96[11:0] ? image_1294 : _GEN_7502; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7504 = 12'h50f == _T_96[11:0] ? image_1295 : _GEN_7503; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7505 = 12'h510 == _T_96[11:0] ? image_1296 : _GEN_7504; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7506 = 12'h511 == _T_96[11:0] ? image_1297 : _GEN_7505; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7507 = 12'h512 == _T_96[11:0] ? image_1298 : _GEN_7506; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7508 = 12'h513 == _T_96[11:0] ? image_1299 : _GEN_7507; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7509 = 12'h514 == _T_96[11:0] ? image_1300 : _GEN_7508; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7510 = 12'h515 == _T_96[11:0] ? image_1301 : _GEN_7509; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7511 = 12'h516 == _T_96[11:0] ? image_1302 : _GEN_7510; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7512 = 12'h517 == _T_96[11:0] ? image_1303 : _GEN_7511; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7513 = 12'h518 == _T_96[11:0] ? image_1304 : _GEN_7512; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7514 = 12'h519 == _T_96[11:0] ? image_1305 : _GEN_7513; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7515 = 12'h51a == _T_96[11:0] ? image_1306 : _GEN_7514; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7516 = 12'h51b == _T_96[11:0] ? image_1307 : _GEN_7515; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7517 = 12'h51c == _T_96[11:0] ? image_1308 : _GEN_7516; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7518 = 12'h51d == _T_96[11:0] ? image_1309 : _GEN_7517; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7519 = 12'h51e == _T_96[11:0] ? image_1310 : _GEN_7518; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7520 = 12'h51f == _T_96[11:0] ? image_1311 : _GEN_7519; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7521 = 12'h520 == _T_96[11:0] ? image_1312 : _GEN_7520; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7522 = 12'h521 == _T_96[11:0] ? image_1313 : _GEN_7521; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7523 = 12'h522 == _T_96[11:0] ? image_1314 : _GEN_7522; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7524 = 12'h523 == _T_96[11:0] ? image_1315 : _GEN_7523; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7525 = 12'h524 == _T_96[11:0] ? image_1316 : _GEN_7524; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7526 = 12'h525 == _T_96[11:0] ? image_1317 : _GEN_7525; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7527 = 12'h526 == _T_96[11:0] ? image_1318 : _GEN_7526; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7528 = 12'h527 == _T_96[11:0] ? image_1319 : _GEN_7527; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7529 = 12'h528 == _T_96[11:0] ? image_1320 : _GEN_7528; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7530 = 12'h529 == _T_96[11:0] ? image_1321 : _GEN_7529; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7531 = 12'h52a == _T_96[11:0] ? image_1322 : _GEN_7530; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7532 = 12'h52b == _T_96[11:0] ? image_1323 : _GEN_7531; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7533 = 12'h52c == _T_96[11:0] ? image_1324 : _GEN_7532; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7534 = 12'h52d == _T_96[11:0] ? image_1325 : _GEN_7533; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7535 = 12'h52e == _T_96[11:0] ? image_1326 : _GEN_7534; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7536 = 12'h52f == _T_96[11:0] ? image_1327 : _GEN_7535; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7537 = 12'h530 == _T_96[11:0] ? image_1328 : _GEN_7536; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7538 = 12'h531 == _T_96[11:0] ? image_1329 : _GEN_7537; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7539 = 12'h532 == _T_96[11:0] ? image_1330 : _GEN_7538; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7540 = 12'h533 == _T_96[11:0] ? image_1331 : _GEN_7539; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7541 = 12'h534 == _T_96[11:0] ? image_1332 : _GEN_7540; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7542 = 12'h535 == _T_96[11:0] ? image_1333 : _GEN_7541; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7543 = 12'h536 == _T_96[11:0] ? image_1334 : _GEN_7542; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7544 = 12'h537 == _T_96[11:0] ? image_1335 : _GEN_7543; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7545 = 12'h538 == _T_96[11:0] ? image_1336 : _GEN_7544; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7546 = 12'h539 == _T_96[11:0] ? image_1337 : _GEN_7545; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7547 = 12'h53a == _T_96[11:0] ? image_1338 : _GEN_7546; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7548 = 12'h53b == _T_96[11:0] ? image_1339 : _GEN_7547; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7549 = 12'h53c == _T_96[11:0] ? image_1340 : _GEN_7548; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7550 = 12'h53d == _T_96[11:0] ? image_1341 : _GEN_7549; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7551 = 12'h53e == _T_96[11:0] ? 4'h0 : _GEN_7550; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7552 = 12'h53f == _T_96[11:0] ? 4'h0 : _GEN_7551; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7553 = 12'h540 == _T_96[11:0] ? image_1344 : _GEN_7552; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7554 = 12'h541 == _T_96[11:0] ? image_1345 : _GEN_7553; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7555 = 12'h542 == _T_96[11:0] ? image_1346 : _GEN_7554; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7556 = 12'h543 == _T_96[11:0] ? image_1347 : _GEN_7555; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7557 = 12'h544 == _T_96[11:0] ? image_1348 : _GEN_7556; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7558 = 12'h545 == _T_96[11:0] ? image_1349 : _GEN_7557; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7559 = 12'h546 == _T_96[11:0] ? image_1350 : _GEN_7558; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7560 = 12'h547 == _T_96[11:0] ? image_1351 : _GEN_7559; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7561 = 12'h548 == _T_96[11:0] ? image_1352 : _GEN_7560; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7562 = 12'h549 == _T_96[11:0] ? image_1353 : _GEN_7561; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7563 = 12'h54a == _T_96[11:0] ? image_1354 : _GEN_7562; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7564 = 12'h54b == _T_96[11:0] ? image_1355 : _GEN_7563; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7565 = 12'h54c == _T_96[11:0] ? image_1356 : _GEN_7564; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7566 = 12'h54d == _T_96[11:0] ? image_1357 : _GEN_7565; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7567 = 12'h54e == _T_96[11:0] ? image_1358 : _GEN_7566; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7568 = 12'h54f == _T_96[11:0] ? image_1359 : _GEN_7567; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7569 = 12'h550 == _T_96[11:0] ? image_1360 : _GEN_7568; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7570 = 12'h551 == _T_96[11:0] ? image_1361 : _GEN_7569; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7571 = 12'h552 == _T_96[11:0] ? image_1362 : _GEN_7570; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7572 = 12'h553 == _T_96[11:0] ? image_1363 : _GEN_7571; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7573 = 12'h554 == _T_96[11:0] ? image_1364 : _GEN_7572; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7574 = 12'h555 == _T_96[11:0] ? image_1365 : _GEN_7573; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7575 = 12'h556 == _T_96[11:0] ? image_1366 : _GEN_7574; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7576 = 12'h557 == _T_96[11:0] ? image_1367 : _GEN_7575; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7577 = 12'h558 == _T_96[11:0] ? image_1368 : _GEN_7576; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7578 = 12'h559 == _T_96[11:0] ? image_1369 : _GEN_7577; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7579 = 12'h55a == _T_96[11:0] ? image_1370 : _GEN_7578; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7580 = 12'h55b == _T_96[11:0] ? image_1371 : _GEN_7579; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7581 = 12'h55c == _T_96[11:0] ? image_1372 : _GEN_7580; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7582 = 12'h55d == _T_96[11:0] ? image_1373 : _GEN_7581; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7583 = 12'h55e == _T_96[11:0] ? image_1374 : _GEN_7582; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7584 = 12'h55f == _T_96[11:0] ? image_1375 : _GEN_7583; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7585 = 12'h560 == _T_96[11:0] ? image_1376 : _GEN_7584; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7586 = 12'h561 == _T_96[11:0] ? image_1377 : _GEN_7585; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7587 = 12'h562 == _T_96[11:0] ? image_1378 : _GEN_7586; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7588 = 12'h563 == _T_96[11:0] ? image_1379 : _GEN_7587; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7589 = 12'h564 == _T_96[11:0] ? image_1380 : _GEN_7588; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7590 = 12'h565 == _T_96[11:0] ? image_1381 : _GEN_7589; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7591 = 12'h566 == _T_96[11:0] ? image_1382 : _GEN_7590; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7592 = 12'h567 == _T_96[11:0] ? image_1383 : _GEN_7591; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7593 = 12'h568 == _T_96[11:0] ? image_1384 : _GEN_7592; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7594 = 12'h569 == _T_96[11:0] ? image_1385 : _GEN_7593; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7595 = 12'h56a == _T_96[11:0] ? image_1386 : _GEN_7594; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7596 = 12'h56b == _T_96[11:0] ? image_1387 : _GEN_7595; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7597 = 12'h56c == _T_96[11:0] ? image_1388 : _GEN_7596; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7598 = 12'h56d == _T_96[11:0] ? image_1389 : _GEN_7597; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7599 = 12'h56e == _T_96[11:0] ? image_1390 : _GEN_7598; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7600 = 12'h56f == _T_96[11:0] ? image_1391 : _GEN_7599; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7601 = 12'h570 == _T_96[11:0] ? image_1392 : _GEN_7600; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7602 = 12'h571 == _T_96[11:0] ? image_1393 : _GEN_7601; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7603 = 12'h572 == _T_96[11:0] ? image_1394 : _GEN_7602; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7604 = 12'h573 == _T_96[11:0] ? image_1395 : _GEN_7603; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7605 = 12'h574 == _T_96[11:0] ? image_1396 : _GEN_7604; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7606 = 12'h575 == _T_96[11:0] ? image_1397 : _GEN_7605; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7607 = 12'h576 == _T_96[11:0] ? image_1398 : _GEN_7606; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7608 = 12'h577 == _T_96[11:0] ? image_1399 : _GEN_7607; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7609 = 12'h578 == _T_96[11:0] ? image_1400 : _GEN_7608; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7610 = 12'h579 == _T_96[11:0] ? image_1401 : _GEN_7609; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7611 = 12'h57a == _T_96[11:0] ? image_1402 : _GEN_7610; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7612 = 12'h57b == _T_96[11:0] ? image_1403 : _GEN_7611; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7613 = 12'h57c == _T_96[11:0] ? image_1404 : _GEN_7612; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7614 = 12'h57d == _T_96[11:0] ? image_1405 : _GEN_7613; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7615 = 12'h57e == _T_96[11:0] ? 4'h0 : _GEN_7614; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7616 = 12'h57f == _T_96[11:0] ? 4'h0 : _GEN_7615; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7617 = 12'h580 == _T_96[11:0] ? image_1408 : _GEN_7616; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7618 = 12'h581 == _T_96[11:0] ? image_1409 : _GEN_7617; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7619 = 12'h582 == _T_96[11:0] ? image_1410 : _GEN_7618; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7620 = 12'h583 == _T_96[11:0] ? image_1411 : _GEN_7619; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7621 = 12'h584 == _T_96[11:0] ? image_1412 : _GEN_7620; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7622 = 12'h585 == _T_96[11:0] ? image_1413 : _GEN_7621; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7623 = 12'h586 == _T_96[11:0] ? image_1414 : _GEN_7622; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7624 = 12'h587 == _T_96[11:0] ? image_1415 : _GEN_7623; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7625 = 12'h588 == _T_96[11:0] ? image_1416 : _GEN_7624; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7626 = 12'h589 == _T_96[11:0] ? image_1417 : _GEN_7625; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7627 = 12'h58a == _T_96[11:0] ? image_1418 : _GEN_7626; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7628 = 12'h58b == _T_96[11:0] ? image_1419 : _GEN_7627; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7629 = 12'h58c == _T_96[11:0] ? image_1420 : _GEN_7628; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7630 = 12'h58d == _T_96[11:0] ? image_1421 : _GEN_7629; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7631 = 12'h58e == _T_96[11:0] ? image_1422 : _GEN_7630; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7632 = 12'h58f == _T_96[11:0] ? image_1423 : _GEN_7631; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7633 = 12'h590 == _T_96[11:0] ? image_1424 : _GEN_7632; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7634 = 12'h591 == _T_96[11:0] ? image_1425 : _GEN_7633; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7635 = 12'h592 == _T_96[11:0] ? image_1426 : _GEN_7634; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7636 = 12'h593 == _T_96[11:0] ? image_1427 : _GEN_7635; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7637 = 12'h594 == _T_96[11:0] ? image_1428 : _GEN_7636; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7638 = 12'h595 == _T_96[11:0] ? image_1429 : _GEN_7637; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7639 = 12'h596 == _T_96[11:0] ? image_1430 : _GEN_7638; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7640 = 12'h597 == _T_96[11:0] ? image_1431 : _GEN_7639; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7641 = 12'h598 == _T_96[11:0] ? image_1432 : _GEN_7640; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7642 = 12'h599 == _T_96[11:0] ? image_1433 : _GEN_7641; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7643 = 12'h59a == _T_96[11:0] ? image_1434 : _GEN_7642; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7644 = 12'h59b == _T_96[11:0] ? image_1435 : _GEN_7643; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7645 = 12'h59c == _T_96[11:0] ? image_1436 : _GEN_7644; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7646 = 12'h59d == _T_96[11:0] ? image_1437 : _GEN_7645; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7647 = 12'h59e == _T_96[11:0] ? image_1438 : _GEN_7646; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7648 = 12'h59f == _T_96[11:0] ? image_1439 : _GEN_7647; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7649 = 12'h5a0 == _T_96[11:0] ? image_1440 : _GEN_7648; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7650 = 12'h5a1 == _T_96[11:0] ? image_1441 : _GEN_7649; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7651 = 12'h5a2 == _T_96[11:0] ? image_1442 : _GEN_7650; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7652 = 12'h5a3 == _T_96[11:0] ? image_1443 : _GEN_7651; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7653 = 12'h5a4 == _T_96[11:0] ? image_1444 : _GEN_7652; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7654 = 12'h5a5 == _T_96[11:0] ? image_1445 : _GEN_7653; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7655 = 12'h5a6 == _T_96[11:0] ? image_1446 : _GEN_7654; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7656 = 12'h5a7 == _T_96[11:0] ? image_1447 : _GEN_7655; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7657 = 12'h5a8 == _T_96[11:0] ? image_1448 : _GEN_7656; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7658 = 12'h5a9 == _T_96[11:0] ? image_1449 : _GEN_7657; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7659 = 12'h5aa == _T_96[11:0] ? image_1450 : _GEN_7658; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7660 = 12'h5ab == _T_96[11:0] ? image_1451 : _GEN_7659; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7661 = 12'h5ac == _T_96[11:0] ? image_1452 : _GEN_7660; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7662 = 12'h5ad == _T_96[11:0] ? image_1453 : _GEN_7661; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7663 = 12'h5ae == _T_96[11:0] ? image_1454 : _GEN_7662; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7664 = 12'h5af == _T_96[11:0] ? image_1455 : _GEN_7663; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7665 = 12'h5b0 == _T_96[11:0] ? image_1456 : _GEN_7664; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7666 = 12'h5b1 == _T_96[11:0] ? image_1457 : _GEN_7665; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7667 = 12'h5b2 == _T_96[11:0] ? image_1458 : _GEN_7666; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7668 = 12'h5b3 == _T_96[11:0] ? image_1459 : _GEN_7667; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7669 = 12'h5b4 == _T_96[11:0] ? image_1460 : _GEN_7668; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7670 = 12'h5b5 == _T_96[11:0] ? image_1461 : _GEN_7669; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7671 = 12'h5b6 == _T_96[11:0] ? image_1462 : _GEN_7670; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7672 = 12'h5b7 == _T_96[11:0] ? image_1463 : _GEN_7671; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7673 = 12'h5b8 == _T_96[11:0] ? image_1464 : _GEN_7672; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7674 = 12'h5b9 == _T_96[11:0] ? image_1465 : _GEN_7673; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7675 = 12'h5ba == _T_96[11:0] ? image_1466 : _GEN_7674; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7676 = 12'h5bb == _T_96[11:0] ? image_1467 : _GEN_7675; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7677 = 12'h5bc == _T_96[11:0] ? image_1468 : _GEN_7676; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7678 = 12'h5bd == _T_96[11:0] ? image_1469 : _GEN_7677; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7679 = 12'h5be == _T_96[11:0] ? 4'h0 : _GEN_7678; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7680 = 12'h5bf == _T_96[11:0] ? 4'h0 : _GEN_7679; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7681 = 12'h5c0 == _T_96[11:0] ? image_1472 : _GEN_7680; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7682 = 12'h5c1 == _T_96[11:0] ? image_1473 : _GEN_7681; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7683 = 12'h5c2 == _T_96[11:0] ? image_1474 : _GEN_7682; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7684 = 12'h5c3 == _T_96[11:0] ? image_1475 : _GEN_7683; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7685 = 12'h5c4 == _T_96[11:0] ? image_1476 : _GEN_7684; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7686 = 12'h5c5 == _T_96[11:0] ? image_1477 : _GEN_7685; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7687 = 12'h5c6 == _T_96[11:0] ? image_1478 : _GEN_7686; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7688 = 12'h5c7 == _T_96[11:0] ? image_1479 : _GEN_7687; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7689 = 12'h5c8 == _T_96[11:0] ? image_1480 : _GEN_7688; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7690 = 12'h5c9 == _T_96[11:0] ? image_1481 : _GEN_7689; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7691 = 12'h5ca == _T_96[11:0] ? image_1482 : _GEN_7690; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7692 = 12'h5cb == _T_96[11:0] ? image_1483 : _GEN_7691; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7693 = 12'h5cc == _T_96[11:0] ? image_1484 : _GEN_7692; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7694 = 12'h5cd == _T_96[11:0] ? image_1485 : _GEN_7693; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7695 = 12'h5ce == _T_96[11:0] ? image_1486 : _GEN_7694; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7696 = 12'h5cf == _T_96[11:0] ? image_1487 : _GEN_7695; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7697 = 12'h5d0 == _T_96[11:0] ? image_1488 : _GEN_7696; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7698 = 12'h5d1 == _T_96[11:0] ? image_1489 : _GEN_7697; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7699 = 12'h5d2 == _T_96[11:0] ? image_1490 : _GEN_7698; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7700 = 12'h5d3 == _T_96[11:0] ? image_1491 : _GEN_7699; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7701 = 12'h5d4 == _T_96[11:0] ? image_1492 : _GEN_7700; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7702 = 12'h5d5 == _T_96[11:0] ? image_1493 : _GEN_7701; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7703 = 12'h5d6 == _T_96[11:0] ? image_1494 : _GEN_7702; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7704 = 12'h5d7 == _T_96[11:0] ? image_1495 : _GEN_7703; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7705 = 12'h5d8 == _T_96[11:0] ? image_1496 : _GEN_7704; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7706 = 12'h5d9 == _T_96[11:0] ? image_1497 : _GEN_7705; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7707 = 12'h5da == _T_96[11:0] ? image_1498 : _GEN_7706; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7708 = 12'h5db == _T_96[11:0] ? image_1499 : _GEN_7707; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7709 = 12'h5dc == _T_96[11:0] ? image_1500 : _GEN_7708; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7710 = 12'h5dd == _T_96[11:0] ? image_1501 : _GEN_7709; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7711 = 12'h5de == _T_96[11:0] ? image_1502 : _GEN_7710; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7712 = 12'h5df == _T_96[11:0] ? image_1503 : _GEN_7711; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7713 = 12'h5e0 == _T_96[11:0] ? image_1504 : _GEN_7712; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7714 = 12'h5e1 == _T_96[11:0] ? image_1505 : _GEN_7713; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7715 = 12'h5e2 == _T_96[11:0] ? image_1506 : _GEN_7714; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7716 = 12'h5e3 == _T_96[11:0] ? image_1507 : _GEN_7715; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7717 = 12'h5e4 == _T_96[11:0] ? image_1508 : _GEN_7716; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7718 = 12'h5e5 == _T_96[11:0] ? image_1509 : _GEN_7717; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7719 = 12'h5e6 == _T_96[11:0] ? image_1510 : _GEN_7718; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7720 = 12'h5e7 == _T_96[11:0] ? image_1511 : _GEN_7719; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7721 = 12'h5e8 == _T_96[11:0] ? image_1512 : _GEN_7720; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7722 = 12'h5e9 == _T_96[11:0] ? image_1513 : _GEN_7721; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7723 = 12'h5ea == _T_96[11:0] ? image_1514 : _GEN_7722; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7724 = 12'h5eb == _T_96[11:0] ? image_1515 : _GEN_7723; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7725 = 12'h5ec == _T_96[11:0] ? image_1516 : _GEN_7724; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7726 = 12'h5ed == _T_96[11:0] ? image_1517 : _GEN_7725; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7727 = 12'h5ee == _T_96[11:0] ? image_1518 : _GEN_7726; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7728 = 12'h5ef == _T_96[11:0] ? image_1519 : _GEN_7727; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7729 = 12'h5f0 == _T_96[11:0] ? image_1520 : _GEN_7728; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7730 = 12'h5f1 == _T_96[11:0] ? image_1521 : _GEN_7729; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7731 = 12'h5f2 == _T_96[11:0] ? image_1522 : _GEN_7730; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7732 = 12'h5f3 == _T_96[11:0] ? image_1523 : _GEN_7731; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7733 = 12'h5f4 == _T_96[11:0] ? image_1524 : _GEN_7732; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7734 = 12'h5f5 == _T_96[11:0] ? image_1525 : _GEN_7733; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7735 = 12'h5f6 == _T_96[11:0] ? image_1526 : _GEN_7734; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7736 = 12'h5f7 == _T_96[11:0] ? image_1527 : _GEN_7735; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7737 = 12'h5f8 == _T_96[11:0] ? image_1528 : _GEN_7736; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7738 = 12'h5f9 == _T_96[11:0] ? image_1529 : _GEN_7737; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7739 = 12'h5fa == _T_96[11:0] ? image_1530 : _GEN_7738; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7740 = 12'h5fb == _T_96[11:0] ? image_1531 : _GEN_7739; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7741 = 12'h5fc == _T_96[11:0] ? image_1532 : _GEN_7740; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7742 = 12'h5fd == _T_96[11:0] ? image_1533 : _GEN_7741; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7743 = 12'h5fe == _T_96[11:0] ? 4'h0 : _GEN_7742; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7744 = 12'h5ff == _T_96[11:0] ? 4'h0 : _GEN_7743; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7745 = 12'h600 == _T_96[11:0] ? image_1536 : _GEN_7744; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7746 = 12'h601 == _T_96[11:0] ? image_1537 : _GEN_7745; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7747 = 12'h602 == _T_96[11:0] ? image_1538 : _GEN_7746; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7748 = 12'h603 == _T_96[11:0] ? image_1539 : _GEN_7747; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7749 = 12'h604 == _T_96[11:0] ? image_1540 : _GEN_7748; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7750 = 12'h605 == _T_96[11:0] ? image_1541 : _GEN_7749; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7751 = 12'h606 == _T_96[11:0] ? image_1542 : _GEN_7750; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7752 = 12'h607 == _T_96[11:0] ? image_1543 : _GEN_7751; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7753 = 12'h608 == _T_96[11:0] ? image_1544 : _GEN_7752; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7754 = 12'h609 == _T_96[11:0] ? image_1545 : _GEN_7753; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7755 = 12'h60a == _T_96[11:0] ? image_1546 : _GEN_7754; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7756 = 12'h60b == _T_96[11:0] ? image_1547 : _GEN_7755; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7757 = 12'h60c == _T_96[11:0] ? image_1548 : _GEN_7756; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7758 = 12'h60d == _T_96[11:0] ? image_1549 : _GEN_7757; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7759 = 12'h60e == _T_96[11:0] ? image_1550 : _GEN_7758; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7760 = 12'h60f == _T_96[11:0] ? image_1551 : _GEN_7759; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7761 = 12'h610 == _T_96[11:0] ? image_1552 : _GEN_7760; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7762 = 12'h611 == _T_96[11:0] ? image_1553 : _GEN_7761; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7763 = 12'h612 == _T_96[11:0] ? image_1554 : _GEN_7762; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7764 = 12'h613 == _T_96[11:0] ? image_1555 : _GEN_7763; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7765 = 12'h614 == _T_96[11:0] ? image_1556 : _GEN_7764; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7766 = 12'h615 == _T_96[11:0] ? image_1557 : _GEN_7765; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7767 = 12'h616 == _T_96[11:0] ? image_1558 : _GEN_7766; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7768 = 12'h617 == _T_96[11:0] ? image_1559 : _GEN_7767; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7769 = 12'h618 == _T_96[11:0] ? image_1560 : _GEN_7768; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7770 = 12'h619 == _T_96[11:0] ? image_1561 : _GEN_7769; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7771 = 12'h61a == _T_96[11:0] ? image_1562 : _GEN_7770; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7772 = 12'h61b == _T_96[11:0] ? image_1563 : _GEN_7771; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7773 = 12'h61c == _T_96[11:0] ? image_1564 : _GEN_7772; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7774 = 12'h61d == _T_96[11:0] ? image_1565 : _GEN_7773; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7775 = 12'h61e == _T_96[11:0] ? image_1566 : _GEN_7774; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7776 = 12'h61f == _T_96[11:0] ? image_1567 : _GEN_7775; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7777 = 12'h620 == _T_96[11:0] ? image_1568 : _GEN_7776; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7778 = 12'h621 == _T_96[11:0] ? image_1569 : _GEN_7777; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7779 = 12'h622 == _T_96[11:0] ? image_1570 : _GEN_7778; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7780 = 12'h623 == _T_96[11:0] ? image_1571 : _GEN_7779; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7781 = 12'h624 == _T_96[11:0] ? image_1572 : _GEN_7780; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7782 = 12'h625 == _T_96[11:0] ? image_1573 : _GEN_7781; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7783 = 12'h626 == _T_96[11:0] ? image_1574 : _GEN_7782; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7784 = 12'h627 == _T_96[11:0] ? image_1575 : _GEN_7783; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7785 = 12'h628 == _T_96[11:0] ? image_1576 : _GEN_7784; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7786 = 12'h629 == _T_96[11:0] ? image_1577 : _GEN_7785; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7787 = 12'h62a == _T_96[11:0] ? image_1578 : _GEN_7786; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7788 = 12'h62b == _T_96[11:0] ? image_1579 : _GEN_7787; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7789 = 12'h62c == _T_96[11:0] ? image_1580 : _GEN_7788; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7790 = 12'h62d == _T_96[11:0] ? image_1581 : _GEN_7789; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7791 = 12'h62e == _T_96[11:0] ? image_1582 : _GEN_7790; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7792 = 12'h62f == _T_96[11:0] ? image_1583 : _GEN_7791; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7793 = 12'h630 == _T_96[11:0] ? image_1584 : _GEN_7792; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7794 = 12'h631 == _T_96[11:0] ? image_1585 : _GEN_7793; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7795 = 12'h632 == _T_96[11:0] ? image_1586 : _GEN_7794; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7796 = 12'h633 == _T_96[11:0] ? image_1587 : _GEN_7795; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7797 = 12'h634 == _T_96[11:0] ? image_1588 : _GEN_7796; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7798 = 12'h635 == _T_96[11:0] ? image_1589 : _GEN_7797; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7799 = 12'h636 == _T_96[11:0] ? image_1590 : _GEN_7798; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7800 = 12'h637 == _T_96[11:0] ? image_1591 : _GEN_7799; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7801 = 12'h638 == _T_96[11:0] ? image_1592 : _GEN_7800; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7802 = 12'h639 == _T_96[11:0] ? image_1593 : _GEN_7801; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7803 = 12'h63a == _T_96[11:0] ? image_1594 : _GEN_7802; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7804 = 12'h63b == _T_96[11:0] ? image_1595 : _GEN_7803; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7805 = 12'h63c == _T_96[11:0] ? image_1596 : _GEN_7804; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7806 = 12'h63d == _T_96[11:0] ? image_1597 : _GEN_7805; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7807 = 12'h63e == _T_96[11:0] ? 4'h0 : _GEN_7806; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7808 = 12'h63f == _T_96[11:0] ? 4'h0 : _GEN_7807; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7809 = 12'h640 == _T_96[11:0] ? image_1600 : _GEN_7808; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7810 = 12'h641 == _T_96[11:0] ? image_1601 : _GEN_7809; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7811 = 12'h642 == _T_96[11:0] ? image_1602 : _GEN_7810; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7812 = 12'h643 == _T_96[11:0] ? image_1603 : _GEN_7811; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7813 = 12'h644 == _T_96[11:0] ? image_1604 : _GEN_7812; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7814 = 12'h645 == _T_96[11:0] ? image_1605 : _GEN_7813; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7815 = 12'h646 == _T_96[11:0] ? image_1606 : _GEN_7814; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7816 = 12'h647 == _T_96[11:0] ? image_1607 : _GEN_7815; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7817 = 12'h648 == _T_96[11:0] ? image_1608 : _GEN_7816; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7818 = 12'h649 == _T_96[11:0] ? image_1609 : _GEN_7817; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7819 = 12'h64a == _T_96[11:0] ? image_1610 : _GEN_7818; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7820 = 12'h64b == _T_96[11:0] ? image_1611 : _GEN_7819; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7821 = 12'h64c == _T_96[11:0] ? image_1612 : _GEN_7820; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7822 = 12'h64d == _T_96[11:0] ? image_1613 : _GEN_7821; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7823 = 12'h64e == _T_96[11:0] ? image_1614 : _GEN_7822; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7824 = 12'h64f == _T_96[11:0] ? image_1615 : _GEN_7823; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7825 = 12'h650 == _T_96[11:0] ? image_1616 : _GEN_7824; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7826 = 12'h651 == _T_96[11:0] ? image_1617 : _GEN_7825; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7827 = 12'h652 == _T_96[11:0] ? image_1618 : _GEN_7826; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7828 = 12'h653 == _T_96[11:0] ? image_1619 : _GEN_7827; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7829 = 12'h654 == _T_96[11:0] ? image_1620 : _GEN_7828; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7830 = 12'h655 == _T_96[11:0] ? image_1621 : _GEN_7829; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7831 = 12'h656 == _T_96[11:0] ? image_1622 : _GEN_7830; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7832 = 12'h657 == _T_96[11:0] ? image_1623 : _GEN_7831; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7833 = 12'h658 == _T_96[11:0] ? image_1624 : _GEN_7832; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7834 = 12'h659 == _T_96[11:0] ? image_1625 : _GEN_7833; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7835 = 12'h65a == _T_96[11:0] ? image_1626 : _GEN_7834; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7836 = 12'h65b == _T_96[11:0] ? image_1627 : _GEN_7835; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7837 = 12'h65c == _T_96[11:0] ? image_1628 : _GEN_7836; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7838 = 12'h65d == _T_96[11:0] ? image_1629 : _GEN_7837; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7839 = 12'h65e == _T_96[11:0] ? image_1630 : _GEN_7838; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7840 = 12'h65f == _T_96[11:0] ? image_1631 : _GEN_7839; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7841 = 12'h660 == _T_96[11:0] ? image_1632 : _GEN_7840; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7842 = 12'h661 == _T_96[11:0] ? image_1633 : _GEN_7841; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7843 = 12'h662 == _T_96[11:0] ? image_1634 : _GEN_7842; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7844 = 12'h663 == _T_96[11:0] ? image_1635 : _GEN_7843; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7845 = 12'h664 == _T_96[11:0] ? image_1636 : _GEN_7844; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7846 = 12'h665 == _T_96[11:0] ? image_1637 : _GEN_7845; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7847 = 12'h666 == _T_96[11:0] ? image_1638 : _GEN_7846; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7848 = 12'h667 == _T_96[11:0] ? image_1639 : _GEN_7847; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7849 = 12'h668 == _T_96[11:0] ? image_1640 : _GEN_7848; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7850 = 12'h669 == _T_96[11:0] ? image_1641 : _GEN_7849; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7851 = 12'h66a == _T_96[11:0] ? image_1642 : _GEN_7850; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7852 = 12'h66b == _T_96[11:0] ? image_1643 : _GEN_7851; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7853 = 12'h66c == _T_96[11:0] ? image_1644 : _GEN_7852; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7854 = 12'h66d == _T_96[11:0] ? image_1645 : _GEN_7853; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7855 = 12'h66e == _T_96[11:0] ? image_1646 : _GEN_7854; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7856 = 12'h66f == _T_96[11:0] ? image_1647 : _GEN_7855; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7857 = 12'h670 == _T_96[11:0] ? image_1648 : _GEN_7856; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7858 = 12'h671 == _T_96[11:0] ? image_1649 : _GEN_7857; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7859 = 12'h672 == _T_96[11:0] ? image_1650 : _GEN_7858; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7860 = 12'h673 == _T_96[11:0] ? image_1651 : _GEN_7859; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7861 = 12'h674 == _T_96[11:0] ? image_1652 : _GEN_7860; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7862 = 12'h675 == _T_96[11:0] ? image_1653 : _GEN_7861; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7863 = 12'h676 == _T_96[11:0] ? image_1654 : _GEN_7862; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7864 = 12'h677 == _T_96[11:0] ? image_1655 : _GEN_7863; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7865 = 12'h678 == _T_96[11:0] ? image_1656 : _GEN_7864; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7866 = 12'h679 == _T_96[11:0] ? image_1657 : _GEN_7865; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7867 = 12'h67a == _T_96[11:0] ? image_1658 : _GEN_7866; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7868 = 12'h67b == _T_96[11:0] ? image_1659 : _GEN_7867; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7869 = 12'h67c == _T_96[11:0] ? image_1660 : _GEN_7868; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7870 = 12'h67d == _T_96[11:0] ? 4'h0 : _GEN_7869; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7871 = 12'h67e == _T_96[11:0] ? 4'h0 : _GEN_7870; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7872 = 12'h67f == _T_96[11:0] ? 4'h0 : _GEN_7871; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7873 = 12'h680 == _T_96[11:0] ? image_1664 : _GEN_7872; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7874 = 12'h681 == _T_96[11:0] ? image_1665 : _GEN_7873; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7875 = 12'h682 == _T_96[11:0] ? image_1666 : _GEN_7874; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7876 = 12'h683 == _T_96[11:0] ? image_1667 : _GEN_7875; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7877 = 12'h684 == _T_96[11:0] ? image_1668 : _GEN_7876; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7878 = 12'h685 == _T_96[11:0] ? image_1669 : _GEN_7877; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7879 = 12'h686 == _T_96[11:0] ? image_1670 : _GEN_7878; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7880 = 12'h687 == _T_96[11:0] ? image_1671 : _GEN_7879; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7881 = 12'h688 == _T_96[11:0] ? image_1672 : _GEN_7880; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7882 = 12'h689 == _T_96[11:0] ? image_1673 : _GEN_7881; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7883 = 12'h68a == _T_96[11:0] ? image_1674 : _GEN_7882; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7884 = 12'h68b == _T_96[11:0] ? image_1675 : _GEN_7883; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7885 = 12'h68c == _T_96[11:0] ? image_1676 : _GEN_7884; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7886 = 12'h68d == _T_96[11:0] ? image_1677 : _GEN_7885; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7887 = 12'h68e == _T_96[11:0] ? image_1678 : _GEN_7886; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7888 = 12'h68f == _T_96[11:0] ? image_1679 : _GEN_7887; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7889 = 12'h690 == _T_96[11:0] ? image_1680 : _GEN_7888; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7890 = 12'h691 == _T_96[11:0] ? image_1681 : _GEN_7889; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7891 = 12'h692 == _T_96[11:0] ? image_1682 : _GEN_7890; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7892 = 12'h693 == _T_96[11:0] ? image_1683 : _GEN_7891; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7893 = 12'h694 == _T_96[11:0] ? image_1684 : _GEN_7892; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7894 = 12'h695 == _T_96[11:0] ? image_1685 : _GEN_7893; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7895 = 12'h696 == _T_96[11:0] ? image_1686 : _GEN_7894; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7896 = 12'h697 == _T_96[11:0] ? image_1687 : _GEN_7895; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7897 = 12'h698 == _T_96[11:0] ? image_1688 : _GEN_7896; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7898 = 12'h699 == _T_96[11:0] ? image_1689 : _GEN_7897; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7899 = 12'h69a == _T_96[11:0] ? image_1690 : _GEN_7898; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7900 = 12'h69b == _T_96[11:0] ? image_1691 : _GEN_7899; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7901 = 12'h69c == _T_96[11:0] ? image_1692 : _GEN_7900; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7902 = 12'h69d == _T_96[11:0] ? image_1693 : _GEN_7901; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7903 = 12'h69e == _T_96[11:0] ? image_1694 : _GEN_7902; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7904 = 12'h69f == _T_96[11:0] ? image_1695 : _GEN_7903; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7905 = 12'h6a0 == _T_96[11:0] ? image_1696 : _GEN_7904; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7906 = 12'h6a1 == _T_96[11:0] ? image_1697 : _GEN_7905; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7907 = 12'h6a2 == _T_96[11:0] ? image_1698 : _GEN_7906; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7908 = 12'h6a3 == _T_96[11:0] ? image_1699 : _GEN_7907; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7909 = 12'h6a4 == _T_96[11:0] ? image_1700 : _GEN_7908; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7910 = 12'h6a5 == _T_96[11:0] ? image_1701 : _GEN_7909; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7911 = 12'h6a6 == _T_96[11:0] ? image_1702 : _GEN_7910; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7912 = 12'h6a7 == _T_96[11:0] ? image_1703 : _GEN_7911; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7913 = 12'h6a8 == _T_96[11:0] ? image_1704 : _GEN_7912; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7914 = 12'h6a9 == _T_96[11:0] ? image_1705 : _GEN_7913; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7915 = 12'h6aa == _T_96[11:0] ? image_1706 : _GEN_7914; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7916 = 12'h6ab == _T_96[11:0] ? image_1707 : _GEN_7915; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7917 = 12'h6ac == _T_96[11:0] ? image_1708 : _GEN_7916; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7918 = 12'h6ad == _T_96[11:0] ? image_1709 : _GEN_7917; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7919 = 12'h6ae == _T_96[11:0] ? image_1710 : _GEN_7918; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7920 = 12'h6af == _T_96[11:0] ? image_1711 : _GEN_7919; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7921 = 12'h6b0 == _T_96[11:0] ? image_1712 : _GEN_7920; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7922 = 12'h6b1 == _T_96[11:0] ? image_1713 : _GEN_7921; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7923 = 12'h6b2 == _T_96[11:0] ? image_1714 : _GEN_7922; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7924 = 12'h6b3 == _T_96[11:0] ? image_1715 : _GEN_7923; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7925 = 12'h6b4 == _T_96[11:0] ? image_1716 : _GEN_7924; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7926 = 12'h6b5 == _T_96[11:0] ? image_1717 : _GEN_7925; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7927 = 12'h6b6 == _T_96[11:0] ? image_1718 : _GEN_7926; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7928 = 12'h6b7 == _T_96[11:0] ? image_1719 : _GEN_7927; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7929 = 12'h6b8 == _T_96[11:0] ? image_1720 : _GEN_7928; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7930 = 12'h6b9 == _T_96[11:0] ? image_1721 : _GEN_7929; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7931 = 12'h6ba == _T_96[11:0] ? image_1722 : _GEN_7930; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7932 = 12'h6bb == _T_96[11:0] ? image_1723 : _GEN_7931; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7933 = 12'h6bc == _T_96[11:0] ? 4'h0 : _GEN_7932; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7934 = 12'h6bd == _T_96[11:0] ? 4'h0 : _GEN_7933; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7935 = 12'h6be == _T_96[11:0] ? 4'h0 : _GEN_7934; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7936 = 12'h6bf == _T_96[11:0] ? 4'h0 : _GEN_7935; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7937 = 12'h6c0 == _T_96[11:0] ? image_1728 : _GEN_7936; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7938 = 12'h6c1 == _T_96[11:0] ? image_1729 : _GEN_7937; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7939 = 12'h6c2 == _T_96[11:0] ? image_1730 : _GEN_7938; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7940 = 12'h6c3 == _T_96[11:0] ? image_1731 : _GEN_7939; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7941 = 12'h6c4 == _T_96[11:0] ? image_1732 : _GEN_7940; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7942 = 12'h6c5 == _T_96[11:0] ? image_1733 : _GEN_7941; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7943 = 12'h6c6 == _T_96[11:0] ? image_1734 : _GEN_7942; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7944 = 12'h6c7 == _T_96[11:0] ? image_1735 : _GEN_7943; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7945 = 12'h6c8 == _T_96[11:0] ? image_1736 : _GEN_7944; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7946 = 12'h6c9 == _T_96[11:0] ? image_1737 : _GEN_7945; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7947 = 12'h6ca == _T_96[11:0] ? image_1738 : _GEN_7946; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7948 = 12'h6cb == _T_96[11:0] ? image_1739 : _GEN_7947; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7949 = 12'h6cc == _T_96[11:0] ? image_1740 : _GEN_7948; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7950 = 12'h6cd == _T_96[11:0] ? image_1741 : _GEN_7949; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7951 = 12'h6ce == _T_96[11:0] ? image_1742 : _GEN_7950; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7952 = 12'h6cf == _T_96[11:0] ? image_1743 : _GEN_7951; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7953 = 12'h6d0 == _T_96[11:0] ? image_1744 : _GEN_7952; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7954 = 12'h6d1 == _T_96[11:0] ? image_1745 : _GEN_7953; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7955 = 12'h6d2 == _T_96[11:0] ? image_1746 : _GEN_7954; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7956 = 12'h6d3 == _T_96[11:0] ? image_1747 : _GEN_7955; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7957 = 12'h6d4 == _T_96[11:0] ? image_1748 : _GEN_7956; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7958 = 12'h6d5 == _T_96[11:0] ? image_1749 : _GEN_7957; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7959 = 12'h6d6 == _T_96[11:0] ? image_1750 : _GEN_7958; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7960 = 12'h6d7 == _T_96[11:0] ? image_1751 : _GEN_7959; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7961 = 12'h6d8 == _T_96[11:0] ? image_1752 : _GEN_7960; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7962 = 12'h6d9 == _T_96[11:0] ? image_1753 : _GEN_7961; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7963 = 12'h6da == _T_96[11:0] ? image_1754 : _GEN_7962; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7964 = 12'h6db == _T_96[11:0] ? image_1755 : _GEN_7963; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7965 = 12'h6dc == _T_96[11:0] ? image_1756 : _GEN_7964; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7966 = 12'h6dd == _T_96[11:0] ? image_1757 : _GEN_7965; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7967 = 12'h6de == _T_96[11:0] ? image_1758 : _GEN_7966; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7968 = 12'h6df == _T_96[11:0] ? image_1759 : _GEN_7967; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7969 = 12'h6e0 == _T_96[11:0] ? image_1760 : _GEN_7968; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7970 = 12'h6e1 == _T_96[11:0] ? image_1761 : _GEN_7969; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7971 = 12'h6e2 == _T_96[11:0] ? image_1762 : _GEN_7970; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7972 = 12'h6e3 == _T_96[11:0] ? image_1763 : _GEN_7971; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7973 = 12'h6e4 == _T_96[11:0] ? image_1764 : _GEN_7972; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7974 = 12'h6e5 == _T_96[11:0] ? image_1765 : _GEN_7973; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7975 = 12'h6e6 == _T_96[11:0] ? image_1766 : _GEN_7974; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7976 = 12'h6e7 == _T_96[11:0] ? image_1767 : _GEN_7975; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7977 = 12'h6e8 == _T_96[11:0] ? image_1768 : _GEN_7976; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7978 = 12'h6e9 == _T_96[11:0] ? image_1769 : _GEN_7977; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7979 = 12'h6ea == _T_96[11:0] ? image_1770 : _GEN_7978; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7980 = 12'h6eb == _T_96[11:0] ? image_1771 : _GEN_7979; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7981 = 12'h6ec == _T_96[11:0] ? image_1772 : _GEN_7980; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7982 = 12'h6ed == _T_96[11:0] ? image_1773 : _GEN_7981; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7983 = 12'h6ee == _T_96[11:0] ? image_1774 : _GEN_7982; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7984 = 12'h6ef == _T_96[11:0] ? image_1775 : _GEN_7983; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7985 = 12'h6f0 == _T_96[11:0] ? image_1776 : _GEN_7984; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7986 = 12'h6f1 == _T_96[11:0] ? image_1777 : _GEN_7985; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7987 = 12'h6f2 == _T_96[11:0] ? image_1778 : _GEN_7986; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7988 = 12'h6f3 == _T_96[11:0] ? image_1779 : _GEN_7987; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7989 = 12'h6f4 == _T_96[11:0] ? image_1780 : _GEN_7988; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7990 = 12'h6f5 == _T_96[11:0] ? image_1781 : _GEN_7989; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7991 = 12'h6f6 == _T_96[11:0] ? image_1782 : _GEN_7990; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7992 = 12'h6f7 == _T_96[11:0] ? image_1783 : _GEN_7991; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7993 = 12'h6f8 == _T_96[11:0] ? image_1784 : _GEN_7992; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7994 = 12'h6f9 == _T_96[11:0] ? image_1785 : _GEN_7993; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7995 = 12'h6fa == _T_96[11:0] ? image_1786 : _GEN_7994; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7996 = 12'h6fb == _T_96[11:0] ? 4'h0 : _GEN_7995; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7997 = 12'h6fc == _T_96[11:0] ? 4'h0 : _GEN_7996; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7998 = 12'h6fd == _T_96[11:0] ? 4'h0 : _GEN_7997; // @[Filter.scala 138:46]
  wire [3:0] _GEN_7999 = 12'h6fe == _T_96[11:0] ? 4'h0 : _GEN_7998; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8000 = 12'h6ff == _T_96[11:0] ? 4'h0 : _GEN_7999; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8001 = 12'h700 == _T_96[11:0] ? 4'h0 : _GEN_8000; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8002 = 12'h701 == _T_96[11:0] ? image_1793 : _GEN_8001; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8003 = 12'h702 == _T_96[11:0] ? image_1794 : _GEN_8002; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8004 = 12'h703 == _T_96[11:0] ? image_1795 : _GEN_8003; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8005 = 12'h704 == _T_96[11:0] ? image_1796 : _GEN_8004; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8006 = 12'h705 == _T_96[11:0] ? image_1797 : _GEN_8005; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8007 = 12'h706 == _T_96[11:0] ? image_1798 : _GEN_8006; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8008 = 12'h707 == _T_96[11:0] ? image_1799 : _GEN_8007; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8009 = 12'h708 == _T_96[11:0] ? image_1800 : _GEN_8008; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8010 = 12'h709 == _T_96[11:0] ? image_1801 : _GEN_8009; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8011 = 12'h70a == _T_96[11:0] ? image_1802 : _GEN_8010; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8012 = 12'h70b == _T_96[11:0] ? image_1803 : _GEN_8011; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8013 = 12'h70c == _T_96[11:0] ? image_1804 : _GEN_8012; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8014 = 12'h70d == _T_96[11:0] ? image_1805 : _GEN_8013; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8015 = 12'h70e == _T_96[11:0] ? image_1806 : _GEN_8014; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8016 = 12'h70f == _T_96[11:0] ? image_1807 : _GEN_8015; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8017 = 12'h710 == _T_96[11:0] ? image_1808 : _GEN_8016; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8018 = 12'h711 == _T_96[11:0] ? image_1809 : _GEN_8017; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8019 = 12'h712 == _T_96[11:0] ? image_1810 : _GEN_8018; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8020 = 12'h713 == _T_96[11:0] ? image_1811 : _GEN_8019; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8021 = 12'h714 == _T_96[11:0] ? image_1812 : _GEN_8020; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8022 = 12'h715 == _T_96[11:0] ? image_1813 : _GEN_8021; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8023 = 12'h716 == _T_96[11:0] ? image_1814 : _GEN_8022; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8024 = 12'h717 == _T_96[11:0] ? image_1815 : _GEN_8023; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8025 = 12'h718 == _T_96[11:0] ? image_1816 : _GEN_8024; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8026 = 12'h719 == _T_96[11:0] ? image_1817 : _GEN_8025; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8027 = 12'h71a == _T_96[11:0] ? image_1818 : _GEN_8026; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8028 = 12'h71b == _T_96[11:0] ? image_1819 : _GEN_8027; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8029 = 12'h71c == _T_96[11:0] ? image_1820 : _GEN_8028; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8030 = 12'h71d == _T_96[11:0] ? image_1821 : _GEN_8029; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8031 = 12'h71e == _T_96[11:0] ? image_1822 : _GEN_8030; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8032 = 12'h71f == _T_96[11:0] ? image_1823 : _GEN_8031; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8033 = 12'h720 == _T_96[11:0] ? image_1824 : _GEN_8032; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8034 = 12'h721 == _T_96[11:0] ? image_1825 : _GEN_8033; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8035 = 12'h722 == _T_96[11:0] ? image_1826 : _GEN_8034; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8036 = 12'h723 == _T_96[11:0] ? image_1827 : _GEN_8035; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8037 = 12'h724 == _T_96[11:0] ? image_1828 : _GEN_8036; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8038 = 12'h725 == _T_96[11:0] ? image_1829 : _GEN_8037; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8039 = 12'h726 == _T_96[11:0] ? image_1830 : _GEN_8038; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8040 = 12'h727 == _T_96[11:0] ? image_1831 : _GEN_8039; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8041 = 12'h728 == _T_96[11:0] ? image_1832 : _GEN_8040; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8042 = 12'h729 == _T_96[11:0] ? image_1833 : _GEN_8041; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8043 = 12'h72a == _T_96[11:0] ? image_1834 : _GEN_8042; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8044 = 12'h72b == _T_96[11:0] ? image_1835 : _GEN_8043; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8045 = 12'h72c == _T_96[11:0] ? image_1836 : _GEN_8044; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8046 = 12'h72d == _T_96[11:0] ? image_1837 : _GEN_8045; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8047 = 12'h72e == _T_96[11:0] ? image_1838 : _GEN_8046; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8048 = 12'h72f == _T_96[11:0] ? image_1839 : _GEN_8047; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8049 = 12'h730 == _T_96[11:0] ? image_1840 : _GEN_8048; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8050 = 12'h731 == _T_96[11:0] ? image_1841 : _GEN_8049; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8051 = 12'h732 == _T_96[11:0] ? image_1842 : _GEN_8050; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8052 = 12'h733 == _T_96[11:0] ? image_1843 : _GEN_8051; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8053 = 12'h734 == _T_96[11:0] ? image_1844 : _GEN_8052; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8054 = 12'h735 == _T_96[11:0] ? image_1845 : _GEN_8053; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8055 = 12'h736 == _T_96[11:0] ? image_1846 : _GEN_8054; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8056 = 12'h737 == _T_96[11:0] ? image_1847 : _GEN_8055; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8057 = 12'h738 == _T_96[11:0] ? image_1848 : _GEN_8056; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8058 = 12'h739 == _T_96[11:0] ? image_1849 : _GEN_8057; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8059 = 12'h73a == _T_96[11:0] ? 4'h0 : _GEN_8058; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8060 = 12'h73b == _T_96[11:0] ? 4'h0 : _GEN_8059; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8061 = 12'h73c == _T_96[11:0] ? 4'h0 : _GEN_8060; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8062 = 12'h73d == _T_96[11:0] ? 4'h0 : _GEN_8061; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8063 = 12'h73e == _T_96[11:0] ? 4'h0 : _GEN_8062; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8064 = 12'h73f == _T_96[11:0] ? 4'h0 : _GEN_8063; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8065 = 12'h740 == _T_96[11:0] ? 4'h0 : _GEN_8064; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8066 = 12'h741 == _T_96[11:0] ? image_1857 : _GEN_8065; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8067 = 12'h742 == _T_96[11:0] ? image_1858 : _GEN_8066; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8068 = 12'h743 == _T_96[11:0] ? image_1859 : _GEN_8067; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8069 = 12'h744 == _T_96[11:0] ? image_1860 : _GEN_8068; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8070 = 12'h745 == _T_96[11:0] ? image_1861 : _GEN_8069; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8071 = 12'h746 == _T_96[11:0] ? image_1862 : _GEN_8070; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8072 = 12'h747 == _T_96[11:0] ? image_1863 : _GEN_8071; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8073 = 12'h748 == _T_96[11:0] ? image_1864 : _GEN_8072; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8074 = 12'h749 == _T_96[11:0] ? image_1865 : _GEN_8073; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8075 = 12'h74a == _T_96[11:0] ? image_1866 : _GEN_8074; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8076 = 12'h74b == _T_96[11:0] ? image_1867 : _GEN_8075; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8077 = 12'h74c == _T_96[11:0] ? image_1868 : _GEN_8076; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8078 = 12'h74d == _T_96[11:0] ? image_1869 : _GEN_8077; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8079 = 12'h74e == _T_96[11:0] ? image_1870 : _GEN_8078; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8080 = 12'h74f == _T_96[11:0] ? image_1871 : _GEN_8079; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8081 = 12'h750 == _T_96[11:0] ? image_1872 : _GEN_8080; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8082 = 12'h751 == _T_96[11:0] ? image_1873 : _GEN_8081; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8083 = 12'h752 == _T_96[11:0] ? image_1874 : _GEN_8082; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8084 = 12'h753 == _T_96[11:0] ? image_1875 : _GEN_8083; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8085 = 12'h754 == _T_96[11:0] ? image_1876 : _GEN_8084; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8086 = 12'h755 == _T_96[11:0] ? image_1877 : _GEN_8085; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8087 = 12'h756 == _T_96[11:0] ? image_1878 : _GEN_8086; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8088 = 12'h757 == _T_96[11:0] ? image_1879 : _GEN_8087; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8089 = 12'h758 == _T_96[11:0] ? image_1880 : _GEN_8088; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8090 = 12'h759 == _T_96[11:0] ? image_1881 : _GEN_8089; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8091 = 12'h75a == _T_96[11:0] ? image_1882 : _GEN_8090; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8092 = 12'h75b == _T_96[11:0] ? image_1883 : _GEN_8091; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8093 = 12'h75c == _T_96[11:0] ? image_1884 : _GEN_8092; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8094 = 12'h75d == _T_96[11:0] ? image_1885 : _GEN_8093; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8095 = 12'h75e == _T_96[11:0] ? image_1886 : _GEN_8094; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8096 = 12'h75f == _T_96[11:0] ? image_1887 : _GEN_8095; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8097 = 12'h760 == _T_96[11:0] ? image_1888 : _GEN_8096; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8098 = 12'h761 == _T_96[11:0] ? image_1889 : _GEN_8097; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8099 = 12'h762 == _T_96[11:0] ? image_1890 : _GEN_8098; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8100 = 12'h763 == _T_96[11:0] ? image_1891 : _GEN_8099; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8101 = 12'h764 == _T_96[11:0] ? image_1892 : _GEN_8100; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8102 = 12'h765 == _T_96[11:0] ? image_1893 : _GEN_8101; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8103 = 12'h766 == _T_96[11:0] ? image_1894 : _GEN_8102; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8104 = 12'h767 == _T_96[11:0] ? image_1895 : _GEN_8103; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8105 = 12'h768 == _T_96[11:0] ? image_1896 : _GEN_8104; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8106 = 12'h769 == _T_96[11:0] ? image_1897 : _GEN_8105; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8107 = 12'h76a == _T_96[11:0] ? image_1898 : _GEN_8106; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8108 = 12'h76b == _T_96[11:0] ? image_1899 : _GEN_8107; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8109 = 12'h76c == _T_96[11:0] ? image_1900 : _GEN_8108; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8110 = 12'h76d == _T_96[11:0] ? image_1901 : _GEN_8109; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8111 = 12'h76e == _T_96[11:0] ? image_1902 : _GEN_8110; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8112 = 12'h76f == _T_96[11:0] ? image_1903 : _GEN_8111; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8113 = 12'h770 == _T_96[11:0] ? image_1904 : _GEN_8112; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8114 = 12'h771 == _T_96[11:0] ? image_1905 : _GEN_8113; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8115 = 12'h772 == _T_96[11:0] ? image_1906 : _GEN_8114; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8116 = 12'h773 == _T_96[11:0] ? image_1907 : _GEN_8115; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8117 = 12'h774 == _T_96[11:0] ? image_1908 : _GEN_8116; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8118 = 12'h775 == _T_96[11:0] ? image_1909 : _GEN_8117; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8119 = 12'h776 == _T_96[11:0] ? image_1910 : _GEN_8118; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8120 = 12'h777 == _T_96[11:0] ? image_1911 : _GEN_8119; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8121 = 12'h778 == _T_96[11:0] ? image_1912 : _GEN_8120; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8122 = 12'h779 == _T_96[11:0] ? image_1913 : _GEN_8121; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8123 = 12'h77a == _T_96[11:0] ? 4'h0 : _GEN_8122; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8124 = 12'h77b == _T_96[11:0] ? 4'h0 : _GEN_8123; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8125 = 12'h77c == _T_96[11:0] ? 4'h0 : _GEN_8124; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8126 = 12'h77d == _T_96[11:0] ? 4'h0 : _GEN_8125; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8127 = 12'h77e == _T_96[11:0] ? 4'h0 : _GEN_8126; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8128 = 12'h77f == _T_96[11:0] ? 4'h0 : _GEN_8127; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8129 = 12'h780 == _T_96[11:0] ? 4'h0 : _GEN_8128; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8130 = 12'h781 == _T_96[11:0] ? image_1921 : _GEN_8129; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8131 = 12'h782 == _T_96[11:0] ? image_1922 : _GEN_8130; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8132 = 12'h783 == _T_96[11:0] ? image_1923 : _GEN_8131; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8133 = 12'h784 == _T_96[11:0] ? image_1924 : _GEN_8132; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8134 = 12'h785 == _T_96[11:0] ? image_1925 : _GEN_8133; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8135 = 12'h786 == _T_96[11:0] ? image_1926 : _GEN_8134; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8136 = 12'h787 == _T_96[11:0] ? image_1927 : _GEN_8135; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8137 = 12'h788 == _T_96[11:0] ? image_1928 : _GEN_8136; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8138 = 12'h789 == _T_96[11:0] ? image_1929 : _GEN_8137; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8139 = 12'h78a == _T_96[11:0] ? image_1930 : _GEN_8138; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8140 = 12'h78b == _T_96[11:0] ? image_1931 : _GEN_8139; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8141 = 12'h78c == _T_96[11:0] ? image_1932 : _GEN_8140; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8142 = 12'h78d == _T_96[11:0] ? image_1933 : _GEN_8141; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8143 = 12'h78e == _T_96[11:0] ? image_1934 : _GEN_8142; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8144 = 12'h78f == _T_96[11:0] ? image_1935 : _GEN_8143; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8145 = 12'h790 == _T_96[11:0] ? image_1936 : _GEN_8144; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8146 = 12'h791 == _T_96[11:0] ? image_1937 : _GEN_8145; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8147 = 12'h792 == _T_96[11:0] ? image_1938 : _GEN_8146; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8148 = 12'h793 == _T_96[11:0] ? image_1939 : _GEN_8147; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8149 = 12'h794 == _T_96[11:0] ? image_1940 : _GEN_8148; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8150 = 12'h795 == _T_96[11:0] ? image_1941 : _GEN_8149; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8151 = 12'h796 == _T_96[11:0] ? image_1942 : _GEN_8150; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8152 = 12'h797 == _T_96[11:0] ? image_1943 : _GEN_8151; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8153 = 12'h798 == _T_96[11:0] ? image_1944 : _GEN_8152; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8154 = 12'h799 == _T_96[11:0] ? image_1945 : _GEN_8153; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8155 = 12'h79a == _T_96[11:0] ? image_1946 : _GEN_8154; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8156 = 12'h79b == _T_96[11:0] ? image_1947 : _GEN_8155; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8157 = 12'h79c == _T_96[11:0] ? image_1948 : _GEN_8156; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8158 = 12'h79d == _T_96[11:0] ? image_1949 : _GEN_8157; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8159 = 12'h79e == _T_96[11:0] ? image_1950 : _GEN_8158; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8160 = 12'h79f == _T_96[11:0] ? image_1951 : _GEN_8159; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8161 = 12'h7a0 == _T_96[11:0] ? image_1952 : _GEN_8160; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8162 = 12'h7a1 == _T_96[11:0] ? image_1953 : _GEN_8161; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8163 = 12'h7a2 == _T_96[11:0] ? image_1954 : _GEN_8162; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8164 = 12'h7a3 == _T_96[11:0] ? image_1955 : _GEN_8163; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8165 = 12'h7a4 == _T_96[11:0] ? image_1956 : _GEN_8164; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8166 = 12'h7a5 == _T_96[11:0] ? image_1957 : _GEN_8165; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8167 = 12'h7a6 == _T_96[11:0] ? image_1958 : _GEN_8166; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8168 = 12'h7a7 == _T_96[11:0] ? image_1959 : _GEN_8167; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8169 = 12'h7a8 == _T_96[11:0] ? image_1960 : _GEN_8168; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8170 = 12'h7a9 == _T_96[11:0] ? image_1961 : _GEN_8169; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8171 = 12'h7aa == _T_96[11:0] ? image_1962 : _GEN_8170; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8172 = 12'h7ab == _T_96[11:0] ? image_1963 : _GEN_8171; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8173 = 12'h7ac == _T_96[11:0] ? image_1964 : _GEN_8172; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8174 = 12'h7ad == _T_96[11:0] ? image_1965 : _GEN_8173; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8175 = 12'h7ae == _T_96[11:0] ? image_1966 : _GEN_8174; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8176 = 12'h7af == _T_96[11:0] ? image_1967 : _GEN_8175; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8177 = 12'h7b0 == _T_96[11:0] ? image_1968 : _GEN_8176; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8178 = 12'h7b1 == _T_96[11:0] ? image_1969 : _GEN_8177; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8179 = 12'h7b2 == _T_96[11:0] ? image_1970 : _GEN_8178; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8180 = 12'h7b3 == _T_96[11:0] ? image_1971 : _GEN_8179; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8181 = 12'h7b4 == _T_96[11:0] ? image_1972 : _GEN_8180; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8182 = 12'h7b5 == _T_96[11:0] ? image_1973 : _GEN_8181; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8183 = 12'h7b6 == _T_96[11:0] ? image_1974 : _GEN_8182; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8184 = 12'h7b7 == _T_96[11:0] ? image_1975 : _GEN_8183; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8185 = 12'h7b8 == _T_96[11:0] ? image_1976 : _GEN_8184; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8186 = 12'h7b9 == _T_96[11:0] ? image_1977 : _GEN_8185; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8187 = 12'h7ba == _T_96[11:0] ? 4'h0 : _GEN_8186; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8188 = 12'h7bb == _T_96[11:0] ? 4'h0 : _GEN_8187; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8189 = 12'h7bc == _T_96[11:0] ? 4'h0 : _GEN_8188; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8190 = 12'h7bd == _T_96[11:0] ? 4'h0 : _GEN_8189; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8191 = 12'h7be == _T_96[11:0] ? 4'h0 : _GEN_8190; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8192 = 12'h7bf == _T_96[11:0] ? 4'h0 : _GEN_8191; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8193 = 12'h7c0 == _T_96[11:0] ? 4'h0 : _GEN_8192; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8194 = 12'h7c1 == _T_96[11:0] ? image_1985 : _GEN_8193; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8195 = 12'h7c2 == _T_96[11:0] ? image_1986 : _GEN_8194; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8196 = 12'h7c3 == _T_96[11:0] ? image_1987 : _GEN_8195; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8197 = 12'h7c4 == _T_96[11:0] ? image_1988 : _GEN_8196; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8198 = 12'h7c5 == _T_96[11:0] ? image_1989 : _GEN_8197; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8199 = 12'h7c6 == _T_96[11:0] ? image_1990 : _GEN_8198; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8200 = 12'h7c7 == _T_96[11:0] ? image_1991 : _GEN_8199; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8201 = 12'h7c8 == _T_96[11:0] ? image_1992 : _GEN_8200; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8202 = 12'h7c9 == _T_96[11:0] ? image_1993 : _GEN_8201; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8203 = 12'h7ca == _T_96[11:0] ? image_1994 : _GEN_8202; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8204 = 12'h7cb == _T_96[11:0] ? image_1995 : _GEN_8203; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8205 = 12'h7cc == _T_96[11:0] ? image_1996 : _GEN_8204; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8206 = 12'h7cd == _T_96[11:0] ? image_1997 : _GEN_8205; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8207 = 12'h7ce == _T_96[11:0] ? image_1998 : _GEN_8206; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8208 = 12'h7cf == _T_96[11:0] ? image_1999 : _GEN_8207; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8209 = 12'h7d0 == _T_96[11:0] ? image_2000 : _GEN_8208; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8210 = 12'h7d1 == _T_96[11:0] ? image_2001 : _GEN_8209; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8211 = 12'h7d2 == _T_96[11:0] ? image_2002 : _GEN_8210; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8212 = 12'h7d3 == _T_96[11:0] ? image_2003 : _GEN_8211; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8213 = 12'h7d4 == _T_96[11:0] ? image_2004 : _GEN_8212; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8214 = 12'h7d5 == _T_96[11:0] ? image_2005 : _GEN_8213; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8215 = 12'h7d6 == _T_96[11:0] ? image_2006 : _GEN_8214; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8216 = 12'h7d7 == _T_96[11:0] ? image_2007 : _GEN_8215; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8217 = 12'h7d8 == _T_96[11:0] ? image_2008 : _GEN_8216; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8218 = 12'h7d9 == _T_96[11:0] ? image_2009 : _GEN_8217; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8219 = 12'h7da == _T_96[11:0] ? image_2010 : _GEN_8218; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8220 = 12'h7db == _T_96[11:0] ? image_2011 : _GEN_8219; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8221 = 12'h7dc == _T_96[11:0] ? image_2012 : _GEN_8220; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8222 = 12'h7dd == _T_96[11:0] ? image_2013 : _GEN_8221; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8223 = 12'h7de == _T_96[11:0] ? image_2014 : _GEN_8222; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8224 = 12'h7df == _T_96[11:0] ? image_2015 : _GEN_8223; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8225 = 12'h7e0 == _T_96[11:0] ? image_2016 : _GEN_8224; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8226 = 12'h7e1 == _T_96[11:0] ? image_2017 : _GEN_8225; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8227 = 12'h7e2 == _T_96[11:0] ? image_2018 : _GEN_8226; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8228 = 12'h7e3 == _T_96[11:0] ? image_2019 : _GEN_8227; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8229 = 12'h7e4 == _T_96[11:0] ? image_2020 : _GEN_8228; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8230 = 12'h7e5 == _T_96[11:0] ? image_2021 : _GEN_8229; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8231 = 12'h7e6 == _T_96[11:0] ? image_2022 : _GEN_8230; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8232 = 12'h7e7 == _T_96[11:0] ? image_2023 : _GEN_8231; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8233 = 12'h7e8 == _T_96[11:0] ? image_2024 : _GEN_8232; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8234 = 12'h7e9 == _T_96[11:0] ? image_2025 : _GEN_8233; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8235 = 12'h7ea == _T_96[11:0] ? image_2026 : _GEN_8234; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8236 = 12'h7eb == _T_96[11:0] ? image_2027 : _GEN_8235; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8237 = 12'h7ec == _T_96[11:0] ? image_2028 : _GEN_8236; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8238 = 12'h7ed == _T_96[11:0] ? image_2029 : _GEN_8237; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8239 = 12'h7ee == _T_96[11:0] ? image_2030 : _GEN_8238; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8240 = 12'h7ef == _T_96[11:0] ? image_2031 : _GEN_8239; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8241 = 12'h7f0 == _T_96[11:0] ? image_2032 : _GEN_8240; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8242 = 12'h7f1 == _T_96[11:0] ? image_2033 : _GEN_8241; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8243 = 12'h7f2 == _T_96[11:0] ? image_2034 : _GEN_8242; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8244 = 12'h7f3 == _T_96[11:0] ? image_2035 : _GEN_8243; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8245 = 12'h7f4 == _T_96[11:0] ? image_2036 : _GEN_8244; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8246 = 12'h7f5 == _T_96[11:0] ? image_2037 : _GEN_8245; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8247 = 12'h7f6 == _T_96[11:0] ? image_2038 : _GEN_8246; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8248 = 12'h7f7 == _T_96[11:0] ? image_2039 : _GEN_8247; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8249 = 12'h7f8 == _T_96[11:0] ? image_2040 : _GEN_8248; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8250 = 12'h7f9 == _T_96[11:0] ? image_2041 : _GEN_8249; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8251 = 12'h7fa == _T_96[11:0] ? 4'h0 : _GEN_8250; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8252 = 12'h7fb == _T_96[11:0] ? 4'h0 : _GEN_8251; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8253 = 12'h7fc == _T_96[11:0] ? 4'h0 : _GEN_8252; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8254 = 12'h7fd == _T_96[11:0] ? 4'h0 : _GEN_8253; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8255 = 12'h7fe == _T_96[11:0] ? 4'h0 : _GEN_8254; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8256 = 12'h7ff == _T_96[11:0] ? 4'h0 : _GEN_8255; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8257 = 12'h800 == _T_96[11:0] ? 4'h0 : _GEN_8256; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8258 = 12'h801 == _T_96[11:0] ? image_2049 : _GEN_8257; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8259 = 12'h802 == _T_96[11:0] ? image_2050 : _GEN_8258; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8260 = 12'h803 == _T_96[11:0] ? image_2051 : _GEN_8259; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8261 = 12'h804 == _T_96[11:0] ? image_2052 : _GEN_8260; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8262 = 12'h805 == _T_96[11:0] ? image_2053 : _GEN_8261; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8263 = 12'h806 == _T_96[11:0] ? image_2054 : _GEN_8262; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8264 = 12'h807 == _T_96[11:0] ? image_2055 : _GEN_8263; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8265 = 12'h808 == _T_96[11:0] ? image_2056 : _GEN_8264; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8266 = 12'h809 == _T_96[11:0] ? image_2057 : _GEN_8265; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8267 = 12'h80a == _T_96[11:0] ? image_2058 : _GEN_8266; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8268 = 12'h80b == _T_96[11:0] ? image_2059 : _GEN_8267; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8269 = 12'h80c == _T_96[11:0] ? image_2060 : _GEN_8268; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8270 = 12'h80d == _T_96[11:0] ? image_2061 : _GEN_8269; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8271 = 12'h80e == _T_96[11:0] ? image_2062 : _GEN_8270; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8272 = 12'h80f == _T_96[11:0] ? image_2063 : _GEN_8271; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8273 = 12'h810 == _T_96[11:0] ? image_2064 : _GEN_8272; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8274 = 12'h811 == _T_96[11:0] ? image_2065 : _GEN_8273; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8275 = 12'h812 == _T_96[11:0] ? image_2066 : _GEN_8274; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8276 = 12'h813 == _T_96[11:0] ? image_2067 : _GEN_8275; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8277 = 12'h814 == _T_96[11:0] ? image_2068 : _GEN_8276; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8278 = 12'h815 == _T_96[11:0] ? image_2069 : _GEN_8277; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8279 = 12'h816 == _T_96[11:0] ? image_2070 : _GEN_8278; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8280 = 12'h817 == _T_96[11:0] ? image_2071 : _GEN_8279; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8281 = 12'h818 == _T_96[11:0] ? image_2072 : _GEN_8280; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8282 = 12'h819 == _T_96[11:0] ? image_2073 : _GEN_8281; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8283 = 12'h81a == _T_96[11:0] ? image_2074 : _GEN_8282; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8284 = 12'h81b == _T_96[11:0] ? image_2075 : _GEN_8283; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8285 = 12'h81c == _T_96[11:0] ? image_2076 : _GEN_8284; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8286 = 12'h81d == _T_96[11:0] ? image_2077 : _GEN_8285; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8287 = 12'h81e == _T_96[11:0] ? image_2078 : _GEN_8286; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8288 = 12'h81f == _T_96[11:0] ? image_2079 : _GEN_8287; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8289 = 12'h820 == _T_96[11:0] ? image_2080 : _GEN_8288; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8290 = 12'h821 == _T_96[11:0] ? image_2081 : _GEN_8289; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8291 = 12'h822 == _T_96[11:0] ? image_2082 : _GEN_8290; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8292 = 12'h823 == _T_96[11:0] ? image_2083 : _GEN_8291; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8293 = 12'h824 == _T_96[11:0] ? image_2084 : _GEN_8292; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8294 = 12'h825 == _T_96[11:0] ? image_2085 : _GEN_8293; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8295 = 12'h826 == _T_96[11:0] ? image_2086 : _GEN_8294; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8296 = 12'h827 == _T_96[11:0] ? image_2087 : _GEN_8295; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8297 = 12'h828 == _T_96[11:0] ? image_2088 : _GEN_8296; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8298 = 12'h829 == _T_96[11:0] ? image_2089 : _GEN_8297; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8299 = 12'h82a == _T_96[11:0] ? image_2090 : _GEN_8298; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8300 = 12'h82b == _T_96[11:0] ? image_2091 : _GEN_8299; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8301 = 12'h82c == _T_96[11:0] ? image_2092 : _GEN_8300; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8302 = 12'h82d == _T_96[11:0] ? image_2093 : _GEN_8301; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8303 = 12'h82e == _T_96[11:0] ? image_2094 : _GEN_8302; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8304 = 12'h82f == _T_96[11:0] ? image_2095 : _GEN_8303; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8305 = 12'h830 == _T_96[11:0] ? image_2096 : _GEN_8304; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8306 = 12'h831 == _T_96[11:0] ? image_2097 : _GEN_8305; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8307 = 12'h832 == _T_96[11:0] ? image_2098 : _GEN_8306; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8308 = 12'h833 == _T_96[11:0] ? image_2099 : _GEN_8307; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8309 = 12'h834 == _T_96[11:0] ? image_2100 : _GEN_8308; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8310 = 12'h835 == _T_96[11:0] ? image_2101 : _GEN_8309; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8311 = 12'h836 == _T_96[11:0] ? image_2102 : _GEN_8310; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8312 = 12'h837 == _T_96[11:0] ? image_2103 : _GEN_8311; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8313 = 12'h838 == _T_96[11:0] ? image_2104 : _GEN_8312; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8314 = 12'h839 == _T_96[11:0] ? image_2105 : _GEN_8313; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8315 = 12'h83a == _T_96[11:0] ? image_2106 : _GEN_8314; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8316 = 12'h83b == _T_96[11:0] ? 4'h0 : _GEN_8315; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8317 = 12'h83c == _T_96[11:0] ? 4'h0 : _GEN_8316; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8318 = 12'h83d == _T_96[11:0] ? 4'h0 : _GEN_8317; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8319 = 12'h83e == _T_96[11:0] ? 4'h0 : _GEN_8318; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8320 = 12'h83f == _T_96[11:0] ? 4'h0 : _GEN_8319; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8321 = 12'h840 == _T_96[11:0] ? 4'h0 : _GEN_8320; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8322 = 12'h841 == _T_96[11:0] ? 4'h0 : _GEN_8321; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8323 = 12'h842 == _T_96[11:0] ? image_2114 : _GEN_8322; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8324 = 12'h843 == _T_96[11:0] ? image_2115 : _GEN_8323; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8325 = 12'h844 == _T_96[11:0] ? image_2116 : _GEN_8324; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8326 = 12'h845 == _T_96[11:0] ? image_2117 : _GEN_8325; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8327 = 12'h846 == _T_96[11:0] ? image_2118 : _GEN_8326; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8328 = 12'h847 == _T_96[11:0] ? image_2119 : _GEN_8327; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8329 = 12'h848 == _T_96[11:0] ? image_2120 : _GEN_8328; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8330 = 12'h849 == _T_96[11:0] ? image_2121 : _GEN_8329; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8331 = 12'h84a == _T_96[11:0] ? image_2122 : _GEN_8330; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8332 = 12'h84b == _T_96[11:0] ? image_2123 : _GEN_8331; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8333 = 12'h84c == _T_96[11:0] ? image_2124 : _GEN_8332; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8334 = 12'h84d == _T_96[11:0] ? image_2125 : _GEN_8333; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8335 = 12'h84e == _T_96[11:0] ? image_2126 : _GEN_8334; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8336 = 12'h84f == _T_96[11:0] ? image_2127 : _GEN_8335; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8337 = 12'h850 == _T_96[11:0] ? image_2128 : _GEN_8336; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8338 = 12'h851 == _T_96[11:0] ? image_2129 : _GEN_8337; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8339 = 12'h852 == _T_96[11:0] ? image_2130 : _GEN_8338; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8340 = 12'h853 == _T_96[11:0] ? image_2131 : _GEN_8339; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8341 = 12'h854 == _T_96[11:0] ? image_2132 : _GEN_8340; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8342 = 12'h855 == _T_96[11:0] ? image_2133 : _GEN_8341; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8343 = 12'h856 == _T_96[11:0] ? image_2134 : _GEN_8342; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8344 = 12'h857 == _T_96[11:0] ? image_2135 : _GEN_8343; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8345 = 12'h858 == _T_96[11:0] ? image_2136 : _GEN_8344; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8346 = 12'h859 == _T_96[11:0] ? image_2137 : _GEN_8345; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8347 = 12'h85a == _T_96[11:0] ? image_2138 : _GEN_8346; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8348 = 12'h85b == _T_96[11:0] ? image_2139 : _GEN_8347; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8349 = 12'h85c == _T_96[11:0] ? image_2140 : _GEN_8348; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8350 = 12'h85d == _T_96[11:0] ? image_2141 : _GEN_8349; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8351 = 12'h85e == _T_96[11:0] ? image_2142 : _GEN_8350; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8352 = 12'h85f == _T_96[11:0] ? image_2143 : _GEN_8351; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8353 = 12'h860 == _T_96[11:0] ? image_2144 : _GEN_8352; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8354 = 12'h861 == _T_96[11:0] ? image_2145 : _GEN_8353; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8355 = 12'h862 == _T_96[11:0] ? image_2146 : _GEN_8354; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8356 = 12'h863 == _T_96[11:0] ? image_2147 : _GEN_8355; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8357 = 12'h864 == _T_96[11:0] ? image_2148 : _GEN_8356; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8358 = 12'h865 == _T_96[11:0] ? image_2149 : _GEN_8357; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8359 = 12'h866 == _T_96[11:0] ? image_2150 : _GEN_8358; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8360 = 12'h867 == _T_96[11:0] ? image_2151 : _GEN_8359; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8361 = 12'h868 == _T_96[11:0] ? image_2152 : _GEN_8360; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8362 = 12'h869 == _T_96[11:0] ? image_2153 : _GEN_8361; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8363 = 12'h86a == _T_96[11:0] ? image_2154 : _GEN_8362; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8364 = 12'h86b == _T_96[11:0] ? image_2155 : _GEN_8363; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8365 = 12'h86c == _T_96[11:0] ? image_2156 : _GEN_8364; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8366 = 12'h86d == _T_96[11:0] ? image_2157 : _GEN_8365; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8367 = 12'h86e == _T_96[11:0] ? image_2158 : _GEN_8366; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8368 = 12'h86f == _T_96[11:0] ? image_2159 : _GEN_8367; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8369 = 12'h870 == _T_96[11:0] ? image_2160 : _GEN_8368; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8370 = 12'h871 == _T_96[11:0] ? image_2161 : _GEN_8369; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8371 = 12'h872 == _T_96[11:0] ? image_2162 : _GEN_8370; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8372 = 12'h873 == _T_96[11:0] ? image_2163 : _GEN_8371; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8373 = 12'h874 == _T_96[11:0] ? image_2164 : _GEN_8372; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8374 = 12'h875 == _T_96[11:0] ? image_2165 : _GEN_8373; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8375 = 12'h876 == _T_96[11:0] ? image_2166 : _GEN_8374; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8376 = 12'h877 == _T_96[11:0] ? image_2167 : _GEN_8375; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8377 = 12'h878 == _T_96[11:0] ? image_2168 : _GEN_8376; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8378 = 12'h879 == _T_96[11:0] ? image_2169 : _GEN_8377; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8379 = 12'h87a == _T_96[11:0] ? image_2170 : _GEN_8378; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8380 = 12'h87b == _T_96[11:0] ? 4'h0 : _GEN_8379; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8381 = 12'h87c == _T_96[11:0] ? 4'h0 : _GEN_8380; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8382 = 12'h87d == _T_96[11:0] ? 4'h0 : _GEN_8381; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8383 = 12'h87e == _T_96[11:0] ? 4'h0 : _GEN_8382; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8384 = 12'h87f == _T_96[11:0] ? 4'h0 : _GEN_8383; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8385 = 12'h880 == _T_96[11:0] ? 4'h0 : _GEN_8384; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8386 = 12'h881 == _T_96[11:0] ? image_2177 : _GEN_8385; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8387 = 12'h882 == _T_96[11:0] ? image_2178 : _GEN_8386; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8388 = 12'h883 == _T_96[11:0] ? image_2179 : _GEN_8387; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8389 = 12'h884 == _T_96[11:0] ? image_2180 : _GEN_8388; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8390 = 12'h885 == _T_96[11:0] ? image_2181 : _GEN_8389; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8391 = 12'h886 == _T_96[11:0] ? image_2182 : _GEN_8390; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8392 = 12'h887 == _T_96[11:0] ? image_2183 : _GEN_8391; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8393 = 12'h888 == _T_96[11:0] ? image_2184 : _GEN_8392; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8394 = 12'h889 == _T_96[11:0] ? image_2185 : _GEN_8393; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8395 = 12'h88a == _T_96[11:0] ? image_2186 : _GEN_8394; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8396 = 12'h88b == _T_96[11:0] ? image_2187 : _GEN_8395; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8397 = 12'h88c == _T_96[11:0] ? image_2188 : _GEN_8396; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8398 = 12'h88d == _T_96[11:0] ? image_2189 : _GEN_8397; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8399 = 12'h88e == _T_96[11:0] ? image_2190 : _GEN_8398; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8400 = 12'h88f == _T_96[11:0] ? image_2191 : _GEN_8399; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8401 = 12'h890 == _T_96[11:0] ? image_2192 : _GEN_8400; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8402 = 12'h891 == _T_96[11:0] ? image_2193 : _GEN_8401; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8403 = 12'h892 == _T_96[11:0] ? image_2194 : _GEN_8402; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8404 = 12'h893 == _T_96[11:0] ? image_2195 : _GEN_8403; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8405 = 12'h894 == _T_96[11:0] ? image_2196 : _GEN_8404; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8406 = 12'h895 == _T_96[11:0] ? image_2197 : _GEN_8405; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8407 = 12'h896 == _T_96[11:0] ? image_2198 : _GEN_8406; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8408 = 12'h897 == _T_96[11:0] ? image_2199 : _GEN_8407; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8409 = 12'h898 == _T_96[11:0] ? image_2200 : _GEN_8408; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8410 = 12'h899 == _T_96[11:0] ? image_2201 : _GEN_8409; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8411 = 12'h89a == _T_96[11:0] ? image_2202 : _GEN_8410; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8412 = 12'h89b == _T_96[11:0] ? image_2203 : _GEN_8411; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8413 = 12'h89c == _T_96[11:0] ? image_2204 : _GEN_8412; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8414 = 12'h89d == _T_96[11:0] ? image_2205 : _GEN_8413; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8415 = 12'h89e == _T_96[11:0] ? image_2206 : _GEN_8414; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8416 = 12'h89f == _T_96[11:0] ? image_2207 : _GEN_8415; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8417 = 12'h8a0 == _T_96[11:0] ? image_2208 : _GEN_8416; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8418 = 12'h8a1 == _T_96[11:0] ? image_2209 : _GEN_8417; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8419 = 12'h8a2 == _T_96[11:0] ? image_2210 : _GEN_8418; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8420 = 12'h8a3 == _T_96[11:0] ? image_2211 : _GEN_8419; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8421 = 12'h8a4 == _T_96[11:0] ? image_2212 : _GEN_8420; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8422 = 12'h8a5 == _T_96[11:0] ? image_2213 : _GEN_8421; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8423 = 12'h8a6 == _T_96[11:0] ? image_2214 : _GEN_8422; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8424 = 12'h8a7 == _T_96[11:0] ? image_2215 : _GEN_8423; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8425 = 12'h8a8 == _T_96[11:0] ? image_2216 : _GEN_8424; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8426 = 12'h8a9 == _T_96[11:0] ? image_2217 : _GEN_8425; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8427 = 12'h8aa == _T_96[11:0] ? image_2218 : _GEN_8426; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8428 = 12'h8ab == _T_96[11:0] ? image_2219 : _GEN_8427; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8429 = 12'h8ac == _T_96[11:0] ? image_2220 : _GEN_8428; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8430 = 12'h8ad == _T_96[11:0] ? image_2221 : _GEN_8429; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8431 = 12'h8ae == _T_96[11:0] ? image_2222 : _GEN_8430; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8432 = 12'h8af == _T_96[11:0] ? image_2223 : _GEN_8431; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8433 = 12'h8b0 == _T_96[11:0] ? image_2224 : _GEN_8432; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8434 = 12'h8b1 == _T_96[11:0] ? image_2225 : _GEN_8433; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8435 = 12'h8b2 == _T_96[11:0] ? image_2226 : _GEN_8434; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8436 = 12'h8b3 == _T_96[11:0] ? image_2227 : _GEN_8435; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8437 = 12'h8b4 == _T_96[11:0] ? image_2228 : _GEN_8436; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8438 = 12'h8b5 == _T_96[11:0] ? image_2229 : _GEN_8437; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8439 = 12'h8b6 == _T_96[11:0] ? image_2230 : _GEN_8438; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8440 = 12'h8b7 == _T_96[11:0] ? image_2231 : _GEN_8439; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8441 = 12'h8b8 == _T_96[11:0] ? image_2232 : _GEN_8440; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8442 = 12'h8b9 == _T_96[11:0] ? image_2233 : _GEN_8441; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8443 = 12'h8ba == _T_96[11:0] ? image_2234 : _GEN_8442; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8444 = 12'h8bb == _T_96[11:0] ? 4'h0 : _GEN_8443; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8445 = 12'h8bc == _T_96[11:0] ? 4'h0 : _GEN_8444; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8446 = 12'h8bd == _T_96[11:0] ? 4'h0 : _GEN_8445; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8447 = 12'h8be == _T_96[11:0] ? 4'h0 : _GEN_8446; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8448 = 12'h8bf == _T_96[11:0] ? 4'h0 : _GEN_8447; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8449 = 12'h8c0 == _T_96[11:0] ? 4'h0 : _GEN_8448; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8450 = 12'h8c1 == _T_96[11:0] ? 4'h0 : _GEN_8449; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8451 = 12'h8c2 == _T_96[11:0] ? 4'h0 : _GEN_8450; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8452 = 12'h8c3 == _T_96[11:0] ? image_2243 : _GEN_8451; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8453 = 12'h8c4 == _T_96[11:0] ? image_2244 : _GEN_8452; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8454 = 12'h8c5 == _T_96[11:0] ? image_2245 : _GEN_8453; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8455 = 12'h8c6 == _T_96[11:0] ? image_2246 : _GEN_8454; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8456 = 12'h8c7 == _T_96[11:0] ? image_2247 : _GEN_8455; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8457 = 12'h8c8 == _T_96[11:0] ? image_2248 : _GEN_8456; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8458 = 12'h8c9 == _T_96[11:0] ? image_2249 : _GEN_8457; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8459 = 12'h8ca == _T_96[11:0] ? image_2250 : _GEN_8458; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8460 = 12'h8cb == _T_96[11:0] ? image_2251 : _GEN_8459; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8461 = 12'h8cc == _T_96[11:0] ? image_2252 : _GEN_8460; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8462 = 12'h8cd == _T_96[11:0] ? image_2253 : _GEN_8461; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8463 = 12'h8ce == _T_96[11:0] ? image_2254 : _GEN_8462; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8464 = 12'h8cf == _T_96[11:0] ? image_2255 : _GEN_8463; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8465 = 12'h8d0 == _T_96[11:0] ? image_2256 : _GEN_8464; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8466 = 12'h8d1 == _T_96[11:0] ? image_2257 : _GEN_8465; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8467 = 12'h8d2 == _T_96[11:0] ? image_2258 : _GEN_8466; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8468 = 12'h8d3 == _T_96[11:0] ? image_2259 : _GEN_8467; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8469 = 12'h8d4 == _T_96[11:0] ? image_2260 : _GEN_8468; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8470 = 12'h8d5 == _T_96[11:0] ? image_2261 : _GEN_8469; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8471 = 12'h8d6 == _T_96[11:0] ? image_2262 : _GEN_8470; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8472 = 12'h8d7 == _T_96[11:0] ? image_2263 : _GEN_8471; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8473 = 12'h8d8 == _T_96[11:0] ? image_2264 : _GEN_8472; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8474 = 12'h8d9 == _T_96[11:0] ? image_2265 : _GEN_8473; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8475 = 12'h8da == _T_96[11:0] ? image_2266 : _GEN_8474; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8476 = 12'h8db == _T_96[11:0] ? image_2267 : _GEN_8475; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8477 = 12'h8dc == _T_96[11:0] ? image_2268 : _GEN_8476; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8478 = 12'h8dd == _T_96[11:0] ? image_2269 : _GEN_8477; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8479 = 12'h8de == _T_96[11:0] ? image_2270 : _GEN_8478; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8480 = 12'h8df == _T_96[11:0] ? image_2271 : _GEN_8479; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8481 = 12'h8e0 == _T_96[11:0] ? image_2272 : _GEN_8480; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8482 = 12'h8e1 == _T_96[11:0] ? image_2273 : _GEN_8481; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8483 = 12'h8e2 == _T_96[11:0] ? image_2274 : _GEN_8482; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8484 = 12'h8e3 == _T_96[11:0] ? image_2275 : _GEN_8483; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8485 = 12'h8e4 == _T_96[11:0] ? image_2276 : _GEN_8484; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8486 = 12'h8e5 == _T_96[11:0] ? image_2277 : _GEN_8485; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8487 = 12'h8e6 == _T_96[11:0] ? image_2278 : _GEN_8486; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8488 = 12'h8e7 == _T_96[11:0] ? image_2279 : _GEN_8487; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8489 = 12'h8e8 == _T_96[11:0] ? image_2280 : _GEN_8488; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8490 = 12'h8e9 == _T_96[11:0] ? image_2281 : _GEN_8489; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8491 = 12'h8ea == _T_96[11:0] ? image_2282 : _GEN_8490; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8492 = 12'h8eb == _T_96[11:0] ? image_2283 : _GEN_8491; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8493 = 12'h8ec == _T_96[11:0] ? image_2284 : _GEN_8492; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8494 = 12'h8ed == _T_96[11:0] ? image_2285 : _GEN_8493; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8495 = 12'h8ee == _T_96[11:0] ? image_2286 : _GEN_8494; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8496 = 12'h8ef == _T_96[11:0] ? image_2287 : _GEN_8495; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8497 = 12'h8f0 == _T_96[11:0] ? image_2288 : _GEN_8496; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8498 = 12'h8f1 == _T_96[11:0] ? image_2289 : _GEN_8497; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8499 = 12'h8f2 == _T_96[11:0] ? image_2290 : _GEN_8498; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8500 = 12'h8f3 == _T_96[11:0] ? image_2291 : _GEN_8499; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8501 = 12'h8f4 == _T_96[11:0] ? image_2292 : _GEN_8500; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8502 = 12'h8f5 == _T_96[11:0] ? image_2293 : _GEN_8501; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8503 = 12'h8f6 == _T_96[11:0] ? image_2294 : _GEN_8502; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8504 = 12'h8f7 == _T_96[11:0] ? image_2295 : _GEN_8503; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8505 = 12'h8f8 == _T_96[11:0] ? image_2296 : _GEN_8504; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8506 = 12'h8f9 == _T_96[11:0] ? image_2297 : _GEN_8505; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8507 = 12'h8fa == _T_96[11:0] ? image_2298 : _GEN_8506; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8508 = 12'h8fb == _T_96[11:0] ? 4'h0 : _GEN_8507; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8509 = 12'h8fc == _T_96[11:0] ? 4'h0 : _GEN_8508; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8510 = 12'h8fd == _T_96[11:0] ? 4'h0 : _GEN_8509; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8511 = 12'h8fe == _T_96[11:0] ? 4'h0 : _GEN_8510; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8512 = 12'h8ff == _T_96[11:0] ? 4'h0 : _GEN_8511; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8513 = 12'h900 == _T_96[11:0] ? 4'h0 : _GEN_8512; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8514 = 12'h901 == _T_96[11:0] ? 4'h0 : _GEN_8513; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8515 = 12'h902 == _T_96[11:0] ? 4'h0 : _GEN_8514; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8516 = 12'h903 == _T_96[11:0] ? image_2307 : _GEN_8515; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8517 = 12'h904 == _T_96[11:0] ? image_2308 : _GEN_8516; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8518 = 12'h905 == _T_96[11:0] ? image_2309 : _GEN_8517; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8519 = 12'h906 == _T_96[11:0] ? image_2310 : _GEN_8518; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8520 = 12'h907 == _T_96[11:0] ? image_2311 : _GEN_8519; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8521 = 12'h908 == _T_96[11:0] ? image_2312 : _GEN_8520; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8522 = 12'h909 == _T_96[11:0] ? image_2313 : _GEN_8521; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8523 = 12'h90a == _T_96[11:0] ? image_2314 : _GEN_8522; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8524 = 12'h90b == _T_96[11:0] ? image_2315 : _GEN_8523; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8525 = 12'h90c == _T_96[11:0] ? image_2316 : _GEN_8524; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8526 = 12'h90d == _T_96[11:0] ? image_2317 : _GEN_8525; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8527 = 12'h90e == _T_96[11:0] ? image_2318 : _GEN_8526; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8528 = 12'h90f == _T_96[11:0] ? image_2319 : _GEN_8527; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8529 = 12'h910 == _T_96[11:0] ? image_2320 : _GEN_8528; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8530 = 12'h911 == _T_96[11:0] ? image_2321 : _GEN_8529; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8531 = 12'h912 == _T_96[11:0] ? image_2322 : _GEN_8530; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8532 = 12'h913 == _T_96[11:0] ? image_2323 : _GEN_8531; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8533 = 12'h914 == _T_96[11:0] ? image_2324 : _GEN_8532; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8534 = 12'h915 == _T_96[11:0] ? image_2325 : _GEN_8533; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8535 = 12'h916 == _T_96[11:0] ? image_2326 : _GEN_8534; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8536 = 12'h917 == _T_96[11:0] ? image_2327 : _GEN_8535; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8537 = 12'h918 == _T_96[11:0] ? image_2328 : _GEN_8536; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8538 = 12'h919 == _T_96[11:0] ? image_2329 : _GEN_8537; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8539 = 12'h91a == _T_96[11:0] ? image_2330 : _GEN_8538; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8540 = 12'h91b == _T_96[11:0] ? image_2331 : _GEN_8539; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8541 = 12'h91c == _T_96[11:0] ? image_2332 : _GEN_8540; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8542 = 12'h91d == _T_96[11:0] ? image_2333 : _GEN_8541; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8543 = 12'h91e == _T_96[11:0] ? image_2334 : _GEN_8542; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8544 = 12'h91f == _T_96[11:0] ? image_2335 : _GEN_8543; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8545 = 12'h920 == _T_96[11:0] ? image_2336 : _GEN_8544; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8546 = 12'h921 == _T_96[11:0] ? image_2337 : _GEN_8545; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8547 = 12'h922 == _T_96[11:0] ? image_2338 : _GEN_8546; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8548 = 12'h923 == _T_96[11:0] ? image_2339 : _GEN_8547; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8549 = 12'h924 == _T_96[11:0] ? image_2340 : _GEN_8548; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8550 = 12'h925 == _T_96[11:0] ? image_2341 : _GEN_8549; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8551 = 12'h926 == _T_96[11:0] ? image_2342 : _GEN_8550; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8552 = 12'h927 == _T_96[11:0] ? image_2343 : _GEN_8551; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8553 = 12'h928 == _T_96[11:0] ? image_2344 : _GEN_8552; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8554 = 12'h929 == _T_96[11:0] ? image_2345 : _GEN_8553; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8555 = 12'h92a == _T_96[11:0] ? image_2346 : _GEN_8554; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8556 = 12'h92b == _T_96[11:0] ? image_2347 : _GEN_8555; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8557 = 12'h92c == _T_96[11:0] ? image_2348 : _GEN_8556; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8558 = 12'h92d == _T_96[11:0] ? image_2349 : _GEN_8557; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8559 = 12'h92e == _T_96[11:0] ? image_2350 : _GEN_8558; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8560 = 12'h92f == _T_96[11:0] ? image_2351 : _GEN_8559; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8561 = 12'h930 == _T_96[11:0] ? image_2352 : _GEN_8560; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8562 = 12'h931 == _T_96[11:0] ? image_2353 : _GEN_8561; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8563 = 12'h932 == _T_96[11:0] ? image_2354 : _GEN_8562; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8564 = 12'h933 == _T_96[11:0] ? image_2355 : _GEN_8563; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8565 = 12'h934 == _T_96[11:0] ? image_2356 : _GEN_8564; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8566 = 12'h935 == _T_96[11:0] ? image_2357 : _GEN_8565; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8567 = 12'h936 == _T_96[11:0] ? image_2358 : _GEN_8566; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8568 = 12'h937 == _T_96[11:0] ? image_2359 : _GEN_8567; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8569 = 12'h938 == _T_96[11:0] ? image_2360 : _GEN_8568; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8570 = 12'h939 == _T_96[11:0] ? image_2361 : _GEN_8569; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8571 = 12'h93a == _T_96[11:0] ? image_2362 : _GEN_8570; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8572 = 12'h93b == _T_96[11:0] ? 4'h0 : _GEN_8571; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8573 = 12'h93c == _T_96[11:0] ? 4'h0 : _GEN_8572; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8574 = 12'h93d == _T_96[11:0] ? 4'h0 : _GEN_8573; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8575 = 12'h93e == _T_96[11:0] ? 4'h0 : _GEN_8574; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8576 = 12'h93f == _T_96[11:0] ? 4'h0 : _GEN_8575; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8577 = 12'h940 == _T_96[11:0] ? 4'h0 : _GEN_8576; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8578 = 12'h941 == _T_96[11:0] ? 4'h0 : _GEN_8577; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8579 = 12'h942 == _T_96[11:0] ? 4'h0 : _GEN_8578; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8580 = 12'h943 == _T_96[11:0] ? 4'h0 : _GEN_8579; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8581 = 12'h944 == _T_96[11:0] ? image_2372 : _GEN_8580; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8582 = 12'h945 == _T_96[11:0] ? image_2373 : _GEN_8581; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8583 = 12'h946 == _T_96[11:0] ? image_2374 : _GEN_8582; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8584 = 12'h947 == _T_96[11:0] ? image_2375 : _GEN_8583; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8585 = 12'h948 == _T_96[11:0] ? image_2376 : _GEN_8584; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8586 = 12'h949 == _T_96[11:0] ? image_2377 : _GEN_8585; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8587 = 12'h94a == _T_96[11:0] ? image_2378 : _GEN_8586; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8588 = 12'h94b == _T_96[11:0] ? image_2379 : _GEN_8587; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8589 = 12'h94c == _T_96[11:0] ? image_2380 : _GEN_8588; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8590 = 12'h94d == _T_96[11:0] ? image_2381 : _GEN_8589; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8591 = 12'h94e == _T_96[11:0] ? image_2382 : _GEN_8590; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8592 = 12'h94f == _T_96[11:0] ? image_2383 : _GEN_8591; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8593 = 12'h950 == _T_96[11:0] ? image_2384 : _GEN_8592; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8594 = 12'h951 == _T_96[11:0] ? image_2385 : _GEN_8593; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8595 = 12'h952 == _T_96[11:0] ? image_2386 : _GEN_8594; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8596 = 12'h953 == _T_96[11:0] ? image_2387 : _GEN_8595; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8597 = 12'h954 == _T_96[11:0] ? image_2388 : _GEN_8596; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8598 = 12'h955 == _T_96[11:0] ? image_2389 : _GEN_8597; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8599 = 12'h956 == _T_96[11:0] ? image_2390 : _GEN_8598; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8600 = 12'h957 == _T_96[11:0] ? image_2391 : _GEN_8599; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8601 = 12'h958 == _T_96[11:0] ? image_2392 : _GEN_8600; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8602 = 12'h959 == _T_96[11:0] ? image_2393 : _GEN_8601; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8603 = 12'h95a == _T_96[11:0] ? image_2394 : _GEN_8602; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8604 = 12'h95b == _T_96[11:0] ? image_2395 : _GEN_8603; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8605 = 12'h95c == _T_96[11:0] ? image_2396 : _GEN_8604; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8606 = 12'h95d == _T_96[11:0] ? image_2397 : _GEN_8605; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8607 = 12'h95e == _T_96[11:0] ? image_2398 : _GEN_8606; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8608 = 12'h95f == _T_96[11:0] ? image_2399 : _GEN_8607; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8609 = 12'h960 == _T_96[11:0] ? image_2400 : _GEN_8608; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8610 = 12'h961 == _T_96[11:0] ? image_2401 : _GEN_8609; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8611 = 12'h962 == _T_96[11:0] ? image_2402 : _GEN_8610; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8612 = 12'h963 == _T_96[11:0] ? image_2403 : _GEN_8611; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8613 = 12'h964 == _T_96[11:0] ? image_2404 : _GEN_8612; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8614 = 12'h965 == _T_96[11:0] ? image_2405 : _GEN_8613; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8615 = 12'h966 == _T_96[11:0] ? image_2406 : _GEN_8614; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8616 = 12'h967 == _T_96[11:0] ? image_2407 : _GEN_8615; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8617 = 12'h968 == _T_96[11:0] ? image_2408 : _GEN_8616; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8618 = 12'h969 == _T_96[11:0] ? image_2409 : _GEN_8617; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8619 = 12'h96a == _T_96[11:0] ? image_2410 : _GEN_8618; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8620 = 12'h96b == _T_96[11:0] ? image_2411 : _GEN_8619; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8621 = 12'h96c == _T_96[11:0] ? image_2412 : _GEN_8620; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8622 = 12'h96d == _T_96[11:0] ? image_2413 : _GEN_8621; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8623 = 12'h96e == _T_96[11:0] ? image_2414 : _GEN_8622; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8624 = 12'h96f == _T_96[11:0] ? image_2415 : _GEN_8623; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8625 = 12'h970 == _T_96[11:0] ? image_2416 : _GEN_8624; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8626 = 12'h971 == _T_96[11:0] ? image_2417 : _GEN_8625; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8627 = 12'h972 == _T_96[11:0] ? image_2418 : _GEN_8626; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8628 = 12'h973 == _T_96[11:0] ? image_2419 : _GEN_8627; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8629 = 12'h974 == _T_96[11:0] ? image_2420 : _GEN_8628; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8630 = 12'h975 == _T_96[11:0] ? image_2421 : _GEN_8629; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8631 = 12'h976 == _T_96[11:0] ? image_2422 : _GEN_8630; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8632 = 12'h977 == _T_96[11:0] ? image_2423 : _GEN_8631; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8633 = 12'h978 == _T_96[11:0] ? image_2424 : _GEN_8632; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8634 = 12'h979 == _T_96[11:0] ? image_2425 : _GEN_8633; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8635 = 12'h97a == _T_96[11:0] ? image_2426 : _GEN_8634; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8636 = 12'h97b == _T_96[11:0] ? 4'h0 : _GEN_8635; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8637 = 12'h97c == _T_96[11:0] ? 4'h0 : _GEN_8636; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8638 = 12'h97d == _T_96[11:0] ? 4'h0 : _GEN_8637; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8639 = 12'h97e == _T_96[11:0] ? 4'h0 : _GEN_8638; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8640 = 12'h97f == _T_96[11:0] ? 4'h0 : _GEN_8639; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8641 = 12'h980 == _T_96[11:0] ? 4'h0 : _GEN_8640; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8642 = 12'h981 == _T_96[11:0] ? 4'h0 : _GEN_8641; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8643 = 12'h982 == _T_96[11:0] ? 4'h0 : _GEN_8642; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8644 = 12'h983 == _T_96[11:0] ? 4'h0 : _GEN_8643; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8645 = 12'h984 == _T_96[11:0] ? 4'h0 : _GEN_8644; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8646 = 12'h985 == _T_96[11:0] ? image_2437 : _GEN_8645; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8647 = 12'h986 == _T_96[11:0] ? image_2438 : _GEN_8646; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8648 = 12'h987 == _T_96[11:0] ? image_2439 : _GEN_8647; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8649 = 12'h988 == _T_96[11:0] ? image_2440 : _GEN_8648; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8650 = 12'h989 == _T_96[11:0] ? image_2441 : _GEN_8649; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8651 = 12'h98a == _T_96[11:0] ? image_2442 : _GEN_8650; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8652 = 12'h98b == _T_96[11:0] ? image_2443 : _GEN_8651; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8653 = 12'h98c == _T_96[11:0] ? image_2444 : _GEN_8652; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8654 = 12'h98d == _T_96[11:0] ? image_2445 : _GEN_8653; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8655 = 12'h98e == _T_96[11:0] ? image_2446 : _GEN_8654; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8656 = 12'h98f == _T_96[11:0] ? image_2447 : _GEN_8655; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8657 = 12'h990 == _T_96[11:0] ? image_2448 : _GEN_8656; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8658 = 12'h991 == _T_96[11:0] ? image_2449 : _GEN_8657; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8659 = 12'h992 == _T_96[11:0] ? image_2450 : _GEN_8658; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8660 = 12'h993 == _T_96[11:0] ? image_2451 : _GEN_8659; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8661 = 12'h994 == _T_96[11:0] ? image_2452 : _GEN_8660; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8662 = 12'h995 == _T_96[11:0] ? image_2453 : _GEN_8661; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8663 = 12'h996 == _T_96[11:0] ? image_2454 : _GEN_8662; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8664 = 12'h997 == _T_96[11:0] ? image_2455 : _GEN_8663; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8665 = 12'h998 == _T_96[11:0] ? image_2456 : _GEN_8664; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8666 = 12'h999 == _T_96[11:0] ? image_2457 : _GEN_8665; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8667 = 12'h99a == _T_96[11:0] ? image_2458 : _GEN_8666; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8668 = 12'h99b == _T_96[11:0] ? image_2459 : _GEN_8667; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8669 = 12'h99c == _T_96[11:0] ? image_2460 : _GEN_8668; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8670 = 12'h99d == _T_96[11:0] ? image_2461 : _GEN_8669; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8671 = 12'h99e == _T_96[11:0] ? image_2462 : _GEN_8670; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8672 = 12'h99f == _T_96[11:0] ? image_2463 : _GEN_8671; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8673 = 12'h9a0 == _T_96[11:0] ? image_2464 : _GEN_8672; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8674 = 12'h9a1 == _T_96[11:0] ? image_2465 : _GEN_8673; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8675 = 12'h9a2 == _T_96[11:0] ? image_2466 : _GEN_8674; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8676 = 12'h9a3 == _T_96[11:0] ? image_2467 : _GEN_8675; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8677 = 12'h9a4 == _T_96[11:0] ? image_2468 : _GEN_8676; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8678 = 12'h9a5 == _T_96[11:0] ? image_2469 : _GEN_8677; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8679 = 12'h9a6 == _T_96[11:0] ? image_2470 : _GEN_8678; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8680 = 12'h9a7 == _T_96[11:0] ? image_2471 : _GEN_8679; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8681 = 12'h9a8 == _T_96[11:0] ? image_2472 : _GEN_8680; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8682 = 12'h9a9 == _T_96[11:0] ? image_2473 : _GEN_8681; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8683 = 12'h9aa == _T_96[11:0] ? image_2474 : _GEN_8682; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8684 = 12'h9ab == _T_96[11:0] ? image_2475 : _GEN_8683; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8685 = 12'h9ac == _T_96[11:0] ? image_2476 : _GEN_8684; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8686 = 12'h9ad == _T_96[11:0] ? image_2477 : _GEN_8685; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8687 = 12'h9ae == _T_96[11:0] ? image_2478 : _GEN_8686; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8688 = 12'h9af == _T_96[11:0] ? image_2479 : _GEN_8687; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8689 = 12'h9b0 == _T_96[11:0] ? image_2480 : _GEN_8688; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8690 = 12'h9b1 == _T_96[11:0] ? image_2481 : _GEN_8689; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8691 = 12'h9b2 == _T_96[11:0] ? image_2482 : _GEN_8690; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8692 = 12'h9b3 == _T_96[11:0] ? image_2483 : _GEN_8691; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8693 = 12'h9b4 == _T_96[11:0] ? image_2484 : _GEN_8692; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8694 = 12'h9b5 == _T_96[11:0] ? image_2485 : _GEN_8693; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8695 = 12'h9b6 == _T_96[11:0] ? image_2486 : _GEN_8694; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8696 = 12'h9b7 == _T_96[11:0] ? image_2487 : _GEN_8695; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8697 = 12'h9b8 == _T_96[11:0] ? image_2488 : _GEN_8696; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8698 = 12'h9b9 == _T_96[11:0] ? image_2489 : _GEN_8697; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8699 = 12'h9ba == _T_96[11:0] ? image_2490 : _GEN_8698; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8700 = 12'h9bb == _T_96[11:0] ? 4'h0 : _GEN_8699; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8701 = 12'h9bc == _T_96[11:0] ? 4'h0 : _GEN_8700; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8702 = 12'h9bd == _T_96[11:0] ? 4'h0 : _GEN_8701; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8703 = 12'h9be == _T_96[11:0] ? 4'h0 : _GEN_8702; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8704 = 12'h9bf == _T_96[11:0] ? 4'h0 : _GEN_8703; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8705 = 12'h9c0 == _T_96[11:0] ? 4'h0 : _GEN_8704; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8706 = 12'h9c1 == _T_96[11:0] ? 4'h0 : _GEN_8705; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8707 = 12'h9c2 == _T_96[11:0] ? 4'h0 : _GEN_8706; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8708 = 12'h9c3 == _T_96[11:0] ? 4'h0 : _GEN_8707; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8709 = 12'h9c4 == _T_96[11:0] ? 4'h0 : _GEN_8708; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8710 = 12'h9c5 == _T_96[11:0] ? 4'h0 : _GEN_8709; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8711 = 12'h9c6 == _T_96[11:0] ? image_2502 : _GEN_8710; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8712 = 12'h9c7 == _T_96[11:0] ? image_2503 : _GEN_8711; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8713 = 12'h9c8 == _T_96[11:0] ? image_2504 : _GEN_8712; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8714 = 12'h9c9 == _T_96[11:0] ? image_2505 : _GEN_8713; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8715 = 12'h9ca == _T_96[11:0] ? image_2506 : _GEN_8714; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8716 = 12'h9cb == _T_96[11:0] ? image_2507 : _GEN_8715; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8717 = 12'h9cc == _T_96[11:0] ? image_2508 : _GEN_8716; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8718 = 12'h9cd == _T_96[11:0] ? image_2509 : _GEN_8717; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8719 = 12'h9ce == _T_96[11:0] ? image_2510 : _GEN_8718; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8720 = 12'h9cf == _T_96[11:0] ? image_2511 : _GEN_8719; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8721 = 12'h9d0 == _T_96[11:0] ? image_2512 : _GEN_8720; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8722 = 12'h9d1 == _T_96[11:0] ? image_2513 : _GEN_8721; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8723 = 12'h9d2 == _T_96[11:0] ? image_2514 : _GEN_8722; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8724 = 12'h9d3 == _T_96[11:0] ? image_2515 : _GEN_8723; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8725 = 12'h9d4 == _T_96[11:0] ? image_2516 : _GEN_8724; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8726 = 12'h9d5 == _T_96[11:0] ? image_2517 : _GEN_8725; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8727 = 12'h9d6 == _T_96[11:0] ? image_2518 : _GEN_8726; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8728 = 12'h9d7 == _T_96[11:0] ? image_2519 : _GEN_8727; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8729 = 12'h9d8 == _T_96[11:0] ? image_2520 : _GEN_8728; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8730 = 12'h9d9 == _T_96[11:0] ? image_2521 : _GEN_8729; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8731 = 12'h9da == _T_96[11:0] ? image_2522 : _GEN_8730; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8732 = 12'h9db == _T_96[11:0] ? image_2523 : _GEN_8731; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8733 = 12'h9dc == _T_96[11:0] ? image_2524 : _GEN_8732; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8734 = 12'h9dd == _T_96[11:0] ? image_2525 : _GEN_8733; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8735 = 12'h9de == _T_96[11:0] ? image_2526 : _GEN_8734; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8736 = 12'h9df == _T_96[11:0] ? image_2527 : _GEN_8735; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8737 = 12'h9e0 == _T_96[11:0] ? image_2528 : _GEN_8736; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8738 = 12'h9e1 == _T_96[11:0] ? image_2529 : _GEN_8737; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8739 = 12'h9e2 == _T_96[11:0] ? image_2530 : _GEN_8738; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8740 = 12'h9e3 == _T_96[11:0] ? image_2531 : _GEN_8739; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8741 = 12'h9e4 == _T_96[11:0] ? image_2532 : _GEN_8740; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8742 = 12'h9e5 == _T_96[11:0] ? image_2533 : _GEN_8741; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8743 = 12'h9e6 == _T_96[11:0] ? image_2534 : _GEN_8742; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8744 = 12'h9e7 == _T_96[11:0] ? image_2535 : _GEN_8743; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8745 = 12'h9e8 == _T_96[11:0] ? image_2536 : _GEN_8744; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8746 = 12'h9e9 == _T_96[11:0] ? image_2537 : _GEN_8745; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8747 = 12'h9ea == _T_96[11:0] ? image_2538 : _GEN_8746; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8748 = 12'h9eb == _T_96[11:0] ? image_2539 : _GEN_8747; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8749 = 12'h9ec == _T_96[11:0] ? image_2540 : _GEN_8748; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8750 = 12'h9ed == _T_96[11:0] ? image_2541 : _GEN_8749; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8751 = 12'h9ee == _T_96[11:0] ? image_2542 : _GEN_8750; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8752 = 12'h9ef == _T_96[11:0] ? image_2543 : _GEN_8751; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8753 = 12'h9f0 == _T_96[11:0] ? image_2544 : _GEN_8752; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8754 = 12'h9f1 == _T_96[11:0] ? image_2545 : _GEN_8753; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8755 = 12'h9f2 == _T_96[11:0] ? image_2546 : _GEN_8754; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8756 = 12'h9f3 == _T_96[11:0] ? image_2547 : _GEN_8755; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8757 = 12'h9f4 == _T_96[11:0] ? image_2548 : _GEN_8756; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8758 = 12'h9f5 == _T_96[11:0] ? image_2549 : _GEN_8757; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8759 = 12'h9f6 == _T_96[11:0] ? image_2550 : _GEN_8758; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8760 = 12'h9f7 == _T_96[11:0] ? image_2551 : _GEN_8759; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8761 = 12'h9f8 == _T_96[11:0] ? image_2552 : _GEN_8760; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8762 = 12'h9f9 == _T_96[11:0] ? image_2553 : _GEN_8761; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8763 = 12'h9fa == _T_96[11:0] ? image_2554 : _GEN_8762; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8764 = 12'h9fb == _T_96[11:0] ? 4'h0 : _GEN_8763; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8765 = 12'h9fc == _T_96[11:0] ? 4'h0 : _GEN_8764; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8766 = 12'h9fd == _T_96[11:0] ? 4'h0 : _GEN_8765; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8767 = 12'h9fe == _T_96[11:0] ? 4'h0 : _GEN_8766; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8768 = 12'h9ff == _T_96[11:0] ? 4'h0 : _GEN_8767; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8769 = 12'ha00 == _T_96[11:0] ? 4'h0 : _GEN_8768; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8770 = 12'ha01 == _T_96[11:0] ? 4'h0 : _GEN_8769; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8771 = 12'ha02 == _T_96[11:0] ? 4'h0 : _GEN_8770; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8772 = 12'ha03 == _T_96[11:0] ? 4'h0 : _GEN_8771; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8773 = 12'ha04 == _T_96[11:0] ? 4'h0 : _GEN_8772; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8774 = 12'ha05 == _T_96[11:0] ? 4'h0 : _GEN_8773; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8775 = 12'ha06 == _T_96[11:0] ? 4'h0 : _GEN_8774; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8776 = 12'ha07 == _T_96[11:0] ? image_2567 : _GEN_8775; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8777 = 12'ha08 == _T_96[11:0] ? image_2568 : _GEN_8776; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8778 = 12'ha09 == _T_96[11:0] ? image_2569 : _GEN_8777; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8779 = 12'ha0a == _T_96[11:0] ? image_2570 : _GEN_8778; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8780 = 12'ha0b == _T_96[11:0] ? image_2571 : _GEN_8779; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8781 = 12'ha0c == _T_96[11:0] ? image_2572 : _GEN_8780; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8782 = 12'ha0d == _T_96[11:0] ? image_2573 : _GEN_8781; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8783 = 12'ha0e == _T_96[11:0] ? image_2574 : _GEN_8782; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8784 = 12'ha0f == _T_96[11:0] ? image_2575 : _GEN_8783; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8785 = 12'ha10 == _T_96[11:0] ? image_2576 : _GEN_8784; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8786 = 12'ha11 == _T_96[11:0] ? image_2577 : _GEN_8785; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8787 = 12'ha12 == _T_96[11:0] ? image_2578 : _GEN_8786; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8788 = 12'ha13 == _T_96[11:0] ? image_2579 : _GEN_8787; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8789 = 12'ha14 == _T_96[11:0] ? image_2580 : _GEN_8788; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8790 = 12'ha15 == _T_96[11:0] ? image_2581 : _GEN_8789; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8791 = 12'ha16 == _T_96[11:0] ? image_2582 : _GEN_8790; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8792 = 12'ha17 == _T_96[11:0] ? image_2583 : _GEN_8791; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8793 = 12'ha18 == _T_96[11:0] ? image_2584 : _GEN_8792; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8794 = 12'ha19 == _T_96[11:0] ? image_2585 : _GEN_8793; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8795 = 12'ha1a == _T_96[11:0] ? image_2586 : _GEN_8794; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8796 = 12'ha1b == _T_96[11:0] ? image_2587 : _GEN_8795; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8797 = 12'ha1c == _T_96[11:0] ? image_2588 : _GEN_8796; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8798 = 12'ha1d == _T_96[11:0] ? image_2589 : _GEN_8797; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8799 = 12'ha1e == _T_96[11:0] ? image_2590 : _GEN_8798; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8800 = 12'ha1f == _T_96[11:0] ? image_2591 : _GEN_8799; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8801 = 12'ha20 == _T_96[11:0] ? image_2592 : _GEN_8800; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8802 = 12'ha21 == _T_96[11:0] ? image_2593 : _GEN_8801; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8803 = 12'ha22 == _T_96[11:0] ? image_2594 : _GEN_8802; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8804 = 12'ha23 == _T_96[11:0] ? image_2595 : _GEN_8803; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8805 = 12'ha24 == _T_96[11:0] ? image_2596 : _GEN_8804; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8806 = 12'ha25 == _T_96[11:0] ? image_2597 : _GEN_8805; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8807 = 12'ha26 == _T_96[11:0] ? image_2598 : _GEN_8806; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8808 = 12'ha27 == _T_96[11:0] ? image_2599 : _GEN_8807; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8809 = 12'ha28 == _T_96[11:0] ? image_2600 : _GEN_8808; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8810 = 12'ha29 == _T_96[11:0] ? image_2601 : _GEN_8809; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8811 = 12'ha2a == _T_96[11:0] ? image_2602 : _GEN_8810; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8812 = 12'ha2b == _T_96[11:0] ? image_2603 : _GEN_8811; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8813 = 12'ha2c == _T_96[11:0] ? image_2604 : _GEN_8812; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8814 = 12'ha2d == _T_96[11:0] ? image_2605 : _GEN_8813; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8815 = 12'ha2e == _T_96[11:0] ? image_2606 : _GEN_8814; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8816 = 12'ha2f == _T_96[11:0] ? image_2607 : _GEN_8815; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8817 = 12'ha30 == _T_96[11:0] ? image_2608 : _GEN_8816; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8818 = 12'ha31 == _T_96[11:0] ? image_2609 : _GEN_8817; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8819 = 12'ha32 == _T_96[11:0] ? image_2610 : _GEN_8818; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8820 = 12'ha33 == _T_96[11:0] ? image_2611 : _GEN_8819; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8821 = 12'ha34 == _T_96[11:0] ? image_2612 : _GEN_8820; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8822 = 12'ha35 == _T_96[11:0] ? image_2613 : _GEN_8821; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8823 = 12'ha36 == _T_96[11:0] ? image_2614 : _GEN_8822; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8824 = 12'ha37 == _T_96[11:0] ? image_2615 : _GEN_8823; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8825 = 12'ha38 == _T_96[11:0] ? image_2616 : _GEN_8824; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8826 = 12'ha39 == _T_96[11:0] ? image_2617 : _GEN_8825; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8827 = 12'ha3a == _T_96[11:0] ? image_2618 : _GEN_8826; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8828 = 12'ha3b == _T_96[11:0] ? 4'h0 : _GEN_8827; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8829 = 12'ha3c == _T_96[11:0] ? 4'h0 : _GEN_8828; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8830 = 12'ha3d == _T_96[11:0] ? 4'h0 : _GEN_8829; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8831 = 12'ha3e == _T_96[11:0] ? 4'h0 : _GEN_8830; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8832 = 12'ha3f == _T_96[11:0] ? 4'h0 : _GEN_8831; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8833 = 12'ha40 == _T_96[11:0] ? 4'h0 : _GEN_8832; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8834 = 12'ha41 == _T_96[11:0] ? 4'h0 : _GEN_8833; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8835 = 12'ha42 == _T_96[11:0] ? 4'h0 : _GEN_8834; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8836 = 12'ha43 == _T_96[11:0] ? 4'h0 : _GEN_8835; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8837 = 12'ha44 == _T_96[11:0] ? 4'h0 : _GEN_8836; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8838 = 12'ha45 == _T_96[11:0] ? 4'h0 : _GEN_8837; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8839 = 12'ha46 == _T_96[11:0] ? 4'h0 : _GEN_8838; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8840 = 12'ha47 == _T_96[11:0] ? 4'h0 : _GEN_8839; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8841 = 12'ha48 == _T_96[11:0] ? image_2632 : _GEN_8840; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8842 = 12'ha49 == _T_96[11:0] ? image_2633 : _GEN_8841; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8843 = 12'ha4a == _T_96[11:0] ? image_2634 : _GEN_8842; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8844 = 12'ha4b == _T_96[11:0] ? image_2635 : _GEN_8843; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8845 = 12'ha4c == _T_96[11:0] ? image_2636 : _GEN_8844; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8846 = 12'ha4d == _T_96[11:0] ? image_2637 : _GEN_8845; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8847 = 12'ha4e == _T_96[11:0] ? image_2638 : _GEN_8846; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8848 = 12'ha4f == _T_96[11:0] ? image_2639 : _GEN_8847; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8849 = 12'ha50 == _T_96[11:0] ? image_2640 : _GEN_8848; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8850 = 12'ha51 == _T_96[11:0] ? image_2641 : _GEN_8849; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8851 = 12'ha52 == _T_96[11:0] ? image_2642 : _GEN_8850; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8852 = 12'ha53 == _T_96[11:0] ? image_2643 : _GEN_8851; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8853 = 12'ha54 == _T_96[11:0] ? image_2644 : _GEN_8852; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8854 = 12'ha55 == _T_96[11:0] ? image_2645 : _GEN_8853; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8855 = 12'ha56 == _T_96[11:0] ? image_2646 : _GEN_8854; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8856 = 12'ha57 == _T_96[11:0] ? image_2647 : _GEN_8855; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8857 = 12'ha58 == _T_96[11:0] ? image_2648 : _GEN_8856; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8858 = 12'ha59 == _T_96[11:0] ? image_2649 : _GEN_8857; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8859 = 12'ha5a == _T_96[11:0] ? image_2650 : _GEN_8858; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8860 = 12'ha5b == _T_96[11:0] ? image_2651 : _GEN_8859; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8861 = 12'ha5c == _T_96[11:0] ? image_2652 : _GEN_8860; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8862 = 12'ha5d == _T_96[11:0] ? image_2653 : _GEN_8861; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8863 = 12'ha5e == _T_96[11:0] ? image_2654 : _GEN_8862; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8864 = 12'ha5f == _T_96[11:0] ? image_2655 : _GEN_8863; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8865 = 12'ha60 == _T_96[11:0] ? image_2656 : _GEN_8864; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8866 = 12'ha61 == _T_96[11:0] ? image_2657 : _GEN_8865; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8867 = 12'ha62 == _T_96[11:0] ? image_2658 : _GEN_8866; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8868 = 12'ha63 == _T_96[11:0] ? image_2659 : _GEN_8867; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8869 = 12'ha64 == _T_96[11:0] ? image_2660 : _GEN_8868; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8870 = 12'ha65 == _T_96[11:0] ? image_2661 : _GEN_8869; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8871 = 12'ha66 == _T_96[11:0] ? image_2662 : _GEN_8870; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8872 = 12'ha67 == _T_96[11:0] ? image_2663 : _GEN_8871; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8873 = 12'ha68 == _T_96[11:0] ? image_2664 : _GEN_8872; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8874 = 12'ha69 == _T_96[11:0] ? image_2665 : _GEN_8873; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8875 = 12'ha6a == _T_96[11:0] ? image_2666 : _GEN_8874; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8876 = 12'ha6b == _T_96[11:0] ? image_2667 : _GEN_8875; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8877 = 12'ha6c == _T_96[11:0] ? image_2668 : _GEN_8876; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8878 = 12'ha6d == _T_96[11:0] ? image_2669 : _GEN_8877; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8879 = 12'ha6e == _T_96[11:0] ? image_2670 : _GEN_8878; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8880 = 12'ha6f == _T_96[11:0] ? image_2671 : _GEN_8879; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8881 = 12'ha70 == _T_96[11:0] ? image_2672 : _GEN_8880; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8882 = 12'ha71 == _T_96[11:0] ? image_2673 : _GEN_8881; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8883 = 12'ha72 == _T_96[11:0] ? image_2674 : _GEN_8882; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8884 = 12'ha73 == _T_96[11:0] ? image_2675 : _GEN_8883; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8885 = 12'ha74 == _T_96[11:0] ? image_2676 : _GEN_8884; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8886 = 12'ha75 == _T_96[11:0] ? image_2677 : _GEN_8885; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8887 = 12'ha76 == _T_96[11:0] ? image_2678 : _GEN_8886; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8888 = 12'ha77 == _T_96[11:0] ? image_2679 : _GEN_8887; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8889 = 12'ha78 == _T_96[11:0] ? image_2680 : _GEN_8888; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8890 = 12'ha79 == _T_96[11:0] ? image_2681 : _GEN_8889; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8891 = 12'ha7a == _T_96[11:0] ? image_2682 : _GEN_8890; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8892 = 12'ha7b == _T_96[11:0] ? 4'h0 : _GEN_8891; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8893 = 12'ha7c == _T_96[11:0] ? 4'h0 : _GEN_8892; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8894 = 12'ha7d == _T_96[11:0] ? 4'h0 : _GEN_8893; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8895 = 12'ha7e == _T_96[11:0] ? 4'h0 : _GEN_8894; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8896 = 12'ha7f == _T_96[11:0] ? 4'h0 : _GEN_8895; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8897 = 12'ha80 == _T_96[11:0] ? 4'h0 : _GEN_8896; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8898 = 12'ha81 == _T_96[11:0] ? 4'h0 : _GEN_8897; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8899 = 12'ha82 == _T_96[11:0] ? 4'h0 : _GEN_8898; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8900 = 12'ha83 == _T_96[11:0] ? 4'h0 : _GEN_8899; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8901 = 12'ha84 == _T_96[11:0] ? 4'h0 : _GEN_8900; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8902 = 12'ha85 == _T_96[11:0] ? 4'h0 : _GEN_8901; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8903 = 12'ha86 == _T_96[11:0] ? 4'h0 : _GEN_8902; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8904 = 12'ha87 == _T_96[11:0] ? 4'h0 : _GEN_8903; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8905 = 12'ha88 == _T_96[11:0] ? 4'h0 : _GEN_8904; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8906 = 12'ha89 == _T_96[11:0] ? image_2697 : _GEN_8905; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8907 = 12'ha8a == _T_96[11:0] ? image_2698 : _GEN_8906; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8908 = 12'ha8b == _T_96[11:0] ? image_2699 : _GEN_8907; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8909 = 12'ha8c == _T_96[11:0] ? image_2700 : _GEN_8908; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8910 = 12'ha8d == _T_96[11:0] ? image_2701 : _GEN_8909; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8911 = 12'ha8e == _T_96[11:0] ? image_2702 : _GEN_8910; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8912 = 12'ha8f == _T_96[11:0] ? image_2703 : _GEN_8911; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8913 = 12'ha90 == _T_96[11:0] ? image_2704 : _GEN_8912; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8914 = 12'ha91 == _T_96[11:0] ? image_2705 : _GEN_8913; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8915 = 12'ha92 == _T_96[11:0] ? image_2706 : _GEN_8914; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8916 = 12'ha93 == _T_96[11:0] ? image_2707 : _GEN_8915; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8917 = 12'ha94 == _T_96[11:0] ? image_2708 : _GEN_8916; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8918 = 12'ha95 == _T_96[11:0] ? image_2709 : _GEN_8917; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8919 = 12'ha96 == _T_96[11:0] ? image_2710 : _GEN_8918; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8920 = 12'ha97 == _T_96[11:0] ? image_2711 : _GEN_8919; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8921 = 12'ha98 == _T_96[11:0] ? image_2712 : _GEN_8920; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8922 = 12'ha99 == _T_96[11:0] ? image_2713 : _GEN_8921; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8923 = 12'ha9a == _T_96[11:0] ? image_2714 : _GEN_8922; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8924 = 12'ha9b == _T_96[11:0] ? image_2715 : _GEN_8923; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8925 = 12'ha9c == _T_96[11:0] ? image_2716 : _GEN_8924; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8926 = 12'ha9d == _T_96[11:0] ? image_2717 : _GEN_8925; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8927 = 12'ha9e == _T_96[11:0] ? image_2718 : _GEN_8926; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8928 = 12'ha9f == _T_96[11:0] ? image_2719 : _GEN_8927; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8929 = 12'haa0 == _T_96[11:0] ? image_2720 : _GEN_8928; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8930 = 12'haa1 == _T_96[11:0] ? image_2721 : _GEN_8929; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8931 = 12'haa2 == _T_96[11:0] ? image_2722 : _GEN_8930; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8932 = 12'haa3 == _T_96[11:0] ? image_2723 : _GEN_8931; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8933 = 12'haa4 == _T_96[11:0] ? image_2724 : _GEN_8932; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8934 = 12'haa5 == _T_96[11:0] ? image_2725 : _GEN_8933; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8935 = 12'haa6 == _T_96[11:0] ? image_2726 : _GEN_8934; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8936 = 12'haa7 == _T_96[11:0] ? image_2727 : _GEN_8935; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8937 = 12'haa8 == _T_96[11:0] ? image_2728 : _GEN_8936; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8938 = 12'haa9 == _T_96[11:0] ? image_2729 : _GEN_8937; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8939 = 12'haaa == _T_96[11:0] ? image_2730 : _GEN_8938; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8940 = 12'haab == _T_96[11:0] ? image_2731 : _GEN_8939; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8941 = 12'haac == _T_96[11:0] ? image_2732 : _GEN_8940; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8942 = 12'haad == _T_96[11:0] ? image_2733 : _GEN_8941; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8943 = 12'haae == _T_96[11:0] ? image_2734 : _GEN_8942; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8944 = 12'haaf == _T_96[11:0] ? image_2735 : _GEN_8943; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8945 = 12'hab0 == _T_96[11:0] ? image_2736 : _GEN_8944; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8946 = 12'hab1 == _T_96[11:0] ? image_2737 : _GEN_8945; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8947 = 12'hab2 == _T_96[11:0] ? image_2738 : _GEN_8946; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8948 = 12'hab3 == _T_96[11:0] ? image_2739 : _GEN_8947; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8949 = 12'hab4 == _T_96[11:0] ? image_2740 : _GEN_8948; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8950 = 12'hab5 == _T_96[11:0] ? image_2741 : _GEN_8949; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8951 = 12'hab6 == _T_96[11:0] ? image_2742 : _GEN_8950; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8952 = 12'hab7 == _T_96[11:0] ? image_2743 : _GEN_8951; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8953 = 12'hab8 == _T_96[11:0] ? image_2744 : _GEN_8952; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8954 = 12'hab9 == _T_96[11:0] ? image_2745 : _GEN_8953; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8955 = 12'haba == _T_96[11:0] ? 4'h0 : _GEN_8954; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8956 = 12'habb == _T_96[11:0] ? 4'h0 : _GEN_8955; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8957 = 12'habc == _T_96[11:0] ? 4'h0 : _GEN_8956; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8958 = 12'habd == _T_96[11:0] ? 4'h0 : _GEN_8957; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8959 = 12'habe == _T_96[11:0] ? 4'h0 : _GEN_8958; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8960 = 12'habf == _T_96[11:0] ? 4'h0 : _GEN_8959; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8961 = 12'hac0 == _T_96[11:0] ? 4'h0 : _GEN_8960; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8962 = 12'hac1 == _T_96[11:0] ? 4'h0 : _GEN_8961; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8963 = 12'hac2 == _T_96[11:0] ? 4'h0 : _GEN_8962; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8964 = 12'hac3 == _T_96[11:0] ? 4'h0 : _GEN_8963; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8965 = 12'hac4 == _T_96[11:0] ? 4'h0 : _GEN_8964; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8966 = 12'hac5 == _T_96[11:0] ? 4'h0 : _GEN_8965; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8967 = 12'hac6 == _T_96[11:0] ? 4'h0 : _GEN_8966; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8968 = 12'hac7 == _T_96[11:0] ? 4'h0 : _GEN_8967; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8969 = 12'hac8 == _T_96[11:0] ? 4'h0 : _GEN_8968; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8970 = 12'hac9 == _T_96[11:0] ? 4'h0 : _GEN_8969; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8971 = 12'haca == _T_96[11:0] ? 4'h0 : _GEN_8970; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8972 = 12'hacb == _T_96[11:0] ? image_2763 : _GEN_8971; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8973 = 12'hacc == _T_96[11:0] ? image_2764 : _GEN_8972; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8974 = 12'hacd == _T_96[11:0] ? image_2765 : _GEN_8973; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8975 = 12'hace == _T_96[11:0] ? image_2766 : _GEN_8974; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8976 = 12'hacf == _T_96[11:0] ? image_2767 : _GEN_8975; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8977 = 12'had0 == _T_96[11:0] ? image_2768 : _GEN_8976; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8978 = 12'had1 == _T_96[11:0] ? image_2769 : _GEN_8977; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8979 = 12'had2 == _T_96[11:0] ? image_2770 : _GEN_8978; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8980 = 12'had3 == _T_96[11:0] ? image_2771 : _GEN_8979; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8981 = 12'had4 == _T_96[11:0] ? image_2772 : _GEN_8980; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8982 = 12'had5 == _T_96[11:0] ? image_2773 : _GEN_8981; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8983 = 12'had6 == _T_96[11:0] ? image_2774 : _GEN_8982; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8984 = 12'had7 == _T_96[11:0] ? image_2775 : _GEN_8983; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8985 = 12'had8 == _T_96[11:0] ? image_2776 : _GEN_8984; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8986 = 12'had9 == _T_96[11:0] ? image_2777 : _GEN_8985; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8987 = 12'hada == _T_96[11:0] ? image_2778 : _GEN_8986; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8988 = 12'hadb == _T_96[11:0] ? image_2779 : _GEN_8987; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8989 = 12'hadc == _T_96[11:0] ? image_2780 : _GEN_8988; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8990 = 12'hadd == _T_96[11:0] ? image_2781 : _GEN_8989; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8991 = 12'hade == _T_96[11:0] ? image_2782 : _GEN_8990; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8992 = 12'hadf == _T_96[11:0] ? image_2783 : _GEN_8991; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8993 = 12'hae0 == _T_96[11:0] ? image_2784 : _GEN_8992; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8994 = 12'hae1 == _T_96[11:0] ? image_2785 : _GEN_8993; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8995 = 12'hae2 == _T_96[11:0] ? image_2786 : _GEN_8994; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8996 = 12'hae3 == _T_96[11:0] ? image_2787 : _GEN_8995; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8997 = 12'hae4 == _T_96[11:0] ? image_2788 : _GEN_8996; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8998 = 12'hae5 == _T_96[11:0] ? image_2789 : _GEN_8997; // @[Filter.scala 138:46]
  wire [3:0] _GEN_8999 = 12'hae6 == _T_96[11:0] ? image_2790 : _GEN_8998; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9000 = 12'hae7 == _T_96[11:0] ? image_2791 : _GEN_8999; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9001 = 12'hae8 == _T_96[11:0] ? image_2792 : _GEN_9000; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9002 = 12'hae9 == _T_96[11:0] ? image_2793 : _GEN_9001; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9003 = 12'haea == _T_96[11:0] ? image_2794 : _GEN_9002; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9004 = 12'haeb == _T_96[11:0] ? image_2795 : _GEN_9003; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9005 = 12'haec == _T_96[11:0] ? image_2796 : _GEN_9004; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9006 = 12'haed == _T_96[11:0] ? image_2797 : _GEN_9005; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9007 = 12'haee == _T_96[11:0] ? image_2798 : _GEN_9006; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9008 = 12'haef == _T_96[11:0] ? image_2799 : _GEN_9007; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9009 = 12'haf0 == _T_96[11:0] ? image_2800 : _GEN_9008; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9010 = 12'haf1 == _T_96[11:0] ? image_2801 : _GEN_9009; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9011 = 12'haf2 == _T_96[11:0] ? image_2802 : _GEN_9010; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9012 = 12'haf3 == _T_96[11:0] ? image_2803 : _GEN_9011; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9013 = 12'haf4 == _T_96[11:0] ? image_2804 : _GEN_9012; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9014 = 12'haf5 == _T_96[11:0] ? image_2805 : _GEN_9013; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9015 = 12'haf6 == _T_96[11:0] ? image_2806 : _GEN_9014; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9016 = 12'haf7 == _T_96[11:0] ? image_2807 : _GEN_9015; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9017 = 12'haf8 == _T_96[11:0] ? image_2808 : _GEN_9016; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9018 = 12'haf9 == _T_96[11:0] ? 4'h0 : _GEN_9017; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9019 = 12'hafa == _T_96[11:0] ? 4'h0 : _GEN_9018; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9020 = 12'hafb == _T_96[11:0] ? 4'h0 : _GEN_9019; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9021 = 12'hafc == _T_96[11:0] ? 4'h0 : _GEN_9020; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9022 = 12'hafd == _T_96[11:0] ? 4'h0 : _GEN_9021; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9023 = 12'hafe == _T_96[11:0] ? 4'h0 : _GEN_9022; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9024 = 12'haff == _T_96[11:0] ? 4'h0 : _GEN_9023; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9025 = 12'hb00 == _T_96[11:0] ? 4'h0 : _GEN_9024; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9026 = 12'hb01 == _T_96[11:0] ? 4'h0 : _GEN_9025; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9027 = 12'hb02 == _T_96[11:0] ? 4'h0 : _GEN_9026; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9028 = 12'hb03 == _T_96[11:0] ? 4'h0 : _GEN_9027; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9029 = 12'hb04 == _T_96[11:0] ? 4'h0 : _GEN_9028; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9030 = 12'hb05 == _T_96[11:0] ? 4'h0 : _GEN_9029; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9031 = 12'hb06 == _T_96[11:0] ? 4'h0 : _GEN_9030; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9032 = 12'hb07 == _T_96[11:0] ? 4'h0 : _GEN_9031; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9033 = 12'hb08 == _T_96[11:0] ? 4'h0 : _GEN_9032; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9034 = 12'hb09 == _T_96[11:0] ? 4'h0 : _GEN_9033; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9035 = 12'hb0a == _T_96[11:0] ? 4'h0 : _GEN_9034; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9036 = 12'hb0b == _T_96[11:0] ? 4'h0 : _GEN_9035; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9037 = 12'hb0c == _T_96[11:0] ? image_2828 : _GEN_9036; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9038 = 12'hb0d == _T_96[11:0] ? image_2829 : _GEN_9037; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9039 = 12'hb0e == _T_96[11:0] ? image_2830 : _GEN_9038; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9040 = 12'hb0f == _T_96[11:0] ? image_2831 : _GEN_9039; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9041 = 12'hb10 == _T_96[11:0] ? image_2832 : _GEN_9040; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9042 = 12'hb11 == _T_96[11:0] ? image_2833 : _GEN_9041; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9043 = 12'hb12 == _T_96[11:0] ? image_2834 : _GEN_9042; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9044 = 12'hb13 == _T_96[11:0] ? image_2835 : _GEN_9043; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9045 = 12'hb14 == _T_96[11:0] ? image_2836 : _GEN_9044; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9046 = 12'hb15 == _T_96[11:0] ? image_2837 : _GEN_9045; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9047 = 12'hb16 == _T_96[11:0] ? image_2838 : _GEN_9046; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9048 = 12'hb17 == _T_96[11:0] ? image_2839 : _GEN_9047; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9049 = 12'hb18 == _T_96[11:0] ? image_2840 : _GEN_9048; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9050 = 12'hb19 == _T_96[11:0] ? image_2841 : _GEN_9049; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9051 = 12'hb1a == _T_96[11:0] ? image_2842 : _GEN_9050; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9052 = 12'hb1b == _T_96[11:0] ? image_2843 : _GEN_9051; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9053 = 12'hb1c == _T_96[11:0] ? image_2844 : _GEN_9052; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9054 = 12'hb1d == _T_96[11:0] ? image_2845 : _GEN_9053; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9055 = 12'hb1e == _T_96[11:0] ? image_2846 : _GEN_9054; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9056 = 12'hb1f == _T_96[11:0] ? image_2847 : _GEN_9055; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9057 = 12'hb20 == _T_96[11:0] ? image_2848 : _GEN_9056; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9058 = 12'hb21 == _T_96[11:0] ? image_2849 : _GEN_9057; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9059 = 12'hb22 == _T_96[11:0] ? image_2850 : _GEN_9058; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9060 = 12'hb23 == _T_96[11:0] ? image_2851 : _GEN_9059; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9061 = 12'hb24 == _T_96[11:0] ? image_2852 : _GEN_9060; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9062 = 12'hb25 == _T_96[11:0] ? image_2853 : _GEN_9061; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9063 = 12'hb26 == _T_96[11:0] ? image_2854 : _GEN_9062; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9064 = 12'hb27 == _T_96[11:0] ? image_2855 : _GEN_9063; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9065 = 12'hb28 == _T_96[11:0] ? image_2856 : _GEN_9064; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9066 = 12'hb29 == _T_96[11:0] ? image_2857 : _GEN_9065; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9067 = 12'hb2a == _T_96[11:0] ? image_2858 : _GEN_9066; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9068 = 12'hb2b == _T_96[11:0] ? image_2859 : _GEN_9067; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9069 = 12'hb2c == _T_96[11:0] ? image_2860 : _GEN_9068; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9070 = 12'hb2d == _T_96[11:0] ? image_2861 : _GEN_9069; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9071 = 12'hb2e == _T_96[11:0] ? image_2862 : _GEN_9070; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9072 = 12'hb2f == _T_96[11:0] ? image_2863 : _GEN_9071; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9073 = 12'hb30 == _T_96[11:0] ? image_2864 : _GEN_9072; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9074 = 12'hb31 == _T_96[11:0] ? image_2865 : _GEN_9073; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9075 = 12'hb32 == _T_96[11:0] ? image_2866 : _GEN_9074; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9076 = 12'hb33 == _T_96[11:0] ? image_2867 : _GEN_9075; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9077 = 12'hb34 == _T_96[11:0] ? image_2868 : _GEN_9076; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9078 = 12'hb35 == _T_96[11:0] ? image_2869 : _GEN_9077; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9079 = 12'hb36 == _T_96[11:0] ? image_2870 : _GEN_9078; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9080 = 12'hb37 == _T_96[11:0] ? image_2871 : _GEN_9079; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9081 = 12'hb38 == _T_96[11:0] ? 4'h0 : _GEN_9080; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9082 = 12'hb39 == _T_96[11:0] ? 4'h0 : _GEN_9081; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9083 = 12'hb3a == _T_96[11:0] ? 4'h0 : _GEN_9082; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9084 = 12'hb3b == _T_96[11:0] ? 4'h0 : _GEN_9083; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9085 = 12'hb3c == _T_96[11:0] ? 4'h0 : _GEN_9084; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9086 = 12'hb3d == _T_96[11:0] ? 4'h0 : _GEN_9085; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9087 = 12'hb3e == _T_96[11:0] ? 4'h0 : _GEN_9086; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9088 = 12'hb3f == _T_96[11:0] ? 4'h0 : _GEN_9087; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9089 = 12'hb40 == _T_96[11:0] ? 4'h0 : _GEN_9088; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9090 = 12'hb41 == _T_96[11:0] ? 4'h0 : _GEN_9089; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9091 = 12'hb42 == _T_96[11:0] ? 4'h0 : _GEN_9090; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9092 = 12'hb43 == _T_96[11:0] ? 4'h0 : _GEN_9091; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9093 = 12'hb44 == _T_96[11:0] ? 4'h0 : _GEN_9092; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9094 = 12'hb45 == _T_96[11:0] ? 4'h0 : _GEN_9093; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9095 = 12'hb46 == _T_96[11:0] ? 4'h0 : _GEN_9094; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9096 = 12'hb47 == _T_96[11:0] ? 4'h0 : _GEN_9095; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9097 = 12'hb48 == _T_96[11:0] ? 4'h0 : _GEN_9096; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9098 = 12'hb49 == _T_96[11:0] ? 4'h0 : _GEN_9097; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9099 = 12'hb4a == _T_96[11:0] ? 4'h0 : _GEN_9098; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9100 = 12'hb4b == _T_96[11:0] ? 4'h0 : _GEN_9099; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9101 = 12'hb4c == _T_96[11:0] ? 4'h0 : _GEN_9100; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9102 = 12'hb4d == _T_96[11:0] ? 4'h0 : _GEN_9101; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9103 = 12'hb4e == _T_96[11:0] ? 4'h0 : _GEN_9102; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9104 = 12'hb4f == _T_96[11:0] ? image_2895 : _GEN_9103; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9105 = 12'hb50 == _T_96[11:0] ? image_2896 : _GEN_9104; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9106 = 12'hb51 == _T_96[11:0] ? image_2897 : _GEN_9105; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9107 = 12'hb52 == _T_96[11:0] ? image_2898 : _GEN_9106; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9108 = 12'hb53 == _T_96[11:0] ? image_2899 : _GEN_9107; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9109 = 12'hb54 == _T_96[11:0] ? image_2900 : _GEN_9108; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9110 = 12'hb55 == _T_96[11:0] ? image_2901 : _GEN_9109; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9111 = 12'hb56 == _T_96[11:0] ? image_2902 : _GEN_9110; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9112 = 12'hb57 == _T_96[11:0] ? image_2903 : _GEN_9111; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9113 = 12'hb58 == _T_96[11:0] ? image_2904 : _GEN_9112; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9114 = 12'hb59 == _T_96[11:0] ? image_2905 : _GEN_9113; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9115 = 12'hb5a == _T_96[11:0] ? image_2906 : _GEN_9114; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9116 = 12'hb5b == _T_96[11:0] ? image_2907 : _GEN_9115; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9117 = 12'hb5c == _T_96[11:0] ? image_2908 : _GEN_9116; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9118 = 12'hb5d == _T_96[11:0] ? image_2909 : _GEN_9117; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9119 = 12'hb5e == _T_96[11:0] ? image_2910 : _GEN_9118; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9120 = 12'hb5f == _T_96[11:0] ? image_2911 : _GEN_9119; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9121 = 12'hb60 == _T_96[11:0] ? image_2912 : _GEN_9120; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9122 = 12'hb61 == _T_96[11:0] ? image_2913 : _GEN_9121; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9123 = 12'hb62 == _T_96[11:0] ? image_2914 : _GEN_9122; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9124 = 12'hb63 == _T_96[11:0] ? image_2915 : _GEN_9123; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9125 = 12'hb64 == _T_96[11:0] ? image_2916 : _GEN_9124; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9126 = 12'hb65 == _T_96[11:0] ? image_2917 : _GEN_9125; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9127 = 12'hb66 == _T_96[11:0] ? image_2918 : _GEN_9126; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9128 = 12'hb67 == _T_96[11:0] ? image_2919 : _GEN_9127; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9129 = 12'hb68 == _T_96[11:0] ? image_2920 : _GEN_9128; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9130 = 12'hb69 == _T_96[11:0] ? image_2921 : _GEN_9129; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9131 = 12'hb6a == _T_96[11:0] ? image_2922 : _GEN_9130; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9132 = 12'hb6b == _T_96[11:0] ? image_2923 : _GEN_9131; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9133 = 12'hb6c == _T_96[11:0] ? image_2924 : _GEN_9132; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9134 = 12'hb6d == _T_96[11:0] ? image_2925 : _GEN_9133; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9135 = 12'hb6e == _T_96[11:0] ? image_2926 : _GEN_9134; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9136 = 12'hb6f == _T_96[11:0] ? image_2927 : _GEN_9135; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9137 = 12'hb70 == _T_96[11:0] ? image_2928 : _GEN_9136; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9138 = 12'hb71 == _T_96[11:0] ? image_2929 : _GEN_9137; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9139 = 12'hb72 == _T_96[11:0] ? image_2930 : _GEN_9138; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9140 = 12'hb73 == _T_96[11:0] ? image_2931 : _GEN_9139; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9141 = 12'hb74 == _T_96[11:0] ? image_2932 : _GEN_9140; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9142 = 12'hb75 == _T_96[11:0] ? image_2933 : _GEN_9141; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9143 = 12'hb76 == _T_96[11:0] ? image_2934 : _GEN_9142; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9144 = 12'hb77 == _T_96[11:0] ? 4'h0 : _GEN_9143; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9145 = 12'hb78 == _T_96[11:0] ? 4'h0 : _GEN_9144; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9146 = 12'hb79 == _T_96[11:0] ? 4'h0 : _GEN_9145; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9147 = 12'hb7a == _T_96[11:0] ? 4'h0 : _GEN_9146; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9148 = 12'hb7b == _T_96[11:0] ? 4'h0 : _GEN_9147; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9149 = 12'hb7c == _T_96[11:0] ? 4'h0 : _GEN_9148; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9150 = 12'hb7d == _T_96[11:0] ? 4'h0 : _GEN_9149; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9151 = 12'hb7e == _T_96[11:0] ? 4'h0 : _GEN_9150; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9152 = 12'hb7f == _T_96[11:0] ? 4'h0 : _GEN_9151; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9153 = 12'hb80 == _T_96[11:0] ? 4'h0 : _GEN_9152; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9154 = 12'hb81 == _T_96[11:0] ? 4'h0 : _GEN_9153; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9155 = 12'hb82 == _T_96[11:0] ? 4'h0 : _GEN_9154; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9156 = 12'hb83 == _T_96[11:0] ? 4'h0 : _GEN_9155; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9157 = 12'hb84 == _T_96[11:0] ? 4'h0 : _GEN_9156; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9158 = 12'hb85 == _T_96[11:0] ? 4'h0 : _GEN_9157; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9159 = 12'hb86 == _T_96[11:0] ? 4'h0 : _GEN_9158; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9160 = 12'hb87 == _T_96[11:0] ? 4'h0 : _GEN_9159; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9161 = 12'hb88 == _T_96[11:0] ? 4'h0 : _GEN_9160; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9162 = 12'hb89 == _T_96[11:0] ? 4'h0 : _GEN_9161; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9163 = 12'hb8a == _T_96[11:0] ? 4'h0 : _GEN_9162; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9164 = 12'hb8b == _T_96[11:0] ? 4'h0 : _GEN_9163; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9165 = 12'hb8c == _T_96[11:0] ? 4'h0 : _GEN_9164; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9166 = 12'hb8d == _T_96[11:0] ? 4'h0 : _GEN_9165; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9167 = 12'hb8e == _T_96[11:0] ? 4'h0 : _GEN_9166; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9168 = 12'hb8f == _T_96[11:0] ? 4'h0 : _GEN_9167; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9169 = 12'hb90 == _T_96[11:0] ? 4'h0 : _GEN_9168; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9170 = 12'hb91 == _T_96[11:0] ? 4'h0 : _GEN_9169; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9171 = 12'hb92 == _T_96[11:0] ? 4'h0 : _GEN_9170; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9172 = 12'hb93 == _T_96[11:0] ? 4'h0 : _GEN_9171; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9173 = 12'hb94 == _T_96[11:0] ? 4'h0 : _GEN_9172; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9174 = 12'hb95 == _T_96[11:0] ? image_2965 : _GEN_9173; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9175 = 12'hb96 == _T_96[11:0] ? image_2966 : _GEN_9174; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9176 = 12'hb97 == _T_96[11:0] ? image_2967 : _GEN_9175; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9177 = 12'hb98 == _T_96[11:0] ? image_2968 : _GEN_9176; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9178 = 12'hb99 == _T_96[11:0] ? image_2969 : _GEN_9177; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9179 = 12'hb9a == _T_96[11:0] ? image_2970 : _GEN_9178; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9180 = 12'hb9b == _T_96[11:0] ? image_2971 : _GEN_9179; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9181 = 12'hb9c == _T_96[11:0] ? image_2972 : _GEN_9180; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9182 = 12'hb9d == _T_96[11:0] ? image_2973 : _GEN_9181; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9183 = 12'hb9e == _T_96[11:0] ? image_2974 : _GEN_9182; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9184 = 12'hb9f == _T_96[11:0] ? image_2975 : _GEN_9183; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9185 = 12'hba0 == _T_96[11:0] ? image_2976 : _GEN_9184; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9186 = 12'hba1 == _T_96[11:0] ? image_2977 : _GEN_9185; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9187 = 12'hba2 == _T_96[11:0] ? image_2978 : _GEN_9186; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9188 = 12'hba3 == _T_96[11:0] ? image_2979 : _GEN_9187; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9189 = 12'hba4 == _T_96[11:0] ? image_2980 : _GEN_9188; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9190 = 12'hba5 == _T_96[11:0] ? image_2981 : _GEN_9189; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9191 = 12'hba6 == _T_96[11:0] ? image_2982 : _GEN_9190; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9192 = 12'hba7 == _T_96[11:0] ? image_2983 : _GEN_9191; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9193 = 12'hba8 == _T_96[11:0] ? image_2984 : _GEN_9192; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9194 = 12'hba9 == _T_96[11:0] ? image_2985 : _GEN_9193; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9195 = 12'hbaa == _T_96[11:0] ? image_2986 : _GEN_9194; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9196 = 12'hbab == _T_96[11:0] ? image_2987 : _GEN_9195; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9197 = 12'hbac == _T_96[11:0] ? image_2988 : _GEN_9196; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9198 = 12'hbad == _T_96[11:0] ? image_2989 : _GEN_9197; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9199 = 12'hbae == _T_96[11:0] ? image_2990 : _GEN_9198; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9200 = 12'hbaf == _T_96[11:0] ? image_2991 : _GEN_9199; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9201 = 12'hbb0 == _T_96[11:0] ? image_2992 : _GEN_9200; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9202 = 12'hbb1 == _T_96[11:0] ? image_2993 : _GEN_9201; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9203 = 12'hbb2 == _T_96[11:0] ? image_2994 : _GEN_9202; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9204 = 12'hbb3 == _T_96[11:0] ? image_2995 : _GEN_9203; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9205 = 12'hbb4 == _T_96[11:0] ? image_2996 : _GEN_9204; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9206 = 12'hbb5 == _T_96[11:0] ? 4'h0 : _GEN_9205; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9207 = 12'hbb6 == _T_96[11:0] ? 4'h0 : _GEN_9206; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9208 = 12'hbb7 == _T_96[11:0] ? 4'h0 : _GEN_9207; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9209 = 12'hbb8 == _T_96[11:0] ? 4'h0 : _GEN_9208; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9210 = 12'hbb9 == _T_96[11:0] ? 4'h0 : _GEN_9209; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9211 = 12'hbba == _T_96[11:0] ? 4'h0 : _GEN_9210; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9212 = 12'hbbb == _T_96[11:0] ? 4'h0 : _GEN_9211; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9213 = 12'hbbc == _T_96[11:0] ? 4'h0 : _GEN_9212; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9214 = 12'hbbd == _T_96[11:0] ? 4'h0 : _GEN_9213; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9215 = 12'hbbe == _T_96[11:0] ? 4'h0 : _GEN_9214; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9216 = 12'hbbf == _T_96[11:0] ? 4'h0 : _GEN_9215; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9217 = 12'hbc0 == _T_96[11:0] ? 4'h0 : _GEN_9216; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9218 = 12'hbc1 == _T_96[11:0] ? 4'h0 : _GEN_9217; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9219 = 12'hbc2 == _T_96[11:0] ? 4'h0 : _GEN_9218; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9220 = 12'hbc3 == _T_96[11:0] ? 4'h0 : _GEN_9219; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9221 = 12'hbc4 == _T_96[11:0] ? 4'h0 : _GEN_9220; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9222 = 12'hbc5 == _T_96[11:0] ? 4'h0 : _GEN_9221; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9223 = 12'hbc6 == _T_96[11:0] ? 4'h0 : _GEN_9222; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9224 = 12'hbc7 == _T_96[11:0] ? 4'h0 : _GEN_9223; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9225 = 12'hbc8 == _T_96[11:0] ? 4'h0 : _GEN_9224; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9226 = 12'hbc9 == _T_96[11:0] ? 4'h0 : _GEN_9225; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9227 = 12'hbca == _T_96[11:0] ? 4'h0 : _GEN_9226; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9228 = 12'hbcb == _T_96[11:0] ? 4'h0 : _GEN_9227; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9229 = 12'hbcc == _T_96[11:0] ? 4'h0 : _GEN_9228; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9230 = 12'hbcd == _T_96[11:0] ? 4'h0 : _GEN_9229; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9231 = 12'hbce == _T_96[11:0] ? 4'h0 : _GEN_9230; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9232 = 12'hbcf == _T_96[11:0] ? 4'h0 : _GEN_9231; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9233 = 12'hbd0 == _T_96[11:0] ? 4'h0 : _GEN_9232; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9234 = 12'hbd1 == _T_96[11:0] ? 4'h0 : _GEN_9233; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9235 = 12'hbd2 == _T_96[11:0] ? 4'h0 : _GEN_9234; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9236 = 12'hbd3 == _T_96[11:0] ? 4'h0 : _GEN_9235; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9237 = 12'hbd4 == _T_96[11:0] ? 4'h0 : _GEN_9236; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9238 = 12'hbd5 == _T_96[11:0] ? 4'h0 : _GEN_9237; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9239 = 12'hbd6 == _T_96[11:0] ? 4'h0 : _GEN_9238; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9240 = 12'hbd7 == _T_96[11:0] ? 4'h0 : _GEN_9239; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9241 = 12'hbd8 == _T_96[11:0] ? 4'h0 : _GEN_9240; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9242 = 12'hbd9 == _T_96[11:0] ? 4'h0 : _GEN_9241; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9243 = 12'hbda == _T_96[11:0] ? 4'h0 : _GEN_9242; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9244 = 12'hbdb == _T_96[11:0] ? image_3035 : _GEN_9243; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9245 = 12'hbdc == _T_96[11:0] ? image_3036 : _GEN_9244; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9246 = 12'hbdd == _T_96[11:0] ? image_3037 : _GEN_9245; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9247 = 12'hbde == _T_96[11:0] ? image_3038 : _GEN_9246; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9248 = 12'hbdf == _T_96[11:0] ? image_3039 : _GEN_9247; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9249 = 12'hbe0 == _T_96[11:0] ? image_3040 : _GEN_9248; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9250 = 12'hbe1 == _T_96[11:0] ? image_3041 : _GEN_9249; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9251 = 12'hbe2 == _T_96[11:0] ? image_3042 : _GEN_9250; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9252 = 12'hbe3 == _T_96[11:0] ? image_3043 : _GEN_9251; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9253 = 12'hbe4 == _T_96[11:0] ? image_3044 : _GEN_9252; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9254 = 12'hbe5 == _T_96[11:0] ? image_3045 : _GEN_9253; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9255 = 12'hbe6 == _T_96[11:0] ? image_3046 : _GEN_9254; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9256 = 12'hbe7 == _T_96[11:0] ? image_3047 : _GEN_9255; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9257 = 12'hbe8 == _T_96[11:0] ? image_3048 : _GEN_9256; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9258 = 12'hbe9 == _T_96[11:0] ? image_3049 : _GEN_9257; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9259 = 12'hbea == _T_96[11:0] ? image_3050 : _GEN_9258; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9260 = 12'hbeb == _T_96[11:0] ? image_3051 : _GEN_9259; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9261 = 12'hbec == _T_96[11:0] ? image_3052 : _GEN_9260; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9262 = 12'hbed == _T_96[11:0] ? image_3053 : _GEN_9261; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9263 = 12'hbee == _T_96[11:0] ? image_3054 : _GEN_9262; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9264 = 12'hbef == _T_96[11:0] ? image_3055 : _GEN_9263; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9265 = 12'hbf0 == _T_96[11:0] ? image_3056 : _GEN_9264; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9266 = 12'hbf1 == _T_96[11:0] ? 4'h0 : _GEN_9265; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9267 = 12'hbf2 == _T_96[11:0] ? 4'h0 : _GEN_9266; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9268 = 12'hbf3 == _T_96[11:0] ? 4'h0 : _GEN_9267; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9269 = 12'hbf4 == _T_96[11:0] ? 4'h0 : _GEN_9268; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9270 = 12'hbf5 == _T_96[11:0] ? 4'h0 : _GEN_9269; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9271 = 12'hbf6 == _T_96[11:0] ? 4'h0 : _GEN_9270; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9272 = 12'hbf7 == _T_96[11:0] ? 4'h0 : _GEN_9271; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9273 = 12'hbf8 == _T_96[11:0] ? 4'h0 : _GEN_9272; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9274 = 12'hbf9 == _T_96[11:0] ? 4'h0 : _GEN_9273; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9275 = 12'hbfa == _T_96[11:0] ? 4'h0 : _GEN_9274; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9276 = 12'hbfb == _T_96[11:0] ? 4'h0 : _GEN_9275; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9277 = 12'hbfc == _T_96[11:0] ? 4'h0 : _GEN_9276; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9278 = 12'hbfd == _T_96[11:0] ? 4'h0 : _GEN_9277; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9279 = 12'hbfe == _T_96[11:0] ? 4'h0 : _GEN_9278; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9280 = 12'hbff == _T_96[11:0] ? 4'h0 : _GEN_9279; // @[Filter.scala 138:46]
  wire [31:0] _T_99 = pixelIndex + 32'h3; // @[Filter.scala 133:29]
  wire [31:0] _T_100 = _T_99 / 32'h40; // @[Filter.scala 133:36]
  wire [31:0] _T_102 = _T_100 + _GEN_24805; // @[Filter.scala 133:51]
  wire [31:0] _T_104 = _T_102 - 32'h1; // @[Filter.scala 133:67]
  wire [31:0] _GEN_3 = _T_99 % 32'h40; // @[Filter.scala 134:36]
  wire [6:0] _T_107 = _GEN_3[6:0]; // @[Filter.scala 134:36]
  wire [6:0] _T_109 = _T_107 + _GEN_24806; // @[Filter.scala 134:51]
  wire [6:0] _T_111 = _T_109 - 7'h1; // @[Filter.scala 134:67]
  wire  _T_113 = _T_104 >= 32'h40; // @[Filter.scala 135:27]
  wire  _T_117 = _T_111 >= 7'h30; // @[Filter.scala 135:59]
  wire  _T_118 = _T_113 | _T_117; // @[Filter.scala 135:54]
  wire [13:0] _T_119 = _T_111 * 7'h40; // @[Filter.scala 138:57]
  wire [31:0] _GEN_24816 = {{18'd0}, _T_119}; // @[Filter.scala 138:72]
  wire [31:0] _T_121 = _GEN_24816 + _T_104; // @[Filter.scala 138:72]
  wire [3:0] _GEN_9294 = 12'hc == _T_121[11:0] ? image_12 : 4'h0; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9295 = 12'hd == _T_121[11:0] ? 4'h0 : _GEN_9294; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9296 = 12'he == _T_121[11:0] ? image_14 : _GEN_9295; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9297 = 12'hf == _T_121[11:0] ? image_15 : _GEN_9296; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9298 = 12'h10 == _T_121[11:0] ? image_16 : _GEN_9297; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9299 = 12'h11 == _T_121[11:0] ? image_17 : _GEN_9298; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9300 = 12'h12 == _T_121[11:0] ? image_18 : _GEN_9299; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9301 = 12'h13 == _T_121[11:0] ? image_19 : _GEN_9300; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9302 = 12'h14 == _T_121[11:0] ? image_20 : _GEN_9301; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9303 = 12'h15 == _T_121[11:0] ? image_21 : _GEN_9302; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9304 = 12'h16 == _T_121[11:0] ? image_22 : _GEN_9303; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9305 = 12'h17 == _T_121[11:0] ? image_23 : _GEN_9304; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9306 = 12'h18 == _T_121[11:0] ? 4'h0 : _GEN_9305; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9307 = 12'h19 == _T_121[11:0] ? 4'h0 : _GEN_9306; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9308 = 12'h1a == _T_121[11:0] ? 4'h0 : _GEN_9307; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9309 = 12'h1b == _T_121[11:0] ? 4'h0 : _GEN_9308; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9310 = 12'h1c == _T_121[11:0] ? 4'h0 : _GEN_9309; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9311 = 12'h1d == _T_121[11:0] ? 4'h0 : _GEN_9310; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9312 = 12'h1e == _T_121[11:0] ? 4'h0 : _GEN_9311; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9313 = 12'h1f == _T_121[11:0] ? 4'h0 : _GEN_9312; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9314 = 12'h20 == _T_121[11:0] ? 4'h0 : _GEN_9313; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9315 = 12'h21 == _T_121[11:0] ? 4'h0 : _GEN_9314; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9316 = 12'h22 == _T_121[11:0] ? 4'h0 : _GEN_9315; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9317 = 12'h23 == _T_121[11:0] ? image_35 : _GEN_9316; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9318 = 12'h24 == _T_121[11:0] ? image_36 : _GEN_9317; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9319 = 12'h25 == _T_121[11:0] ? image_37 : _GEN_9318; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9320 = 12'h26 == _T_121[11:0] ? image_38 : _GEN_9319; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9321 = 12'h27 == _T_121[11:0] ? image_39 : _GEN_9320; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9322 = 12'h28 == _T_121[11:0] ? image_40 : _GEN_9321; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9323 = 12'h29 == _T_121[11:0] ? image_41 : _GEN_9322; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9324 = 12'h2a == _T_121[11:0] ? image_42 : _GEN_9323; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9325 = 12'h2b == _T_121[11:0] ? 4'h0 : _GEN_9324; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9326 = 12'h2c == _T_121[11:0] ? 4'h0 : _GEN_9325; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9327 = 12'h2d == _T_121[11:0] ? 4'h0 : _GEN_9326; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9328 = 12'h2e == _T_121[11:0] ? 4'h0 : _GEN_9327; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9329 = 12'h2f == _T_121[11:0] ? 4'h0 : _GEN_9328; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9330 = 12'h30 == _T_121[11:0] ? 4'h0 : _GEN_9329; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9331 = 12'h31 == _T_121[11:0] ? 4'h0 : _GEN_9330; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9332 = 12'h32 == _T_121[11:0] ? 4'h0 : _GEN_9331; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9333 = 12'h33 == _T_121[11:0] ? 4'h0 : _GEN_9332; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9334 = 12'h34 == _T_121[11:0] ? 4'h0 : _GEN_9333; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9335 = 12'h35 == _T_121[11:0] ? 4'h0 : _GEN_9334; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9336 = 12'h36 == _T_121[11:0] ? 4'h0 : _GEN_9335; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9337 = 12'h37 == _T_121[11:0] ? 4'h0 : _GEN_9336; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9338 = 12'h38 == _T_121[11:0] ? 4'h0 : _GEN_9337; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9339 = 12'h39 == _T_121[11:0] ? 4'h0 : _GEN_9338; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9340 = 12'h3a == _T_121[11:0] ? 4'h0 : _GEN_9339; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9341 = 12'h3b == _T_121[11:0] ? 4'h0 : _GEN_9340; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9342 = 12'h3c == _T_121[11:0] ? 4'h0 : _GEN_9341; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9343 = 12'h3d == _T_121[11:0] ? 4'h0 : _GEN_9342; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9344 = 12'h3e == _T_121[11:0] ? 4'h0 : _GEN_9343; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9345 = 12'h3f == _T_121[11:0] ? 4'h0 : _GEN_9344; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9346 = 12'h40 == _T_121[11:0] ? 4'h0 : _GEN_9345; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9347 = 12'h41 == _T_121[11:0] ? 4'h0 : _GEN_9346; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9348 = 12'h42 == _T_121[11:0] ? 4'h0 : _GEN_9347; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9349 = 12'h43 == _T_121[11:0] ? 4'h0 : _GEN_9348; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9350 = 12'h44 == _T_121[11:0] ? 4'h0 : _GEN_9349; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9351 = 12'h45 == _T_121[11:0] ? 4'h0 : _GEN_9350; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9352 = 12'h46 == _T_121[11:0] ? 4'h0 : _GEN_9351; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9353 = 12'h47 == _T_121[11:0] ? 4'h0 : _GEN_9352; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9354 = 12'h48 == _T_121[11:0] ? 4'h0 : _GEN_9353; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9355 = 12'h49 == _T_121[11:0] ? 4'h0 : _GEN_9354; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9356 = 12'h4a == _T_121[11:0] ? 4'h0 : _GEN_9355; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9357 = 12'h4b == _T_121[11:0] ? image_75 : _GEN_9356; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9358 = 12'h4c == _T_121[11:0] ? image_76 : _GEN_9357; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9359 = 12'h4d == _T_121[11:0] ? image_77 : _GEN_9358; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9360 = 12'h4e == _T_121[11:0] ? image_78 : _GEN_9359; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9361 = 12'h4f == _T_121[11:0] ? image_79 : _GEN_9360; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9362 = 12'h50 == _T_121[11:0] ? image_80 : _GEN_9361; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9363 = 12'h51 == _T_121[11:0] ? image_81 : _GEN_9362; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9364 = 12'h52 == _T_121[11:0] ? image_82 : _GEN_9363; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9365 = 12'h53 == _T_121[11:0] ? image_83 : _GEN_9364; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9366 = 12'h54 == _T_121[11:0] ? image_84 : _GEN_9365; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9367 = 12'h55 == _T_121[11:0] ? image_85 : _GEN_9366; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9368 = 12'h56 == _T_121[11:0] ? image_86 : _GEN_9367; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9369 = 12'h57 == _T_121[11:0] ? image_87 : _GEN_9368; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9370 = 12'h58 == _T_121[11:0] ? image_88 : _GEN_9369; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9371 = 12'h59 == _T_121[11:0] ? image_89 : _GEN_9370; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9372 = 12'h5a == _T_121[11:0] ? image_90 : _GEN_9371; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9373 = 12'h5b == _T_121[11:0] ? 4'h0 : _GEN_9372; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9374 = 12'h5c == _T_121[11:0] ? 4'h0 : _GEN_9373; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9375 = 12'h5d == _T_121[11:0] ? image_93 : _GEN_9374; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9376 = 12'h5e == _T_121[11:0] ? 4'h0 : _GEN_9375; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9377 = 12'h5f == _T_121[11:0] ? image_95 : _GEN_9376; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9378 = 12'h60 == _T_121[11:0] ? image_96 : _GEN_9377; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9379 = 12'h61 == _T_121[11:0] ? image_97 : _GEN_9378; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9380 = 12'h62 == _T_121[11:0] ? image_98 : _GEN_9379; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9381 = 12'h63 == _T_121[11:0] ? image_99 : _GEN_9380; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9382 = 12'h64 == _T_121[11:0] ? image_100 : _GEN_9381; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9383 = 12'h65 == _T_121[11:0] ? image_101 : _GEN_9382; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9384 = 12'h66 == _T_121[11:0] ? image_102 : _GEN_9383; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9385 = 12'h67 == _T_121[11:0] ? image_103 : _GEN_9384; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9386 = 12'h68 == _T_121[11:0] ? image_104 : _GEN_9385; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9387 = 12'h69 == _T_121[11:0] ? image_105 : _GEN_9386; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9388 = 12'h6a == _T_121[11:0] ? image_106 : _GEN_9387; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9389 = 12'h6b == _T_121[11:0] ? image_107 : _GEN_9388; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9390 = 12'h6c == _T_121[11:0] ? image_108 : _GEN_9389; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9391 = 12'h6d == _T_121[11:0] ? 4'h0 : _GEN_9390; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9392 = 12'h6e == _T_121[11:0] ? 4'h0 : _GEN_9391; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9393 = 12'h6f == _T_121[11:0] ? 4'h0 : _GEN_9392; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9394 = 12'h70 == _T_121[11:0] ? 4'h0 : _GEN_9393; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9395 = 12'h71 == _T_121[11:0] ? 4'h0 : _GEN_9394; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9396 = 12'h72 == _T_121[11:0] ? 4'h0 : _GEN_9395; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9397 = 12'h73 == _T_121[11:0] ? 4'h0 : _GEN_9396; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9398 = 12'h74 == _T_121[11:0] ? 4'h0 : _GEN_9397; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9399 = 12'h75 == _T_121[11:0] ? 4'h0 : _GEN_9398; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9400 = 12'h76 == _T_121[11:0] ? 4'h0 : _GEN_9399; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9401 = 12'h77 == _T_121[11:0] ? 4'h0 : _GEN_9400; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9402 = 12'h78 == _T_121[11:0] ? 4'h0 : _GEN_9401; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9403 = 12'h79 == _T_121[11:0] ? 4'h0 : _GEN_9402; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9404 = 12'h7a == _T_121[11:0] ? 4'h0 : _GEN_9403; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9405 = 12'h7b == _T_121[11:0] ? 4'h0 : _GEN_9404; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9406 = 12'h7c == _T_121[11:0] ? 4'h0 : _GEN_9405; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9407 = 12'h7d == _T_121[11:0] ? 4'h0 : _GEN_9406; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9408 = 12'h7e == _T_121[11:0] ? 4'h0 : _GEN_9407; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9409 = 12'h7f == _T_121[11:0] ? 4'h0 : _GEN_9408; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9410 = 12'h80 == _T_121[11:0] ? 4'h0 : _GEN_9409; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9411 = 12'h81 == _T_121[11:0] ? 4'h0 : _GEN_9410; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9412 = 12'h82 == _T_121[11:0] ? 4'h0 : _GEN_9411; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9413 = 12'h83 == _T_121[11:0] ? 4'h0 : _GEN_9412; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9414 = 12'h84 == _T_121[11:0] ? 4'h0 : _GEN_9413; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9415 = 12'h85 == _T_121[11:0] ? 4'h0 : _GEN_9414; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9416 = 12'h86 == _T_121[11:0] ? 4'h0 : _GEN_9415; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9417 = 12'h87 == _T_121[11:0] ? 4'h0 : _GEN_9416; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9418 = 12'h88 == _T_121[11:0] ? image_136 : _GEN_9417; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9419 = 12'h89 == _T_121[11:0] ? image_137 : _GEN_9418; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9420 = 12'h8a == _T_121[11:0] ? image_138 : _GEN_9419; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9421 = 12'h8b == _T_121[11:0] ? image_139 : _GEN_9420; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9422 = 12'h8c == _T_121[11:0] ? image_140 : _GEN_9421; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9423 = 12'h8d == _T_121[11:0] ? image_141 : _GEN_9422; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9424 = 12'h8e == _T_121[11:0] ? image_142 : _GEN_9423; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9425 = 12'h8f == _T_121[11:0] ? image_143 : _GEN_9424; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9426 = 12'h90 == _T_121[11:0] ? image_144 : _GEN_9425; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9427 = 12'h91 == _T_121[11:0] ? image_145 : _GEN_9426; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9428 = 12'h92 == _T_121[11:0] ? image_146 : _GEN_9427; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9429 = 12'h93 == _T_121[11:0] ? image_147 : _GEN_9428; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9430 = 12'h94 == _T_121[11:0] ? image_148 : _GEN_9429; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9431 = 12'h95 == _T_121[11:0] ? image_149 : _GEN_9430; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9432 = 12'h96 == _T_121[11:0] ? image_150 : _GEN_9431; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9433 = 12'h97 == _T_121[11:0] ? image_151 : _GEN_9432; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9434 = 12'h98 == _T_121[11:0] ? image_152 : _GEN_9433; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9435 = 12'h99 == _T_121[11:0] ? image_153 : _GEN_9434; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9436 = 12'h9a == _T_121[11:0] ? image_154 : _GEN_9435; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9437 = 12'h9b == _T_121[11:0] ? image_155 : _GEN_9436; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9438 = 12'h9c == _T_121[11:0] ? 4'h0 : _GEN_9437; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9439 = 12'h9d == _T_121[11:0] ? image_157 : _GEN_9438; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9440 = 12'h9e == _T_121[11:0] ? image_158 : _GEN_9439; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9441 = 12'h9f == _T_121[11:0] ? image_159 : _GEN_9440; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9442 = 12'ha0 == _T_121[11:0] ? image_160 : _GEN_9441; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9443 = 12'ha1 == _T_121[11:0] ? image_161 : _GEN_9442; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9444 = 12'ha2 == _T_121[11:0] ? image_162 : _GEN_9443; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9445 = 12'ha3 == _T_121[11:0] ? image_163 : _GEN_9444; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9446 = 12'ha4 == _T_121[11:0] ? image_164 : _GEN_9445; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9447 = 12'ha5 == _T_121[11:0] ? image_165 : _GEN_9446; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9448 = 12'ha6 == _T_121[11:0] ? image_166 : _GEN_9447; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9449 = 12'ha7 == _T_121[11:0] ? image_167 : _GEN_9448; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9450 = 12'ha8 == _T_121[11:0] ? image_168 : _GEN_9449; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9451 = 12'ha9 == _T_121[11:0] ? image_169 : _GEN_9450; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9452 = 12'haa == _T_121[11:0] ? image_170 : _GEN_9451; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9453 = 12'hab == _T_121[11:0] ? image_171 : _GEN_9452; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9454 = 12'hac == _T_121[11:0] ? image_172 : _GEN_9453; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9455 = 12'had == _T_121[11:0] ? image_173 : _GEN_9454; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9456 = 12'hae == _T_121[11:0] ? image_174 : _GEN_9455; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9457 = 12'haf == _T_121[11:0] ? image_175 : _GEN_9456; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9458 = 12'hb0 == _T_121[11:0] ? image_176 : _GEN_9457; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9459 = 12'hb1 == _T_121[11:0] ? image_177 : _GEN_9458; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9460 = 12'hb2 == _T_121[11:0] ? image_178 : _GEN_9459; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9461 = 12'hb3 == _T_121[11:0] ? image_179 : _GEN_9460; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9462 = 12'hb4 == _T_121[11:0] ? 4'h0 : _GEN_9461; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9463 = 12'hb5 == _T_121[11:0] ? 4'h0 : _GEN_9462; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9464 = 12'hb6 == _T_121[11:0] ? 4'h0 : _GEN_9463; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9465 = 12'hb7 == _T_121[11:0] ? 4'h0 : _GEN_9464; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9466 = 12'hb8 == _T_121[11:0] ? 4'h0 : _GEN_9465; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9467 = 12'hb9 == _T_121[11:0] ? 4'h0 : _GEN_9466; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9468 = 12'hba == _T_121[11:0] ? 4'h0 : _GEN_9467; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9469 = 12'hbb == _T_121[11:0] ? 4'h0 : _GEN_9468; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9470 = 12'hbc == _T_121[11:0] ? 4'h0 : _GEN_9469; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9471 = 12'hbd == _T_121[11:0] ? 4'h0 : _GEN_9470; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9472 = 12'hbe == _T_121[11:0] ? 4'h0 : _GEN_9471; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9473 = 12'hbf == _T_121[11:0] ? 4'h0 : _GEN_9472; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9474 = 12'hc0 == _T_121[11:0] ? 4'h0 : _GEN_9473; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9475 = 12'hc1 == _T_121[11:0] ? 4'h0 : _GEN_9474; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9476 = 12'hc2 == _T_121[11:0] ? 4'h0 : _GEN_9475; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9477 = 12'hc3 == _T_121[11:0] ? 4'h0 : _GEN_9476; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9478 = 12'hc4 == _T_121[11:0] ? 4'h0 : _GEN_9477; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9479 = 12'hc5 == _T_121[11:0] ? 4'h0 : _GEN_9478; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9480 = 12'hc6 == _T_121[11:0] ? 4'h0 : _GEN_9479; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9481 = 12'hc7 == _T_121[11:0] ? image_199 : _GEN_9480; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9482 = 12'hc8 == _T_121[11:0] ? image_200 : _GEN_9481; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9483 = 12'hc9 == _T_121[11:0] ? image_201 : _GEN_9482; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9484 = 12'hca == _T_121[11:0] ? image_202 : _GEN_9483; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9485 = 12'hcb == _T_121[11:0] ? image_203 : _GEN_9484; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9486 = 12'hcc == _T_121[11:0] ? image_204 : _GEN_9485; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9487 = 12'hcd == _T_121[11:0] ? image_205 : _GEN_9486; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9488 = 12'hce == _T_121[11:0] ? image_206 : _GEN_9487; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9489 = 12'hcf == _T_121[11:0] ? image_207 : _GEN_9488; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9490 = 12'hd0 == _T_121[11:0] ? image_208 : _GEN_9489; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9491 = 12'hd1 == _T_121[11:0] ? image_209 : _GEN_9490; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9492 = 12'hd2 == _T_121[11:0] ? image_210 : _GEN_9491; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9493 = 12'hd3 == _T_121[11:0] ? image_211 : _GEN_9492; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9494 = 12'hd4 == _T_121[11:0] ? image_212 : _GEN_9493; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9495 = 12'hd5 == _T_121[11:0] ? image_213 : _GEN_9494; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9496 = 12'hd6 == _T_121[11:0] ? image_214 : _GEN_9495; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9497 = 12'hd7 == _T_121[11:0] ? image_215 : _GEN_9496; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9498 = 12'hd8 == _T_121[11:0] ? image_216 : _GEN_9497; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9499 = 12'hd9 == _T_121[11:0] ? image_217 : _GEN_9498; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9500 = 12'hda == _T_121[11:0] ? image_218 : _GEN_9499; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9501 = 12'hdb == _T_121[11:0] ? image_219 : _GEN_9500; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9502 = 12'hdc == _T_121[11:0] ? image_220 : _GEN_9501; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9503 = 12'hdd == _T_121[11:0] ? image_221 : _GEN_9502; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9504 = 12'hde == _T_121[11:0] ? image_222 : _GEN_9503; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9505 = 12'hdf == _T_121[11:0] ? image_223 : _GEN_9504; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9506 = 12'he0 == _T_121[11:0] ? image_224 : _GEN_9505; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9507 = 12'he1 == _T_121[11:0] ? image_225 : _GEN_9506; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9508 = 12'he2 == _T_121[11:0] ? image_226 : _GEN_9507; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9509 = 12'he3 == _T_121[11:0] ? image_227 : _GEN_9508; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9510 = 12'he4 == _T_121[11:0] ? image_228 : _GEN_9509; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9511 = 12'he5 == _T_121[11:0] ? image_229 : _GEN_9510; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9512 = 12'he6 == _T_121[11:0] ? image_230 : _GEN_9511; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9513 = 12'he7 == _T_121[11:0] ? image_231 : _GEN_9512; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9514 = 12'he8 == _T_121[11:0] ? image_232 : _GEN_9513; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9515 = 12'he9 == _T_121[11:0] ? image_233 : _GEN_9514; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9516 = 12'hea == _T_121[11:0] ? image_234 : _GEN_9515; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9517 = 12'heb == _T_121[11:0] ? image_235 : _GEN_9516; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9518 = 12'hec == _T_121[11:0] ? image_236 : _GEN_9517; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9519 = 12'hed == _T_121[11:0] ? image_237 : _GEN_9518; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9520 = 12'hee == _T_121[11:0] ? image_238 : _GEN_9519; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9521 = 12'hef == _T_121[11:0] ? image_239 : _GEN_9520; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9522 = 12'hf0 == _T_121[11:0] ? image_240 : _GEN_9521; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9523 = 12'hf1 == _T_121[11:0] ? image_241 : _GEN_9522; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9524 = 12'hf2 == _T_121[11:0] ? image_242 : _GEN_9523; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9525 = 12'hf3 == _T_121[11:0] ? image_243 : _GEN_9524; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9526 = 12'hf4 == _T_121[11:0] ? image_244 : _GEN_9525; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9527 = 12'hf5 == _T_121[11:0] ? image_245 : _GEN_9526; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9528 = 12'hf6 == _T_121[11:0] ? image_246 : _GEN_9527; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9529 = 12'hf7 == _T_121[11:0] ? 4'h0 : _GEN_9528; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9530 = 12'hf8 == _T_121[11:0] ? 4'h0 : _GEN_9529; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9531 = 12'hf9 == _T_121[11:0] ? 4'h0 : _GEN_9530; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9532 = 12'hfa == _T_121[11:0] ? 4'h0 : _GEN_9531; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9533 = 12'hfb == _T_121[11:0] ? 4'h0 : _GEN_9532; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9534 = 12'hfc == _T_121[11:0] ? 4'h0 : _GEN_9533; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9535 = 12'hfd == _T_121[11:0] ? 4'h0 : _GEN_9534; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9536 = 12'hfe == _T_121[11:0] ? 4'h0 : _GEN_9535; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9537 = 12'hff == _T_121[11:0] ? 4'h0 : _GEN_9536; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9538 = 12'h100 == _T_121[11:0] ? 4'h0 : _GEN_9537; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9539 = 12'h101 == _T_121[11:0] ? 4'h0 : _GEN_9538; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9540 = 12'h102 == _T_121[11:0] ? 4'h0 : _GEN_9539; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9541 = 12'h103 == _T_121[11:0] ? 4'h0 : _GEN_9540; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9542 = 12'h104 == _T_121[11:0] ? 4'h0 : _GEN_9541; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9543 = 12'h105 == _T_121[11:0] ? 4'h0 : _GEN_9542; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9544 = 12'h106 == _T_121[11:0] ? image_262 : _GEN_9543; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9545 = 12'h107 == _T_121[11:0] ? image_263 : _GEN_9544; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9546 = 12'h108 == _T_121[11:0] ? image_264 : _GEN_9545; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9547 = 12'h109 == _T_121[11:0] ? image_265 : _GEN_9546; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9548 = 12'h10a == _T_121[11:0] ? image_266 : _GEN_9547; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9549 = 12'h10b == _T_121[11:0] ? image_267 : _GEN_9548; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9550 = 12'h10c == _T_121[11:0] ? image_268 : _GEN_9549; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9551 = 12'h10d == _T_121[11:0] ? image_269 : _GEN_9550; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9552 = 12'h10e == _T_121[11:0] ? image_270 : _GEN_9551; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9553 = 12'h10f == _T_121[11:0] ? image_271 : _GEN_9552; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9554 = 12'h110 == _T_121[11:0] ? image_272 : _GEN_9553; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9555 = 12'h111 == _T_121[11:0] ? image_273 : _GEN_9554; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9556 = 12'h112 == _T_121[11:0] ? image_274 : _GEN_9555; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9557 = 12'h113 == _T_121[11:0] ? image_275 : _GEN_9556; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9558 = 12'h114 == _T_121[11:0] ? image_276 : _GEN_9557; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9559 = 12'h115 == _T_121[11:0] ? image_277 : _GEN_9558; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9560 = 12'h116 == _T_121[11:0] ? image_278 : _GEN_9559; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9561 = 12'h117 == _T_121[11:0] ? image_279 : _GEN_9560; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9562 = 12'h118 == _T_121[11:0] ? image_280 : _GEN_9561; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9563 = 12'h119 == _T_121[11:0] ? image_281 : _GEN_9562; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9564 = 12'h11a == _T_121[11:0] ? image_282 : _GEN_9563; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9565 = 12'h11b == _T_121[11:0] ? image_283 : _GEN_9564; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9566 = 12'h11c == _T_121[11:0] ? image_284 : _GEN_9565; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9567 = 12'h11d == _T_121[11:0] ? image_285 : _GEN_9566; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9568 = 12'h11e == _T_121[11:0] ? image_286 : _GEN_9567; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9569 = 12'h11f == _T_121[11:0] ? image_287 : _GEN_9568; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9570 = 12'h120 == _T_121[11:0] ? image_288 : _GEN_9569; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9571 = 12'h121 == _T_121[11:0] ? image_289 : _GEN_9570; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9572 = 12'h122 == _T_121[11:0] ? image_290 : _GEN_9571; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9573 = 12'h123 == _T_121[11:0] ? image_291 : _GEN_9572; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9574 = 12'h124 == _T_121[11:0] ? image_292 : _GEN_9573; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9575 = 12'h125 == _T_121[11:0] ? image_293 : _GEN_9574; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9576 = 12'h126 == _T_121[11:0] ? image_294 : _GEN_9575; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9577 = 12'h127 == _T_121[11:0] ? image_295 : _GEN_9576; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9578 = 12'h128 == _T_121[11:0] ? image_296 : _GEN_9577; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9579 = 12'h129 == _T_121[11:0] ? image_297 : _GEN_9578; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9580 = 12'h12a == _T_121[11:0] ? image_298 : _GEN_9579; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9581 = 12'h12b == _T_121[11:0] ? image_299 : _GEN_9580; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9582 = 12'h12c == _T_121[11:0] ? image_300 : _GEN_9581; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9583 = 12'h12d == _T_121[11:0] ? image_301 : _GEN_9582; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9584 = 12'h12e == _T_121[11:0] ? image_302 : _GEN_9583; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9585 = 12'h12f == _T_121[11:0] ? image_303 : _GEN_9584; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9586 = 12'h130 == _T_121[11:0] ? image_304 : _GEN_9585; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9587 = 12'h131 == _T_121[11:0] ? image_305 : _GEN_9586; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9588 = 12'h132 == _T_121[11:0] ? image_306 : _GEN_9587; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9589 = 12'h133 == _T_121[11:0] ? image_307 : _GEN_9588; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9590 = 12'h134 == _T_121[11:0] ? image_308 : _GEN_9589; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9591 = 12'h135 == _T_121[11:0] ? image_309 : _GEN_9590; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9592 = 12'h136 == _T_121[11:0] ? image_310 : _GEN_9591; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9593 = 12'h137 == _T_121[11:0] ? image_311 : _GEN_9592; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9594 = 12'h138 == _T_121[11:0] ? image_312 : _GEN_9593; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9595 = 12'h139 == _T_121[11:0] ? image_313 : _GEN_9594; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9596 = 12'h13a == _T_121[11:0] ? image_314 : _GEN_9595; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9597 = 12'h13b == _T_121[11:0] ? image_315 : _GEN_9596; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9598 = 12'h13c == _T_121[11:0] ? 4'h0 : _GEN_9597; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9599 = 12'h13d == _T_121[11:0] ? 4'h0 : _GEN_9598; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9600 = 12'h13e == _T_121[11:0] ? 4'h0 : _GEN_9599; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9601 = 12'h13f == _T_121[11:0] ? 4'h0 : _GEN_9600; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9602 = 12'h140 == _T_121[11:0] ? 4'h0 : _GEN_9601; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9603 = 12'h141 == _T_121[11:0] ? 4'h0 : _GEN_9602; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9604 = 12'h142 == _T_121[11:0] ? 4'h0 : _GEN_9603; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9605 = 12'h143 == _T_121[11:0] ? 4'h0 : _GEN_9604; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9606 = 12'h144 == _T_121[11:0] ? 4'h0 : _GEN_9605; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9607 = 12'h145 == _T_121[11:0] ? image_325 : _GEN_9606; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9608 = 12'h146 == _T_121[11:0] ? image_326 : _GEN_9607; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9609 = 12'h147 == _T_121[11:0] ? image_327 : _GEN_9608; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9610 = 12'h148 == _T_121[11:0] ? image_328 : _GEN_9609; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9611 = 12'h149 == _T_121[11:0] ? image_329 : _GEN_9610; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9612 = 12'h14a == _T_121[11:0] ? image_330 : _GEN_9611; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9613 = 12'h14b == _T_121[11:0] ? image_331 : _GEN_9612; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9614 = 12'h14c == _T_121[11:0] ? image_332 : _GEN_9613; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9615 = 12'h14d == _T_121[11:0] ? image_333 : _GEN_9614; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9616 = 12'h14e == _T_121[11:0] ? image_334 : _GEN_9615; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9617 = 12'h14f == _T_121[11:0] ? image_335 : _GEN_9616; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9618 = 12'h150 == _T_121[11:0] ? image_336 : _GEN_9617; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9619 = 12'h151 == _T_121[11:0] ? image_337 : _GEN_9618; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9620 = 12'h152 == _T_121[11:0] ? image_338 : _GEN_9619; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9621 = 12'h153 == _T_121[11:0] ? image_339 : _GEN_9620; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9622 = 12'h154 == _T_121[11:0] ? image_340 : _GEN_9621; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9623 = 12'h155 == _T_121[11:0] ? image_341 : _GEN_9622; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9624 = 12'h156 == _T_121[11:0] ? image_342 : _GEN_9623; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9625 = 12'h157 == _T_121[11:0] ? image_343 : _GEN_9624; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9626 = 12'h158 == _T_121[11:0] ? image_344 : _GEN_9625; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9627 = 12'h159 == _T_121[11:0] ? image_345 : _GEN_9626; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9628 = 12'h15a == _T_121[11:0] ? image_346 : _GEN_9627; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9629 = 12'h15b == _T_121[11:0] ? image_347 : _GEN_9628; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9630 = 12'h15c == _T_121[11:0] ? image_348 : _GEN_9629; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9631 = 12'h15d == _T_121[11:0] ? image_349 : _GEN_9630; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9632 = 12'h15e == _T_121[11:0] ? image_350 : _GEN_9631; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9633 = 12'h15f == _T_121[11:0] ? image_351 : _GEN_9632; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9634 = 12'h160 == _T_121[11:0] ? image_352 : _GEN_9633; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9635 = 12'h161 == _T_121[11:0] ? image_353 : _GEN_9634; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9636 = 12'h162 == _T_121[11:0] ? image_354 : _GEN_9635; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9637 = 12'h163 == _T_121[11:0] ? image_355 : _GEN_9636; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9638 = 12'h164 == _T_121[11:0] ? image_356 : _GEN_9637; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9639 = 12'h165 == _T_121[11:0] ? image_357 : _GEN_9638; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9640 = 12'h166 == _T_121[11:0] ? image_358 : _GEN_9639; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9641 = 12'h167 == _T_121[11:0] ? image_359 : _GEN_9640; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9642 = 12'h168 == _T_121[11:0] ? image_360 : _GEN_9641; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9643 = 12'h169 == _T_121[11:0] ? image_361 : _GEN_9642; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9644 = 12'h16a == _T_121[11:0] ? image_362 : _GEN_9643; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9645 = 12'h16b == _T_121[11:0] ? image_363 : _GEN_9644; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9646 = 12'h16c == _T_121[11:0] ? image_364 : _GEN_9645; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9647 = 12'h16d == _T_121[11:0] ? image_365 : _GEN_9646; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9648 = 12'h16e == _T_121[11:0] ? image_366 : _GEN_9647; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9649 = 12'h16f == _T_121[11:0] ? image_367 : _GEN_9648; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9650 = 12'h170 == _T_121[11:0] ? image_368 : _GEN_9649; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9651 = 12'h171 == _T_121[11:0] ? image_369 : _GEN_9650; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9652 = 12'h172 == _T_121[11:0] ? image_370 : _GEN_9651; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9653 = 12'h173 == _T_121[11:0] ? image_371 : _GEN_9652; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9654 = 12'h174 == _T_121[11:0] ? image_372 : _GEN_9653; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9655 = 12'h175 == _T_121[11:0] ? image_373 : _GEN_9654; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9656 = 12'h176 == _T_121[11:0] ? image_374 : _GEN_9655; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9657 = 12'h177 == _T_121[11:0] ? image_375 : _GEN_9656; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9658 = 12'h178 == _T_121[11:0] ? image_376 : _GEN_9657; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9659 = 12'h179 == _T_121[11:0] ? image_377 : _GEN_9658; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9660 = 12'h17a == _T_121[11:0] ? image_378 : _GEN_9659; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9661 = 12'h17b == _T_121[11:0] ? image_379 : _GEN_9660; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9662 = 12'h17c == _T_121[11:0] ? 4'h0 : _GEN_9661; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9663 = 12'h17d == _T_121[11:0] ? 4'h0 : _GEN_9662; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9664 = 12'h17e == _T_121[11:0] ? 4'h0 : _GEN_9663; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9665 = 12'h17f == _T_121[11:0] ? 4'h0 : _GEN_9664; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9666 = 12'h180 == _T_121[11:0] ? 4'h0 : _GEN_9665; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9667 = 12'h181 == _T_121[11:0] ? 4'h0 : _GEN_9666; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9668 = 12'h182 == _T_121[11:0] ? 4'h0 : _GEN_9667; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9669 = 12'h183 == _T_121[11:0] ? 4'h0 : _GEN_9668; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9670 = 12'h184 == _T_121[11:0] ? image_388 : _GEN_9669; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9671 = 12'h185 == _T_121[11:0] ? image_389 : _GEN_9670; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9672 = 12'h186 == _T_121[11:0] ? image_390 : _GEN_9671; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9673 = 12'h187 == _T_121[11:0] ? image_391 : _GEN_9672; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9674 = 12'h188 == _T_121[11:0] ? image_392 : _GEN_9673; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9675 = 12'h189 == _T_121[11:0] ? image_393 : _GEN_9674; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9676 = 12'h18a == _T_121[11:0] ? image_394 : _GEN_9675; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9677 = 12'h18b == _T_121[11:0] ? image_395 : _GEN_9676; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9678 = 12'h18c == _T_121[11:0] ? image_396 : _GEN_9677; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9679 = 12'h18d == _T_121[11:0] ? image_397 : _GEN_9678; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9680 = 12'h18e == _T_121[11:0] ? image_398 : _GEN_9679; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9681 = 12'h18f == _T_121[11:0] ? image_399 : _GEN_9680; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9682 = 12'h190 == _T_121[11:0] ? image_400 : _GEN_9681; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9683 = 12'h191 == _T_121[11:0] ? image_401 : _GEN_9682; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9684 = 12'h192 == _T_121[11:0] ? image_402 : _GEN_9683; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9685 = 12'h193 == _T_121[11:0] ? image_403 : _GEN_9684; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9686 = 12'h194 == _T_121[11:0] ? image_404 : _GEN_9685; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9687 = 12'h195 == _T_121[11:0] ? image_405 : _GEN_9686; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9688 = 12'h196 == _T_121[11:0] ? image_406 : _GEN_9687; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9689 = 12'h197 == _T_121[11:0] ? image_407 : _GEN_9688; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9690 = 12'h198 == _T_121[11:0] ? image_408 : _GEN_9689; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9691 = 12'h199 == _T_121[11:0] ? image_409 : _GEN_9690; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9692 = 12'h19a == _T_121[11:0] ? image_410 : _GEN_9691; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9693 = 12'h19b == _T_121[11:0] ? image_411 : _GEN_9692; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9694 = 12'h19c == _T_121[11:0] ? image_412 : _GEN_9693; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9695 = 12'h19d == _T_121[11:0] ? image_413 : _GEN_9694; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9696 = 12'h19e == _T_121[11:0] ? image_414 : _GEN_9695; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9697 = 12'h19f == _T_121[11:0] ? image_415 : _GEN_9696; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9698 = 12'h1a0 == _T_121[11:0] ? image_416 : _GEN_9697; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9699 = 12'h1a1 == _T_121[11:0] ? image_417 : _GEN_9698; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9700 = 12'h1a2 == _T_121[11:0] ? image_418 : _GEN_9699; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9701 = 12'h1a3 == _T_121[11:0] ? image_419 : _GEN_9700; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9702 = 12'h1a4 == _T_121[11:0] ? image_420 : _GEN_9701; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9703 = 12'h1a5 == _T_121[11:0] ? image_421 : _GEN_9702; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9704 = 12'h1a6 == _T_121[11:0] ? image_422 : _GEN_9703; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9705 = 12'h1a7 == _T_121[11:0] ? image_423 : _GEN_9704; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9706 = 12'h1a8 == _T_121[11:0] ? image_424 : _GEN_9705; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9707 = 12'h1a9 == _T_121[11:0] ? image_425 : _GEN_9706; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9708 = 12'h1aa == _T_121[11:0] ? image_426 : _GEN_9707; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9709 = 12'h1ab == _T_121[11:0] ? image_427 : _GEN_9708; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9710 = 12'h1ac == _T_121[11:0] ? image_428 : _GEN_9709; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9711 = 12'h1ad == _T_121[11:0] ? image_429 : _GEN_9710; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9712 = 12'h1ae == _T_121[11:0] ? image_430 : _GEN_9711; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9713 = 12'h1af == _T_121[11:0] ? image_431 : _GEN_9712; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9714 = 12'h1b0 == _T_121[11:0] ? image_432 : _GEN_9713; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9715 = 12'h1b1 == _T_121[11:0] ? image_433 : _GEN_9714; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9716 = 12'h1b2 == _T_121[11:0] ? image_434 : _GEN_9715; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9717 = 12'h1b3 == _T_121[11:0] ? image_435 : _GEN_9716; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9718 = 12'h1b4 == _T_121[11:0] ? image_436 : _GEN_9717; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9719 = 12'h1b5 == _T_121[11:0] ? image_437 : _GEN_9718; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9720 = 12'h1b6 == _T_121[11:0] ? image_438 : _GEN_9719; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9721 = 12'h1b7 == _T_121[11:0] ? image_439 : _GEN_9720; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9722 = 12'h1b8 == _T_121[11:0] ? image_440 : _GEN_9721; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9723 = 12'h1b9 == _T_121[11:0] ? image_441 : _GEN_9722; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9724 = 12'h1ba == _T_121[11:0] ? image_442 : _GEN_9723; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9725 = 12'h1bb == _T_121[11:0] ? image_443 : _GEN_9724; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9726 = 12'h1bc == _T_121[11:0] ? image_444 : _GEN_9725; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9727 = 12'h1bd == _T_121[11:0] ? 4'h0 : _GEN_9726; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9728 = 12'h1be == _T_121[11:0] ? 4'h0 : _GEN_9727; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9729 = 12'h1bf == _T_121[11:0] ? 4'h0 : _GEN_9728; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9730 = 12'h1c0 == _T_121[11:0] ? 4'h0 : _GEN_9729; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9731 = 12'h1c1 == _T_121[11:0] ? 4'h0 : _GEN_9730; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9732 = 12'h1c2 == _T_121[11:0] ? 4'h0 : _GEN_9731; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9733 = 12'h1c3 == _T_121[11:0] ? image_451 : _GEN_9732; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9734 = 12'h1c4 == _T_121[11:0] ? image_452 : _GEN_9733; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9735 = 12'h1c5 == _T_121[11:0] ? image_453 : _GEN_9734; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9736 = 12'h1c6 == _T_121[11:0] ? image_454 : _GEN_9735; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9737 = 12'h1c7 == _T_121[11:0] ? image_455 : _GEN_9736; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9738 = 12'h1c8 == _T_121[11:0] ? image_456 : _GEN_9737; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9739 = 12'h1c9 == _T_121[11:0] ? image_457 : _GEN_9738; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9740 = 12'h1ca == _T_121[11:0] ? image_458 : _GEN_9739; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9741 = 12'h1cb == _T_121[11:0] ? image_459 : _GEN_9740; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9742 = 12'h1cc == _T_121[11:0] ? image_460 : _GEN_9741; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9743 = 12'h1cd == _T_121[11:0] ? image_461 : _GEN_9742; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9744 = 12'h1ce == _T_121[11:0] ? image_462 : _GEN_9743; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9745 = 12'h1cf == _T_121[11:0] ? image_463 : _GEN_9744; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9746 = 12'h1d0 == _T_121[11:0] ? image_464 : _GEN_9745; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9747 = 12'h1d1 == _T_121[11:0] ? image_465 : _GEN_9746; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9748 = 12'h1d2 == _T_121[11:0] ? image_466 : _GEN_9747; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9749 = 12'h1d3 == _T_121[11:0] ? image_467 : _GEN_9748; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9750 = 12'h1d4 == _T_121[11:0] ? image_468 : _GEN_9749; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9751 = 12'h1d5 == _T_121[11:0] ? image_469 : _GEN_9750; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9752 = 12'h1d6 == _T_121[11:0] ? image_470 : _GEN_9751; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9753 = 12'h1d7 == _T_121[11:0] ? image_471 : _GEN_9752; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9754 = 12'h1d8 == _T_121[11:0] ? image_472 : _GEN_9753; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9755 = 12'h1d9 == _T_121[11:0] ? image_473 : _GEN_9754; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9756 = 12'h1da == _T_121[11:0] ? image_474 : _GEN_9755; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9757 = 12'h1db == _T_121[11:0] ? image_475 : _GEN_9756; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9758 = 12'h1dc == _T_121[11:0] ? image_476 : _GEN_9757; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9759 = 12'h1dd == _T_121[11:0] ? image_477 : _GEN_9758; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9760 = 12'h1de == _T_121[11:0] ? image_478 : _GEN_9759; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9761 = 12'h1df == _T_121[11:0] ? image_479 : _GEN_9760; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9762 = 12'h1e0 == _T_121[11:0] ? image_480 : _GEN_9761; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9763 = 12'h1e1 == _T_121[11:0] ? image_481 : _GEN_9762; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9764 = 12'h1e2 == _T_121[11:0] ? image_482 : _GEN_9763; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9765 = 12'h1e3 == _T_121[11:0] ? image_483 : _GEN_9764; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9766 = 12'h1e4 == _T_121[11:0] ? image_484 : _GEN_9765; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9767 = 12'h1e5 == _T_121[11:0] ? image_485 : _GEN_9766; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9768 = 12'h1e6 == _T_121[11:0] ? image_486 : _GEN_9767; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9769 = 12'h1e7 == _T_121[11:0] ? image_487 : _GEN_9768; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9770 = 12'h1e8 == _T_121[11:0] ? image_488 : _GEN_9769; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9771 = 12'h1e9 == _T_121[11:0] ? image_489 : _GEN_9770; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9772 = 12'h1ea == _T_121[11:0] ? image_490 : _GEN_9771; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9773 = 12'h1eb == _T_121[11:0] ? image_491 : _GEN_9772; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9774 = 12'h1ec == _T_121[11:0] ? image_492 : _GEN_9773; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9775 = 12'h1ed == _T_121[11:0] ? image_493 : _GEN_9774; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9776 = 12'h1ee == _T_121[11:0] ? image_494 : _GEN_9775; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9777 = 12'h1ef == _T_121[11:0] ? image_495 : _GEN_9776; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9778 = 12'h1f0 == _T_121[11:0] ? image_496 : _GEN_9777; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9779 = 12'h1f1 == _T_121[11:0] ? image_497 : _GEN_9778; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9780 = 12'h1f2 == _T_121[11:0] ? image_498 : _GEN_9779; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9781 = 12'h1f3 == _T_121[11:0] ? image_499 : _GEN_9780; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9782 = 12'h1f4 == _T_121[11:0] ? image_500 : _GEN_9781; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9783 = 12'h1f5 == _T_121[11:0] ? image_501 : _GEN_9782; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9784 = 12'h1f6 == _T_121[11:0] ? image_502 : _GEN_9783; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9785 = 12'h1f7 == _T_121[11:0] ? image_503 : _GEN_9784; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9786 = 12'h1f8 == _T_121[11:0] ? image_504 : _GEN_9785; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9787 = 12'h1f9 == _T_121[11:0] ? image_505 : _GEN_9786; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9788 = 12'h1fa == _T_121[11:0] ? image_506 : _GEN_9787; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9789 = 12'h1fb == _T_121[11:0] ? image_507 : _GEN_9788; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9790 = 12'h1fc == _T_121[11:0] ? image_508 : _GEN_9789; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9791 = 12'h1fd == _T_121[11:0] ? image_509 : _GEN_9790; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9792 = 12'h1fe == _T_121[11:0] ? 4'h0 : _GEN_9791; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9793 = 12'h1ff == _T_121[11:0] ? 4'h0 : _GEN_9792; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9794 = 12'h200 == _T_121[11:0] ? 4'h0 : _GEN_9793; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9795 = 12'h201 == _T_121[11:0] ? 4'h0 : _GEN_9794; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9796 = 12'h202 == _T_121[11:0] ? 4'h0 : _GEN_9795; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9797 = 12'h203 == _T_121[11:0] ? image_515 : _GEN_9796; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9798 = 12'h204 == _T_121[11:0] ? image_516 : _GEN_9797; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9799 = 12'h205 == _T_121[11:0] ? image_517 : _GEN_9798; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9800 = 12'h206 == _T_121[11:0] ? image_518 : _GEN_9799; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9801 = 12'h207 == _T_121[11:0] ? image_519 : _GEN_9800; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9802 = 12'h208 == _T_121[11:0] ? image_520 : _GEN_9801; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9803 = 12'h209 == _T_121[11:0] ? image_521 : _GEN_9802; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9804 = 12'h20a == _T_121[11:0] ? image_522 : _GEN_9803; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9805 = 12'h20b == _T_121[11:0] ? image_523 : _GEN_9804; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9806 = 12'h20c == _T_121[11:0] ? image_524 : _GEN_9805; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9807 = 12'h20d == _T_121[11:0] ? image_525 : _GEN_9806; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9808 = 12'h20e == _T_121[11:0] ? image_526 : _GEN_9807; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9809 = 12'h20f == _T_121[11:0] ? image_527 : _GEN_9808; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9810 = 12'h210 == _T_121[11:0] ? image_528 : _GEN_9809; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9811 = 12'h211 == _T_121[11:0] ? image_529 : _GEN_9810; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9812 = 12'h212 == _T_121[11:0] ? image_530 : _GEN_9811; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9813 = 12'h213 == _T_121[11:0] ? image_531 : _GEN_9812; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9814 = 12'h214 == _T_121[11:0] ? image_532 : _GEN_9813; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9815 = 12'h215 == _T_121[11:0] ? image_533 : _GEN_9814; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9816 = 12'h216 == _T_121[11:0] ? image_534 : _GEN_9815; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9817 = 12'h217 == _T_121[11:0] ? image_535 : _GEN_9816; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9818 = 12'h218 == _T_121[11:0] ? image_536 : _GEN_9817; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9819 = 12'h219 == _T_121[11:0] ? image_537 : _GEN_9818; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9820 = 12'h21a == _T_121[11:0] ? image_538 : _GEN_9819; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9821 = 12'h21b == _T_121[11:0] ? image_539 : _GEN_9820; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9822 = 12'h21c == _T_121[11:0] ? image_540 : _GEN_9821; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9823 = 12'h21d == _T_121[11:0] ? image_541 : _GEN_9822; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9824 = 12'h21e == _T_121[11:0] ? image_542 : _GEN_9823; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9825 = 12'h21f == _T_121[11:0] ? image_543 : _GEN_9824; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9826 = 12'h220 == _T_121[11:0] ? image_544 : _GEN_9825; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9827 = 12'h221 == _T_121[11:0] ? image_545 : _GEN_9826; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9828 = 12'h222 == _T_121[11:0] ? image_546 : _GEN_9827; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9829 = 12'h223 == _T_121[11:0] ? image_547 : _GEN_9828; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9830 = 12'h224 == _T_121[11:0] ? image_548 : _GEN_9829; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9831 = 12'h225 == _T_121[11:0] ? image_549 : _GEN_9830; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9832 = 12'h226 == _T_121[11:0] ? image_550 : _GEN_9831; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9833 = 12'h227 == _T_121[11:0] ? image_551 : _GEN_9832; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9834 = 12'h228 == _T_121[11:0] ? image_552 : _GEN_9833; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9835 = 12'h229 == _T_121[11:0] ? image_553 : _GEN_9834; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9836 = 12'h22a == _T_121[11:0] ? image_554 : _GEN_9835; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9837 = 12'h22b == _T_121[11:0] ? image_555 : _GEN_9836; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9838 = 12'h22c == _T_121[11:0] ? image_556 : _GEN_9837; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9839 = 12'h22d == _T_121[11:0] ? image_557 : _GEN_9838; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9840 = 12'h22e == _T_121[11:0] ? image_558 : _GEN_9839; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9841 = 12'h22f == _T_121[11:0] ? image_559 : _GEN_9840; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9842 = 12'h230 == _T_121[11:0] ? image_560 : _GEN_9841; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9843 = 12'h231 == _T_121[11:0] ? image_561 : _GEN_9842; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9844 = 12'h232 == _T_121[11:0] ? image_562 : _GEN_9843; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9845 = 12'h233 == _T_121[11:0] ? image_563 : _GEN_9844; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9846 = 12'h234 == _T_121[11:0] ? image_564 : _GEN_9845; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9847 = 12'h235 == _T_121[11:0] ? image_565 : _GEN_9846; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9848 = 12'h236 == _T_121[11:0] ? image_566 : _GEN_9847; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9849 = 12'h237 == _T_121[11:0] ? 4'h0 : _GEN_9848; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9850 = 12'h238 == _T_121[11:0] ? 4'h0 : _GEN_9849; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9851 = 12'h239 == _T_121[11:0] ? 4'h0 : _GEN_9850; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9852 = 12'h23a == _T_121[11:0] ? 4'h0 : _GEN_9851; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9853 = 12'h23b == _T_121[11:0] ? image_571 : _GEN_9852; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9854 = 12'h23c == _T_121[11:0] ? image_572 : _GEN_9853; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9855 = 12'h23d == _T_121[11:0] ? image_573 : _GEN_9854; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9856 = 12'h23e == _T_121[11:0] ? image_574 : _GEN_9855; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9857 = 12'h23f == _T_121[11:0] ? 4'h0 : _GEN_9856; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9858 = 12'h240 == _T_121[11:0] ? 4'h0 : _GEN_9857; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9859 = 12'h241 == _T_121[11:0] ? 4'h0 : _GEN_9858; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9860 = 12'h242 == _T_121[11:0] ? image_578 : _GEN_9859; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9861 = 12'h243 == _T_121[11:0] ? image_579 : _GEN_9860; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9862 = 12'h244 == _T_121[11:0] ? image_580 : _GEN_9861; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9863 = 12'h245 == _T_121[11:0] ? image_581 : _GEN_9862; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9864 = 12'h246 == _T_121[11:0] ? image_582 : _GEN_9863; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9865 = 12'h247 == _T_121[11:0] ? image_583 : _GEN_9864; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9866 = 12'h248 == _T_121[11:0] ? image_584 : _GEN_9865; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9867 = 12'h249 == _T_121[11:0] ? image_585 : _GEN_9866; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9868 = 12'h24a == _T_121[11:0] ? image_586 : _GEN_9867; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9869 = 12'h24b == _T_121[11:0] ? image_587 : _GEN_9868; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9870 = 12'h24c == _T_121[11:0] ? image_588 : _GEN_9869; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9871 = 12'h24d == _T_121[11:0] ? image_589 : _GEN_9870; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9872 = 12'h24e == _T_121[11:0] ? image_590 : _GEN_9871; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9873 = 12'h24f == _T_121[11:0] ? image_591 : _GEN_9872; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9874 = 12'h250 == _T_121[11:0] ? image_592 : _GEN_9873; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9875 = 12'h251 == _T_121[11:0] ? image_593 : _GEN_9874; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9876 = 12'h252 == _T_121[11:0] ? image_594 : _GEN_9875; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9877 = 12'h253 == _T_121[11:0] ? image_595 : _GEN_9876; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9878 = 12'h254 == _T_121[11:0] ? image_596 : _GEN_9877; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9879 = 12'h255 == _T_121[11:0] ? image_597 : _GEN_9878; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9880 = 12'h256 == _T_121[11:0] ? image_598 : _GEN_9879; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9881 = 12'h257 == _T_121[11:0] ? image_599 : _GEN_9880; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9882 = 12'h258 == _T_121[11:0] ? image_600 : _GEN_9881; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9883 = 12'h259 == _T_121[11:0] ? image_601 : _GEN_9882; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9884 = 12'h25a == _T_121[11:0] ? image_602 : _GEN_9883; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9885 = 12'h25b == _T_121[11:0] ? image_603 : _GEN_9884; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9886 = 12'h25c == _T_121[11:0] ? image_604 : _GEN_9885; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9887 = 12'h25d == _T_121[11:0] ? image_605 : _GEN_9886; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9888 = 12'h25e == _T_121[11:0] ? image_606 : _GEN_9887; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9889 = 12'h25f == _T_121[11:0] ? image_607 : _GEN_9888; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9890 = 12'h260 == _T_121[11:0] ? 4'h0 : _GEN_9889; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9891 = 12'h261 == _T_121[11:0] ? 4'h0 : _GEN_9890; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9892 = 12'h262 == _T_121[11:0] ? 4'h0 : _GEN_9891; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9893 = 12'h263 == _T_121[11:0] ? 4'h0 : _GEN_9892; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9894 = 12'h264 == _T_121[11:0] ? 4'h0 : _GEN_9893; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9895 = 12'h265 == _T_121[11:0] ? 4'h0 : _GEN_9894; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9896 = 12'h266 == _T_121[11:0] ? image_614 : _GEN_9895; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9897 = 12'h267 == _T_121[11:0] ? image_615 : _GEN_9896; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9898 = 12'h268 == _T_121[11:0] ? image_616 : _GEN_9897; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9899 = 12'h269 == _T_121[11:0] ? image_617 : _GEN_9898; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9900 = 12'h26a == _T_121[11:0] ? image_618 : _GEN_9899; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9901 = 12'h26b == _T_121[11:0] ? image_619 : _GEN_9900; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9902 = 12'h26c == _T_121[11:0] ? image_620 : _GEN_9901; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9903 = 12'h26d == _T_121[11:0] ? image_621 : _GEN_9902; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9904 = 12'h26e == _T_121[11:0] ? image_622 : _GEN_9903; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9905 = 12'h26f == _T_121[11:0] ? image_623 : _GEN_9904; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9906 = 12'h270 == _T_121[11:0] ? image_624 : _GEN_9905; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9907 = 12'h271 == _T_121[11:0] ? image_625 : _GEN_9906; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9908 = 12'h272 == _T_121[11:0] ? image_626 : _GEN_9907; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9909 = 12'h273 == _T_121[11:0] ? image_627 : _GEN_9908; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9910 = 12'h274 == _T_121[11:0] ? image_628 : _GEN_9909; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9911 = 12'h275 == _T_121[11:0] ? 4'h0 : _GEN_9910; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9912 = 12'h276 == _T_121[11:0] ? 4'h0 : _GEN_9911; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9913 = 12'h277 == _T_121[11:0] ? 4'h0 : _GEN_9912; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9914 = 12'h278 == _T_121[11:0] ? 4'h0 : _GEN_9913; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9915 = 12'h279 == _T_121[11:0] ? 4'h0 : _GEN_9914; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9916 = 12'h27a == _T_121[11:0] ? 4'h0 : _GEN_9915; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9917 = 12'h27b == _T_121[11:0] ? 4'h0 : _GEN_9916; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9918 = 12'h27c == _T_121[11:0] ? image_636 : _GEN_9917; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9919 = 12'h27d == _T_121[11:0] ? image_637 : _GEN_9918; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9920 = 12'h27e == _T_121[11:0] ? image_638 : _GEN_9919; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9921 = 12'h27f == _T_121[11:0] ? image_639 : _GEN_9920; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9922 = 12'h280 == _T_121[11:0] ? 4'h0 : _GEN_9921; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9923 = 12'h281 == _T_121[11:0] ? 4'h0 : _GEN_9922; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9924 = 12'h282 == _T_121[11:0] ? image_642 : _GEN_9923; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9925 = 12'h283 == _T_121[11:0] ? image_643 : _GEN_9924; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9926 = 12'h284 == _T_121[11:0] ? image_644 : _GEN_9925; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9927 = 12'h285 == _T_121[11:0] ? image_645 : _GEN_9926; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9928 = 12'h286 == _T_121[11:0] ? image_646 : _GEN_9927; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9929 = 12'h287 == _T_121[11:0] ? image_647 : _GEN_9928; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9930 = 12'h288 == _T_121[11:0] ? image_648 : _GEN_9929; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9931 = 12'h289 == _T_121[11:0] ? image_649 : _GEN_9930; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9932 = 12'h28a == _T_121[11:0] ? image_650 : _GEN_9931; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9933 = 12'h28b == _T_121[11:0] ? image_651 : _GEN_9932; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9934 = 12'h28c == _T_121[11:0] ? image_652 : _GEN_9933; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9935 = 12'h28d == _T_121[11:0] ? image_653 : _GEN_9934; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9936 = 12'h28e == _T_121[11:0] ? image_654 : _GEN_9935; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9937 = 12'h28f == _T_121[11:0] ? image_655 : _GEN_9936; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9938 = 12'h290 == _T_121[11:0] ? image_656 : _GEN_9937; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9939 = 12'h291 == _T_121[11:0] ? image_657 : _GEN_9938; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9940 = 12'h292 == _T_121[11:0] ? image_658 : _GEN_9939; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9941 = 12'h293 == _T_121[11:0] ? image_659 : _GEN_9940; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9942 = 12'h294 == _T_121[11:0] ? image_660 : _GEN_9941; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9943 = 12'h295 == _T_121[11:0] ? image_661 : _GEN_9942; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9944 = 12'h296 == _T_121[11:0] ? image_662 : _GEN_9943; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9945 = 12'h297 == _T_121[11:0] ? image_663 : _GEN_9944; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9946 = 12'h298 == _T_121[11:0] ? image_664 : _GEN_9945; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9947 = 12'h299 == _T_121[11:0] ? image_665 : _GEN_9946; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9948 = 12'h29a == _T_121[11:0] ? image_666 : _GEN_9947; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9949 = 12'h29b == _T_121[11:0] ? image_667 : _GEN_9948; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9950 = 12'h29c == _T_121[11:0] ? image_668 : _GEN_9949; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9951 = 12'h29d == _T_121[11:0] ? image_669 : _GEN_9950; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9952 = 12'h29e == _T_121[11:0] ? image_670 : _GEN_9951; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9953 = 12'h29f == _T_121[11:0] ? 4'h0 : _GEN_9952; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9954 = 12'h2a0 == _T_121[11:0] ? 4'h0 : _GEN_9953; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9955 = 12'h2a1 == _T_121[11:0] ? 4'h0 : _GEN_9954; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9956 = 12'h2a2 == _T_121[11:0] ? 4'h0 : _GEN_9955; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9957 = 12'h2a3 == _T_121[11:0] ? 4'h0 : _GEN_9956; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9958 = 12'h2a4 == _T_121[11:0] ? 4'h0 : _GEN_9957; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9959 = 12'h2a5 == _T_121[11:0] ? 4'h0 : _GEN_9958; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9960 = 12'h2a6 == _T_121[11:0] ? 4'h0 : _GEN_9959; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9961 = 12'h2a7 == _T_121[11:0] ? image_679 : _GEN_9960; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9962 = 12'h2a8 == _T_121[11:0] ? image_680 : _GEN_9961; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9963 = 12'h2a9 == _T_121[11:0] ? image_681 : _GEN_9962; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9964 = 12'h2aa == _T_121[11:0] ? image_682 : _GEN_9963; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9965 = 12'h2ab == _T_121[11:0] ? image_683 : _GEN_9964; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9966 = 12'h2ac == _T_121[11:0] ? image_684 : _GEN_9965; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9967 = 12'h2ad == _T_121[11:0] ? image_685 : _GEN_9966; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9968 = 12'h2ae == _T_121[11:0] ? image_686 : _GEN_9967; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9969 = 12'h2af == _T_121[11:0] ? image_687 : _GEN_9968; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9970 = 12'h2b0 == _T_121[11:0] ? image_688 : _GEN_9969; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9971 = 12'h2b1 == _T_121[11:0] ? image_689 : _GEN_9970; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9972 = 12'h2b2 == _T_121[11:0] ? image_690 : _GEN_9971; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9973 = 12'h2b3 == _T_121[11:0] ? image_691 : _GEN_9972; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9974 = 12'h2b4 == _T_121[11:0] ? image_692 : _GEN_9973; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9975 = 12'h2b5 == _T_121[11:0] ? image_693 : _GEN_9974; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9976 = 12'h2b6 == _T_121[11:0] ? image_694 : _GEN_9975; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9977 = 12'h2b7 == _T_121[11:0] ? image_695 : _GEN_9976; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9978 = 12'h2b8 == _T_121[11:0] ? image_696 : _GEN_9977; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9979 = 12'h2b9 == _T_121[11:0] ? image_697 : _GEN_9978; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9980 = 12'h2ba == _T_121[11:0] ? image_698 : _GEN_9979; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9981 = 12'h2bb == _T_121[11:0] ? 4'h0 : _GEN_9980; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9982 = 12'h2bc == _T_121[11:0] ? 4'h0 : _GEN_9981; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9983 = 12'h2bd == _T_121[11:0] ? image_701 : _GEN_9982; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9984 = 12'h2be == _T_121[11:0] ? image_702 : _GEN_9983; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9985 = 12'h2bf == _T_121[11:0] ? image_703 : _GEN_9984; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9986 = 12'h2c0 == _T_121[11:0] ? 4'h0 : _GEN_9985; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9987 = 12'h2c1 == _T_121[11:0] ? image_705 : _GEN_9986; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9988 = 12'h2c2 == _T_121[11:0] ? image_706 : _GEN_9987; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9989 = 12'h2c3 == _T_121[11:0] ? image_707 : _GEN_9988; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9990 = 12'h2c4 == _T_121[11:0] ? image_708 : _GEN_9989; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9991 = 12'h2c5 == _T_121[11:0] ? image_709 : _GEN_9990; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9992 = 12'h2c6 == _T_121[11:0] ? image_710 : _GEN_9991; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9993 = 12'h2c7 == _T_121[11:0] ? image_711 : _GEN_9992; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9994 = 12'h2c8 == _T_121[11:0] ? image_712 : _GEN_9993; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9995 = 12'h2c9 == _T_121[11:0] ? image_713 : _GEN_9994; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9996 = 12'h2ca == _T_121[11:0] ? image_714 : _GEN_9995; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9997 = 12'h2cb == _T_121[11:0] ? image_715 : _GEN_9996; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9998 = 12'h2cc == _T_121[11:0] ? image_716 : _GEN_9997; // @[Filter.scala 138:46]
  wire [3:0] _GEN_9999 = 12'h2cd == _T_121[11:0] ? image_717 : _GEN_9998; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10000 = 12'h2ce == _T_121[11:0] ? image_718 : _GEN_9999; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10001 = 12'h2cf == _T_121[11:0] ? image_719 : _GEN_10000; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10002 = 12'h2d0 == _T_121[11:0] ? image_720 : _GEN_10001; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10003 = 12'h2d1 == _T_121[11:0] ? image_721 : _GEN_10002; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10004 = 12'h2d2 == _T_121[11:0] ? image_722 : _GEN_10003; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10005 = 12'h2d3 == _T_121[11:0] ? image_723 : _GEN_10004; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10006 = 12'h2d4 == _T_121[11:0] ? image_724 : _GEN_10005; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10007 = 12'h2d5 == _T_121[11:0] ? image_725 : _GEN_10006; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10008 = 12'h2d6 == _T_121[11:0] ? image_726 : _GEN_10007; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10009 = 12'h2d7 == _T_121[11:0] ? image_727 : _GEN_10008; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10010 = 12'h2d8 == _T_121[11:0] ? image_728 : _GEN_10009; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10011 = 12'h2d9 == _T_121[11:0] ? image_729 : _GEN_10010; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10012 = 12'h2da == _T_121[11:0] ? image_730 : _GEN_10011; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10013 = 12'h2db == _T_121[11:0] ? image_731 : _GEN_10012; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10014 = 12'h2dc == _T_121[11:0] ? image_732 : _GEN_10013; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10015 = 12'h2dd == _T_121[11:0] ? image_733 : _GEN_10014; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10016 = 12'h2de == _T_121[11:0] ? image_734 : _GEN_10015; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10017 = 12'h2df == _T_121[11:0] ? 4'h0 : _GEN_10016; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10018 = 12'h2e0 == _T_121[11:0] ? image_736 : _GEN_10017; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10019 = 12'h2e1 == _T_121[11:0] ? image_737 : _GEN_10018; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10020 = 12'h2e2 == _T_121[11:0] ? 4'h0 : _GEN_10019; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10021 = 12'h2e3 == _T_121[11:0] ? image_739 : _GEN_10020; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10022 = 12'h2e4 == _T_121[11:0] ? image_740 : _GEN_10021; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10023 = 12'h2e5 == _T_121[11:0] ? image_741 : _GEN_10022; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10024 = 12'h2e6 == _T_121[11:0] ? 4'h0 : _GEN_10023; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10025 = 12'h2e7 == _T_121[11:0] ? 4'h0 : _GEN_10024; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10026 = 12'h2e8 == _T_121[11:0] ? image_744 : _GEN_10025; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10027 = 12'h2e9 == _T_121[11:0] ? image_745 : _GEN_10026; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10028 = 12'h2ea == _T_121[11:0] ? image_746 : _GEN_10027; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10029 = 12'h2eb == _T_121[11:0] ? image_747 : _GEN_10028; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10030 = 12'h2ec == _T_121[11:0] ? image_748 : _GEN_10029; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10031 = 12'h2ed == _T_121[11:0] ? image_749 : _GEN_10030; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10032 = 12'h2ee == _T_121[11:0] ? image_750 : _GEN_10031; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10033 = 12'h2ef == _T_121[11:0] ? image_751 : _GEN_10032; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10034 = 12'h2f0 == _T_121[11:0] ? image_752 : _GEN_10033; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10035 = 12'h2f1 == _T_121[11:0] ? image_753 : _GEN_10034; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10036 = 12'h2f2 == _T_121[11:0] ? image_754 : _GEN_10035; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10037 = 12'h2f3 == _T_121[11:0] ? image_755 : _GEN_10036; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10038 = 12'h2f4 == _T_121[11:0] ? image_756 : _GEN_10037; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10039 = 12'h2f5 == _T_121[11:0] ? 4'h0 : _GEN_10038; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10040 = 12'h2f6 == _T_121[11:0] ? image_758 : _GEN_10039; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10041 = 12'h2f7 == _T_121[11:0] ? 4'h0 : _GEN_10040; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10042 = 12'h2f8 == _T_121[11:0] ? image_760 : _GEN_10041; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10043 = 12'h2f9 == _T_121[11:0] ? image_761 : _GEN_10042; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10044 = 12'h2fa == _T_121[11:0] ? image_762 : _GEN_10043; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10045 = 12'h2fb == _T_121[11:0] ? image_763 : _GEN_10044; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10046 = 12'h2fc == _T_121[11:0] ? 4'h0 : _GEN_10045; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10047 = 12'h2fd == _T_121[11:0] ? image_765 : _GEN_10046; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10048 = 12'h2fe == _T_121[11:0] ? image_766 : _GEN_10047; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10049 = 12'h2ff == _T_121[11:0] ? image_767 : _GEN_10048; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10050 = 12'h300 == _T_121[11:0] ? image_768 : _GEN_10049; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10051 = 12'h301 == _T_121[11:0] ? image_769 : _GEN_10050; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10052 = 12'h302 == _T_121[11:0] ? image_770 : _GEN_10051; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10053 = 12'h303 == _T_121[11:0] ? image_771 : _GEN_10052; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10054 = 12'h304 == _T_121[11:0] ? image_772 : _GEN_10053; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10055 = 12'h305 == _T_121[11:0] ? image_773 : _GEN_10054; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10056 = 12'h306 == _T_121[11:0] ? image_774 : _GEN_10055; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10057 = 12'h307 == _T_121[11:0] ? image_775 : _GEN_10056; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10058 = 12'h308 == _T_121[11:0] ? image_776 : _GEN_10057; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10059 = 12'h309 == _T_121[11:0] ? image_777 : _GEN_10058; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10060 = 12'h30a == _T_121[11:0] ? image_778 : _GEN_10059; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10061 = 12'h30b == _T_121[11:0] ? image_779 : _GEN_10060; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10062 = 12'h30c == _T_121[11:0] ? image_780 : _GEN_10061; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10063 = 12'h30d == _T_121[11:0] ? image_781 : _GEN_10062; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10064 = 12'h30e == _T_121[11:0] ? image_782 : _GEN_10063; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10065 = 12'h30f == _T_121[11:0] ? image_783 : _GEN_10064; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10066 = 12'h310 == _T_121[11:0] ? image_784 : _GEN_10065; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10067 = 12'h311 == _T_121[11:0] ? image_785 : _GEN_10066; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10068 = 12'h312 == _T_121[11:0] ? image_786 : _GEN_10067; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10069 = 12'h313 == _T_121[11:0] ? image_787 : _GEN_10068; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10070 = 12'h314 == _T_121[11:0] ? image_788 : _GEN_10069; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10071 = 12'h315 == _T_121[11:0] ? image_789 : _GEN_10070; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10072 = 12'h316 == _T_121[11:0] ? image_790 : _GEN_10071; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10073 = 12'h317 == _T_121[11:0] ? image_791 : _GEN_10072; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10074 = 12'h318 == _T_121[11:0] ? image_792 : _GEN_10073; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10075 = 12'h319 == _T_121[11:0] ? image_793 : _GEN_10074; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10076 = 12'h31a == _T_121[11:0] ? image_794 : _GEN_10075; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10077 = 12'h31b == _T_121[11:0] ? image_795 : _GEN_10076; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10078 = 12'h31c == _T_121[11:0] ? image_796 : _GEN_10077; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10079 = 12'h31d == _T_121[11:0] ? image_797 : _GEN_10078; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10080 = 12'h31e == _T_121[11:0] ? 4'h0 : _GEN_10079; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10081 = 12'h31f == _T_121[11:0] ? 4'h0 : _GEN_10080; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10082 = 12'h320 == _T_121[11:0] ? image_800 : _GEN_10081; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10083 = 12'h321 == _T_121[11:0] ? image_801 : _GEN_10082; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10084 = 12'h322 == _T_121[11:0] ? image_802 : _GEN_10083; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10085 = 12'h323 == _T_121[11:0] ? image_803 : _GEN_10084; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10086 = 12'h324 == _T_121[11:0] ? image_804 : _GEN_10085; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10087 = 12'h325 == _T_121[11:0] ? image_805 : _GEN_10086; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10088 = 12'h326 == _T_121[11:0] ? image_806 : _GEN_10087; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10089 = 12'h327 == _T_121[11:0] ? 4'h0 : _GEN_10088; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10090 = 12'h328 == _T_121[11:0] ? image_808 : _GEN_10089; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10091 = 12'h329 == _T_121[11:0] ? image_809 : _GEN_10090; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10092 = 12'h32a == _T_121[11:0] ? image_810 : _GEN_10091; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10093 = 12'h32b == _T_121[11:0] ? image_811 : _GEN_10092; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10094 = 12'h32c == _T_121[11:0] ? image_812 : _GEN_10093; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10095 = 12'h32d == _T_121[11:0] ? image_813 : _GEN_10094; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10096 = 12'h32e == _T_121[11:0] ? image_814 : _GEN_10095; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10097 = 12'h32f == _T_121[11:0] ? image_815 : _GEN_10096; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10098 = 12'h330 == _T_121[11:0] ? image_816 : _GEN_10097; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10099 = 12'h331 == _T_121[11:0] ? image_817 : _GEN_10098; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10100 = 12'h332 == _T_121[11:0] ? image_818 : _GEN_10099; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10101 = 12'h333 == _T_121[11:0] ? image_819 : _GEN_10100; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10102 = 12'h334 == _T_121[11:0] ? image_820 : _GEN_10101; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10103 = 12'h335 == _T_121[11:0] ? 4'h0 : _GEN_10102; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10104 = 12'h336 == _T_121[11:0] ? image_822 : _GEN_10103; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10105 = 12'h337 == _T_121[11:0] ? image_823 : _GEN_10104; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10106 = 12'h338 == _T_121[11:0] ? image_824 : _GEN_10105; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10107 = 12'h339 == _T_121[11:0] ? image_825 : _GEN_10106; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10108 = 12'h33a == _T_121[11:0] ? image_826 : _GEN_10107; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10109 = 12'h33b == _T_121[11:0] ? 4'h0 : _GEN_10108; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10110 = 12'h33c == _T_121[11:0] ? image_828 : _GEN_10109; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10111 = 12'h33d == _T_121[11:0] ? image_829 : _GEN_10110; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10112 = 12'h33e == _T_121[11:0] ? image_830 : _GEN_10111; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10113 = 12'h33f == _T_121[11:0] ? image_831 : _GEN_10112; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10114 = 12'h340 == _T_121[11:0] ? 4'h0 : _GEN_10113; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10115 = 12'h341 == _T_121[11:0] ? image_833 : _GEN_10114; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10116 = 12'h342 == _T_121[11:0] ? image_834 : _GEN_10115; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10117 = 12'h343 == _T_121[11:0] ? image_835 : _GEN_10116; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10118 = 12'h344 == _T_121[11:0] ? image_836 : _GEN_10117; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10119 = 12'h345 == _T_121[11:0] ? image_837 : _GEN_10118; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10120 = 12'h346 == _T_121[11:0] ? image_838 : _GEN_10119; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10121 = 12'h347 == _T_121[11:0] ? image_839 : _GEN_10120; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10122 = 12'h348 == _T_121[11:0] ? image_840 : _GEN_10121; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10123 = 12'h349 == _T_121[11:0] ? image_841 : _GEN_10122; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10124 = 12'h34a == _T_121[11:0] ? image_842 : _GEN_10123; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10125 = 12'h34b == _T_121[11:0] ? image_843 : _GEN_10124; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10126 = 12'h34c == _T_121[11:0] ? image_844 : _GEN_10125; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10127 = 12'h34d == _T_121[11:0] ? image_845 : _GEN_10126; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10128 = 12'h34e == _T_121[11:0] ? image_846 : _GEN_10127; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10129 = 12'h34f == _T_121[11:0] ? image_847 : _GEN_10128; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10130 = 12'h350 == _T_121[11:0] ? image_848 : _GEN_10129; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10131 = 12'h351 == _T_121[11:0] ? image_849 : _GEN_10130; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10132 = 12'h352 == _T_121[11:0] ? image_850 : _GEN_10131; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10133 = 12'h353 == _T_121[11:0] ? image_851 : _GEN_10132; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10134 = 12'h354 == _T_121[11:0] ? image_852 : _GEN_10133; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10135 = 12'h355 == _T_121[11:0] ? image_853 : _GEN_10134; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10136 = 12'h356 == _T_121[11:0] ? image_854 : _GEN_10135; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10137 = 12'h357 == _T_121[11:0] ? image_855 : _GEN_10136; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10138 = 12'h358 == _T_121[11:0] ? image_856 : _GEN_10137; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10139 = 12'h359 == _T_121[11:0] ? image_857 : _GEN_10138; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10140 = 12'h35a == _T_121[11:0] ? image_858 : _GEN_10139; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10141 = 12'h35b == _T_121[11:0] ? image_859 : _GEN_10140; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10142 = 12'h35c == _T_121[11:0] ? image_860 : _GEN_10141; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10143 = 12'h35d == _T_121[11:0] ? image_861 : _GEN_10142; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10144 = 12'h35e == _T_121[11:0] ? image_862 : _GEN_10143; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10145 = 12'h35f == _T_121[11:0] ? 4'h0 : _GEN_10144; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10146 = 12'h360 == _T_121[11:0] ? 4'h0 : _GEN_10145; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10147 = 12'h361 == _T_121[11:0] ? image_865 : _GEN_10146; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10148 = 12'h362 == _T_121[11:0] ? image_866 : _GEN_10147; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10149 = 12'h363 == _T_121[11:0] ? image_867 : _GEN_10148; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10150 = 12'h364 == _T_121[11:0] ? image_868 : _GEN_10149; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10151 = 12'h365 == _T_121[11:0] ? image_869 : _GEN_10150; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10152 = 12'h366 == _T_121[11:0] ? 4'h0 : _GEN_10151; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10153 = 12'h367 == _T_121[11:0] ? 4'h0 : _GEN_10152; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10154 = 12'h368 == _T_121[11:0] ? image_872 : _GEN_10153; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10155 = 12'h369 == _T_121[11:0] ? image_873 : _GEN_10154; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10156 = 12'h36a == _T_121[11:0] ? image_874 : _GEN_10155; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10157 = 12'h36b == _T_121[11:0] ? image_875 : _GEN_10156; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10158 = 12'h36c == _T_121[11:0] ? image_876 : _GEN_10157; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10159 = 12'h36d == _T_121[11:0] ? image_877 : _GEN_10158; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10160 = 12'h36e == _T_121[11:0] ? image_878 : _GEN_10159; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10161 = 12'h36f == _T_121[11:0] ? image_879 : _GEN_10160; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10162 = 12'h370 == _T_121[11:0] ? image_880 : _GEN_10161; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10163 = 12'h371 == _T_121[11:0] ? image_881 : _GEN_10162; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10164 = 12'h372 == _T_121[11:0] ? image_882 : _GEN_10163; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10165 = 12'h373 == _T_121[11:0] ? image_883 : _GEN_10164; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10166 = 12'h374 == _T_121[11:0] ? image_884 : _GEN_10165; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10167 = 12'h375 == _T_121[11:0] ? image_885 : _GEN_10166; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10168 = 12'h376 == _T_121[11:0] ? 4'h0 : _GEN_10167; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10169 = 12'h377 == _T_121[11:0] ? 4'h0 : _GEN_10168; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10170 = 12'h378 == _T_121[11:0] ? 4'h0 : _GEN_10169; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10171 = 12'h379 == _T_121[11:0] ? 4'h0 : _GEN_10170; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10172 = 12'h37a == _T_121[11:0] ? 4'h0 : _GEN_10171; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10173 = 12'h37b == _T_121[11:0] ? image_891 : _GEN_10172; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10174 = 12'h37c == _T_121[11:0] ? image_892 : _GEN_10173; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10175 = 12'h37d == _T_121[11:0] ? image_893 : _GEN_10174; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10176 = 12'h37e == _T_121[11:0] ? image_894 : _GEN_10175; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10177 = 12'h37f == _T_121[11:0] ? image_895 : _GEN_10176; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10178 = 12'h380 == _T_121[11:0] ? 4'h0 : _GEN_10177; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10179 = 12'h381 == _T_121[11:0] ? image_897 : _GEN_10178; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10180 = 12'h382 == _T_121[11:0] ? image_898 : _GEN_10179; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10181 = 12'h383 == _T_121[11:0] ? image_899 : _GEN_10180; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10182 = 12'h384 == _T_121[11:0] ? image_900 : _GEN_10181; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10183 = 12'h385 == _T_121[11:0] ? image_901 : _GEN_10182; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10184 = 12'h386 == _T_121[11:0] ? image_902 : _GEN_10183; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10185 = 12'h387 == _T_121[11:0] ? image_903 : _GEN_10184; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10186 = 12'h388 == _T_121[11:0] ? image_904 : _GEN_10185; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10187 = 12'h389 == _T_121[11:0] ? image_905 : _GEN_10186; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10188 = 12'h38a == _T_121[11:0] ? image_906 : _GEN_10187; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10189 = 12'h38b == _T_121[11:0] ? image_907 : _GEN_10188; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10190 = 12'h38c == _T_121[11:0] ? image_908 : _GEN_10189; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10191 = 12'h38d == _T_121[11:0] ? image_909 : _GEN_10190; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10192 = 12'h38e == _T_121[11:0] ? image_910 : _GEN_10191; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10193 = 12'h38f == _T_121[11:0] ? image_911 : _GEN_10192; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10194 = 12'h390 == _T_121[11:0] ? image_912 : _GEN_10193; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10195 = 12'h391 == _T_121[11:0] ? image_913 : _GEN_10194; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10196 = 12'h392 == _T_121[11:0] ? image_914 : _GEN_10195; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10197 = 12'h393 == _T_121[11:0] ? image_915 : _GEN_10196; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10198 = 12'h394 == _T_121[11:0] ? image_916 : _GEN_10197; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10199 = 12'h395 == _T_121[11:0] ? image_917 : _GEN_10198; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10200 = 12'h396 == _T_121[11:0] ? image_918 : _GEN_10199; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10201 = 12'h397 == _T_121[11:0] ? image_919 : _GEN_10200; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10202 = 12'h398 == _T_121[11:0] ? image_920 : _GEN_10201; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10203 = 12'h399 == _T_121[11:0] ? image_921 : _GEN_10202; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10204 = 12'h39a == _T_121[11:0] ? image_922 : _GEN_10203; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10205 = 12'h39b == _T_121[11:0] ? image_923 : _GEN_10204; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10206 = 12'h39c == _T_121[11:0] ? image_924 : _GEN_10205; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10207 = 12'h39d == _T_121[11:0] ? image_925 : _GEN_10206; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10208 = 12'h39e == _T_121[11:0] ? image_926 : _GEN_10207; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10209 = 12'h39f == _T_121[11:0] ? image_927 : _GEN_10208; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10210 = 12'h3a0 == _T_121[11:0] ? 4'h0 : _GEN_10209; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10211 = 12'h3a1 == _T_121[11:0] ? image_929 : _GEN_10210; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10212 = 12'h3a2 == _T_121[11:0] ? image_930 : _GEN_10211; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10213 = 12'h3a3 == _T_121[11:0] ? 4'h0 : _GEN_10212; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10214 = 12'h3a4 == _T_121[11:0] ? 4'h0 : _GEN_10213; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10215 = 12'h3a5 == _T_121[11:0] ? 4'h0 : _GEN_10214; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10216 = 12'h3a6 == _T_121[11:0] ? 4'h0 : _GEN_10215; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10217 = 12'h3a7 == _T_121[11:0] ? image_935 : _GEN_10216; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10218 = 12'h3a8 == _T_121[11:0] ? image_936 : _GEN_10217; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10219 = 12'h3a9 == _T_121[11:0] ? image_937 : _GEN_10218; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10220 = 12'h3aa == _T_121[11:0] ? image_938 : _GEN_10219; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10221 = 12'h3ab == _T_121[11:0] ? image_939 : _GEN_10220; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10222 = 12'h3ac == _T_121[11:0] ? image_940 : _GEN_10221; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10223 = 12'h3ad == _T_121[11:0] ? image_941 : _GEN_10222; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10224 = 12'h3ae == _T_121[11:0] ? image_942 : _GEN_10223; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10225 = 12'h3af == _T_121[11:0] ? image_943 : _GEN_10224; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10226 = 12'h3b0 == _T_121[11:0] ? image_944 : _GEN_10225; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10227 = 12'h3b1 == _T_121[11:0] ? image_945 : _GEN_10226; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10228 = 12'h3b2 == _T_121[11:0] ? image_946 : _GEN_10227; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10229 = 12'h3b3 == _T_121[11:0] ? image_947 : _GEN_10228; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10230 = 12'h3b4 == _T_121[11:0] ? image_948 : _GEN_10229; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10231 = 12'h3b5 == _T_121[11:0] ? image_949 : _GEN_10230; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10232 = 12'h3b6 == _T_121[11:0] ? image_950 : _GEN_10231; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10233 = 12'h3b7 == _T_121[11:0] ? image_951 : _GEN_10232; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10234 = 12'h3b8 == _T_121[11:0] ? image_952 : _GEN_10233; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10235 = 12'h3b9 == _T_121[11:0] ? image_953 : _GEN_10234; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10236 = 12'h3ba == _T_121[11:0] ? image_954 : _GEN_10235; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10237 = 12'h3bb == _T_121[11:0] ? image_955 : _GEN_10236; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10238 = 12'h3bc == _T_121[11:0] ? image_956 : _GEN_10237; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10239 = 12'h3bd == _T_121[11:0] ? image_957 : _GEN_10238; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10240 = 12'h3be == _T_121[11:0] ? image_958 : _GEN_10239; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10241 = 12'h3bf == _T_121[11:0] ? image_959 : _GEN_10240; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10242 = 12'h3c0 == _T_121[11:0] ? 4'h0 : _GEN_10241; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10243 = 12'h3c1 == _T_121[11:0] ? image_961 : _GEN_10242; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10244 = 12'h3c2 == _T_121[11:0] ? image_962 : _GEN_10243; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10245 = 12'h3c3 == _T_121[11:0] ? image_963 : _GEN_10244; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10246 = 12'h3c4 == _T_121[11:0] ? image_964 : _GEN_10245; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10247 = 12'h3c5 == _T_121[11:0] ? image_965 : _GEN_10246; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10248 = 12'h3c6 == _T_121[11:0] ? image_966 : _GEN_10247; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10249 = 12'h3c7 == _T_121[11:0] ? image_967 : _GEN_10248; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10250 = 12'h3c8 == _T_121[11:0] ? image_968 : _GEN_10249; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10251 = 12'h3c9 == _T_121[11:0] ? image_969 : _GEN_10250; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10252 = 12'h3ca == _T_121[11:0] ? image_970 : _GEN_10251; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10253 = 12'h3cb == _T_121[11:0] ? image_971 : _GEN_10252; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10254 = 12'h3cc == _T_121[11:0] ? image_972 : _GEN_10253; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10255 = 12'h3cd == _T_121[11:0] ? image_973 : _GEN_10254; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10256 = 12'h3ce == _T_121[11:0] ? image_974 : _GEN_10255; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10257 = 12'h3cf == _T_121[11:0] ? image_975 : _GEN_10256; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10258 = 12'h3d0 == _T_121[11:0] ? image_976 : _GEN_10257; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10259 = 12'h3d1 == _T_121[11:0] ? image_977 : _GEN_10258; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10260 = 12'h3d2 == _T_121[11:0] ? image_978 : _GEN_10259; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10261 = 12'h3d3 == _T_121[11:0] ? image_979 : _GEN_10260; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10262 = 12'h3d4 == _T_121[11:0] ? image_980 : _GEN_10261; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10263 = 12'h3d5 == _T_121[11:0] ? image_981 : _GEN_10262; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10264 = 12'h3d6 == _T_121[11:0] ? image_982 : _GEN_10263; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10265 = 12'h3d7 == _T_121[11:0] ? image_983 : _GEN_10264; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10266 = 12'h3d8 == _T_121[11:0] ? image_984 : _GEN_10265; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10267 = 12'h3d9 == _T_121[11:0] ? image_985 : _GEN_10266; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10268 = 12'h3da == _T_121[11:0] ? image_986 : _GEN_10267; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10269 = 12'h3db == _T_121[11:0] ? image_987 : _GEN_10268; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10270 = 12'h3dc == _T_121[11:0] ? image_988 : _GEN_10269; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10271 = 12'h3dd == _T_121[11:0] ? image_989 : _GEN_10270; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10272 = 12'h3de == _T_121[11:0] ? image_990 : _GEN_10271; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10273 = 12'h3df == _T_121[11:0] ? image_991 : _GEN_10272; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10274 = 12'h3e0 == _T_121[11:0] ? image_992 : _GEN_10273; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10275 = 12'h3e1 == _T_121[11:0] ? 4'h0 : _GEN_10274; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10276 = 12'h3e2 == _T_121[11:0] ? 4'h0 : _GEN_10275; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10277 = 12'h3e3 == _T_121[11:0] ? 4'h0 : _GEN_10276; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10278 = 12'h3e4 == _T_121[11:0] ? 4'h0 : _GEN_10277; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10279 = 12'h3e5 == _T_121[11:0] ? image_997 : _GEN_10278; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10280 = 12'h3e6 == _T_121[11:0] ? image_998 : _GEN_10279; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10281 = 12'h3e7 == _T_121[11:0] ? image_999 : _GEN_10280; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10282 = 12'h3e8 == _T_121[11:0] ? image_1000 : _GEN_10281; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10283 = 12'h3e9 == _T_121[11:0] ? image_1001 : _GEN_10282; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10284 = 12'h3ea == _T_121[11:0] ? image_1002 : _GEN_10283; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10285 = 12'h3eb == _T_121[11:0] ? image_1003 : _GEN_10284; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10286 = 12'h3ec == _T_121[11:0] ? image_1004 : _GEN_10285; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10287 = 12'h3ed == _T_121[11:0] ? image_1005 : _GEN_10286; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10288 = 12'h3ee == _T_121[11:0] ? image_1006 : _GEN_10287; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10289 = 12'h3ef == _T_121[11:0] ? image_1007 : _GEN_10288; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10290 = 12'h3f0 == _T_121[11:0] ? image_1008 : _GEN_10289; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10291 = 12'h3f1 == _T_121[11:0] ? image_1009 : _GEN_10290; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10292 = 12'h3f2 == _T_121[11:0] ? image_1010 : _GEN_10291; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10293 = 12'h3f3 == _T_121[11:0] ? image_1011 : _GEN_10292; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10294 = 12'h3f4 == _T_121[11:0] ? image_1012 : _GEN_10293; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10295 = 12'h3f5 == _T_121[11:0] ? image_1013 : _GEN_10294; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10296 = 12'h3f6 == _T_121[11:0] ? image_1014 : _GEN_10295; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10297 = 12'h3f7 == _T_121[11:0] ? image_1015 : _GEN_10296; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10298 = 12'h3f8 == _T_121[11:0] ? image_1016 : _GEN_10297; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10299 = 12'h3f9 == _T_121[11:0] ? image_1017 : _GEN_10298; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10300 = 12'h3fa == _T_121[11:0] ? image_1018 : _GEN_10299; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10301 = 12'h3fb == _T_121[11:0] ? image_1019 : _GEN_10300; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10302 = 12'h3fc == _T_121[11:0] ? image_1020 : _GEN_10301; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10303 = 12'h3fd == _T_121[11:0] ? 4'h0 : _GEN_10302; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10304 = 12'h3fe == _T_121[11:0] ? 4'h0 : _GEN_10303; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10305 = 12'h3ff == _T_121[11:0] ? 4'h0 : _GEN_10304; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10306 = 12'h400 == _T_121[11:0] ? image_1024 : _GEN_10305; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10307 = 12'h401 == _T_121[11:0] ? image_1025 : _GEN_10306; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10308 = 12'h402 == _T_121[11:0] ? image_1026 : _GEN_10307; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10309 = 12'h403 == _T_121[11:0] ? image_1027 : _GEN_10308; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10310 = 12'h404 == _T_121[11:0] ? image_1028 : _GEN_10309; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10311 = 12'h405 == _T_121[11:0] ? image_1029 : _GEN_10310; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10312 = 12'h406 == _T_121[11:0] ? image_1030 : _GEN_10311; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10313 = 12'h407 == _T_121[11:0] ? image_1031 : _GEN_10312; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10314 = 12'h408 == _T_121[11:0] ? image_1032 : _GEN_10313; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10315 = 12'h409 == _T_121[11:0] ? image_1033 : _GEN_10314; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10316 = 12'h40a == _T_121[11:0] ? image_1034 : _GEN_10315; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10317 = 12'h40b == _T_121[11:0] ? image_1035 : _GEN_10316; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10318 = 12'h40c == _T_121[11:0] ? image_1036 : _GEN_10317; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10319 = 12'h40d == _T_121[11:0] ? image_1037 : _GEN_10318; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10320 = 12'h40e == _T_121[11:0] ? image_1038 : _GEN_10319; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10321 = 12'h40f == _T_121[11:0] ? image_1039 : _GEN_10320; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10322 = 12'h410 == _T_121[11:0] ? image_1040 : _GEN_10321; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10323 = 12'h411 == _T_121[11:0] ? image_1041 : _GEN_10322; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10324 = 12'h412 == _T_121[11:0] ? image_1042 : _GEN_10323; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10325 = 12'h413 == _T_121[11:0] ? image_1043 : _GEN_10324; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10326 = 12'h414 == _T_121[11:0] ? image_1044 : _GEN_10325; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10327 = 12'h415 == _T_121[11:0] ? image_1045 : _GEN_10326; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10328 = 12'h416 == _T_121[11:0] ? image_1046 : _GEN_10327; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10329 = 12'h417 == _T_121[11:0] ? image_1047 : _GEN_10328; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10330 = 12'h418 == _T_121[11:0] ? image_1048 : _GEN_10329; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10331 = 12'h419 == _T_121[11:0] ? image_1049 : _GEN_10330; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10332 = 12'h41a == _T_121[11:0] ? image_1050 : _GEN_10331; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10333 = 12'h41b == _T_121[11:0] ? image_1051 : _GEN_10332; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10334 = 12'h41c == _T_121[11:0] ? image_1052 : _GEN_10333; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10335 = 12'h41d == _T_121[11:0] ? image_1053 : _GEN_10334; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10336 = 12'h41e == _T_121[11:0] ? image_1054 : _GEN_10335; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10337 = 12'h41f == _T_121[11:0] ? image_1055 : _GEN_10336; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10338 = 12'h420 == _T_121[11:0] ? image_1056 : _GEN_10337; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10339 = 12'h421 == _T_121[11:0] ? image_1057 : _GEN_10338; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10340 = 12'h422 == _T_121[11:0] ? image_1058 : _GEN_10339; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10341 = 12'h423 == _T_121[11:0] ? image_1059 : _GEN_10340; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10342 = 12'h424 == _T_121[11:0] ? image_1060 : _GEN_10341; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10343 = 12'h425 == _T_121[11:0] ? image_1061 : _GEN_10342; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10344 = 12'h426 == _T_121[11:0] ? image_1062 : _GEN_10343; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10345 = 12'h427 == _T_121[11:0] ? image_1063 : _GEN_10344; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10346 = 12'h428 == _T_121[11:0] ? image_1064 : _GEN_10345; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10347 = 12'h429 == _T_121[11:0] ? image_1065 : _GEN_10346; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10348 = 12'h42a == _T_121[11:0] ? image_1066 : _GEN_10347; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10349 = 12'h42b == _T_121[11:0] ? image_1067 : _GEN_10348; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10350 = 12'h42c == _T_121[11:0] ? image_1068 : _GEN_10349; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10351 = 12'h42d == _T_121[11:0] ? image_1069 : _GEN_10350; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10352 = 12'h42e == _T_121[11:0] ? image_1070 : _GEN_10351; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10353 = 12'h42f == _T_121[11:0] ? image_1071 : _GEN_10352; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10354 = 12'h430 == _T_121[11:0] ? image_1072 : _GEN_10353; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10355 = 12'h431 == _T_121[11:0] ? image_1073 : _GEN_10354; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10356 = 12'h432 == _T_121[11:0] ? image_1074 : _GEN_10355; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10357 = 12'h433 == _T_121[11:0] ? image_1075 : _GEN_10356; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10358 = 12'h434 == _T_121[11:0] ? image_1076 : _GEN_10357; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10359 = 12'h435 == _T_121[11:0] ? image_1077 : _GEN_10358; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10360 = 12'h436 == _T_121[11:0] ? image_1078 : _GEN_10359; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10361 = 12'h437 == _T_121[11:0] ? image_1079 : _GEN_10360; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10362 = 12'h438 == _T_121[11:0] ? image_1080 : _GEN_10361; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10363 = 12'h439 == _T_121[11:0] ? image_1081 : _GEN_10362; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10364 = 12'h43a == _T_121[11:0] ? image_1082 : _GEN_10363; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10365 = 12'h43b == _T_121[11:0] ? image_1083 : _GEN_10364; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10366 = 12'h43c == _T_121[11:0] ? image_1084 : _GEN_10365; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10367 = 12'h43d == _T_121[11:0] ? image_1085 : _GEN_10366; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10368 = 12'h43e == _T_121[11:0] ? 4'h0 : _GEN_10367; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10369 = 12'h43f == _T_121[11:0] ? 4'h0 : _GEN_10368; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10370 = 12'h440 == _T_121[11:0] ? image_1088 : _GEN_10369; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10371 = 12'h441 == _T_121[11:0] ? image_1089 : _GEN_10370; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10372 = 12'h442 == _T_121[11:0] ? image_1090 : _GEN_10371; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10373 = 12'h443 == _T_121[11:0] ? image_1091 : _GEN_10372; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10374 = 12'h444 == _T_121[11:0] ? image_1092 : _GEN_10373; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10375 = 12'h445 == _T_121[11:0] ? image_1093 : _GEN_10374; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10376 = 12'h446 == _T_121[11:0] ? image_1094 : _GEN_10375; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10377 = 12'h447 == _T_121[11:0] ? image_1095 : _GEN_10376; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10378 = 12'h448 == _T_121[11:0] ? image_1096 : _GEN_10377; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10379 = 12'h449 == _T_121[11:0] ? image_1097 : _GEN_10378; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10380 = 12'h44a == _T_121[11:0] ? image_1098 : _GEN_10379; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10381 = 12'h44b == _T_121[11:0] ? image_1099 : _GEN_10380; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10382 = 12'h44c == _T_121[11:0] ? image_1100 : _GEN_10381; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10383 = 12'h44d == _T_121[11:0] ? image_1101 : _GEN_10382; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10384 = 12'h44e == _T_121[11:0] ? image_1102 : _GEN_10383; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10385 = 12'h44f == _T_121[11:0] ? image_1103 : _GEN_10384; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10386 = 12'h450 == _T_121[11:0] ? image_1104 : _GEN_10385; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10387 = 12'h451 == _T_121[11:0] ? image_1105 : _GEN_10386; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10388 = 12'h452 == _T_121[11:0] ? image_1106 : _GEN_10387; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10389 = 12'h453 == _T_121[11:0] ? image_1107 : _GEN_10388; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10390 = 12'h454 == _T_121[11:0] ? image_1108 : _GEN_10389; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10391 = 12'h455 == _T_121[11:0] ? image_1109 : _GEN_10390; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10392 = 12'h456 == _T_121[11:0] ? image_1110 : _GEN_10391; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10393 = 12'h457 == _T_121[11:0] ? image_1111 : _GEN_10392; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10394 = 12'h458 == _T_121[11:0] ? image_1112 : _GEN_10393; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10395 = 12'h459 == _T_121[11:0] ? image_1113 : _GEN_10394; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10396 = 12'h45a == _T_121[11:0] ? image_1114 : _GEN_10395; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10397 = 12'h45b == _T_121[11:0] ? image_1115 : _GEN_10396; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10398 = 12'h45c == _T_121[11:0] ? image_1116 : _GEN_10397; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10399 = 12'h45d == _T_121[11:0] ? image_1117 : _GEN_10398; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10400 = 12'h45e == _T_121[11:0] ? image_1118 : _GEN_10399; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10401 = 12'h45f == _T_121[11:0] ? image_1119 : _GEN_10400; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10402 = 12'h460 == _T_121[11:0] ? image_1120 : _GEN_10401; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10403 = 12'h461 == _T_121[11:0] ? image_1121 : _GEN_10402; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10404 = 12'h462 == _T_121[11:0] ? image_1122 : _GEN_10403; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10405 = 12'h463 == _T_121[11:0] ? image_1123 : _GEN_10404; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10406 = 12'h464 == _T_121[11:0] ? image_1124 : _GEN_10405; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10407 = 12'h465 == _T_121[11:0] ? image_1125 : _GEN_10406; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10408 = 12'h466 == _T_121[11:0] ? image_1126 : _GEN_10407; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10409 = 12'h467 == _T_121[11:0] ? image_1127 : _GEN_10408; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10410 = 12'h468 == _T_121[11:0] ? image_1128 : _GEN_10409; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10411 = 12'h469 == _T_121[11:0] ? image_1129 : _GEN_10410; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10412 = 12'h46a == _T_121[11:0] ? image_1130 : _GEN_10411; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10413 = 12'h46b == _T_121[11:0] ? image_1131 : _GEN_10412; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10414 = 12'h46c == _T_121[11:0] ? image_1132 : _GEN_10413; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10415 = 12'h46d == _T_121[11:0] ? image_1133 : _GEN_10414; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10416 = 12'h46e == _T_121[11:0] ? image_1134 : _GEN_10415; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10417 = 12'h46f == _T_121[11:0] ? image_1135 : _GEN_10416; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10418 = 12'h470 == _T_121[11:0] ? image_1136 : _GEN_10417; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10419 = 12'h471 == _T_121[11:0] ? image_1137 : _GEN_10418; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10420 = 12'h472 == _T_121[11:0] ? image_1138 : _GEN_10419; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10421 = 12'h473 == _T_121[11:0] ? image_1139 : _GEN_10420; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10422 = 12'h474 == _T_121[11:0] ? image_1140 : _GEN_10421; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10423 = 12'h475 == _T_121[11:0] ? image_1141 : _GEN_10422; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10424 = 12'h476 == _T_121[11:0] ? image_1142 : _GEN_10423; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10425 = 12'h477 == _T_121[11:0] ? image_1143 : _GEN_10424; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10426 = 12'h478 == _T_121[11:0] ? image_1144 : _GEN_10425; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10427 = 12'h479 == _T_121[11:0] ? image_1145 : _GEN_10426; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10428 = 12'h47a == _T_121[11:0] ? image_1146 : _GEN_10427; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10429 = 12'h47b == _T_121[11:0] ? image_1147 : _GEN_10428; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10430 = 12'h47c == _T_121[11:0] ? image_1148 : _GEN_10429; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10431 = 12'h47d == _T_121[11:0] ? 4'h0 : _GEN_10430; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10432 = 12'h47e == _T_121[11:0] ? 4'h0 : _GEN_10431; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10433 = 12'h47f == _T_121[11:0] ? 4'h0 : _GEN_10432; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10434 = 12'h480 == _T_121[11:0] ? image_1152 : _GEN_10433; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10435 = 12'h481 == _T_121[11:0] ? image_1153 : _GEN_10434; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10436 = 12'h482 == _T_121[11:0] ? image_1154 : _GEN_10435; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10437 = 12'h483 == _T_121[11:0] ? image_1155 : _GEN_10436; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10438 = 12'h484 == _T_121[11:0] ? image_1156 : _GEN_10437; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10439 = 12'h485 == _T_121[11:0] ? image_1157 : _GEN_10438; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10440 = 12'h486 == _T_121[11:0] ? image_1158 : _GEN_10439; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10441 = 12'h487 == _T_121[11:0] ? image_1159 : _GEN_10440; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10442 = 12'h488 == _T_121[11:0] ? image_1160 : _GEN_10441; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10443 = 12'h489 == _T_121[11:0] ? image_1161 : _GEN_10442; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10444 = 12'h48a == _T_121[11:0] ? image_1162 : _GEN_10443; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10445 = 12'h48b == _T_121[11:0] ? image_1163 : _GEN_10444; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10446 = 12'h48c == _T_121[11:0] ? image_1164 : _GEN_10445; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10447 = 12'h48d == _T_121[11:0] ? image_1165 : _GEN_10446; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10448 = 12'h48e == _T_121[11:0] ? image_1166 : _GEN_10447; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10449 = 12'h48f == _T_121[11:0] ? image_1167 : _GEN_10448; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10450 = 12'h490 == _T_121[11:0] ? image_1168 : _GEN_10449; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10451 = 12'h491 == _T_121[11:0] ? image_1169 : _GEN_10450; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10452 = 12'h492 == _T_121[11:0] ? image_1170 : _GEN_10451; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10453 = 12'h493 == _T_121[11:0] ? image_1171 : _GEN_10452; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10454 = 12'h494 == _T_121[11:0] ? image_1172 : _GEN_10453; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10455 = 12'h495 == _T_121[11:0] ? image_1173 : _GEN_10454; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10456 = 12'h496 == _T_121[11:0] ? image_1174 : _GEN_10455; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10457 = 12'h497 == _T_121[11:0] ? image_1175 : _GEN_10456; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10458 = 12'h498 == _T_121[11:0] ? image_1176 : _GEN_10457; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10459 = 12'h499 == _T_121[11:0] ? image_1177 : _GEN_10458; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10460 = 12'h49a == _T_121[11:0] ? image_1178 : _GEN_10459; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10461 = 12'h49b == _T_121[11:0] ? image_1179 : _GEN_10460; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10462 = 12'h49c == _T_121[11:0] ? image_1180 : _GEN_10461; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10463 = 12'h49d == _T_121[11:0] ? image_1181 : _GEN_10462; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10464 = 12'h49e == _T_121[11:0] ? image_1182 : _GEN_10463; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10465 = 12'h49f == _T_121[11:0] ? image_1183 : _GEN_10464; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10466 = 12'h4a0 == _T_121[11:0] ? image_1184 : _GEN_10465; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10467 = 12'h4a1 == _T_121[11:0] ? image_1185 : _GEN_10466; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10468 = 12'h4a2 == _T_121[11:0] ? image_1186 : _GEN_10467; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10469 = 12'h4a3 == _T_121[11:0] ? image_1187 : _GEN_10468; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10470 = 12'h4a4 == _T_121[11:0] ? image_1188 : _GEN_10469; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10471 = 12'h4a5 == _T_121[11:0] ? image_1189 : _GEN_10470; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10472 = 12'h4a6 == _T_121[11:0] ? image_1190 : _GEN_10471; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10473 = 12'h4a7 == _T_121[11:0] ? image_1191 : _GEN_10472; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10474 = 12'h4a8 == _T_121[11:0] ? image_1192 : _GEN_10473; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10475 = 12'h4a9 == _T_121[11:0] ? image_1193 : _GEN_10474; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10476 = 12'h4aa == _T_121[11:0] ? image_1194 : _GEN_10475; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10477 = 12'h4ab == _T_121[11:0] ? image_1195 : _GEN_10476; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10478 = 12'h4ac == _T_121[11:0] ? image_1196 : _GEN_10477; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10479 = 12'h4ad == _T_121[11:0] ? image_1197 : _GEN_10478; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10480 = 12'h4ae == _T_121[11:0] ? image_1198 : _GEN_10479; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10481 = 12'h4af == _T_121[11:0] ? image_1199 : _GEN_10480; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10482 = 12'h4b0 == _T_121[11:0] ? image_1200 : _GEN_10481; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10483 = 12'h4b1 == _T_121[11:0] ? image_1201 : _GEN_10482; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10484 = 12'h4b2 == _T_121[11:0] ? image_1202 : _GEN_10483; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10485 = 12'h4b3 == _T_121[11:0] ? image_1203 : _GEN_10484; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10486 = 12'h4b4 == _T_121[11:0] ? image_1204 : _GEN_10485; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10487 = 12'h4b5 == _T_121[11:0] ? image_1205 : _GEN_10486; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10488 = 12'h4b6 == _T_121[11:0] ? image_1206 : _GEN_10487; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10489 = 12'h4b7 == _T_121[11:0] ? image_1207 : _GEN_10488; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10490 = 12'h4b8 == _T_121[11:0] ? image_1208 : _GEN_10489; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10491 = 12'h4b9 == _T_121[11:0] ? 4'h0 : _GEN_10490; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10492 = 12'h4ba == _T_121[11:0] ? 4'h0 : _GEN_10491; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10493 = 12'h4bb == _T_121[11:0] ? 4'h0 : _GEN_10492; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10494 = 12'h4bc == _T_121[11:0] ? 4'h0 : _GEN_10493; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10495 = 12'h4bd == _T_121[11:0] ? 4'h0 : _GEN_10494; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10496 = 12'h4be == _T_121[11:0] ? 4'h0 : _GEN_10495; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10497 = 12'h4bf == _T_121[11:0] ? 4'h0 : _GEN_10496; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10498 = 12'h4c0 == _T_121[11:0] ? image_1216 : _GEN_10497; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10499 = 12'h4c1 == _T_121[11:0] ? image_1217 : _GEN_10498; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10500 = 12'h4c2 == _T_121[11:0] ? image_1218 : _GEN_10499; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10501 = 12'h4c3 == _T_121[11:0] ? image_1219 : _GEN_10500; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10502 = 12'h4c4 == _T_121[11:0] ? image_1220 : _GEN_10501; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10503 = 12'h4c5 == _T_121[11:0] ? image_1221 : _GEN_10502; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10504 = 12'h4c6 == _T_121[11:0] ? image_1222 : _GEN_10503; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10505 = 12'h4c7 == _T_121[11:0] ? image_1223 : _GEN_10504; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10506 = 12'h4c8 == _T_121[11:0] ? image_1224 : _GEN_10505; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10507 = 12'h4c9 == _T_121[11:0] ? image_1225 : _GEN_10506; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10508 = 12'h4ca == _T_121[11:0] ? image_1226 : _GEN_10507; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10509 = 12'h4cb == _T_121[11:0] ? image_1227 : _GEN_10508; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10510 = 12'h4cc == _T_121[11:0] ? image_1228 : _GEN_10509; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10511 = 12'h4cd == _T_121[11:0] ? image_1229 : _GEN_10510; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10512 = 12'h4ce == _T_121[11:0] ? image_1230 : _GEN_10511; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10513 = 12'h4cf == _T_121[11:0] ? image_1231 : _GEN_10512; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10514 = 12'h4d0 == _T_121[11:0] ? image_1232 : _GEN_10513; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10515 = 12'h4d1 == _T_121[11:0] ? image_1233 : _GEN_10514; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10516 = 12'h4d2 == _T_121[11:0] ? image_1234 : _GEN_10515; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10517 = 12'h4d3 == _T_121[11:0] ? image_1235 : _GEN_10516; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10518 = 12'h4d4 == _T_121[11:0] ? image_1236 : _GEN_10517; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10519 = 12'h4d5 == _T_121[11:0] ? image_1237 : _GEN_10518; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10520 = 12'h4d6 == _T_121[11:0] ? image_1238 : _GEN_10519; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10521 = 12'h4d7 == _T_121[11:0] ? image_1239 : _GEN_10520; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10522 = 12'h4d8 == _T_121[11:0] ? image_1240 : _GEN_10521; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10523 = 12'h4d9 == _T_121[11:0] ? image_1241 : _GEN_10522; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10524 = 12'h4da == _T_121[11:0] ? image_1242 : _GEN_10523; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10525 = 12'h4db == _T_121[11:0] ? image_1243 : _GEN_10524; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10526 = 12'h4dc == _T_121[11:0] ? image_1244 : _GEN_10525; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10527 = 12'h4dd == _T_121[11:0] ? image_1245 : _GEN_10526; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10528 = 12'h4de == _T_121[11:0] ? image_1246 : _GEN_10527; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10529 = 12'h4df == _T_121[11:0] ? image_1247 : _GEN_10528; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10530 = 12'h4e0 == _T_121[11:0] ? image_1248 : _GEN_10529; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10531 = 12'h4e1 == _T_121[11:0] ? image_1249 : _GEN_10530; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10532 = 12'h4e2 == _T_121[11:0] ? image_1250 : _GEN_10531; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10533 = 12'h4e3 == _T_121[11:0] ? image_1251 : _GEN_10532; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10534 = 12'h4e4 == _T_121[11:0] ? image_1252 : _GEN_10533; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10535 = 12'h4e5 == _T_121[11:0] ? image_1253 : _GEN_10534; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10536 = 12'h4e6 == _T_121[11:0] ? image_1254 : _GEN_10535; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10537 = 12'h4e7 == _T_121[11:0] ? image_1255 : _GEN_10536; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10538 = 12'h4e8 == _T_121[11:0] ? image_1256 : _GEN_10537; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10539 = 12'h4e9 == _T_121[11:0] ? image_1257 : _GEN_10538; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10540 = 12'h4ea == _T_121[11:0] ? image_1258 : _GEN_10539; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10541 = 12'h4eb == _T_121[11:0] ? image_1259 : _GEN_10540; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10542 = 12'h4ec == _T_121[11:0] ? image_1260 : _GEN_10541; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10543 = 12'h4ed == _T_121[11:0] ? image_1261 : _GEN_10542; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10544 = 12'h4ee == _T_121[11:0] ? image_1262 : _GEN_10543; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10545 = 12'h4ef == _T_121[11:0] ? image_1263 : _GEN_10544; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10546 = 12'h4f0 == _T_121[11:0] ? image_1264 : _GEN_10545; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10547 = 12'h4f1 == _T_121[11:0] ? image_1265 : _GEN_10546; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10548 = 12'h4f2 == _T_121[11:0] ? image_1266 : _GEN_10547; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10549 = 12'h4f3 == _T_121[11:0] ? image_1267 : _GEN_10548; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10550 = 12'h4f4 == _T_121[11:0] ? image_1268 : _GEN_10549; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10551 = 12'h4f5 == _T_121[11:0] ? image_1269 : _GEN_10550; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10552 = 12'h4f6 == _T_121[11:0] ? image_1270 : _GEN_10551; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10553 = 12'h4f7 == _T_121[11:0] ? image_1271 : _GEN_10552; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10554 = 12'h4f8 == _T_121[11:0] ? image_1272 : _GEN_10553; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10555 = 12'h4f9 == _T_121[11:0] ? image_1273 : _GEN_10554; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10556 = 12'h4fa == _T_121[11:0] ? image_1274 : _GEN_10555; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10557 = 12'h4fb == _T_121[11:0] ? image_1275 : _GEN_10556; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10558 = 12'h4fc == _T_121[11:0] ? 4'h0 : _GEN_10557; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10559 = 12'h4fd == _T_121[11:0] ? 4'h0 : _GEN_10558; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10560 = 12'h4fe == _T_121[11:0] ? 4'h0 : _GEN_10559; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10561 = 12'h4ff == _T_121[11:0] ? 4'h0 : _GEN_10560; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10562 = 12'h500 == _T_121[11:0] ? image_1280 : _GEN_10561; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10563 = 12'h501 == _T_121[11:0] ? image_1281 : _GEN_10562; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10564 = 12'h502 == _T_121[11:0] ? image_1282 : _GEN_10563; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10565 = 12'h503 == _T_121[11:0] ? image_1283 : _GEN_10564; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10566 = 12'h504 == _T_121[11:0] ? image_1284 : _GEN_10565; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10567 = 12'h505 == _T_121[11:0] ? image_1285 : _GEN_10566; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10568 = 12'h506 == _T_121[11:0] ? image_1286 : _GEN_10567; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10569 = 12'h507 == _T_121[11:0] ? image_1287 : _GEN_10568; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10570 = 12'h508 == _T_121[11:0] ? image_1288 : _GEN_10569; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10571 = 12'h509 == _T_121[11:0] ? image_1289 : _GEN_10570; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10572 = 12'h50a == _T_121[11:0] ? image_1290 : _GEN_10571; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10573 = 12'h50b == _T_121[11:0] ? image_1291 : _GEN_10572; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10574 = 12'h50c == _T_121[11:0] ? image_1292 : _GEN_10573; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10575 = 12'h50d == _T_121[11:0] ? image_1293 : _GEN_10574; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10576 = 12'h50e == _T_121[11:0] ? image_1294 : _GEN_10575; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10577 = 12'h50f == _T_121[11:0] ? image_1295 : _GEN_10576; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10578 = 12'h510 == _T_121[11:0] ? image_1296 : _GEN_10577; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10579 = 12'h511 == _T_121[11:0] ? image_1297 : _GEN_10578; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10580 = 12'h512 == _T_121[11:0] ? image_1298 : _GEN_10579; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10581 = 12'h513 == _T_121[11:0] ? image_1299 : _GEN_10580; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10582 = 12'h514 == _T_121[11:0] ? image_1300 : _GEN_10581; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10583 = 12'h515 == _T_121[11:0] ? image_1301 : _GEN_10582; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10584 = 12'h516 == _T_121[11:0] ? image_1302 : _GEN_10583; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10585 = 12'h517 == _T_121[11:0] ? image_1303 : _GEN_10584; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10586 = 12'h518 == _T_121[11:0] ? image_1304 : _GEN_10585; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10587 = 12'h519 == _T_121[11:0] ? image_1305 : _GEN_10586; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10588 = 12'h51a == _T_121[11:0] ? image_1306 : _GEN_10587; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10589 = 12'h51b == _T_121[11:0] ? image_1307 : _GEN_10588; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10590 = 12'h51c == _T_121[11:0] ? image_1308 : _GEN_10589; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10591 = 12'h51d == _T_121[11:0] ? image_1309 : _GEN_10590; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10592 = 12'h51e == _T_121[11:0] ? image_1310 : _GEN_10591; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10593 = 12'h51f == _T_121[11:0] ? image_1311 : _GEN_10592; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10594 = 12'h520 == _T_121[11:0] ? image_1312 : _GEN_10593; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10595 = 12'h521 == _T_121[11:0] ? image_1313 : _GEN_10594; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10596 = 12'h522 == _T_121[11:0] ? image_1314 : _GEN_10595; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10597 = 12'h523 == _T_121[11:0] ? image_1315 : _GEN_10596; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10598 = 12'h524 == _T_121[11:0] ? image_1316 : _GEN_10597; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10599 = 12'h525 == _T_121[11:0] ? image_1317 : _GEN_10598; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10600 = 12'h526 == _T_121[11:0] ? image_1318 : _GEN_10599; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10601 = 12'h527 == _T_121[11:0] ? image_1319 : _GEN_10600; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10602 = 12'h528 == _T_121[11:0] ? image_1320 : _GEN_10601; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10603 = 12'h529 == _T_121[11:0] ? image_1321 : _GEN_10602; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10604 = 12'h52a == _T_121[11:0] ? image_1322 : _GEN_10603; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10605 = 12'h52b == _T_121[11:0] ? image_1323 : _GEN_10604; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10606 = 12'h52c == _T_121[11:0] ? image_1324 : _GEN_10605; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10607 = 12'h52d == _T_121[11:0] ? image_1325 : _GEN_10606; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10608 = 12'h52e == _T_121[11:0] ? image_1326 : _GEN_10607; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10609 = 12'h52f == _T_121[11:0] ? image_1327 : _GEN_10608; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10610 = 12'h530 == _T_121[11:0] ? image_1328 : _GEN_10609; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10611 = 12'h531 == _T_121[11:0] ? image_1329 : _GEN_10610; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10612 = 12'h532 == _T_121[11:0] ? image_1330 : _GEN_10611; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10613 = 12'h533 == _T_121[11:0] ? image_1331 : _GEN_10612; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10614 = 12'h534 == _T_121[11:0] ? image_1332 : _GEN_10613; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10615 = 12'h535 == _T_121[11:0] ? image_1333 : _GEN_10614; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10616 = 12'h536 == _T_121[11:0] ? image_1334 : _GEN_10615; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10617 = 12'h537 == _T_121[11:0] ? image_1335 : _GEN_10616; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10618 = 12'h538 == _T_121[11:0] ? image_1336 : _GEN_10617; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10619 = 12'h539 == _T_121[11:0] ? image_1337 : _GEN_10618; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10620 = 12'h53a == _T_121[11:0] ? image_1338 : _GEN_10619; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10621 = 12'h53b == _T_121[11:0] ? image_1339 : _GEN_10620; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10622 = 12'h53c == _T_121[11:0] ? image_1340 : _GEN_10621; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10623 = 12'h53d == _T_121[11:0] ? image_1341 : _GEN_10622; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10624 = 12'h53e == _T_121[11:0] ? 4'h0 : _GEN_10623; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10625 = 12'h53f == _T_121[11:0] ? 4'h0 : _GEN_10624; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10626 = 12'h540 == _T_121[11:0] ? image_1344 : _GEN_10625; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10627 = 12'h541 == _T_121[11:0] ? image_1345 : _GEN_10626; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10628 = 12'h542 == _T_121[11:0] ? image_1346 : _GEN_10627; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10629 = 12'h543 == _T_121[11:0] ? image_1347 : _GEN_10628; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10630 = 12'h544 == _T_121[11:0] ? image_1348 : _GEN_10629; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10631 = 12'h545 == _T_121[11:0] ? image_1349 : _GEN_10630; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10632 = 12'h546 == _T_121[11:0] ? image_1350 : _GEN_10631; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10633 = 12'h547 == _T_121[11:0] ? image_1351 : _GEN_10632; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10634 = 12'h548 == _T_121[11:0] ? image_1352 : _GEN_10633; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10635 = 12'h549 == _T_121[11:0] ? image_1353 : _GEN_10634; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10636 = 12'h54a == _T_121[11:0] ? image_1354 : _GEN_10635; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10637 = 12'h54b == _T_121[11:0] ? image_1355 : _GEN_10636; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10638 = 12'h54c == _T_121[11:0] ? image_1356 : _GEN_10637; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10639 = 12'h54d == _T_121[11:0] ? image_1357 : _GEN_10638; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10640 = 12'h54e == _T_121[11:0] ? image_1358 : _GEN_10639; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10641 = 12'h54f == _T_121[11:0] ? image_1359 : _GEN_10640; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10642 = 12'h550 == _T_121[11:0] ? image_1360 : _GEN_10641; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10643 = 12'h551 == _T_121[11:0] ? image_1361 : _GEN_10642; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10644 = 12'h552 == _T_121[11:0] ? image_1362 : _GEN_10643; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10645 = 12'h553 == _T_121[11:0] ? image_1363 : _GEN_10644; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10646 = 12'h554 == _T_121[11:0] ? image_1364 : _GEN_10645; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10647 = 12'h555 == _T_121[11:0] ? image_1365 : _GEN_10646; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10648 = 12'h556 == _T_121[11:0] ? image_1366 : _GEN_10647; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10649 = 12'h557 == _T_121[11:0] ? image_1367 : _GEN_10648; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10650 = 12'h558 == _T_121[11:0] ? image_1368 : _GEN_10649; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10651 = 12'h559 == _T_121[11:0] ? image_1369 : _GEN_10650; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10652 = 12'h55a == _T_121[11:0] ? image_1370 : _GEN_10651; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10653 = 12'h55b == _T_121[11:0] ? image_1371 : _GEN_10652; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10654 = 12'h55c == _T_121[11:0] ? image_1372 : _GEN_10653; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10655 = 12'h55d == _T_121[11:0] ? image_1373 : _GEN_10654; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10656 = 12'h55e == _T_121[11:0] ? image_1374 : _GEN_10655; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10657 = 12'h55f == _T_121[11:0] ? image_1375 : _GEN_10656; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10658 = 12'h560 == _T_121[11:0] ? image_1376 : _GEN_10657; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10659 = 12'h561 == _T_121[11:0] ? image_1377 : _GEN_10658; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10660 = 12'h562 == _T_121[11:0] ? image_1378 : _GEN_10659; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10661 = 12'h563 == _T_121[11:0] ? image_1379 : _GEN_10660; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10662 = 12'h564 == _T_121[11:0] ? image_1380 : _GEN_10661; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10663 = 12'h565 == _T_121[11:0] ? image_1381 : _GEN_10662; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10664 = 12'h566 == _T_121[11:0] ? image_1382 : _GEN_10663; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10665 = 12'h567 == _T_121[11:0] ? image_1383 : _GEN_10664; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10666 = 12'h568 == _T_121[11:0] ? image_1384 : _GEN_10665; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10667 = 12'h569 == _T_121[11:0] ? image_1385 : _GEN_10666; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10668 = 12'h56a == _T_121[11:0] ? image_1386 : _GEN_10667; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10669 = 12'h56b == _T_121[11:0] ? image_1387 : _GEN_10668; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10670 = 12'h56c == _T_121[11:0] ? image_1388 : _GEN_10669; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10671 = 12'h56d == _T_121[11:0] ? image_1389 : _GEN_10670; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10672 = 12'h56e == _T_121[11:0] ? image_1390 : _GEN_10671; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10673 = 12'h56f == _T_121[11:0] ? image_1391 : _GEN_10672; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10674 = 12'h570 == _T_121[11:0] ? image_1392 : _GEN_10673; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10675 = 12'h571 == _T_121[11:0] ? image_1393 : _GEN_10674; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10676 = 12'h572 == _T_121[11:0] ? image_1394 : _GEN_10675; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10677 = 12'h573 == _T_121[11:0] ? image_1395 : _GEN_10676; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10678 = 12'h574 == _T_121[11:0] ? image_1396 : _GEN_10677; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10679 = 12'h575 == _T_121[11:0] ? image_1397 : _GEN_10678; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10680 = 12'h576 == _T_121[11:0] ? image_1398 : _GEN_10679; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10681 = 12'h577 == _T_121[11:0] ? image_1399 : _GEN_10680; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10682 = 12'h578 == _T_121[11:0] ? image_1400 : _GEN_10681; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10683 = 12'h579 == _T_121[11:0] ? image_1401 : _GEN_10682; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10684 = 12'h57a == _T_121[11:0] ? image_1402 : _GEN_10683; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10685 = 12'h57b == _T_121[11:0] ? image_1403 : _GEN_10684; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10686 = 12'h57c == _T_121[11:0] ? image_1404 : _GEN_10685; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10687 = 12'h57d == _T_121[11:0] ? image_1405 : _GEN_10686; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10688 = 12'h57e == _T_121[11:0] ? 4'h0 : _GEN_10687; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10689 = 12'h57f == _T_121[11:0] ? 4'h0 : _GEN_10688; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10690 = 12'h580 == _T_121[11:0] ? image_1408 : _GEN_10689; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10691 = 12'h581 == _T_121[11:0] ? image_1409 : _GEN_10690; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10692 = 12'h582 == _T_121[11:0] ? image_1410 : _GEN_10691; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10693 = 12'h583 == _T_121[11:0] ? image_1411 : _GEN_10692; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10694 = 12'h584 == _T_121[11:0] ? image_1412 : _GEN_10693; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10695 = 12'h585 == _T_121[11:0] ? image_1413 : _GEN_10694; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10696 = 12'h586 == _T_121[11:0] ? image_1414 : _GEN_10695; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10697 = 12'h587 == _T_121[11:0] ? image_1415 : _GEN_10696; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10698 = 12'h588 == _T_121[11:0] ? image_1416 : _GEN_10697; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10699 = 12'h589 == _T_121[11:0] ? image_1417 : _GEN_10698; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10700 = 12'h58a == _T_121[11:0] ? image_1418 : _GEN_10699; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10701 = 12'h58b == _T_121[11:0] ? image_1419 : _GEN_10700; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10702 = 12'h58c == _T_121[11:0] ? image_1420 : _GEN_10701; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10703 = 12'h58d == _T_121[11:0] ? image_1421 : _GEN_10702; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10704 = 12'h58e == _T_121[11:0] ? image_1422 : _GEN_10703; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10705 = 12'h58f == _T_121[11:0] ? image_1423 : _GEN_10704; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10706 = 12'h590 == _T_121[11:0] ? image_1424 : _GEN_10705; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10707 = 12'h591 == _T_121[11:0] ? image_1425 : _GEN_10706; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10708 = 12'h592 == _T_121[11:0] ? image_1426 : _GEN_10707; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10709 = 12'h593 == _T_121[11:0] ? image_1427 : _GEN_10708; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10710 = 12'h594 == _T_121[11:0] ? image_1428 : _GEN_10709; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10711 = 12'h595 == _T_121[11:0] ? image_1429 : _GEN_10710; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10712 = 12'h596 == _T_121[11:0] ? image_1430 : _GEN_10711; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10713 = 12'h597 == _T_121[11:0] ? image_1431 : _GEN_10712; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10714 = 12'h598 == _T_121[11:0] ? image_1432 : _GEN_10713; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10715 = 12'h599 == _T_121[11:0] ? image_1433 : _GEN_10714; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10716 = 12'h59a == _T_121[11:0] ? image_1434 : _GEN_10715; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10717 = 12'h59b == _T_121[11:0] ? image_1435 : _GEN_10716; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10718 = 12'h59c == _T_121[11:0] ? image_1436 : _GEN_10717; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10719 = 12'h59d == _T_121[11:0] ? image_1437 : _GEN_10718; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10720 = 12'h59e == _T_121[11:0] ? image_1438 : _GEN_10719; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10721 = 12'h59f == _T_121[11:0] ? image_1439 : _GEN_10720; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10722 = 12'h5a0 == _T_121[11:0] ? image_1440 : _GEN_10721; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10723 = 12'h5a1 == _T_121[11:0] ? image_1441 : _GEN_10722; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10724 = 12'h5a2 == _T_121[11:0] ? image_1442 : _GEN_10723; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10725 = 12'h5a3 == _T_121[11:0] ? image_1443 : _GEN_10724; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10726 = 12'h5a4 == _T_121[11:0] ? image_1444 : _GEN_10725; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10727 = 12'h5a5 == _T_121[11:0] ? image_1445 : _GEN_10726; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10728 = 12'h5a6 == _T_121[11:0] ? image_1446 : _GEN_10727; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10729 = 12'h5a7 == _T_121[11:0] ? image_1447 : _GEN_10728; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10730 = 12'h5a8 == _T_121[11:0] ? image_1448 : _GEN_10729; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10731 = 12'h5a9 == _T_121[11:0] ? image_1449 : _GEN_10730; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10732 = 12'h5aa == _T_121[11:0] ? image_1450 : _GEN_10731; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10733 = 12'h5ab == _T_121[11:0] ? image_1451 : _GEN_10732; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10734 = 12'h5ac == _T_121[11:0] ? image_1452 : _GEN_10733; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10735 = 12'h5ad == _T_121[11:0] ? image_1453 : _GEN_10734; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10736 = 12'h5ae == _T_121[11:0] ? image_1454 : _GEN_10735; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10737 = 12'h5af == _T_121[11:0] ? image_1455 : _GEN_10736; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10738 = 12'h5b0 == _T_121[11:0] ? image_1456 : _GEN_10737; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10739 = 12'h5b1 == _T_121[11:0] ? image_1457 : _GEN_10738; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10740 = 12'h5b2 == _T_121[11:0] ? image_1458 : _GEN_10739; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10741 = 12'h5b3 == _T_121[11:0] ? image_1459 : _GEN_10740; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10742 = 12'h5b4 == _T_121[11:0] ? image_1460 : _GEN_10741; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10743 = 12'h5b5 == _T_121[11:0] ? image_1461 : _GEN_10742; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10744 = 12'h5b6 == _T_121[11:0] ? image_1462 : _GEN_10743; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10745 = 12'h5b7 == _T_121[11:0] ? image_1463 : _GEN_10744; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10746 = 12'h5b8 == _T_121[11:0] ? image_1464 : _GEN_10745; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10747 = 12'h5b9 == _T_121[11:0] ? image_1465 : _GEN_10746; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10748 = 12'h5ba == _T_121[11:0] ? image_1466 : _GEN_10747; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10749 = 12'h5bb == _T_121[11:0] ? image_1467 : _GEN_10748; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10750 = 12'h5bc == _T_121[11:0] ? image_1468 : _GEN_10749; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10751 = 12'h5bd == _T_121[11:0] ? image_1469 : _GEN_10750; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10752 = 12'h5be == _T_121[11:0] ? 4'h0 : _GEN_10751; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10753 = 12'h5bf == _T_121[11:0] ? 4'h0 : _GEN_10752; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10754 = 12'h5c0 == _T_121[11:0] ? image_1472 : _GEN_10753; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10755 = 12'h5c1 == _T_121[11:0] ? image_1473 : _GEN_10754; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10756 = 12'h5c2 == _T_121[11:0] ? image_1474 : _GEN_10755; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10757 = 12'h5c3 == _T_121[11:0] ? image_1475 : _GEN_10756; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10758 = 12'h5c4 == _T_121[11:0] ? image_1476 : _GEN_10757; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10759 = 12'h5c5 == _T_121[11:0] ? image_1477 : _GEN_10758; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10760 = 12'h5c6 == _T_121[11:0] ? image_1478 : _GEN_10759; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10761 = 12'h5c7 == _T_121[11:0] ? image_1479 : _GEN_10760; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10762 = 12'h5c8 == _T_121[11:0] ? image_1480 : _GEN_10761; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10763 = 12'h5c9 == _T_121[11:0] ? image_1481 : _GEN_10762; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10764 = 12'h5ca == _T_121[11:0] ? image_1482 : _GEN_10763; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10765 = 12'h5cb == _T_121[11:0] ? image_1483 : _GEN_10764; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10766 = 12'h5cc == _T_121[11:0] ? image_1484 : _GEN_10765; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10767 = 12'h5cd == _T_121[11:0] ? image_1485 : _GEN_10766; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10768 = 12'h5ce == _T_121[11:0] ? image_1486 : _GEN_10767; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10769 = 12'h5cf == _T_121[11:0] ? image_1487 : _GEN_10768; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10770 = 12'h5d0 == _T_121[11:0] ? image_1488 : _GEN_10769; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10771 = 12'h5d1 == _T_121[11:0] ? image_1489 : _GEN_10770; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10772 = 12'h5d2 == _T_121[11:0] ? image_1490 : _GEN_10771; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10773 = 12'h5d3 == _T_121[11:0] ? image_1491 : _GEN_10772; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10774 = 12'h5d4 == _T_121[11:0] ? image_1492 : _GEN_10773; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10775 = 12'h5d5 == _T_121[11:0] ? image_1493 : _GEN_10774; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10776 = 12'h5d6 == _T_121[11:0] ? image_1494 : _GEN_10775; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10777 = 12'h5d7 == _T_121[11:0] ? image_1495 : _GEN_10776; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10778 = 12'h5d8 == _T_121[11:0] ? image_1496 : _GEN_10777; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10779 = 12'h5d9 == _T_121[11:0] ? image_1497 : _GEN_10778; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10780 = 12'h5da == _T_121[11:0] ? image_1498 : _GEN_10779; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10781 = 12'h5db == _T_121[11:0] ? image_1499 : _GEN_10780; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10782 = 12'h5dc == _T_121[11:0] ? image_1500 : _GEN_10781; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10783 = 12'h5dd == _T_121[11:0] ? image_1501 : _GEN_10782; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10784 = 12'h5de == _T_121[11:0] ? image_1502 : _GEN_10783; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10785 = 12'h5df == _T_121[11:0] ? image_1503 : _GEN_10784; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10786 = 12'h5e0 == _T_121[11:0] ? image_1504 : _GEN_10785; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10787 = 12'h5e1 == _T_121[11:0] ? image_1505 : _GEN_10786; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10788 = 12'h5e2 == _T_121[11:0] ? image_1506 : _GEN_10787; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10789 = 12'h5e3 == _T_121[11:0] ? image_1507 : _GEN_10788; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10790 = 12'h5e4 == _T_121[11:0] ? image_1508 : _GEN_10789; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10791 = 12'h5e5 == _T_121[11:0] ? image_1509 : _GEN_10790; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10792 = 12'h5e6 == _T_121[11:0] ? image_1510 : _GEN_10791; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10793 = 12'h5e7 == _T_121[11:0] ? image_1511 : _GEN_10792; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10794 = 12'h5e8 == _T_121[11:0] ? image_1512 : _GEN_10793; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10795 = 12'h5e9 == _T_121[11:0] ? image_1513 : _GEN_10794; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10796 = 12'h5ea == _T_121[11:0] ? image_1514 : _GEN_10795; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10797 = 12'h5eb == _T_121[11:0] ? image_1515 : _GEN_10796; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10798 = 12'h5ec == _T_121[11:0] ? image_1516 : _GEN_10797; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10799 = 12'h5ed == _T_121[11:0] ? image_1517 : _GEN_10798; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10800 = 12'h5ee == _T_121[11:0] ? image_1518 : _GEN_10799; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10801 = 12'h5ef == _T_121[11:0] ? image_1519 : _GEN_10800; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10802 = 12'h5f0 == _T_121[11:0] ? image_1520 : _GEN_10801; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10803 = 12'h5f1 == _T_121[11:0] ? image_1521 : _GEN_10802; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10804 = 12'h5f2 == _T_121[11:0] ? image_1522 : _GEN_10803; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10805 = 12'h5f3 == _T_121[11:0] ? image_1523 : _GEN_10804; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10806 = 12'h5f4 == _T_121[11:0] ? image_1524 : _GEN_10805; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10807 = 12'h5f5 == _T_121[11:0] ? image_1525 : _GEN_10806; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10808 = 12'h5f6 == _T_121[11:0] ? image_1526 : _GEN_10807; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10809 = 12'h5f7 == _T_121[11:0] ? image_1527 : _GEN_10808; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10810 = 12'h5f8 == _T_121[11:0] ? image_1528 : _GEN_10809; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10811 = 12'h5f9 == _T_121[11:0] ? image_1529 : _GEN_10810; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10812 = 12'h5fa == _T_121[11:0] ? image_1530 : _GEN_10811; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10813 = 12'h5fb == _T_121[11:0] ? image_1531 : _GEN_10812; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10814 = 12'h5fc == _T_121[11:0] ? image_1532 : _GEN_10813; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10815 = 12'h5fd == _T_121[11:0] ? image_1533 : _GEN_10814; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10816 = 12'h5fe == _T_121[11:0] ? 4'h0 : _GEN_10815; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10817 = 12'h5ff == _T_121[11:0] ? 4'h0 : _GEN_10816; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10818 = 12'h600 == _T_121[11:0] ? image_1536 : _GEN_10817; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10819 = 12'h601 == _T_121[11:0] ? image_1537 : _GEN_10818; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10820 = 12'h602 == _T_121[11:0] ? image_1538 : _GEN_10819; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10821 = 12'h603 == _T_121[11:0] ? image_1539 : _GEN_10820; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10822 = 12'h604 == _T_121[11:0] ? image_1540 : _GEN_10821; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10823 = 12'h605 == _T_121[11:0] ? image_1541 : _GEN_10822; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10824 = 12'h606 == _T_121[11:0] ? image_1542 : _GEN_10823; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10825 = 12'h607 == _T_121[11:0] ? image_1543 : _GEN_10824; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10826 = 12'h608 == _T_121[11:0] ? image_1544 : _GEN_10825; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10827 = 12'h609 == _T_121[11:0] ? image_1545 : _GEN_10826; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10828 = 12'h60a == _T_121[11:0] ? image_1546 : _GEN_10827; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10829 = 12'h60b == _T_121[11:0] ? image_1547 : _GEN_10828; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10830 = 12'h60c == _T_121[11:0] ? image_1548 : _GEN_10829; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10831 = 12'h60d == _T_121[11:0] ? image_1549 : _GEN_10830; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10832 = 12'h60e == _T_121[11:0] ? image_1550 : _GEN_10831; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10833 = 12'h60f == _T_121[11:0] ? image_1551 : _GEN_10832; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10834 = 12'h610 == _T_121[11:0] ? image_1552 : _GEN_10833; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10835 = 12'h611 == _T_121[11:0] ? image_1553 : _GEN_10834; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10836 = 12'h612 == _T_121[11:0] ? image_1554 : _GEN_10835; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10837 = 12'h613 == _T_121[11:0] ? image_1555 : _GEN_10836; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10838 = 12'h614 == _T_121[11:0] ? image_1556 : _GEN_10837; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10839 = 12'h615 == _T_121[11:0] ? image_1557 : _GEN_10838; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10840 = 12'h616 == _T_121[11:0] ? image_1558 : _GEN_10839; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10841 = 12'h617 == _T_121[11:0] ? image_1559 : _GEN_10840; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10842 = 12'h618 == _T_121[11:0] ? image_1560 : _GEN_10841; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10843 = 12'h619 == _T_121[11:0] ? image_1561 : _GEN_10842; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10844 = 12'h61a == _T_121[11:0] ? image_1562 : _GEN_10843; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10845 = 12'h61b == _T_121[11:0] ? image_1563 : _GEN_10844; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10846 = 12'h61c == _T_121[11:0] ? image_1564 : _GEN_10845; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10847 = 12'h61d == _T_121[11:0] ? image_1565 : _GEN_10846; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10848 = 12'h61e == _T_121[11:0] ? image_1566 : _GEN_10847; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10849 = 12'h61f == _T_121[11:0] ? image_1567 : _GEN_10848; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10850 = 12'h620 == _T_121[11:0] ? image_1568 : _GEN_10849; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10851 = 12'h621 == _T_121[11:0] ? image_1569 : _GEN_10850; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10852 = 12'h622 == _T_121[11:0] ? image_1570 : _GEN_10851; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10853 = 12'h623 == _T_121[11:0] ? image_1571 : _GEN_10852; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10854 = 12'h624 == _T_121[11:0] ? image_1572 : _GEN_10853; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10855 = 12'h625 == _T_121[11:0] ? image_1573 : _GEN_10854; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10856 = 12'h626 == _T_121[11:0] ? image_1574 : _GEN_10855; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10857 = 12'h627 == _T_121[11:0] ? image_1575 : _GEN_10856; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10858 = 12'h628 == _T_121[11:0] ? image_1576 : _GEN_10857; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10859 = 12'h629 == _T_121[11:0] ? image_1577 : _GEN_10858; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10860 = 12'h62a == _T_121[11:0] ? image_1578 : _GEN_10859; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10861 = 12'h62b == _T_121[11:0] ? image_1579 : _GEN_10860; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10862 = 12'h62c == _T_121[11:0] ? image_1580 : _GEN_10861; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10863 = 12'h62d == _T_121[11:0] ? image_1581 : _GEN_10862; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10864 = 12'h62e == _T_121[11:0] ? image_1582 : _GEN_10863; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10865 = 12'h62f == _T_121[11:0] ? image_1583 : _GEN_10864; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10866 = 12'h630 == _T_121[11:0] ? image_1584 : _GEN_10865; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10867 = 12'h631 == _T_121[11:0] ? image_1585 : _GEN_10866; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10868 = 12'h632 == _T_121[11:0] ? image_1586 : _GEN_10867; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10869 = 12'h633 == _T_121[11:0] ? image_1587 : _GEN_10868; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10870 = 12'h634 == _T_121[11:0] ? image_1588 : _GEN_10869; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10871 = 12'h635 == _T_121[11:0] ? image_1589 : _GEN_10870; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10872 = 12'h636 == _T_121[11:0] ? image_1590 : _GEN_10871; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10873 = 12'h637 == _T_121[11:0] ? image_1591 : _GEN_10872; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10874 = 12'h638 == _T_121[11:0] ? image_1592 : _GEN_10873; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10875 = 12'h639 == _T_121[11:0] ? image_1593 : _GEN_10874; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10876 = 12'h63a == _T_121[11:0] ? image_1594 : _GEN_10875; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10877 = 12'h63b == _T_121[11:0] ? image_1595 : _GEN_10876; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10878 = 12'h63c == _T_121[11:0] ? image_1596 : _GEN_10877; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10879 = 12'h63d == _T_121[11:0] ? image_1597 : _GEN_10878; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10880 = 12'h63e == _T_121[11:0] ? 4'h0 : _GEN_10879; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10881 = 12'h63f == _T_121[11:0] ? 4'h0 : _GEN_10880; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10882 = 12'h640 == _T_121[11:0] ? image_1600 : _GEN_10881; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10883 = 12'h641 == _T_121[11:0] ? image_1601 : _GEN_10882; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10884 = 12'h642 == _T_121[11:0] ? image_1602 : _GEN_10883; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10885 = 12'h643 == _T_121[11:0] ? image_1603 : _GEN_10884; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10886 = 12'h644 == _T_121[11:0] ? image_1604 : _GEN_10885; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10887 = 12'h645 == _T_121[11:0] ? image_1605 : _GEN_10886; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10888 = 12'h646 == _T_121[11:0] ? image_1606 : _GEN_10887; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10889 = 12'h647 == _T_121[11:0] ? image_1607 : _GEN_10888; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10890 = 12'h648 == _T_121[11:0] ? image_1608 : _GEN_10889; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10891 = 12'h649 == _T_121[11:0] ? image_1609 : _GEN_10890; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10892 = 12'h64a == _T_121[11:0] ? image_1610 : _GEN_10891; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10893 = 12'h64b == _T_121[11:0] ? image_1611 : _GEN_10892; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10894 = 12'h64c == _T_121[11:0] ? image_1612 : _GEN_10893; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10895 = 12'h64d == _T_121[11:0] ? image_1613 : _GEN_10894; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10896 = 12'h64e == _T_121[11:0] ? image_1614 : _GEN_10895; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10897 = 12'h64f == _T_121[11:0] ? image_1615 : _GEN_10896; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10898 = 12'h650 == _T_121[11:0] ? image_1616 : _GEN_10897; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10899 = 12'h651 == _T_121[11:0] ? image_1617 : _GEN_10898; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10900 = 12'h652 == _T_121[11:0] ? image_1618 : _GEN_10899; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10901 = 12'h653 == _T_121[11:0] ? image_1619 : _GEN_10900; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10902 = 12'h654 == _T_121[11:0] ? image_1620 : _GEN_10901; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10903 = 12'h655 == _T_121[11:0] ? image_1621 : _GEN_10902; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10904 = 12'h656 == _T_121[11:0] ? image_1622 : _GEN_10903; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10905 = 12'h657 == _T_121[11:0] ? image_1623 : _GEN_10904; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10906 = 12'h658 == _T_121[11:0] ? image_1624 : _GEN_10905; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10907 = 12'h659 == _T_121[11:0] ? image_1625 : _GEN_10906; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10908 = 12'h65a == _T_121[11:0] ? image_1626 : _GEN_10907; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10909 = 12'h65b == _T_121[11:0] ? image_1627 : _GEN_10908; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10910 = 12'h65c == _T_121[11:0] ? image_1628 : _GEN_10909; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10911 = 12'h65d == _T_121[11:0] ? image_1629 : _GEN_10910; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10912 = 12'h65e == _T_121[11:0] ? image_1630 : _GEN_10911; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10913 = 12'h65f == _T_121[11:0] ? image_1631 : _GEN_10912; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10914 = 12'h660 == _T_121[11:0] ? image_1632 : _GEN_10913; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10915 = 12'h661 == _T_121[11:0] ? image_1633 : _GEN_10914; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10916 = 12'h662 == _T_121[11:0] ? image_1634 : _GEN_10915; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10917 = 12'h663 == _T_121[11:0] ? image_1635 : _GEN_10916; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10918 = 12'h664 == _T_121[11:0] ? image_1636 : _GEN_10917; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10919 = 12'h665 == _T_121[11:0] ? image_1637 : _GEN_10918; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10920 = 12'h666 == _T_121[11:0] ? image_1638 : _GEN_10919; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10921 = 12'h667 == _T_121[11:0] ? image_1639 : _GEN_10920; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10922 = 12'h668 == _T_121[11:0] ? image_1640 : _GEN_10921; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10923 = 12'h669 == _T_121[11:0] ? image_1641 : _GEN_10922; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10924 = 12'h66a == _T_121[11:0] ? image_1642 : _GEN_10923; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10925 = 12'h66b == _T_121[11:0] ? image_1643 : _GEN_10924; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10926 = 12'h66c == _T_121[11:0] ? image_1644 : _GEN_10925; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10927 = 12'h66d == _T_121[11:0] ? image_1645 : _GEN_10926; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10928 = 12'h66e == _T_121[11:0] ? image_1646 : _GEN_10927; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10929 = 12'h66f == _T_121[11:0] ? image_1647 : _GEN_10928; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10930 = 12'h670 == _T_121[11:0] ? image_1648 : _GEN_10929; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10931 = 12'h671 == _T_121[11:0] ? image_1649 : _GEN_10930; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10932 = 12'h672 == _T_121[11:0] ? image_1650 : _GEN_10931; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10933 = 12'h673 == _T_121[11:0] ? image_1651 : _GEN_10932; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10934 = 12'h674 == _T_121[11:0] ? image_1652 : _GEN_10933; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10935 = 12'h675 == _T_121[11:0] ? image_1653 : _GEN_10934; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10936 = 12'h676 == _T_121[11:0] ? image_1654 : _GEN_10935; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10937 = 12'h677 == _T_121[11:0] ? image_1655 : _GEN_10936; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10938 = 12'h678 == _T_121[11:0] ? image_1656 : _GEN_10937; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10939 = 12'h679 == _T_121[11:0] ? image_1657 : _GEN_10938; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10940 = 12'h67a == _T_121[11:0] ? image_1658 : _GEN_10939; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10941 = 12'h67b == _T_121[11:0] ? image_1659 : _GEN_10940; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10942 = 12'h67c == _T_121[11:0] ? image_1660 : _GEN_10941; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10943 = 12'h67d == _T_121[11:0] ? 4'h0 : _GEN_10942; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10944 = 12'h67e == _T_121[11:0] ? 4'h0 : _GEN_10943; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10945 = 12'h67f == _T_121[11:0] ? 4'h0 : _GEN_10944; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10946 = 12'h680 == _T_121[11:0] ? image_1664 : _GEN_10945; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10947 = 12'h681 == _T_121[11:0] ? image_1665 : _GEN_10946; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10948 = 12'h682 == _T_121[11:0] ? image_1666 : _GEN_10947; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10949 = 12'h683 == _T_121[11:0] ? image_1667 : _GEN_10948; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10950 = 12'h684 == _T_121[11:0] ? image_1668 : _GEN_10949; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10951 = 12'h685 == _T_121[11:0] ? image_1669 : _GEN_10950; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10952 = 12'h686 == _T_121[11:0] ? image_1670 : _GEN_10951; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10953 = 12'h687 == _T_121[11:0] ? image_1671 : _GEN_10952; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10954 = 12'h688 == _T_121[11:0] ? image_1672 : _GEN_10953; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10955 = 12'h689 == _T_121[11:0] ? image_1673 : _GEN_10954; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10956 = 12'h68a == _T_121[11:0] ? image_1674 : _GEN_10955; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10957 = 12'h68b == _T_121[11:0] ? image_1675 : _GEN_10956; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10958 = 12'h68c == _T_121[11:0] ? image_1676 : _GEN_10957; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10959 = 12'h68d == _T_121[11:0] ? image_1677 : _GEN_10958; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10960 = 12'h68e == _T_121[11:0] ? image_1678 : _GEN_10959; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10961 = 12'h68f == _T_121[11:0] ? image_1679 : _GEN_10960; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10962 = 12'h690 == _T_121[11:0] ? image_1680 : _GEN_10961; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10963 = 12'h691 == _T_121[11:0] ? image_1681 : _GEN_10962; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10964 = 12'h692 == _T_121[11:0] ? image_1682 : _GEN_10963; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10965 = 12'h693 == _T_121[11:0] ? image_1683 : _GEN_10964; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10966 = 12'h694 == _T_121[11:0] ? image_1684 : _GEN_10965; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10967 = 12'h695 == _T_121[11:0] ? image_1685 : _GEN_10966; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10968 = 12'h696 == _T_121[11:0] ? image_1686 : _GEN_10967; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10969 = 12'h697 == _T_121[11:0] ? image_1687 : _GEN_10968; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10970 = 12'h698 == _T_121[11:0] ? image_1688 : _GEN_10969; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10971 = 12'h699 == _T_121[11:0] ? image_1689 : _GEN_10970; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10972 = 12'h69a == _T_121[11:0] ? image_1690 : _GEN_10971; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10973 = 12'h69b == _T_121[11:0] ? image_1691 : _GEN_10972; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10974 = 12'h69c == _T_121[11:0] ? image_1692 : _GEN_10973; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10975 = 12'h69d == _T_121[11:0] ? image_1693 : _GEN_10974; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10976 = 12'h69e == _T_121[11:0] ? image_1694 : _GEN_10975; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10977 = 12'h69f == _T_121[11:0] ? image_1695 : _GEN_10976; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10978 = 12'h6a0 == _T_121[11:0] ? image_1696 : _GEN_10977; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10979 = 12'h6a1 == _T_121[11:0] ? image_1697 : _GEN_10978; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10980 = 12'h6a2 == _T_121[11:0] ? image_1698 : _GEN_10979; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10981 = 12'h6a3 == _T_121[11:0] ? image_1699 : _GEN_10980; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10982 = 12'h6a4 == _T_121[11:0] ? image_1700 : _GEN_10981; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10983 = 12'h6a5 == _T_121[11:0] ? image_1701 : _GEN_10982; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10984 = 12'h6a6 == _T_121[11:0] ? image_1702 : _GEN_10983; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10985 = 12'h6a7 == _T_121[11:0] ? image_1703 : _GEN_10984; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10986 = 12'h6a8 == _T_121[11:0] ? image_1704 : _GEN_10985; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10987 = 12'h6a9 == _T_121[11:0] ? image_1705 : _GEN_10986; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10988 = 12'h6aa == _T_121[11:0] ? image_1706 : _GEN_10987; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10989 = 12'h6ab == _T_121[11:0] ? image_1707 : _GEN_10988; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10990 = 12'h6ac == _T_121[11:0] ? image_1708 : _GEN_10989; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10991 = 12'h6ad == _T_121[11:0] ? image_1709 : _GEN_10990; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10992 = 12'h6ae == _T_121[11:0] ? image_1710 : _GEN_10991; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10993 = 12'h6af == _T_121[11:0] ? image_1711 : _GEN_10992; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10994 = 12'h6b0 == _T_121[11:0] ? image_1712 : _GEN_10993; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10995 = 12'h6b1 == _T_121[11:0] ? image_1713 : _GEN_10994; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10996 = 12'h6b2 == _T_121[11:0] ? image_1714 : _GEN_10995; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10997 = 12'h6b3 == _T_121[11:0] ? image_1715 : _GEN_10996; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10998 = 12'h6b4 == _T_121[11:0] ? image_1716 : _GEN_10997; // @[Filter.scala 138:46]
  wire [3:0] _GEN_10999 = 12'h6b5 == _T_121[11:0] ? image_1717 : _GEN_10998; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11000 = 12'h6b6 == _T_121[11:0] ? image_1718 : _GEN_10999; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11001 = 12'h6b7 == _T_121[11:0] ? image_1719 : _GEN_11000; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11002 = 12'h6b8 == _T_121[11:0] ? image_1720 : _GEN_11001; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11003 = 12'h6b9 == _T_121[11:0] ? image_1721 : _GEN_11002; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11004 = 12'h6ba == _T_121[11:0] ? image_1722 : _GEN_11003; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11005 = 12'h6bb == _T_121[11:0] ? image_1723 : _GEN_11004; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11006 = 12'h6bc == _T_121[11:0] ? 4'h0 : _GEN_11005; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11007 = 12'h6bd == _T_121[11:0] ? 4'h0 : _GEN_11006; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11008 = 12'h6be == _T_121[11:0] ? 4'h0 : _GEN_11007; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11009 = 12'h6bf == _T_121[11:0] ? 4'h0 : _GEN_11008; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11010 = 12'h6c0 == _T_121[11:0] ? image_1728 : _GEN_11009; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11011 = 12'h6c1 == _T_121[11:0] ? image_1729 : _GEN_11010; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11012 = 12'h6c2 == _T_121[11:0] ? image_1730 : _GEN_11011; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11013 = 12'h6c3 == _T_121[11:0] ? image_1731 : _GEN_11012; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11014 = 12'h6c4 == _T_121[11:0] ? image_1732 : _GEN_11013; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11015 = 12'h6c5 == _T_121[11:0] ? image_1733 : _GEN_11014; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11016 = 12'h6c6 == _T_121[11:0] ? image_1734 : _GEN_11015; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11017 = 12'h6c7 == _T_121[11:0] ? image_1735 : _GEN_11016; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11018 = 12'h6c8 == _T_121[11:0] ? image_1736 : _GEN_11017; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11019 = 12'h6c9 == _T_121[11:0] ? image_1737 : _GEN_11018; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11020 = 12'h6ca == _T_121[11:0] ? image_1738 : _GEN_11019; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11021 = 12'h6cb == _T_121[11:0] ? image_1739 : _GEN_11020; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11022 = 12'h6cc == _T_121[11:0] ? image_1740 : _GEN_11021; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11023 = 12'h6cd == _T_121[11:0] ? image_1741 : _GEN_11022; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11024 = 12'h6ce == _T_121[11:0] ? image_1742 : _GEN_11023; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11025 = 12'h6cf == _T_121[11:0] ? image_1743 : _GEN_11024; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11026 = 12'h6d0 == _T_121[11:0] ? image_1744 : _GEN_11025; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11027 = 12'h6d1 == _T_121[11:0] ? image_1745 : _GEN_11026; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11028 = 12'h6d2 == _T_121[11:0] ? image_1746 : _GEN_11027; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11029 = 12'h6d3 == _T_121[11:0] ? image_1747 : _GEN_11028; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11030 = 12'h6d4 == _T_121[11:0] ? image_1748 : _GEN_11029; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11031 = 12'h6d5 == _T_121[11:0] ? image_1749 : _GEN_11030; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11032 = 12'h6d6 == _T_121[11:0] ? image_1750 : _GEN_11031; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11033 = 12'h6d7 == _T_121[11:0] ? image_1751 : _GEN_11032; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11034 = 12'h6d8 == _T_121[11:0] ? image_1752 : _GEN_11033; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11035 = 12'h6d9 == _T_121[11:0] ? image_1753 : _GEN_11034; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11036 = 12'h6da == _T_121[11:0] ? image_1754 : _GEN_11035; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11037 = 12'h6db == _T_121[11:0] ? image_1755 : _GEN_11036; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11038 = 12'h6dc == _T_121[11:0] ? image_1756 : _GEN_11037; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11039 = 12'h6dd == _T_121[11:0] ? image_1757 : _GEN_11038; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11040 = 12'h6de == _T_121[11:0] ? image_1758 : _GEN_11039; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11041 = 12'h6df == _T_121[11:0] ? image_1759 : _GEN_11040; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11042 = 12'h6e0 == _T_121[11:0] ? image_1760 : _GEN_11041; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11043 = 12'h6e1 == _T_121[11:0] ? image_1761 : _GEN_11042; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11044 = 12'h6e2 == _T_121[11:0] ? image_1762 : _GEN_11043; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11045 = 12'h6e3 == _T_121[11:0] ? image_1763 : _GEN_11044; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11046 = 12'h6e4 == _T_121[11:0] ? image_1764 : _GEN_11045; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11047 = 12'h6e5 == _T_121[11:0] ? image_1765 : _GEN_11046; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11048 = 12'h6e6 == _T_121[11:0] ? image_1766 : _GEN_11047; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11049 = 12'h6e7 == _T_121[11:0] ? image_1767 : _GEN_11048; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11050 = 12'h6e8 == _T_121[11:0] ? image_1768 : _GEN_11049; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11051 = 12'h6e9 == _T_121[11:0] ? image_1769 : _GEN_11050; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11052 = 12'h6ea == _T_121[11:0] ? image_1770 : _GEN_11051; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11053 = 12'h6eb == _T_121[11:0] ? image_1771 : _GEN_11052; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11054 = 12'h6ec == _T_121[11:0] ? image_1772 : _GEN_11053; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11055 = 12'h6ed == _T_121[11:0] ? image_1773 : _GEN_11054; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11056 = 12'h6ee == _T_121[11:0] ? image_1774 : _GEN_11055; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11057 = 12'h6ef == _T_121[11:0] ? image_1775 : _GEN_11056; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11058 = 12'h6f0 == _T_121[11:0] ? image_1776 : _GEN_11057; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11059 = 12'h6f1 == _T_121[11:0] ? image_1777 : _GEN_11058; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11060 = 12'h6f2 == _T_121[11:0] ? image_1778 : _GEN_11059; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11061 = 12'h6f3 == _T_121[11:0] ? image_1779 : _GEN_11060; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11062 = 12'h6f4 == _T_121[11:0] ? image_1780 : _GEN_11061; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11063 = 12'h6f5 == _T_121[11:0] ? image_1781 : _GEN_11062; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11064 = 12'h6f6 == _T_121[11:0] ? image_1782 : _GEN_11063; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11065 = 12'h6f7 == _T_121[11:0] ? image_1783 : _GEN_11064; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11066 = 12'h6f8 == _T_121[11:0] ? image_1784 : _GEN_11065; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11067 = 12'h6f9 == _T_121[11:0] ? image_1785 : _GEN_11066; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11068 = 12'h6fa == _T_121[11:0] ? image_1786 : _GEN_11067; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11069 = 12'h6fb == _T_121[11:0] ? 4'h0 : _GEN_11068; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11070 = 12'h6fc == _T_121[11:0] ? 4'h0 : _GEN_11069; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11071 = 12'h6fd == _T_121[11:0] ? 4'h0 : _GEN_11070; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11072 = 12'h6fe == _T_121[11:0] ? 4'h0 : _GEN_11071; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11073 = 12'h6ff == _T_121[11:0] ? 4'h0 : _GEN_11072; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11074 = 12'h700 == _T_121[11:0] ? 4'h0 : _GEN_11073; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11075 = 12'h701 == _T_121[11:0] ? image_1793 : _GEN_11074; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11076 = 12'h702 == _T_121[11:0] ? image_1794 : _GEN_11075; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11077 = 12'h703 == _T_121[11:0] ? image_1795 : _GEN_11076; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11078 = 12'h704 == _T_121[11:0] ? image_1796 : _GEN_11077; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11079 = 12'h705 == _T_121[11:0] ? image_1797 : _GEN_11078; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11080 = 12'h706 == _T_121[11:0] ? image_1798 : _GEN_11079; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11081 = 12'h707 == _T_121[11:0] ? image_1799 : _GEN_11080; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11082 = 12'h708 == _T_121[11:0] ? image_1800 : _GEN_11081; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11083 = 12'h709 == _T_121[11:0] ? image_1801 : _GEN_11082; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11084 = 12'h70a == _T_121[11:0] ? image_1802 : _GEN_11083; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11085 = 12'h70b == _T_121[11:0] ? image_1803 : _GEN_11084; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11086 = 12'h70c == _T_121[11:0] ? image_1804 : _GEN_11085; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11087 = 12'h70d == _T_121[11:0] ? image_1805 : _GEN_11086; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11088 = 12'h70e == _T_121[11:0] ? image_1806 : _GEN_11087; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11089 = 12'h70f == _T_121[11:0] ? image_1807 : _GEN_11088; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11090 = 12'h710 == _T_121[11:0] ? image_1808 : _GEN_11089; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11091 = 12'h711 == _T_121[11:0] ? image_1809 : _GEN_11090; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11092 = 12'h712 == _T_121[11:0] ? image_1810 : _GEN_11091; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11093 = 12'h713 == _T_121[11:0] ? image_1811 : _GEN_11092; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11094 = 12'h714 == _T_121[11:0] ? image_1812 : _GEN_11093; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11095 = 12'h715 == _T_121[11:0] ? image_1813 : _GEN_11094; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11096 = 12'h716 == _T_121[11:0] ? image_1814 : _GEN_11095; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11097 = 12'h717 == _T_121[11:0] ? image_1815 : _GEN_11096; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11098 = 12'h718 == _T_121[11:0] ? image_1816 : _GEN_11097; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11099 = 12'h719 == _T_121[11:0] ? image_1817 : _GEN_11098; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11100 = 12'h71a == _T_121[11:0] ? image_1818 : _GEN_11099; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11101 = 12'h71b == _T_121[11:0] ? image_1819 : _GEN_11100; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11102 = 12'h71c == _T_121[11:0] ? image_1820 : _GEN_11101; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11103 = 12'h71d == _T_121[11:0] ? image_1821 : _GEN_11102; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11104 = 12'h71e == _T_121[11:0] ? image_1822 : _GEN_11103; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11105 = 12'h71f == _T_121[11:0] ? image_1823 : _GEN_11104; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11106 = 12'h720 == _T_121[11:0] ? image_1824 : _GEN_11105; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11107 = 12'h721 == _T_121[11:0] ? image_1825 : _GEN_11106; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11108 = 12'h722 == _T_121[11:0] ? image_1826 : _GEN_11107; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11109 = 12'h723 == _T_121[11:0] ? image_1827 : _GEN_11108; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11110 = 12'h724 == _T_121[11:0] ? image_1828 : _GEN_11109; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11111 = 12'h725 == _T_121[11:0] ? image_1829 : _GEN_11110; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11112 = 12'h726 == _T_121[11:0] ? image_1830 : _GEN_11111; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11113 = 12'h727 == _T_121[11:0] ? image_1831 : _GEN_11112; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11114 = 12'h728 == _T_121[11:0] ? image_1832 : _GEN_11113; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11115 = 12'h729 == _T_121[11:0] ? image_1833 : _GEN_11114; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11116 = 12'h72a == _T_121[11:0] ? image_1834 : _GEN_11115; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11117 = 12'h72b == _T_121[11:0] ? image_1835 : _GEN_11116; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11118 = 12'h72c == _T_121[11:0] ? image_1836 : _GEN_11117; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11119 = 12'h72d == _T_121[11:0] ? image_1837 : _GEN_11118; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11120 = 12'h72e == _T_121[11:0] ? image_1838 : _GEN_11119; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11121 = 12'h72f == _T_121[11:0] ? image_1839 : _GEN_11120; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11122 = 12'h730 == _T_121[11:0] ? image_1840 : _GEN_11121; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11123 = 12'h731 == _T_121[11:0] ? image_1841 : _GEN_11122; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11124 = 12'h732 == _T_121[11:0] ? image_1842 : _GEN_11123; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11125 = 12'h733 == _T_121[11:0] ? image_1843 : _GEN_11124; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11126 = 12'h734 == _T_121[11:0] ? image_1844 : _GEN_11125; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11127 = 12'h735 == _T_121[11:0] ? image_1845 : _GEN_11126; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11128 = 12'h736 == _T_121[11:0] ? image_1846 : _GEN_11127; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11129 = 12'h737 == _T_121[11:0] ? image_1847 : _GEN_11128; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11130 = 12'h738 == _T_121[11:0] ? image_1848 : _GEN_11129; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11131 = 12'h739 == _T_121[11:0] ? image_1849 : _GEN_11130; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11132 = 12'h73a == _T_121[11:0] ? 4'h0 : _GEN_11131; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11133 = 12'h73b == _T_121[11:0] ? 4'h0 : _GEN_11132; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11134 = 12'h73c == _T_121[11:0] ? 4'h0 : _GEN_11133; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11135 = 12'h73d == _T_121[11:0] ? 4'h0 : _GEN_11134; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11136 = 12'h73e == _T_121[11:0] ? 4'h0 : _GEN_11135; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11137 = 12'h73f == _T_121[11:0] ? 4'h0 : _GEN_11136; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11138 = 12'h740 == _T_121[11:0] ? 4'h0 : _GEN_11137; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11139 = 12'h741 == _T_121[11:0] ? image_1857 : _GEN_11138; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11140 = 12'h742 == _T_121[11:0] ? image_1858 : _GEN_11139; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11141 = 12'h743 == _T_121[11:0] ? image_1859 : _GEN_11140; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11142 = 12'h744 == _T_121[11:0] ? image_1860 : _GEN_11141; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11143 = 12'h745 == _T_121[11:0] ? image_1861 : _GEN_11142; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11144 = 12'h746 == _T_121[11:0] ? image_1862 : _GEN_11143; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11145 = 12'h747 == _T_121[11:0] ? image_1863 : _GEN_11144; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11146 = 12'h748 == _T_121[11:0] ? image_1864 : _GEN_11145; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11147 = 12'h749 == _T_121[11:0] ? image_1865 : _GEN_11146; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11148 = 12'h74a == _T_121[11:0] ? image_1866 : _GEN_11147; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11149 = 12'h74b == _T_121[11:0] ? image_1867 : _GEN_11148; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11150 = 12'h74c == _T_121[11:0] ? image_1868 : _GEN_11149; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11151 = 12'h74d == _T_121[11:0] ? image_1869 : _GEN_11150; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11152 = 12'h74e == _T_121[11:0] ? image_1870 : _GEN_11151; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11153 = 12'h74f == _T_121[11:0] ? image_1871 : _GEN_11152; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11154 = 12'h750 == _T_121[11:0] ? image_1872 : _GEN_11153; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11155 = 12'h751 == _T_121[11:0] ? image_1873 : _GEN_11154; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11156 = 12'h752 == _T_121[11:0] ? image_1874 : _GEN_11155; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11157 = 12'h753 == _T_121[11:0] ? image_1875 : _GEN_11156; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11158 = 12'h754 == _T_121[11:0] ? image_1876 : _GEN_11157; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11159 = 12'h755 == _T_121[11:0] ? image_1877 : _GEN_11158; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11160 = 12'h756 == _T_121[11:0] ? image_1878 : _GEN_11159; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11161 = 12'h757 == _T_121[11:0] ? image_1879 : _GEN_11160; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11162 = 12'h758 == _T_121[11:0] ? image_1880 : _GEN_11161; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11163 = 12'h759 == _T_121[11:0] ? image_1881 : _GEN_11162; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11164 = 12'h75a == _T_121[11:0] ? image_1882 : _GEN_11163; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11165 = 12'h75b == _T_121[11:0] ? image_1883 : _GEN_11164; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11166 = 12'h75c == _T_121[11:0] ? image_1884 : _GEN_11165; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11167 = 12'h75d == _T_121[11:0] ? image_1885 : _GEN_11166; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11168 = 12'h75e == _T_121[11:0] ? image_1886 : _GEN_11167; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11169 = 12'h75f == _T_121[11:0] ? image_1887 : _GEN_11168; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11170 = 12'h760 == _T_121[11:0] ? image_1888 : _GEN_11169; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11171 = 12'h761 == _T_121[11:0] ? image_1889 : _GEN_11170; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11172 = 12'h762 == _T_121[11:0] ? image_1890 : _GEN_11171; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11173 = 12'h763 == _T_121[11:0] ? image_1891 : _GEN_11172; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11174 = 12'h764 == _T_121[11:0] ? image_1892 : _GEN_11173; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11175 = 12'h765 == _T_121[11:0] ? image_1893 : _GEN_11174; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11176 = 12'h766 == _T_121[11:0] ? image_1894 : _GEN_11175; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11177 = 12'h767 == _T_121[11:0] ? image_1895 : _GEN_11176; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11178 = 12'h768 == _T_121[11:0] ? image_1896 : _GEN_11177; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11179 = 12'h769 == _T_121[11:0] ? image_1897 : _GEN_11178; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11180 = 12'h76a == _T_121[11:0] ? image_1898 : _GEN_11179; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11181 = 12'h76b == _T_121[11:0] ? image_1899 : _GEN_11180; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11182 = 12'h76c == _T_121[11:0] ? image_1900 : _GEN_11181; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11183 = 12'h76d == _T_121[11:0] ? image_1901 : _GEN_11182; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11184 = 12'h76e == _T_121[11:0] ? image_1902 : _GEN_11183; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11185 = 12'h76f == _T_121[11:0] ? image_1903 : _GEN_11184; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11186 = 12'h770 == _T_121[11:0] ? image_1904 : _GEN_11185; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11187 = 12'h771 == _T_121[11:0] ? image_1905 : _GEN_11186; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11188 = 12'h772 == _T_121[11:0] ? image_1906 : _GEN_11187; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11189 = 12'h773 == _T_121[11:0] ? image_1907 : _GEN_11188; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11190 = 12'h774 == _T_121[11:0] ? image_1908 : _GEN_11189; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11191 = 12'h775 == _T_121[11:0] ? image_1909 : _GEN_11190; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11192 = 12'h776 == _T_121[11:0] ? image_1910 : _GEN_11191; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11193 = 12'h777 == _T_121[11:0] ? image_1911 : _GEN_11192; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11194 = 12'h778 == _T_121[11:0] ? image_1912 : _GEN_11193; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11195 = 12'h779 == _T_121[11:0] ? image_1913 : _GEN_11194; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11196 = 12'h77a == _T_121[11:0] ? 4'h0 : _GEN_11195; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11197 = 12'h77b == _T_121[11:0] ? 4'h0 : _GEN_11196; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11198 = 12'h77c == _T_121[11:0] ? 4'h0 : _GEN_11197; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11199 = 12'h77d == _T_121[11:0] ? 4'h0 : _GEN_11198; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11200 = 12'h77e == _T_121[11:0] ? 4'h0 : _GEN_11199; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11201 = 12'h77f == _T_121[11:0] ? 4'h0 : _GEN_11200; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11202 = 12'h780 == _T_121[11:0] ? 4'h0 : _GEN_11201; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11203 = 12'h781 == _T_121[11:0] ? image_1921 : _GEN_11202; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11204 = 12'h782 == _T_121[11:0] ? image_1922 : _GEN_11203; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11205 = 12'h783 == _T_121[11:0] ? image_1923 : _GEN_11204; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11206 = 12'h784 == _T_121[11:0] ? image_1924 : _GEN_11205; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11207 = 12'h785 == _T_121[11:0] ? image_1925 : _GEN_11206; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11208 = 12'h786 == _T_121[11:0] ? image_1926 : _GEN_11207; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11209 = 12'h787 == _T_121[11:0] ? image_1927 : _GEN_11208; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11210 = 12'h788 == _T_121[11:0] ? image_1928 : _GEN_11209; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11211 = 12'h789 == _T_121[11:0] ? image_1929 : _GEN_11210; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11212 = 12'h78a == _T_121[11:0] ? image_1930 : _GEN_11211; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11213 = 12'h78b == _T_121[11:0] ? image_1931 : _GEN_11212; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11214 = 12'h78c == _T_121[11:0] ? image_1932 : _GEN_11213; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11215 = 12'h78d == _T_121[11:0] ? image_1933 : _GEN_11214; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11216 = 12'h78e == _T_121[11:0] ? image_1934 : _GEN_11215; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11217 = 12'h78f == _T_121[11:0] ? image_1935 : _GEN_11216; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11218 = 12'h790 == _T_121[11:0] ? image_1936 : _GEN_11217; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11219 = 12'h791 == _T_121[11:0] ? image_1937 : _GEN_11218; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11220 = 12'h792 == _T_121[11:0] ? image_1938 : _GEN_11219; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11221 = 12'h793 == _T_121[11:0] ? image_1939 : _GEN_11220; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11222 = 12'h794 == _T_121[11:0] ? image_1940 : _GEN_11221; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11223 = 12'h795 == _T_121[11:0] ? image_1941 : _GEN_11222; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11224 = 12'h796 == _T_121[11:0] ? image_1942 : _GEN_11223; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11225 = 12'h797 == _T_121[11:0] ? image_1943 : _GEN_11224; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11226 = 12'h798 == _T_121[11:0] ? image_1944 : _GEN_11225; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11227 = 12'h799 == _T_121[11:0] ? image_1945 : _GEN_11226; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11228 = 12'h79a == _T_121[11:0] ? image_1946 : _GEN_11227; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11229 = 12'h79b == _T_121[11:0] ? image_1947 : _GEN_11228; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11230 = 12'h79c == _T_121[11:0] ? image_1948 : _GEN_11229; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11231 = 12'h79d == _T_121[11:0] ? image_1949 : _GEN_11230; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11232 = 12'h79e == _T_121[11:0] ? image_1950 : _GEN_11231; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11233 = 12'h79f == _T_121[11:0] ? image_1951 : _GEN_11232; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11234 = 12'h7a0 == _T_121[11:0] ? image_1952 : _GEN_11233; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11235 = 12'h7a1 == _T_121[11:0] ? image_1953 : _GEN_11234; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11236 = 12'h7a2 == _T_121[11:0] ? image_1954 : _GEN_11235; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11237 = 12'h7a3 == _T_121[11:0] ? image_1955 : _GEN_11236; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11238 = 12'h7a4 == _T_121[11:0] ? image_1956 : _GEN_11237; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11239 = 12'h7a5 == _T_121[11:0] ? image_1957 : _GEN_11238; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11240 = 12'h7a6 == _T_121[11:0] ? image_1958 : _GEN_11239; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11241 = 12'h7a7 == _T_121[11:0] ? image_1959 : _GEN_11240; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11242 = 12'h7a8 == _T_121[11:0] ? image_1960 : _GEN_11241; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11243 = 12'h7a9 == _T_121[11:0] ? image_1961 : _GEN_11242; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11244 = 12'h7aa == _T_121[11:0] ? image_1962 : _GEN_11243; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11245 = 12'h7ab == _T_121[11:0] ? image_1963 : _GEN_11244; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11246 = 12'h7ac == _T_121[11:0] ? image_1964 : _GEN_11245; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11247 = 12'h7ad == _T_121[11:0] ? image_1965 : _GEN_11246; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11248 = 12'h7ae == _T_121[11:0] ? image_1966 : _GEN_11247; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11249 = 12'h7af == _T_121[11:0] ? image_1967 : _GEN_11248; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11250 = 12'h7b0 == _T_121[11:0] ? image_1968 : _GEN_11249; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11251 = 12'h7b1 == _T_121[11:0] ? image_1969 : _GEN_11250; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11252 = 12'h7b2 == _T_121[11:0] ? image_1970 : _GEN_11251; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11253 = 12'h7b3 == _T_121[11:0] ? image_1971 : _GEN_11252; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11254 = 12'h7b4 == _T_121[11:0] ? image_1972 : _GEN_11253; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11255 = 12'h7b5 == _T_121[11:0] ? image_1973 : _GEN_11254; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11256 = 12'h7b6 == _T_121[11:0] ? image_1974 : _GEN_11255; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11257 = 12'h7b7 == _T_121[11:0] ? image_1975 : _GEN_11256; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11258 = 12'h7b8 == _T_121[11:0] ? image_1976 : _GEN_11257; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11259 = 12'h7b9 == _T_121[11:0] ? image_1977 : _GEN_11258; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11260 = 12'h7ba == _T_121[11:0] ? 4'h0 : _GEN_11259; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11261 = 12'h7bb == _T_121[11:0] ? 4'h0 : _GEN_11260; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11262 = 12'h7bc == _T_121[11:0] ? 4'h0 : _GEN_11261; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11263 = 12'h7bd == _T_121[11:0] ? 4'h0 : _GEN_11262; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11264 = 12'h7be == _T_121[11:0] ? 4'h0 : _GEN_11263; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11265 = 12'h7bf == _T_121[11:0] ? 4'h0 : _GEN_11264; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11266 = 12'h7c0 == _T_121[11:0] ? 4'h0 : _GEN_11265; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11267 = 12'h7c1 == _T_121[11:0] ? image_1985 : _GEN_11266; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11268 = 12'h7c2 == _T_121[11:0] ? image_1986 : _GEN_11267; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11269 = 12'h7c3 == _T_121[11:0] ? image_1987 : _GEN_11268; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11270 = 12'h7c4 == _T_121[11:0] ? image_1988 : _GEN_11269; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11271 = 12'h7c5 == _T_121[11:0] ? image_1989 : _GEN_11270; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11272 = 12'h7c6 == _T_121[11:0] ? image_1990 : _GEN_11271; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11273 = 12'h7c7 == _T_121[11:0] ? image_1991 : _GEN_11272; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11274 = 12'h7c8 == _T_121[11:0] ? image_1992 : _GEN_11273; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11275 = 12'h7c9 == _T_121[11:0] ? image_1993 : _GEN_11274; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11276 = 12'h7ca == _T_121[11:0] ? image_1994 : _GEN_11275; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11277 = 12'h7cb == _T_121[11:0] ? image_1995 : _GEN_11276; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11278 = 12'h7cc == _T_121[11:0] ? image_1996 : _GEN_11277; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11279 = 12'h7cd == _T_121[11:0] ? image_1997 : _GEN_11278; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11280 = 12'h7ce == _T_121[11:0] ? image_1998 : _GEN_11279; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11281 = 12'h7cf == _T_121[11:0] ? image_1999 : _GEN_11280; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11282 = 12'h7d0 == _T_121[11:0] ? image_2000 : _GEN_11281; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11283 = 12'h7d1 == _T_121[11:0] ? image_2001 : _GEN_11282; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11284 = 12'h7d2 == _T_121[11:0] ? image_2002 : _GEN_11283; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11285 = 12'h7d3 == _T_121[11:0] ? image_2003 : _GEN_11284; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11286 = 12'h7d4 == _T_121[11:0] ? image_2004 : _GEN_11285; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11287 = 12'h7d5 == _T_121[11:0] ? image_2005 : _GEN_11286; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11288 = 12'h7d6 == _T_121[11:0] ? image_2006 : _GEN_11287; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11289 = 12'h7d7 == _T_121[11:0] ? image_2007 : _GEN_11288; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11290 = 12'h7d8 == _T_121[11:0] ? image_2008 : _GEN_11289; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11291 = 12'h7d9 == _T_121[11:0] ? image_2009 : _GEN_11290; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11292 = 12'h7da == _T_121[11:0] ? image_2010 : _GEN_11291; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11293 = 12'h7db == _T_121[11:0] ? image_2011 : _GEN_11292; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11294 = 12'h7dc == _T_121[11:0] ? image_2012 : _GEN_11293; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11295 = 12'h7dd == _T_121[11:0] ? image_2013 : _GEN_11294; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11296 = 12'h7de == _T_121[11:0] ? image_2014 : _GEN_11295; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11297 = 12'h7df == _T_121[11:0] ? image_2015 : _GEN_11296; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11298 = 12'h7e0 == _T_121[11:0] ? image_2016 : _GEN_11297; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11299 = 12'h7e1 == _T_121[11:0] ? image_2017 : _GEN_11298; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11300 = 12'h7e2 == _T_121[11:0] ? image_2018 : _GEN_11299; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11301 = 12'h7e3 == _T_121[11:0] ? image_2019 : _GEN_11300; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11302 = 12'h7e4 == _T_121[11:0] ? image_2020 : _GEN_11301; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11303 = 12'h7e5 == _T_121[11:0] ? image_2021 : _GEN_11302; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11304 = 12'h7e6 == _T_121[11:0] ? image_2022 : _GEN_11303; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11305 = 12'h7e7 == _T_121[11:0] ? image_2023 : _GEN_11304; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11306 = 12'h7e8 == _T_121[11:0] ? image_2024 : _GEN_11305; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11307 = 12'h7e9 == _T_121[11:0] ? image_2025 : _GEN_11306; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11308 = 12'h7ea == _T_121[11:0] ? image_2026 : _GEN_11307; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11309 = 12'h7eb == _T_121[11:0] ? image_2027 : _GEN_11308; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11310 = 12'h7ec == _T_121[11:0] ? image_2028 : _GEN_11309; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11311 = 12'h7ed == _T_121[11:0] ? image_2029 : _GEN_11310; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11312 = 12'h7ee == _T_121[11:0] ? image_2030 : _GEN_11311; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11313 = 12'h7ef == _T_121[11:0] ? image_2031 : _GEN_11312; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11314 = 12'h7f0 == _T_121[11:0] ? image_2032 : _GEN_11313; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11315 = 12'h7f1 == _T_121[11:0] ? image_2033 : _GEN_11314; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11316 = 12'h7f2 == _T_121[11:0] ? image_2034 : _GEN_11315; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11317 = 12'h7f3 == _T_121[11:0] ? image_2035 : _GEN_11316; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11318 = 12'h7f4 == _T_121[11:0] ? image_2036 : _GEN_11317; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11319 = 12'h7f5 == _T_121[11:0] ? image_2037 : _GEN_11318; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11320 = 12'h7f6 == _T_121[11:0] ? image_2038 : _GEN_11319; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11321 = 12'h7f7 == _T_121[11:0] ? image_2039 : _GEN_11320; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11322 = 12'h7f8 == _T_121[11:0] ? image_2040 : _GEN_11321; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11323 = 12'h7f9 == _T_121[11:0] ? image_2041 : _GEN_11322; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11324 = 12'h7fa == _T_121[11:0] ? 4'h0 : _GEN_11323; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11325 = 12'h7fb == _T_121[11:0] ? 4'h0 : _GEN_11324; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11326 = 12'h7fc == _T_121[11:0] ? 4'h0 : _GEN_11325; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11327 = 12'h7fd == _T_121[11:0] ? 4'h0 : _GEN_11326; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11328 = 12'h7fe == _T_121[11:0] ? 4'h0 : _GEN_11327; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11329 = 12'h7ff == _T_121[11:0] ? 4'h0 : _GEN_11328; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11330 = 12'h800 == _T_121[11:0] ? 4'h0 : _GEN_11329; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11331 = 12'h801 == _T_121[11:0] ? image_2049 : _GEN_11330; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11332 = 12'h802 == _T_121[11:0] ? image_2050 : _GEN_11331; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11333 = 12'h803 == _T_121[11:0] ? image_2051 : _GEN_11332; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11334 = 12'h804 == _T_121[11:0] ? image_2052 : _GEN_11333; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11335 = 12'h805 == _T_121[11:0] ? image_2053 : _GEN_11334; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11336 = 12'h806 == _T_121[11:0] ? image_2054 : _GEN_11335; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11337 = 12'h807 == _T_121[11:0] ? image_2055 : _GEN_11336; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11338 = 12'h808 == _T_121[11:0] ? image_2056 : _GEN_11337; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11339 = 12'h809 == _T_121[11:0] ? image_2057 : _GEN_11338; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11340 = 12'h80a == _T_121[11:0] ? image_2058 : _GEN_11339; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11341 = 12'h80b == _T_121[11:0] ? image_2059 : _GEN_11340; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11342 = 12'h80c == _T_121[11:0] ? image_2060 : _GEN_11341; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11343 = 12'h80d == _T_121[11:0] ? image_2061 : _GEN_11342; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11344 = 12'h80e == _T_121[11:0] ? image_2062 : _GEN_11343; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11345 = 12'h80f == _T_121[11:0] ? image_2063 : _GEN_11344; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11346 = 12'h810 == _T_121[11:0] ? image_2064 : _GEN_11345; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11347 = 12'h811 == _T_121[11:0] ? image_2065 : _GEN_11346; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11348 = 12'h812 == _T_121[11:0] ? image_2066 : _GEN_11347; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11349 = 12'h813 == _T_121[11:0] ? image_2067 : _GEN_11348; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11350 = 12'h814 == _T_121[11:0] ? image_2068 : _GEN_11349; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11351 = 12'h815 == _T_121[11:0] ? image_2069 : _GEN_11350; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11352 = 12'h816 == _T_121[11:0] ? image_2070 : _GEN_11351; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11353 = 12'h817 == _T_121[11:0] ? image_2071 : _GEN_11352; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11354 = 12'h818 == _T_121[11:0] ? image_2072 : _GEN_11353; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11355 = 12'h819 == _T_121[11:0] ? image_2073 : _GEN_11354; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11356 = 12'h81a == _T_121[11:0] ? image_2074 : _GEN_11355; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11357 = 12'h81b == _T_121[11:0] ? image_2075 : _GEN_11356; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11358 = 12'h81c == _T_121[11:0] ? image_2076 : _GEN_11357; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11359 = 12'h81d == _T_121[11:0] ? image_2077 : _GEN_11358; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11360 = 12'h81e == _T_121[11:0] ? image_2078 : _GEN_11359; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11361 = 12'h81f == _T_121[11:0] ? image_2079 : _GEN_11360; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11362 = 12'h820 == _T_121[11:0] ? image_2080 : _GEN_11361; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11363 = 12'h821 == _T_121[11:0] ? image_2081 : _GEN_11362; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11364 = 12'h822 == _T_121[11:0] ? image_2082 : _GEN_11363; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11365 = 12'h823 == _T_121[11:0] ? image_2083 : _GEN_11364; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11366 = 12'h824 == _T_121[11:0] ? image_2084 : _GEN_11365; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11367 = 12'h825 == _T_121[11:0] ? image_2085 : _GEN_11366; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11368 = 12'h826 == _T_121[11:0] ? image_2086 : _GEN_11367; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11369 = 12'h827 == _T_121[11:0] ? image_2087 : _GEN_11368; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11370 = 12'h828 == _T_121[11:0] ? image_2088 : _GEN_11369; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11371 = 12'h829 == _T_121[11:0] ? image_2089 : _GEN_11370; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11372 = 12'h82a == _T_121[11:0] ? image_2090 : _GEN_11371; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11373 = 12'h82b == _T_121[11:0] ? image_2091 : _GEN_11372; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11374 = 12'h82c == _T_121[11:0] ? image_2092 : _GEN_11373; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11375 = 12'h82d == _T_121[11:0] ? image_2093 : _GEN_11374; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11376 = 12'h82e == _T_121[11:0] ? image_2094 : _GEN_11375; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11377 = 12'h82f == _T_121[11:0] ? image_2095 : _GEN_11376; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11378 = 12'h830 == _T_121[11:0] ? image_2096 : _GEN_11377; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11379 = 12'h831 == _T_121[11:0] ? image_2097 : _GEN_11378; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11380 = 12'h832 == _T_121[11:0] ? image_2098 : _GEN_11379; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11381 = 12'h833 == _T_121[11:0] ? image_2099 : _GEN_11380; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11382 = 12'h834 == _T_121[11:0] ? image_2100 : _GEN_11381; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11383 = 12'h835 == _T_121[11:0] ? image_2101 : _GEN_11382; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11384 = 12'h836 == _T_121[11:0] ? image_2102 : _GEN_11383; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11385 = 12'h837 == _T_121[11:0] ? image_2103 : _GEN_11384; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11386 = 12'h838 == _T_121[11:0] ? image_2104 : _GEN_11385; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11387 = 12'h839 == _T_121[11:0] ? image_2105 : _GEN_11386; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11388 = 12'h83a == _T_121[11:0] ? image_2106 : _GEN_11387; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11389 = 12'h83b == _T_121[11:0] ? 4'h0 : _GEN_11388; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11390 = 12'h83c == _T_121[11:0] ? 4'h0 : _GEN_11389; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11391 = 12'h83d == _T_121[11:0] ? 4'h0 : _GEN_11390; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11392 = 12'h83e == _T_121[11:0] ? 4'h0 : _GEN_11391; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11393 = 12'h83f == _T_121[11:0] ? 4'h0 : _GEN_11392; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11394 = 12'h840 == _T_121[11:0] ? 4'h0 : _GEN_11393; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11395 = 12'h841 == _T_121[11:0] ? 4'h0 : _GEN_11394; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11396 = 12'h842 == _T_121[11:0] ? image_2114 : _GEN_11395; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11397 = 12'h843 == _T_121[11:0] ? image_2115 : _GEN_11396; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11398 = 12'h844 == _T_121[11:0] ? image_2116 : _GEN_11397; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11399 = 12'h845 == _T_121[11:0] ? image_2117 : _GEN_11398; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11400 = 12'h846 == _T_121[11:0] ? image_2118 : _GEN_11399; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11401 = 12'h847 == _T_121[11:0] ? image_2119 : _GEN_11400; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11402 = 12'h848 == _T_121[11:0] ? image_2120 : _GEN_11401; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11403 = 12'h849 == _T_121[11:0] ? image_2121 : _GEN_11402; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11404 = 12'h84a == _T_121[11:0] ? image_2122 : _GEN_11403; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11405 = 12'h84b == _T_121[11:0] ? image_2123 : _GEN_11404; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11406 = 12'h84c == _T_121[11:0] ? image_2124 : _GEN_11405; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11407 = 12'h84d == _T_121[11:0] ? image_2125 : _GEN_11406; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11408 = 12'h84e == _T_121[11:0] ? image_2126 : _GEN_11407; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11409 = 12'h84f == _T_121[11:0] ? image_2127 : _GEN_11408; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11410 = 12'h850 == _T_121[11:0] ? image_2128 : _GEN_11409; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11411 = 12'h851 == _T_121[11:0] ? image_2129 : _GEN_11410; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11412 = 12'h852 == _T_121[11:0] ? image_2130 : _GEN_11411; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11413 = 12'h853 == _T_121[11:0] ? image_2131 : _GEN_11412; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11414 = 12'h854 == _T_121[11:0] ? image_2132 : _GEN_11413; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11415 = 12'h855 == _T_121[11:0] ? image_2133 : _GEN_11414; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11416 = 12'h856 == _T_121[11:0] ? image_2134 : _GEN_11415; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11417 = 12'h857 == _T_121[11:0] ? image_2135 : _GEN_11416; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11418 = 12'h858 == _T_121[11:0] ? image_2136 : _GEN_11417; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11419 = 12'h859 == _T_121[11:0] ? image_2137 : _GEN_11418; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11420 = 12'h85a == _T_121[11:0] ? image_2138 : _GEN_11419; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11421 = 12'h85b == _T_121[11:0] ? image_2139 : _GEN_11420; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11422 = 12'h85c == _T_121[11:0] ? image_2140 : _GEN_11421; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11423 = 12'h85d == _T_121[11:0] ? image_2141 : _GEN_11422; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11424 = 12'h85e == _T_121[11:0] ? image_2142 : _GEN_11423; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11425 = 12'h85f == _T_121[11:0] ? image_2143 : _GEN_11424; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11426 = 12'h860 == _T_121[11:0] ? image_2144 : _GEN_11425; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11427 = 12'h861 == _T_121[11:0] ? image_2145 : _GEN_11426; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11428 = 12'h862 == _T_121[11:0] ? image_2146 : _GEN_11427; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11429 = 12'h863 == _T_121[11:0] ? image_2147 : _GEN_11428; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11430 = 12'h864 == _T_121[11:0] ? image_2148 : _GEN_11429; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11431 = 12'h865 == _T_121[11:0] ? image_2149 : _GEN_11430; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11432 = 12'h866 == _T_121[11:0] ? image_2150 : _GEN_11431; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11433 = 12'h867 == _T_121[11:0] ? image_2151 : _GEN_11432; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11434 = 12'h868 == _T_121[11:0] ? image_2152 : _GEN_11433; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11435 = 12'h869 == _T_121[11:0] ? image_2153 : _GEN_11434; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11436 = 12'h86a == _T_121[11:0] ? image_2154 : _GEN_11435; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11437 = 12'h86b == _T_121[11:0] ? image_2155 : _GEN_11436; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11438 = 12'h86c == _T_121[11:0] ? image_2156 : _GEN_11437; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11439 = 12'h86d == _T_121[11:0] ? image_2157 : _GEN_11438; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11440 = 12'h86e == _T_121[11:0] ? image_2158 : _GEN_11439; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11441 = 12'h86f == _T_121[11:0] ? image_2159 : _GEN_11440; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11442 = 12'h870 == _T_121[11:0] ? image_2160 : _GEN_11441; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11443 = 12'h871 == _T_121[11:0] ? image_2161 : _GEN_11442; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11444 = 12'h872 == _T_121[11:0] ? image_2162 : _GEN_11443; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11445 = 12'h873 == _T_121[11:0] ? image_2163 : _GEN_11444; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11446 = 12'h874 == _T_121[11:0] ? image_2164 : _GEN_11445; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11447 = 12'h875 == _T_121[11:0] ? image_2165 : _GEN_11446; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11448 = 12'h876 == _T_121[11:0] ? image_2166 : _GEN_11447; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11449 = 12'h877 == _T_121[11:0] ? image_2167 : _GEN_11448; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11450 = 12'h878 == _T_121[11:0] ? image_2168 : _GEN_11449; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11451 = 12'h879 == _T_121[11:0] ? image_2169 : _GEN_11450; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11452 = 12'h87a == _T_121[11:0] ? image_2170 : _GEN_11451; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11453 = 12'h87b == _T_121[11:0] ? 4'h0 : _GEN_11452; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11454 = 12'h87c == _T_121[11:0] ? 4'h0 : _GEN_11453; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11455 = 12'h87d == _T_121[11:0] ? 4'h0 : _GEN_11454; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11456 = 12'h87e == _T_121[11:0] ? 4'h0 : _GEN_11455; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11457 = 12'h87f == _T_121[11:0] ? 4'h0 : _GEN_11456; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11458 = 12'h880 == _T_121[11:0] ? 4'h0 : _GEN_11457; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11459 = 12'h881 == _T_121[11:0] ? image_2177 : _GEN_11458; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11460 = 12'h882 == _T_121[11:0] ? image_2178 : _GEN_11459; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11461 = 12'h883 == _T_121[11:0] ? image_2179 : _GEN_11460; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11462 = 12'h884 == _T_121[11:0] ? image_2180 : _GEN_11461; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11463 = 12'h885 == _T_121[11:0] ? image_2181 : _GEN_11462; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11464 = 12'h886 == _T_121[11:0] ? image_2182 : _GEN_11463; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11465 = 12'h887 == _T_121[11:0] ? image_2183 : _GEN_11464; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11466 = 12'h888 == _T_121[11:0] ? image_2184 : _GEN_11465; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11467 = 12'h889 == _T_121[11:0] ? image_2185 : _GEN_11466; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11468 = 12'h88a == _T_121[11:0] ? image_2186 : _GEN_11467; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11469 = 12'h88b == _T_121[11:0] ? image_2187 : _GEN_11468; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11470 = 12'h88c == _T_121[11:0] ? image_2188 : _GEN_11469; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11471 = 12'h88d == _T_121[11:0] ? image_2189 : _GEN_11470; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11472 = 12'h88e == _T_121[11:0] ? image_2190 : _GEN_11471; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11473 = 12'h88f == _T_121[11:0] ? image_2191 : _GEN_11472; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11474 = 12'h890 == _T_121[11:0] ? image_2192 : _GEN_11473; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11475 = 12'h891 == _T_121[11:0] ? image_2193 : _GEN_11474; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11476 = 12'h892 == _T_121[11:0] ? image_2194 : _GEN_11475; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11477 = 12'h893 == _T_121[11:0] ? image_2195 : _GEN_11476; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11478 = 12'h894 == _T_121[11:0] ? image_2196 : _GEN_11477; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11479 = 12'h895 == _T_121[11:0] ? image_2197 : _GEN_11478; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11480 = 12'h896 == _T_121[11:0] ? image_2198 : _GEN_11479; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11481 = 12'h897 == _T_121[11:0] ? image_2199 : _GEN_11480; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11482 = 12'h898 == _T_121[11:0] ? image_2200 : _GEN_11481; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11483 = 12'h899 == _T_121[11:0] ? image_2201 : _GEN_11482; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11484 = 12'h89a == _T_121[11:0] ? image_2202 : _GEN_11483; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11485 = 12'h89b == _T_121[11:0] ? image_2203 : _GEN_11484; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11486 = 12'h89c == _T_121[11:0] ? image_2204 : _GEN_11485; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11487 = 12'h89d == _T_121[11:0] ? image_2205 : _GEN_11486; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11488 = 12'h89e == _T_121[11:0] ? image_2206 : _GEN_11487; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11489 = 12'h89f == _T_121[11:0] ? image_2207 : _GEN_11488; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11490 = 12'h8a0 == _T_121[11:0] ? image_2208 : _GEN_11489; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11491 = 12'h8a1 == _T_121[11:0] ? image_2209 : _GEN_11490; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11492 = 12'h8a2 == _T_121[11:0] ? image_2210 : _GEN_11491; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11493 = 12'h8a3 == _T_121[11:0] ? image_2211 : _GEN_11492; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11494 = 12'h8a4 == _T_121[11:0] ? image_2212 : _GEN_11493; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11495 = 12'h8a5 == _T_121[11:0] ? image_2213 : _GEN_11494; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11496 = 12'h8a6 == _T_121[11:0] ? image_2214 : _GEN_11495; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11497 = 12'h8a7 == _T_121[11:0] ? image_2215 : _GEN_11496; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11498 = 12'h8a8 == _T_121[11:0] ? image_2216 : _GEN_11497; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11499 = 12'h8a9 == _T_121[11:0] ? image_2217 : _GEN_11498; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11500 = 12'h8aa == _T_121[11:0] ? image_2218 : _GEN_11499; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11501 = 12'h8ab == _T_121[11:0] ? image_2219 : _GEN_11500; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11502 = 12'h8ac == _T_121[11:0] ? image_2220 : _GEN_11501; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11503 = 12'h8ad == _T_121[11:0] ? image_2221 : _GEN_11502; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11504 = 12'h8ae == _T_121[11:0] ? image_2222 : _GEN_11503; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11505 = 12'h8af == _T_121[11:0] ? image_2223 : _GEN_11504; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11506 = 12'h8b0 == _T_121[11:0] ? image_2224 : _GEN_11505; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11507 = 12'h8b1 == _T_121[11:0] ? image_2225 : _GEN_11506; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11508 = 12'h8b2 == _T_121[11:0] ? image_2226 : _GEN_11507; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11509 = 12'h8b3 == _T_121[11:0] ? image_2227 : _GEN_11508; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11510 = 12'h8b4 == _T_121[11:0] ? image_2228 : _GEN_11509; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11511 = 12'h8b5 == _T_121[11:0] ? image_2229 : _GEN_11510; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11512 = 12'h8b6 == _T_121[11:0] ? image_2230 : _GEN_11511; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11513 = 12'h8b7 == _T_121[11:0] ? image_2231 : _GEN_11512; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11514 = 12'h8b8 == _T_121[11:0] ? image_2232 : _GEN_11513; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11515 = 12'h8b9 == _T_121[11:0] ? image_2233 : _GEN_11514; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11516 = 12'h8ba == _T_121[11:0] ? image_2234 : _GEN_11515; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11517 = 12'h8bb == _T_121[11:0] ? 4'h0 : _GEN_11516; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11518 = 12'h8bc == _T_121[11:0] ? 4'h0 : _GEN_11517; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11519 = 12'h8bd == _T_121[11:0] ? 4'h0 : _GEN_11518; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11520 = 12'h8be == _T_121[11:0] ? 4'h0 : _GEN_11519; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11521 = 12'h8bf == _T_121[11:0] ? 4'h0 : _GEN_11520; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11522 = 12'h8c0 == _T_121[11:0] ? 4'h0 : _GEN_11521; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11523 = 12'h8c1 == _T_121[11:0] ? 4'h0 : _GEN_11522; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11524 = 12'h8c2 == _T_121[11:0] ? 4'h0 : _GEN_11523; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11525 = 12'h8c3 == _T_121[11:0] ? image_2243 : _GEN_11524; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11526 = 12'h8c4 == _T_121[11:0] ? image_2244 : _GEN_11525; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11527 = 12'h8c5 == _T_121[11:0] ? image_2245 : _GEN_11526; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11528 = 12'h8c6 == _T_121[11:0] ? image_2246 : _GEN_11527; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11529 = 12'h8c7 == _T_121[11:0] ? image_2247 : _GEN_11528; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11530 = 12'h8c8 == _T_121[11:0] ? image_2248 : _GEN_11529; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11531 = 12'h8c9 == _T_121[11:0] ? image_2249 : _GEN_11530; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11532 = 12'h8ca == _T_121[11:0] ? image_2250 : _GEN_11531; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11533 = 12'h8cb == _T_121[11:0] ? image_2251 : _GEN_11532; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11534 = 12'h8cc == _T_121[11:0] ? image_2252 : _GEN_11533; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11535 = 12'h8cd == _T_121[11:0] ? image_2253 : _GEN_11534; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11536 = 12'h8ce == _T_121[11:0] ? image_2254 : _GEN_11535; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11537 = 12'h8cf == _T_121[11:0] ? image_2255 : _GEN_11536; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11538 = 12'h8d0 == _T_121[11:0] ? image_2256 : _GEN_11537; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11539 = 12'h8d1 == _T_121[11:0] ? image_2257 : _GEN_11538; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11540 = 12'h8d2 == _T_121[11:0] ? image_2258 : _GEN_11539; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11541 = 12'h8d3 == _T_121[11:0] ? image_2259 : _GEN_11540; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11542 = 12'h8d4 == _T_121[11:0] ? image_2260 : _GEN_11541; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11543 = 12'h8d5 == _T_121[11:0] ? image_2261 : _GEN_11542; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11544 = 12'h8d6 == _T_121[11:0] ? image_2262 : _GEN_11543; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11545 = 12'h8d7 == _T_121[11:0] ? image_2263 : _GEN_11544; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11546 = 12'h8d8 == _T_121[11:0] ? image_2264 : _GEN_11545; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11547 = 12'h8d9 == _T_121[11:0] ? image_2265 : _GEN_11546; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11548 = 12'h8da == _T_121[11:0] ? image_2266 : _GEN_11547; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11549 = 12'h8db == _T_121[11:0] ? image_2267 : _GEN_11548; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11550 = 12'h8dc == _T_121[11:0] ? image_2268 : _GEN_11549; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11551 = 12'h8dd == _T_121[11:0] ? image_2269 : _GEN_11550; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11552 = 12'h8de == _T_121[11:0] ? image_2270 : _GEN_11551; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11553 = 12'h8df == _T_121[11:0] ? image_2271 : _GEN_11552; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11554 = 12'h8e0 == _T_121[11:0] ? image_2272 : _GEN_11553; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11555 = 12'h8e1 == _T_121[11:0] ? image_2273 : _GEN_11554; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11556 = 12'h8e2 == _T_121[11:0] ? image_2274 : _GEN_11555; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11557 = 12'h8e3 == _T_121[11:0] ? image_2275 : _GEN_11556; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11558 = 12'h8e4 == _T_121[11:0] ? image_2276 : _GEN_11557; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11559 = 12'h8e5 == _T_121[11:0] ? image_2277 : _GEN_11558; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11560 = 12'h8e6 == _T_121[11:0] ? image_2278 : _GEN_11559; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11561 = 12'h8e7 == _T_121[11:0] ? image_2279 : _GEN_11560; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11562 = 12'h8e8 == _T_121[11:0] ? image_2280 : _GEN_11561; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11563 = 12'h8e9 == _T_121[11:0] ? image_2281 : _GEN_11562; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11564 = 12'h8ea == _T_121[11:0] ? image_2282 : _GEN_11563; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11565 = 12'h8eb == _T_121[11:0] ? image_2283 : _GEN_11564; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11566 = 12'h8ec == _T_121[11:0] ? image_2284 : _GEN_11565; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11567 = 12'h8ed == _T_121[11:0] ? image_2285 : _GEN_11566; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11568 = 12'h8ee == _T_121[11:0] ? image_2286 : _GEN_11567; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11569 = 12'h8ef == _T_121[11:0] ? image_2287 : _GEN_11568; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11570 = 12'h8f0 == _T_121[11:0] ? image_2288 : _GEN_11569; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11571 = 12'h8f1 == _T_121[11:0] ? image_2289 : _GEN_11570; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11572 = 12'h8f2 == _T_121[11:0] ? image_2290 : _GEN_11571; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11573 = 12'h8f3 == _T_121[11:0] ? image_2291 : _GEN_11572; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11574 = 12'h8f4 == _T_121[11:0] ? image_2292 : _GEN_11573; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11575 = 12'h8f5 == _T_121[11:0] ? image_2293 : _GEN_11574; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11576 = 12'h8f6 == _T_121[11:0] ? image_2294 : _GEN_11575; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11577 = 12'h8f7 == _T_121[11:0] ? image_2295 : _GEN_11576; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11578 = 12'h8f8 == _T_121[11:0] ? image_2296 : _GEN_11577; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11579 = 12'h8f9 == _T_121[11:0] ? image_2297 : _GEN_11578; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11580 = 12'h8fa == _T_121[11:0] ? image_2298 : _GEN_11579; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11581 = 12'h8fb == _T_121[11:0] ? 4'h0 : _GEN_11580; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11582 = 12'h8fc == _T_121[11:0] ? 4'h0 : _GEN_11581; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11583 = 12'h8fd == _T_121[11:0] ? 4'h0 : _GEN_11582; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11584 = 12'h8fe == _T_121[11:0] ? 4'h0 : _GEN_11583; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11585 = 12'h8ff == _T_121[11:0] ? 4'h0 : _GEN_11584; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11586 = 12'h900 == _T_121[11:0] ? 4'h0 : _GEN_11585; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11587 = 12'h901 == _T_121[11:0] ? 4'h0 : _GEN_11586; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11588 = 12'h902 == _T_121[11:0] ? 4'h0 : _GEN_11587; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11589 = 12'h903 == _T_121[11:0] ? image_2307 : _GEN_11588; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11590 = 12'h904 == _T_121[11:0] ? image_2308 : _GEN_11589; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11591 = 12'h905 == _T_121[11:0] ? image_2309 : _GEN_11590; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11592 = 12'h906 == _T_121[11:0] ? image_2310 : _GEN_11591; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11593 = 12'h907 == _T_121[11:0] ? image_2311 : _GEN_11592; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11594 = 12'h908 == _T_121[11:0] ? image_2312 : _GEN_11593; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11595 = 12'h909 == _T_121[11:0] ? image_2313 : _GEN_11594; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11596 = 12'h90a == _T_121[11:0] ? image_2314 : _GEN_11595; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11597 = 12'h90b == _T_121[11:0] ? image_2315 : _GEN_11596; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11598 = 12'h90c == _T_121[11:0] ? image_2316 : _GEN_11597; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11599 = 12'h90d == _T_121[11:0] ? image_2317 : _GEN_11598; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11600 = 12'h90e == _T_121[11:0] ? image_2318 : _GEN_11599; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11601 = 12'h90f == _T_121[11:0] ? image_2319 : _GEN_11600; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11602 = 12'h910 == _T_121[11:0] ? image_2320 : _GEN_11601; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11603 = 12'h911 == _T_121[11:0] ? image_2321 : _GEN_11602; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11604 = 12'h912 == _T_121[11:0] ? image_2322 : _GEN_11603; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11605 = 12'h913 == _T_121[11:0] ? image_2323 : _GEN_11604; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11606 = 12'h914 == _T_121[11:0] ? image_2324 : _GEN_11605; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11607 = 12'h915 == _T_121[11:0] ? image_2325 : _GEN_11606; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11608 = 12'h916 == _T_121[11:0] ? image_2326 : _GEN_11607; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11609 = 12'h917 == _T_121[11:0] ? image_2327 : _GEN_11608; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11610 = 12'h918 == _T_121[11:0] ? image_2328 : _GEN_11609; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11611 = 12'h919 == _T_121[11:0] ? image_2329 : _GEN_11610; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11612 = 12'h91a == _T_121[11:0] ? image_2330 : _GEN_11611; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11613 = 12'h91b == _T_121[11:0] ? image_2331 : _GEN_11612; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11614 = 12'h91c == _T_121[11:0] ? image_2332 : _GEN_11613; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11615 = 12'h91d == _T_121[11:0] ? image_2333 : _GEN_11614; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11616 = 12'h91e == _T_121[11:0] ? image_2334 : _GEN_11615; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11617 = 12'h91f == _T_121[11:0] ? image_2335 : _GEN_11616; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11618 = 12'h920 == _T_121[11:0] ? image_2336 : _GEN_11617; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11619 = 12'h921 == _T_121[11:0] ? image_2337 : _GEN_11618; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11620 = 12'h922 == _T_121[11:0] ? image_2338 : _GEN_11619; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11621 = 12'h923 == _T_121[11:0] ? image_2339 : _GEN_11620; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11622 = 12'h924 == _T_121[11:0] ? image_2340 : _GEN_11621; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11623 = 12'h925 == _T_121[11:0] ? image_2341 : _GEN_11622; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11624 = 12'h926 == _T_121[11:0] ? image_2342 : _GEN_11623; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11625 = 12'h927 == _T_121[11:0] ? image_2343 : _GEN_11624; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11626 = 12'h928 == _T_121[11:0] ? image_2344 : _GEN_11625; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11627 = 12'h929 == _T_121[11:0] ? image_2345 : _GEN_11626; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11628 = 12'h92a == _T_121[11:0] ? image_2346 : _GEN_11627; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11629 = 12'h92b == _T_121[11:0] ? image_2347 : _GEN_11628; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11630 = 12'h92c == _T_121[11:0] ? image_2348 : _GEN_11629; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11631 = 12'h92d == _T_121[11:0] ? image_2349 : _GEN_11630; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11632 = 12'h92e == _T_121[11:0] ? image_2350 : _GEN_11631; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11633 = 12'h92f == _T_121[11:0] ? image_2351 : _GEN_11632; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11634 = 12'h930 == _T_121[11:0] ? image_2352 : _GEN_11633; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11635 = 12'h931 == _T_121[11:0] ? image_2353 : _GEN_11634; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11636 = 12'h932 == _T_121[11:0] ? image_2354 : _GEN_11635; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11637 = 12'h933 == _T_121[11:0] ? image_2355 : _GEN_11636; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11638 = 12'h934 == _T_121[11:0] ? image_2356 : _GEN_11637; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11639 = 12'h935 == _T_121[11:0] ? image_2357 : _GEN_11638; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11640 = 12'h936 == _T_121[11:0] ? image_2358 : _GEN_11639; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11641 = 12'h937 == _T_121[11:0] ? image_2359 : _GEN_11640; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11642 = 12'h938 == _T_121[11:0] ? image_2360 : _GEN_11641; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11643 = 12'h939 == _T_121[11:0] ? image_2361 : _GEN_11642; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11644 = 12'h93a == _T_121[11:0] ? image_2362 : _GEN_11643; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11645 = 12'h93b == _T_121[11:0] ? 4'h0 : _GEN_11644; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11646 = 12'h93c == _T_121[11:0] ? 4'h0 : _GEN_11645; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11647 = 12'h93d == _T_121[11:0] ? 4'h0 : _GEN_11646; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11648 = 12'h93e == _T_121[11:0] ? 4'h0 : _GEN_11647; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11649 = 12'h93f == _T_121[11:0] ? 4'h0 : _GEN_11648; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11650 = 12'h940 == _T_121[11:0] ? 4'h0 : _GEN_11649; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11651 = 12'h941 == _T_121[11:0] ? 4'h0 : _GEN_11650; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11652 = 12'h942 == _T_121[11:0] ? 4'h0 : _GEN_11651; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11653 = 12'h943 == _T_121[11:0] ? 4'h0 : _GEN_11652; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11654 = 12'h944 == _T_121[11:0] ? image_2372 : _GEN_11653; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11655 = 12'h945 == _T_121[11:0] ? image_2373 : _GEN_11654; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11656 = 12'h946 == _T_121[11:0] ? image_2374 : _GEN_11655; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11657 = 12'h947 == _T_121[11:0] ? image_2375 : _GEN_11656; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11658 = 12'h948 == _T_121[11:0] ? image_2376 : _GEN_11657; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11659 = 12'h949 == _T_121[11:0] ? image_2377 : _GEN_11658; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11660 = 12'h94a == _T_121[11:0] ? image_2378 : _GEN_11659; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11661 = 12'h94b == _T_121[11:0] ? image_2379 : _GEN_11660; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11662 = 12'h94c == _T_121[11:0] ? image_2380 : _GEN_11661; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11663 = 12'h94d == _T_121[11:0] ? image_2381 : _GEN_11662; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11664 = 12'h94e == _T_121[11:0] ? image_2382 : _GEN_11663; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11665 = 12'h94f == _T_121[11:0] ? image_2383 : _GEN_11664; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11666 = 12'h950 == _T_121[11:0] ? image_2384 : _GEN_11665; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11667 = 12'h951 == _T_121[11:0] ? image_2385 : _GEN_11666; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11668 = 12'h952 == _T_121[11:0] ? image_2386 : _GEN_11667; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11669 = 12'h953 == _T_121[11:0] ? image_2387 : _GEN_11668; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11670 = 12'h954 == _T_121[11:0] ? image_2388 : _GEN_11669; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11671 = 12'h955 == _T_121[11:0] ? image_2389 : _GEN_11670; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11672 = 12'h956 == _T_121[11:0] ? image_2390 : _GEN_11671; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11673 = 12'h957 == _T_121[11:0] ? image_2391 : _GEN_11672; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11674 = 12'h958 == _T_121[11:0] ? image_2392 : _GEN_11673; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11675 = 12'h959 == _T_121[11:0] ? image_2393 : _GEN_11674; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11676 = 12'h95a == _T_121[11:0] ? image_2394 : _GEN_11675; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11677 = 12'h95b == _T_121[11:0] ? image_2395 : _GEN_11676; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11678 = 12'h95c == _T_121[11:0] ? image_2396 : _GEN_11677; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11679 = 12'h95d == _T_121[11:0] ? image_2397 : _GEN_11678; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11680 = 12'h95e == _T_121[11:0] ? image_2398 : _GEN_11679; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11681 = 12'h95f == _T_121[11:0] ? image_2399 : _GEN_11680; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11682 = 12'h960 == _T_121[11:0] ? image_2400 : _GEN_11681; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11683 = 12'h961 == _T_121[11:0] ? image_2401 : _GEN_11682; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11684 = 12'h962 == _T_121[11:0] ? image_2402 : _GEN_11683; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11685 = 12'h963 == _T_121[11:0] ? image_2403 : _GEN_11684; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11686 = 12'h964 == _T_121[11:0] ? image_2404 : _GEN_11685; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11687 = 12'h965 == _T_121[11:0] ? image_2405 : _GEN_11686; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11688 = 12'h966 == _T_121[11:0] ? image_2406 : _GEN_11687; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11689 = 12'h967 == _T_121[11:0] ? image_2407 : _GEN_11688; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11690 = 12'h968 == _T_121[11:0] ? image_2408 : _GEN_11689; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11691 = 12'h969 == _T_121[11:0] ? image_2409 : _GEN_11690; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11692 = 12'h96a == _T_121[11:0] ? image_2410 : _GEN_11691; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11693 = 12'h96b == _T_121[11:0] ? image_2411 : _GEN_11692; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11694 = 12'h96c == _T_121[11:0] ? image_2412 : _GEN_11693; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11695 = 12'h96d == _T_121[11:0] ? image_2413 : _GEN_11694; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11696 = 12'h96e == _T_121[11:0] ? image_2414 : _GEN_11695; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11697 = 12'h96f == _T_121[11:0] ? image_2415 : _GEN_11696; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11698 = 12'h970 == _T_121[11:0] ? image_2416 : _GEN_11697; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11699 = 12'h971 == _T_121[11:0] ? image_2417 : _GEN_11698; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11700 = 12'h972 == _T_121[11:0] ? image_2418 : _GEN_11699; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11701 = 12'h973 == _T_121[11:0] ? image_2419 : _GEN_11700; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11702 = 12'h974 == _T_121[11:0] ? image_2420 : _GEN_11701; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11703 = 12'h975 == _T_121[11:0] ? image_2421 : _GEN_11702; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11704 = 12'h976 == _T_121[11:0] ? image_2422 : _GEN_11703; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11705 = 12'h977 == _T_121[11:0] ? image_2423 : _GEN_11704; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11706 = 12'h978 == _T_121[11:0] ? image_2424 : _GEN_11705; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11707 = 12'h979 == _T_121[11:0] ? image_2425 : _GEN_11706; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11708 = 12'h97a == _T_121[11:0] ? image_2426 : _GEN_11707; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11709 = 12'h97b == _T_121[11:0] ? 4'h0 : _GEN_11708; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11710 = 12'h97c == _T_121[11:0] ? 4'h0 : _GEN_11709; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11711 = 12'h97d == _T_121[11:0] ? 4'h0 : _GEN_11710; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11712 = 12'h97e == _T_121[11:0] ? 4'h0 : _GEN_11711; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11713 = 12'h97f == _T_121[11:0] ? 4'h0 : _GEN_11712; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11714 = 12'h980 == _T_121[11:0] ? 4'h0 : _GEN_11713; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11715 = 12'h981 == _T_121[11:0] ? 4'h0 : _GEN_11714; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11716 = 12'h982 == _T_121[11:0] ? 4'h0 : _GEN_11715; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11717 = 12'h983 == _T_121[11:0] ? 4'h0 : _GEN_11716; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11718 = 12'h984 == _T_121[11:0] ? 4'h0 : _GEN_11717; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11719 = 12'h985 == _T_121[11:0] ? image_2437 : _GEN_11718; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11720 = 12'h986 == _T_121[11:0] ? image_2438 : _GEN_11719; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11721 = 12'h987 == _T_121[11:0] ? image_2439 : _GEN_11720; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11722 = 12'h988 == _T_121[11:0] ? image_2440 : _GEN_11721; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11723 = 12'h989 == _T_121[11:0] ? image_2441 : _GEN_11722; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11724 = 12'h98a == _T_121[11:0] ? image_2442 : _GEN_11723; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11725 = 12'h98b == _T_121[11:0] ? image_2443 : _GEN_11724; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11726 = 12'h98c == _T_121[11:0] ? image_2444 : _GEN_11725; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11727 = 12'h98d == _T_121[11:0] ? image_2445 : _GEN_11726; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11728 = 12'h98e == _T_121[11:0] ? image_2446 : _GEN_11727; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11729 = 12'h98f == _T_121[11:0] ? image_2447 : _GEN_11728; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11730 = 12'h990 == _T_121[11:0] ? image_2448 : _GEN_11729; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11731 = 12'h991 == _T_121[11:0] ? image_2449 : _GEN_11730; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11732 = 12'h992 == _T_121[11:0] ? image_2450 : _GEN_11731; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11733 = 12'h993 == _T_121[11:0] ? image_2451 : _GEN_11732; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11734 = 12'h994 == _T_121[11:0] ? image_2452 : _GEN_11733; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11735 = 12'h995 == _T_121[11:0] ? image_2453 : _GEN_11734; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11736 = 12'h996 == _T_121[11:0] ? image_2454 : _GEN_11735; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11737 = 12'h997 == _T_121[11:0] ? image_2455 : _GEN_11736; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11738 = 12'h998 == _T_121[11:0] ? image_2456 : _GEN_11737; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11739 = 12'h999 == _T_121[11:0] ? image_2457 : _GEN_11738; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11740 = 12'h99a == _T_121[11:0] ? image_2458 : _GEN_11739; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11741 = 12'h99b == _T_121[11:0] ? image_2459 : _GEN_11740; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11742 = 12'h99c == _T_121[11:0] ? image_2460 : _GEN_11741; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11743 = 12'h99d == _T_121[11:0] ? image_2461 : _GEN_11742; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11744 = 12'h99e == _T_121[11:0] ? image_2462 : _GEN_11743; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11745 = 12'h99f == _T_121[11:0] ? image_2463 : _GEN_11744; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11746 = 12'h9a0 == _T_121[11:0] ? image_2464 : _GEN_11745; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11747 = 12'h9a1 == _T_121[11:0] ? image_2465 : _GEN_11746; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11748 = 12'h9a2 == _T_121[11:0] ? image_2466 : _GEN_11747; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11749 = 12'h9a3 == _T_121[11:0] ? image_2467 : _GEN_11748; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11750 = 12'h9a4 == _T_121[11:0] ? image_2468 : _GEN_11749; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11751 = 12'h9a5 == _T_121[11:0] ? image_2469 : _GEN_11750; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11752 = 12'h9a6 == _T_121[11:0] ? image_2470 : _GEN_11751; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11753 = 12'h9a7 == _T_121[11:0] ? image_2471 : _GEN_11752; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11754 = 12'h9a8 == _T_121[11:0] ? image_2472 : _GEN_11753; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11755 = 12'h9a9 == _T_121[11:0] ? image_2473 : _GEN_11754; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11756 = 12'h9aa == _T_121[11:0] ? image_2474 : _GEN_11755; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11757 = 12'h9ab == _T_121[11:0] ? image_2475 : _GEN_11756; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11758 = 12'h9ac == _T_121[11:0] ? image_2476 : _GEN_11757; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11759 = 12'h9ad == _T_121[11:0] ? image_2477 : _GEN_11758; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11760 = 12'h9ae == _T_121[11:0] ? image_2478 : _GEN_11759; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11761 = 12'h9af == _T_121[11:0] ? image_2479 : _GEN_11760; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11762 = 12'h9b0 == _T_121[11:0] ? image_2480 : _GEN_11761; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11763 = 12'h9b1 == _T_121[11:0] ? image_2481 : _GEN_11762; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11764 = 12'h9b2 == _T_121[11:0] ? image_2482 : _GEN_11763; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11765 = 12'h9b3 == _T_121[11:0] ? image_2483 : _GEN_11764; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11766 = 12'h9b4 == _T_121[11:0] ? image_2484 : _GEN_11765; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11767 = 12'h9b5 == _T_121[11:0] ? image_2485 : _GEN_11766; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11768 = 12'h9b6 == _T_121[11:0] ? image_2486 : _GEN_11767; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11769 = 12'h9b7 == _T_121[11:0] ? image_2487 : _GEN_11768; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11770 = 12'h9b8 == _T_121[11:0] ? image_2488 : _GEN_11769; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11771 = 12'h9b9 == _T_121[11:0] ? image_2489 : _GEN_11770; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11772 = 12'h9ba == _T_121[11:0] ? image_2490 : _GEN_11771; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11773 = 12'h9bb == _T_121[11:0] ? 4'h0 : _GEN_11772; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11774 = 12'h9bc == _T_121[11:0] ? 4'h0 : _GEN_11773; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11775 = 12'h9bd == _T_121[11:0] ? 4'h0 : _GEN_11774; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11776 = 12'h9be == _T_121[11:0] ? 4'h0 : _GEN_11775; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11777 = 12'h9bf == _T_121[11:0] ? 4'h0 : _GEN_11776; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11778 = 12'h9c0 == _T_121[11:0] ? 4'h0 : _GEN_11777; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11779 = 12'h9c1 == _T_121[11:0] ? 4'h0 : _GEN_11778; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11780 = 12'h9c2 == _T_121[11:0] ? 4'h0 : _GEN_11779; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11781 = 12'h9c3 == _T_121[11:0] ? 4'h0 : _GEN_11780; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11782 = 12'h9c4 == _T_121[11:0] ? 4'h0 : _GEN_11781; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11783 = 12'h9c5 == _T_121[11:0] ? 4'h0 : _GEN_11782; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11784 = 12'h9c6 == _T_121[11:0] ? image_2502 : _GEN_11783; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11785 = 12'h9c7 == _T_121[11:0] ? image_2503 : _GEN_11784; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11786 = 12'h9c8 == _T_121[11:0] ? image_2504 : _GEN_11785; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11787 = 12'h9c9 == _T_121[11:0] ? image_2505 : _GEN_11786; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11788 = 12'h9ca == _T_121[11:0] ? image_2506 : _GEN_11787; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11789 = 12'h9cb == _T_121[11:0] ? image_2507 : _GEN_11788; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11790 = 12'h9cc == _T_121[11:0] ? image_2508 : _GEN_11789; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11791 = 12'h9cd == _T_121[11:0] ? image_2509 : _GEN_11790; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11792 = 12'h9ce == _T_121[11:0] ? image_2510 : _GEN_11791; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11793 = 12'h9cf == _T_121[11:0] ? image_2511 : _GEN_11792; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11794 = 12'h9d0 == _T_121[11:0] ? image_2512 : _GEN_11793; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11795 = 12'h9d1 == _T_121[11:0] ? image_2513 : _GEN_11794; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11796 = 12'h9d2 == _T_121[11:0] ? image_2514 : _GEN_11795; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11797 = 12'h9d3 == _T_121[11:0] ? image_2515 : _GEN_11796; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11798 = 12'h9d4 == _T_121[11:0] ? image_2516 : _GEN_11797; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11799 = 12'h9d5 == _T_121[11:0] ? image_2517 : _GEN_11798; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11800 = 12'h9d6 == _T_121[11:0] ? image_2518 : _GEN_11799; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11801 = 12'h9d7 == _T_121[11:0] ? image_2519 : _GEN_11800; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11802 = 12'h9d8 == _T_121[11:0] ? image_2520 : _GEN_11801; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11803 = 12'h9d9 == _T_121[11:0] ? image_2521 : _GEN_11802; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11804 = 12'h9da == _T_121[11:0] ? image_2522 : _GEN_11803; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11805 = 12'h9db == _T_121[11:0] ? image_2523 : _GEN_11804; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11806 = 12'h9dc == _T_121[11:0] ? image_2524 : _GEN_11805; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11807 = 12'h9dd == _T_121[11:0] ? image_2525 : _GEN_11806; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11808 = 12'h9de == _T_121[11:0] ? image_2526 : _GEN_11807; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11809 = 12'h9df == _T_121[11:0] ? image_2527 : _GEN_11808; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11810 = 12'h9e0 == _T_121[11:0] ? image_2528 : _GEN_11809; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11811 = 12'h9e1 == _T_121[11:0] ? image_2529 : _GEN_11810; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11812 = 12'h9e2 == _T_121[11:0] ? image_2530 : _GEN_11811; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11813 = 12'h9e3 == _T_121[11:0] ? image_2531 : _GEN_11812; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11814 = 12'h9e4 == _T_121[11:0] ? image_2532 : _GEN_11813; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11815 = 12'h9e5 == _T_121[11:0] ? image_2533 : _GEN_11814; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11816 = 12'h9e6 == _T_121[11:0] ? image_2534 : _GEN_11815; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11817 = 12'h9e7 == _T_121[11:0] ? image_2535 : _GEN_11816; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11818 = 12'h9e8 == _T_121[11:0] ? image_2536 : _GEN_11817; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11819 = 12'h9e9 == _T_121[11:0] ? image_2537 : _GEN_11818; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11820 = 12'h9ea == _T_121[11:0] ? image_2538 : _GEN_11819; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11821 = 12'h9eb == _T_121[11:0] ? image_2539 : _GEN_11820; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11822 = 12'h9ec == _T_121[11:0] ? image_2540 : _GEN_11821; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11823 = 12'h9ed == _T_121[11:0] ? image_2541 : _GEN_11822; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11824 = 12'h9ee == _T_121[11:0] ? image_2542 : _GEN_11823; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11825 = 12'h9ef == _T_121[11:0] ? image_2543 : _GEN_11824; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11826 = 12'h9f0 == _T_121[11:0] ? image_2544 : _GEN_11825; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11827 = 12'h9f1 == _T_121[11:0] ? image_2545 : _GEN_11826; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11828 = 12'h9f2 == _T_121[11:0] ? image_2546 : _GEN_11827; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11829 = 12'h9f3 == _T_121[11:0] ? image_2547 : _GEN_11828; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11830 = 12'h9f4 == _T_121[11:0] ? image_2548 : _GEN_11829; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11831 = 12'h9f5 == _T_121[11:0] ? image_2549 : _GEN_11830; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11832 = 12'h9f6 == _T_121[11:0] ? image_2550 : _GEN_11831; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11833 = 12'h9f7 == _T_121[11:0] ? image_2551 : _GEN_11832; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11834 = 12'h9f8 == _T_121[11:0] ? image_2552 : _GEN_11833; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11835 = 12'h9f9 == _T_121[11:0] ? image_2553 : _GEN_11834; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11836 = 12'h9fa == _T_121[11:0] ? image_2554 : _GEN_11835; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11837 = 12'h9fb == _T_121[11:0] ? 4'h0 : _GEN_11836; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11838 = 12'h9fc == _T_121[11:0] ? 4'h0 : _GEN_11837; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11839 = 12'h9fd == _T_121[11:0] ? 4'h0 : _GEN_11838; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11840 = 12'h9fe == _T_121[11:0] ? 4'h0 : _GEN_11839; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11841 = 12'h9ff == _T_121[11:0] ? 4'h0 : _GEN_11840; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11842 = 12'ha00 == _T_121[11:0] ? 4'h0 : _GEN_11841; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11843 = 12'ha01 == _T_121[11:0] ? 4'h0 : _GEN_11842; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11844 = 12'ha02 == _T_121[11:0] ? 4'h0 : _GEN_11843; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11845 = 12'ha03 == _T_121[11:0] ? 4'h0 : _GEN_11844; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11846 = 12'ha04 == _T_121[11:0] ? 4'h0 : _GEN_11845; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11847 = 12'ha05 == _T_121[11:0] ? 4'h0 : _GEN_11846; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11848 = 12'ha06 == _T_121[11:0] ? 4'h0 : _GEN_11847; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11849 = 12'ha07 == _T_121[11:0] ? image_2567 : _GEN_11848; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11850 = 12'ha08 == _T_121[11:0] ? image_2568 : _GEN_11849; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11851 = 12'ha09 == _T_121[11:0] ? image_2569 : _GEN_11850; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11852 = 12'ha0a == _T_121[11:0] ? image_2570 : _GEN_11851; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11853 = 12'ha0b == _T_121[11:0] ? image_2571 : _GEN_11852; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11854 = 12'ha0c == _T_121[11:0] ? image_2572 : _GEN_11853; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11855 = 12'ha0d == _T_121[11:0] ? image_2573 : _GEN_11854; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11856 = 12'ha0e == _T_121[11:0] ? image_2574 : _GEN_11855; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11857 = 12'ha0f == _T_121[11:0] ? image_2575 : _GEN_11856; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11858 = 12'ha10 == _T_121[11:0] ? image_2576 : _GEN_11857; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11859 = 12'ha11 == _T_121[11:0] ? image_2577 : _GEN_11858; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11860 = 12'ha12 == _T_121[11:0] ? image_2578 : _GEN_11859; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11861 = 12'ha13 == _T_121[11:0] ? image_2579 : _GEN_11860; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11862 = 12'ha14 == _T_121[11:0] ? image_2580 : _GEN_11861; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11863 = 12'ha15 == _T_121[11:0] ? image_2581 : _GEN_11862; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11864 = 12'ha16 == _T_121[11:0] ? image_2582 : _GEN_11863; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11865 = 12'ha17 == _T_121[11:0] ? image_2583 : _GEN_11864; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11866 = 12'ha18 == _T_121[11:0] ? image_2584 : _GEN_11865; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11867 = 12'ha19 == _T_121[11:0] ? image_2585 : _GEN_11866; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11868 = 12'ha1a == _T_121[11:0] ? image_2586 : _GEN_11867; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11869 = 12'ha1b == _T_121[11:0] ? image_2587 : _GEN_11868; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11870 = 12'ha1c == _T_121[11:0] ? image_2588 : _GEN_11869; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11871 = 12'ha1d == _T_121[11:0] ? image_2589 : _GEN_11870; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11872 = 12'ha1e == _T_121[11:0] ? image_2590 : _GEN_11871; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11873 = 12'ha1f == _T_121[11:0] ? image_2591 : _GEN_11872; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11874 = 12'ha20 == _T_121[11:0] ? image_2592 : _GEN_11873; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11875 = 12'ha21 == _T_121[11:0] ? image_2593 : _GEN_11874; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11876 = 12'ha22 == _T_121[11:0] ? image_2594 : _GEN_11875; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11877 = 12'ha23 == _T_121[11:0] ? image_2595 : _GEN_11876; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11878 = 12'ha24 == _T_121[11:0] ? image_2596 : _GEN_11877; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11879 = 12'ha25 == _T_121[11:0] ? image_2597 : _GEN_11878; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11880 = 12'ha26 == _T_121[11:0] ? image_2598 : _GEN_11879; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11881 = 12'ha27 == _T_121[11:0] ? image_2599 : _GEN_11880; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11882 = 12'ha28 == _T_121[11:0] ? image_2600 : _GEN_11881; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11883 = 12'ha29 == _T_121[11:0] ? image_2601 : _GEN_11882; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11884 = 12'ha2a == _T_121[11:0] ? image_2602 : _GEN_11883; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11885 = 12'ha2b == _T_121[11:0] ? image_2603 : _GEN_11884; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11886 = 12'ha2c == _T_121[11:0] ? image_2604 : _GEN_11885; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11887 = 12'ha2d == _T_121[11:0] ? image_2605 : _GEN_11886; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11888 = 12'ha2e == _T_121[11:0] ? image_2606 : _GEN_11887; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11889 = 12'ha2f == _T_121[11:0] ? image_2607 : _GEN_11888; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11890 = 12'ha30 == _T_121[11:0] ? image_2608 : _GEN_11889; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11891 = 12'ha31 == _T_121[11:0] ? image_2609 : _GEN_11890; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11892 = 12'ha32 == _T_121[11:0] ? image_2610 : _GEN_11891; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11893 = 12'ha33 == _T_121[11:0] ? image_2611 : _GEN_11892; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11894 = 12'ha34 == _T_121[11:0] ? image_2612 : _GEN_11893; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11895 = 12'ha35 == _T_121[11:0] ? image_2613 : _GEN_11894; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11896 = 12'ha36 == _T_121[11:0] ? image_2614 : _GEN_11895; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11897 = 12'ha37 == _T_121[11:0] ? image_2615 : _GEN_11896; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11898 = 12'ha38 == _T_121[11:0] ? image_2616 : _GEN_11897; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11899 = 12'ha39 == _T_121[11:0] ? image_2617 : _GEN_11898; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11900 = 12'ha3a == _T_121[11:0] ? image_2618 : _GEN_11899; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11901 = 12'ha3b == _T_121[11:0] ? 4'h0 : _GEN_11900; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11902 = 12'ha3c == _T_121[11:0] ? 4'h0 : _GEN_11901; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11903 = 12'ha3d == _T_121[11:0] ? 4'h0 : _GEN_11902; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11904 = 12'ha3e == _T_121[11:0] ? 4'h0 : _GEN_11903; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11905 = 12'ha3f == _T_121[11:0] ? 4'h0 : _GEN_11904; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11906 = 12'ha40 == _T_121[11:0] ? 4'h0 : _GEN_11905; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11907 = 12'ha41 == _T_121[11:0] ? 4'h0 : _GEN_11906; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11908 = 12'ha42 == _T_121[11:0] ? 4'h0 : _GEN_11907; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11909 = 12'ha43 == _T_121[11:0] ? 4'h0 : _GEN_11908; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11910 = 12'ha44 == _T_121[11:0] ? 4'h0 : _GEN_11909; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11911 = 12'ha45 == _T_121[11:0] ? 4'h0 : _GEN_11910; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11912 = 12'ha46 == _T_121[11:0] ? 4'h0 : _GEN_11911; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11913 = 12'ha47 == _T_121[11:0] ? 4'h0 : _GEN_11912; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11914 = 12'ha48 == _T_121[11:0] ? image_2632 : _GEN_11913; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11915 = 12'ha49 == _T_121[11:0] ? image_2633 : _GEN_11914; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11916 = 12'ha4a == _T_121[11:0] ? image_2634 : _GEN_11915; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11917 = 12'ha4b == _T_121[11:0] ? image_2635 : _GEN_11916; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11918 = 12'ha4c == _T_121[11:0] ? image_2636 : _GEN_11917; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11919 = 12'ha4d == _T_121[11:0] ? image_2637 : _GEN_11918; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11920 = 12'ha4e == _T_121[11:0] ? image_2638 : _GEN_11919; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11921 = 12'ha4f == _T_121[11:0] ? image_2639 : _GEN_11920; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11922 = 12'ha50 == _T_121[11:0] ? image_2640 : _GEN_11921; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11923 = 12'ha51 == _T_121[11:0] ? image_2641 : _GEN_11922; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11924 = 12'ha52 == _T_121[11:0] ? image_2642 : _GEN_11923; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11925 = 12'ha53 == _T_121[11:0] ? image_2643 : _GEN_11924; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11926 = 12'ha54 == _T_121[11:0] ? image_2644 : _GEN_11925; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11927 = 12'ha55 == _T_121[11:0] ? image_2645 : _GEN_11926; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11928 = 12'ha56 == _T_121[11:0] ? image_2646 : _GEN_11927; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11929 = 12'ha57 == _T_121[11:0] ? image_2647 : _GEN_11928; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11930 = 12'ha58 == _T_121[11:0] ? image_2648 : _GEN_11929; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11931 = 12'ha59 == _T_121[11:0] ? image_2649 : _GEN_11930; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11932 = 12'ha5a == _T_121[11:0] ? image_2650 : _GEN_11931; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11933 = 12'ha5b == _T_121[11:0] ? image_2651 : _GEN_11932; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11934 = 12'ha5c == _T_121[11:0] ? image_2652 : _GEN_11933; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11935 = 12'ha5d == _T_121[11:0] ? image_2653 : _GEN_11934; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11936 = 12'ha5e == _T_121[11:0] ? image_2654 : _GEN_11935; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11937 = 12'ha5f == _T_121[11:0] ? image_2655 : _GEN_11936; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11938 = 12'ha60 == _T_121[11:0] ? image_2656 : _GEN_11937; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11939 = 12'ha61 == _T_121[11:0] ? image_2657 : _GEN_11938; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11940 = 12'ha62 == _T_121[11:0] ? image_2658 : _GEN_11939; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11941 = 12'ha63 == _T_121[11:0] ? image_2659 : _GEN_11940; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11942 = 12'ha64 == _T_121[11:0] ? image_2660 : _GEN_11941; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11943 = 12'ha65 == _T_121[11:0] ? image_2661 : _GEN_11942; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11944 = 12'ha66 == _T_121[11:0] ? image_2662 : _GEN_11943; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11945 = 12'ha67 == _T_121[11:0] ? image_2663 : _GEN_11944; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11946 = 12'ha68 == _T_121[11:0] ? image_2664 : _GEN_11945; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11947 = 12'ha69 == _T_121[11:0] ? image_2665 : _GEN_11946; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11948 = 12'ha6a == _T_121[11:0] ? image_2666 : _GEN_11947; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11949 = 12'ha6b == _T_121[11:0] ? image_2667 : _GEN_11948; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11950 = 12'ha6c == _T_121[11:0] ? image_2668 : _GEN_11949; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11951 = 12'ha6d == _T_121[11:0] ? image_2669 : _GEN_11950; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11952 = 12'ha6e == _T_121[11:0] ? image_2670 : _GEN_11951; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11953 = 12'ha6f == _T_121[11:0] ? image_2671 : _GEN_11952; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11954 = 12'ha70 == _T_121[11:0] ? image_2672 : _GEN_11953; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11955 = 12'ha71 == _T_121[11:0] ? image_2673 : _GEN_11954; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11956 = 12'ha72 == _T_121[11:0] ? image_2674 : _GEN_11955; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11957 = 12'ha73 == _T_121[11:0] ? image_2675 : _GEN_11956; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11958 = 12'ha74 == _T_121[11:0] ? image_2676 : _GEN_11957; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11959 = 12'ha75 == _T_121[11:0] ? image_2677 : _GEN_11958; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11960 = 12'ha76 == _T_121[11:0] ? image_2678 : _GEN_11959; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11961 = 12'ha77 == _T_121[11:0] ? image_2679 : _GEN_11960; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11962 = 12'ha78 == _T_121[11:0] ? image_2680 : _GEN_11961; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11963 = 12'ha79 == _T_121[11:0] ? image_2681 : _GEN_11962; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11964 = 12'ha7a == _T_121[11:0] ? image_2682 : _GEN_11963; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11965 = 12'ha7b == _T_121[11:0] ? 4'h0 : _GEN_11964; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11966 = 12'ha7c == _T_121[11:0] ? 4'h0 : _GEN_11965; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11967 = 12'ha7d == _T_121[11:0] ? 4'h0 : _GEN_11966; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11968 = 12'ha7e == _T_121[11:0] ? 4'h0 : _GEN_11967; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11969 = 12'ha7f == _T_121[11:0] ? 4'h0 : _GEN_11968; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11970 = 12'ha80 == _T_121[11:0] ? 4'h0 : _GEN_11969; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11971 = 12'ha81 == _T_121[11:0] ? 4'h0 : _GEN_11970; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11972 = 12'ha82 == _T_121[11:0] ? 4'h0 : _GEN_11971; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11973 = 12'ha83 == _T_121[11:0] ? 4'h0 : _GEN_11972; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11974 = 12'ha84 == _T_121[11:0] ? 4'h0 : _GEN_11973; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11975 = 12'ha85 == _T_121[11:0] ? 4'h0 : _GEN_11974; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11976 = 12'ha86 == _T_121[11:0] ? 4'h0 : _GEN_11975; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11977 = 12'ha87 == _T_121[11:0] ? 4'h0 : _GEN_11976; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11978 = 12'ha88 == _T_121[11:0] ? 4'h0 : _GEN_11977; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11979 = 12'ha89 == _T_121[11:0] ? image_2697 : _GEN_11978; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11980 = 12'ha8a == _T_121[11:0] ? image_2698 : _GEN_11979; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11981 = 12'ha8b == _T_121[11:0] ? image_2699 : _GEN_11980; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11982 = 12'ha8c == _T_121[11:0] ? image_2700 : _GEN_11981; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11983 = 12'ha8d == _T_121[11:0] ? image_2701 : _GEN_11982; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11984 = 12'ha8e == _T_121[11:0] ? image_2702 : _GEN_11983; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11985 = 12'ha8f == _T_121[11:0] ? image_2703 : _GEN_11984; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11986 = 12'ha90 == _T_121[11:0] ? image_2704 : _GEN_11985; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11987 = 12'ha91 == _T_121[11:0] ? image_2705 : _GEN_11986; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11988 = 12'ha92 == _T_121[11:0] ? image_2706 : _GEN_11987; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11989 = 12'ha93 == _T_121[11:0] ? image_2707 : _GEN_11988; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11990 = 12'ha94 == _T_121[11:0] ? image_2708 : _GEN_11989; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11991 = 12'ha95 == _T_121[11:0] ? image_2709 : _GEN_11990; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11992 = 12'ha96 == _T_121[11:0] ? image_2710 : _GEN_11991; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11993 = 12'ha97 == _T_121[11:0] ? image_2711 : _GEN_11992; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11994 = 12'ha98 == _T_121[11:0] ? image_2712 : _GEN_11993; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11995 = 12'ha99 == _T_121[11:0] ? image_2713 : _GEN_11994; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11996 = 12'ha9a == _T_121[11:0] ? image_2714 : _GEN_11995; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11997 = 12'ha9b == _T_121[11:0] ? image_2715 : _GEN_11996; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11998 = 12'ha9c == _T_121[11:0] ? image_2716 : _GEN_11997; // @[Filter.scala 138:46]
  wire [3:0] _GEN_11999 = 12'ha9d == _T_121[11:0] ? image_2717 : _GEN_11998; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12000 = 12'ha9e == _T_121[11:0] ? image_2718 : _GEN_11999; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12001 = 12'ha9f == _T_121[11:0] ? image_2719 : _GEN_12000; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12002 = 12'haa0 == _T_121[11:0] ? image_2720 : _GEN_12001; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12003 = 12'haa1 == _T_121[11:0] ? image_2721 : _GEN_12002; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12004 = 12'haa2 == _T_121[11:0] ? image_2722 : _GEN_12003; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12005 = 12'haa3 == _T_121[11:0] ? image_2723 : _GEN_12004; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12006 = 12'haa4 == _T_121[11:0] ? image_2724 : _GEN_12005; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12007 = 12'haa5 == _T_121[11:0] ? image_2725 : _GEN_12006; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12008 = 12'haa6 == _T_121[11:0] ? image_2726 : _GEN_12007; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12009 = 12'haa7 == _T_121[11:0] ? image_2727 : _GEN_12008; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12010 = 12'haa8 == _T_121[11:0] ? image_2728 : _GEN_12009; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12011 = 12'haa9 == _T_121[11:0] ? image_2729 : _GEN_12010; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12012 = 12'haaa == _T_121[11:0] ? image_2730 : _GEN_12011; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12013 = 12'haab == _T_121[11:0] ? image_2731 : _GEN_12012; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12014 = 12'haac == _T_121[11:0] ? image_2732 : _GEN_12013; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12015 = 12'haad == _T_121[11:0] ? image_2733 : _GEN_12014; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12016 = 12'haae == _T_121[11:0] ? image_2734 : _GEN_12015; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12017 = 12'haaf == _T_121[11:0] ? image_2735 : _GEN_12016; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12018 = 12'hab0 == _T_121[11:0] ? image_2736 : _GEN_12017; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12019 = 12'hab1 == _T_121[11:0] ? image_2737 : _GEN_12018; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12020 = 12'hab2 == _T_121[11:0] ? image_2738 : _GEN_12019; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12021 = 12'hab3 == _T_121[11:0] ? image_2739 : _GEN_12020; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12022 = 12'hab4 == _T_121[11:0] ? image_2740 : _GEN_12021; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12023 = 12'hab5 == _T_121[11:0] ? image_2741 : _GEN_12022; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12024 = 12'hab6 == _T_121[11:0] ? image_2742 : _GEN_12023; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12025 = 12'hab7 == _T_121[11:0] ? image_2743 : _GEN_12024; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12026 = 12'hab8 == _T_121[11:0] ? image_2744 : _GEN_12025; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12027 = 12'hab9 == _T_121[11:0] ? image_2745 : _GEN_12026; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12028 = 12'haba == _T_121[11:0] ? 4'h0 : _GEN_12027; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12029 = 12'habb == _T_121[11:0] ? 4'h0 : _GEN_12028; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12030 = 12'habc == _T_121[11:0] ? 4'h0 : _GEN_12029; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12031 = 12'habd == _T_121[11:0] ? 4'h0 : _GEN_12030; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12032 = 12'habe == _T_121[11:0] ? 4'h0 : _GEN_12031; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12033 = 12'habf == _T_121[11:0] ? 4'h0 : _GEN_12032; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12034 = 12'hac0 == _T_121[11:0] ? 4'h0 : _GEN_12033; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12035 = 12'hac1 == _T_121[11:0] ? 4'h0 : _GEN_12034; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12036 = 12'hac2 == _T_121[11:0] ? 4'h0 : _GEN_12035; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12037 = 12'hac3 == _T_121[11:0] ? 4'h0 : _GEN_12036; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12038 = 12'hac4 == _T_121[11:0] ? 4'h0 : _GEN_12037; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12039 = 12'hac5 == _T_121[11:0] ? 4'h0 : _GEN_12038; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12040 = 12'hac6 == _T_121[11:0] ? 4'h0 : _GEN_12039; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12041 = 12'hac7 == _T_121[11:0] ? 4'h0 : _GEN_12040; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12042 = 12'hac8 == _T_121[11:0] ? 4'h0 : _GEN_12041; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12043 = 12'hac9 == _T_121[11:0] ? 4'h0 : _GEN_12042; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12044 = 12'haca == _T_121[11:0] ? 4'h0 : _GEN_12043; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12045 = 12'hacb == _T_121[11:0] ? image_2763 : _GEN_12044; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12046 = 12'hacc == _T_121[11:0] ? image_2764 : _GEN_12045; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12047 = 12'hacd == _T_121[11:0] ? image_2765 : _GEN_12046; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12048 = 12'hace == _T_121[11:0] ? image_2766 : _GEN_12047; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12049 = 12'hacf == _T_121[11:0] ? image_2767 : _GEN_12048; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12050 = 12'had0 == _T_121[11:0] ? image_2768 : _GEN_12049; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12051 = 12'had1 == _T_121[11:0] ? image_2769 : _GEN_12050; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12052 = 12'had2 == _T_121[11:0] ? image_2770 : _GEN_12051; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12053 = 12'had3 == _T_121[11:0] ? image_2771 : _GEN_12052; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12054 = 12'had4 == _T_121[11:0] ? image_2772 : _GEN_12053; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12055 = 12'had5 == _T_121[11:0] ? image_2773 : _GEN_12054; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12056 = 12'had6 == _T_121[11:0] ? image_2774 : _GEN_12055; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12057 = 12'had7 == _T_121[11:0] ? image_2775 : _GEN_12056; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12058 = 12'had8 == _T_121[11:0] ? image_2776 : _GEN_12057; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12059 = 12'had9 == _T_121[11:0] ? image_2777 : _GEN_12058; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12060 = 12'hada == _T_121[11:0] ? image_2778 : _GEN_12059; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12061 = 12'hadb == _T_121[11:0] ? image_2779 : _GEN_12060; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12062 = 12'hadc == _T_121[11:0] ? image_2780 : _GEN_12061; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12063 = 12'hadd == _T_121[11:0] ? image_2781 : _GEN_12062; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12064 = 12'hade == _T_121[11:0] ? image_2782 : _GEN_12063; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12065 = 12'hadf == _T_121[11:0] ? image_2783 : _GEN_12064; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12066 = 12'hae0 == _T_121[11:0] ? image_2784 : _GEN_12065; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12067 = 12'hae1 == _T_121[11:0] ? image_2785 : _GEN_12066; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12068 = 12'hae2 == _T_121[11:0] ? image_2786 : _GEN_12067; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12069 = 12'hae3 == _T_121[11:0] ? image_2787 : _GEN_12068; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12070 = 12'hae4 == _T_121[11:0] ? image_2788 : _GEN_12069; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12071 = 12'hae5 == _T_121[11:0] ? image_2789 : _GEN_12070; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12072 = 12'hae6 == _T_121[11:0] ? image_2790 : _GEN_12071; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12073 = 12'hae7 == _T_121[11:0] ? image_2791 : _GEN_12072; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12074 = 12'hae8 == _T_121[11:0] ? image_2792 : _GEN_12073; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12075 = 12'hae9 == _T_121[11:0] ? image_2793 : _GEN_12074; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12076 = 12'haea == _T_121[11:0] ? image_2794 : _GEN_12075; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12077 = 12'haeb == _T_121[11:0] ? image_2795 : _GEN_12076; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12078 = 12'haec == _T_121[11:0] ? image_2796 : _GEN_12077; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12079 = 12'haed == _T_121[11:0] ? image_2797 : _GEN_12078; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12080 = 12'haee == _T_121[11:0] ? image_2798 : _GEN_12079; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12081 = 12'haef == _T_121[11:0] ? image_2799 : _GEN_12080; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12082 = 12'haf0 == _T_121[11:0] ? image_2800 : _GEN_12081; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12083 = 12'haf1 == _T_121[11:0] ? image_2801 : _GEN_12082; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12084 = 12'haf2 == _T_121[11:0] ? image_2802 : _GEN_12083; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12085 = 12'haf3 == _T_121[11:0] ? image_2803 : _GEN_12084; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12086 = 12'haf4 == _T_121[11:0] ? image_2804 : _GEN_12085; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12087 = 12'haf5 == _T_121[11:0] ? image_2805 : _GEN_12086; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12088 = 12'haf6 == _T_121[11:0] ? image_2806 : _GEN_12087; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12089 = 12'haf7 == _T_121[11:0] ? image_2807 : _GEN_12088; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12090 = 12'haf8 == _T_121[11:0] ? image_2808 : _GEN_12089; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12091 = 12'haf9 == _T_121[11:0] ? 4'h0 : _GEN_12090; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12092 = 12'hafa == _T_121[11:0] ? 4'h0 : _GEN_12091; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12093 = 12'hafb == _T_121[11:0] ? 4'h0 : _GEN_12092; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12094 = 12'hafc == _T_121[11:0] ? 4'h0 : _GEN_12093; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12095 = 12'hafd == _T_121[11:0] ? 4'h0 : _GEN_12094; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12096 = 12'hafe == _T_121[11:0] ? 4'h0 : _GEN_12095; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12097 = 12'haff == _T_121[11:0] ? 4'h0 : _GEN_12096; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12098 = 12'hb00 == _T_121[11:0] ? 4'h0 : _GEN_12097; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12099 = 12'hb01 == _T_121[11:0] ? 4'h0 : _GEN_12098; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12100 = 12'hb02 == _T_121[11:0] ? 4'h0 : _GEN_12099; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12101 = 12'hb03 == _T_121[11:0] ? 4'h0 : _GEN_12100; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12102 = 12'hb04 == _T_121[11:0] ? 4'h0 : _GEN_12101; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12103 = 12'hb05 == _T_121[11:0] ? 4'h0 : _GEN_12102; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12104 = 12'hb06 == _T_121[11:0] ? 4'h0 : _GEN_12103; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12105 = 12'hb07 == _T_121[11:0] ? 4'h0 : _GEN_12104; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12106 = 12'hb08 == _T_121[11:0] ? 4'h0 : _GEN_12105; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12107 = 12'hb09 == _T_121[11:0] ? 4'h0 : _GEN_12106; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12108 = 12'hb0a == _T_121[11:0] ? 4'h0 : _GEN_12107; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12109 = 12'hb0b == _T_121[11:0] ? 4'h0 : _GEN_12108; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12110 = 12'hb0c == _T_121[11:0] ? image_2828 : _GEN_12109; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12111 = 12'hb0d == _T_121[11:0] ? image_2829 : _GEN_12110; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12112 = 12'hb0e == _T_121[11:0] ? image_2830 : _GEN_12111; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12113 = 12'hb0f == _T_121[11:0] ? image_2831 : _GEN_12112; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12114 = 12'hb10 == _T_121[11:0] ? image_2832 : _GEN_12113; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12115 = 12'hb11 == _T_121[11:0] ? image_2833 : _GEN_12114; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12116 = 12'hb12 == _T_121[11:0] ? image_2834 : _GEN_12115; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12117 = 12'hb13 == _T_121[11:0] ? image_2835 : _GEN_12116; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12118 = 12'hb14 == _T_121[11:0] ? image_2836 : _GEN_12117; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12119 = 12'hb15 == _T_121[11:0] ? image_2837 : _GEN_12118; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12120 = 12'hb16 == _T_121[11:0] ? image_2838 : _GEN_12119; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12121 = 12'hb17 == _T_121[11:0] ? image_2839 : _GEN_12120; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12122 = 12'hb18 == _T_121[11:0] ? image_2840 : _GEN_12121; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12123 = 12'hb19 == _T_121[11:0] ? image_2841 : _GEN_12122; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12124 = 12'hb1a == _T_121[11:0] ? image_2842 : _GEN_12123; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12125 = 12'hb1b == _T_121[11:0] ? image_2843 : _GEN_12124; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12126 = 12'hb1c == _T_121[11:0] ? image_2844 : _GEN_12125; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12127 = 12'hb1d == _T_121[11:0] ? image_2845 : _GEN_12126; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12128 = 12'hb1e == _T_121[11:0] ? image_2846 : _GEN_12127; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12129 = 12'hb1f == _T_121[11:0] ? image_2847 : _GEN_12128; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12130 = 12'hb20 == _T_121[11:0] ? image_2848 : _GEN_12129; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12131 = 12'hb21 == _T_121[11:0] ? image_2849 : _GEN_12130; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12132 = 12'hb22 == _T_121[11:0] ? image_2850 : _GEN_12131; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12133 = 12'hb23 == _T_121[11:0] ? image_2851 : _GEN_12132; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12134 = 12'hb24 == _T_121[11:0] ? image_2852 : _GEN_12133; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12135 = 12'hb25 == _T_121[11:0] ? image_2853 : _GEN_12134; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12136 = 12'hb26 == _T_121[11:0] ? image_2854 : _GEN_12135; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12137 = 12'hb27 == _T_121[11:0] ? image_2855 : _GEN_12136; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12138 = 12'hb28 == _T_121[11:0] ? image_2856 : _GEN_12137; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12139 = 12'hb29 == _T_121[11:0] ? image_2857 : _GEN_12138; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12140 = 12'hb2a == _T_121[11:0] ? image_2858 : _GEN_12139; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12141 = 12'hb2b == _T_121[11:0] ? image_2859 : _GEN_12140; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12142 = 12'hb2c == _T_121[11:0] ? image_2860 : _GEN_12141; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12143 = 12'hb2d == _T_121[11:0] ? image_2861 : _GEN_12142; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12144 = 12'hb2e == _T_121[11:0] ? image_2862 : _GEN_12143; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12145 = 12'hb2f == _T_121[11:0] ? image_2863 : _GEN_12144; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12146 = 12'hb30 == _T_121[11:0] ? image_2864 : _GEN_12145; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12147 = 12'hb31 == _T_121[11:0] ? image_2865 : _GEN_12146; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12148 = 12'hb32 == _T_121[11:0] ? image_2866 : _GEN_12147; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12149 = 12'hb33 == _T_121[11:0] ? image_2867 : _GEN_12148; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12150 = 12'hb34 == _T_121[11:0] ? image_2868 : _GEN_12149; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12151 = 12'hb35 == _T_121[11:0] ? image_2869 : _GEN_12150; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12152 = 12'hb36 == _T_121[11:0] ? image_2870 : _GEN_12151; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12153 = 12'hb37 == _T_121[11:0] ? image_2871 : _GEN_12152; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12154 = 12'hb38 == _T_121[11:0] ? 4'h0 : _GEN_12153; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12155 = 12'hb39 == _T_121[11:0] ? 4'h0 : _GEN_12154; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12156 = 12'hb3a == _T_121[11:0] ? 4'h0 : _GEN_12155; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12157 = 12'hb3b == _T_121[11:0] ? 4'h0 : _GEN_12156; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12158 = 12'hb3c == _T_121[11:0] ? 4'h0 : _GEN_12157; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12159 = 12'hb3d == _T_121[11:0] ? 4'h0 : _GEN_12158; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12160 = 12'hb3e == _T_121[11:0] ? 4'h0 : _GEN_12159; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12161 = 12'hb3f == _T_121[11:0] ? 4'h0 : _GEN_12160; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12162 = 12'hb40 == _T_121[11:0] ? 4'h0 : _GEN_12161; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12163 = 12'hb41 == _T_121[11:0] ? 4'h0 : _GEN_12162; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12164 = 12'hb42 == _T_121[11:0] ? 4'h0 : _GEN_12163; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12165 = 12'hb43 == _T_121[11:0] ? 4'h0 : _GEN_12164; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12166 = 12'hb44 == _T_121[11:0] ? 4'h0 : _GEN_12165; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12167 = 12'hb45 == _T_121[11:0] ? 4'h0 : _GEN_12166; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12168 = 12'hb46 == _T_121[11:0] ? 4'h0 : _GEN_12167; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12169 = 12'hb47 == _T_121[11:0] ? 4'h0 : _GEN_12168; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12170 = 12'hb48 == _T_121[11:0] ? 4'h0 : _GEN_12169; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12171 = 12'hb49 == _T_121[11:0] ? 4'h0 : _GEN_12170; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12172 = 12'hb4a == _T_121[11:0] ? 4'h0 : _GEN_12171; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12173 = 12'hb4b == _T_121[11:0] ? 4'h0 : _GEN_12172; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12174 = 12'hb4c == _T_121[11:0] ? 4'h0 : _GEN_12173; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12175 = 12'hb4d == _T_121[11:0] ? 4'h0 : _GEN_12174; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12176 = 12'hb4e == _T_121[11:0] ? 4'h0 : _GEN_12175; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12177 = 12'hb4f == _T_121[11:0] ? image_2895 : _GEN_12176; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12178 = 12'hb50 == _T_121[11:0] ? image_2896 : _GEN_12177; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12179 = 12'hb51 == _T_121[11:0] ? image_2897 : _GEN_12178; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12180 = 12'hb52 == _T_121[11:0] ? image_2898 : _GEN_12179; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12181 = 12'hb53 == _T_121[11:0] ? image_2899 : _GEN_12180; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12182 = 12'hb54 == _T_121[11:0] ? image_2900 : _GEN_12181; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12183 = 12'hb55 == _T_121[11:0] ? image_2901 : _GEN_12182; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12184 = 12'hb56 == _T_121[11:0] ? image_2902 : _GEN_12183; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12185 = 12'hb57 == _T_121[11:0] ? image_2903 : _GEN_12184; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12186 = 12'hb58 == _T_121[11:0] ? image_2904 : _GEN_12185; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12187 = 12'hb59 == _T_121[11:0] ? image_2905 : _GEN_12186; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12188 = 12'hb5a == _T_121[11:0] ? image_2906 : _GEN_12187; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12189 = 12'hb5b == _T_121[11:0] ? image_2907 : _GEN_12188; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12190 = 12'hb5c == _T_121[11:0] ? image_2908 : _GEN_12189; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12191 = 12'hb5d == _T_121[11:0] ? image_2909 : _GEN_12190; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12192 = 12'hb5e == _T_121[11:0] ? image_2910 : _GEN_12191; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12193 = 12'hb5f == _T_121[11:0] ? image_2911 : _GEN_12192; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12194 = 12'hb60 == _T_121[11:0] ? image_2912 : _GEN_12193; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12195 = 12'hb61 == _T_121[11:0] ? image_2913 : _GEN_12194; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12196 = 12'hb62 == _T_121[11:0] ? image_2914 : _GEN_12195; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12197 = 12'hb63 == _T_121[11:0] ? image_2915 : _GEN_12196; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12198 = 12'hb64 == _T_121[11:0] ? image_2916 : _GEN_12197; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12199 = 12'hb65 == _T_121[11:0] ? image_2917 : _GEN_12198; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12200 = 12'hb66 == _T_121[11:0] ? image_2918 : _GEN_12199; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12201 = 12'hb67 == _T_121[11:0] ? image_2919 : _GEN_12200; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12202 = 12'hb68 == _T_121[11:0] ? image_2920 : _GEN_12201; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12203 = 12'hb69 == _T_121[11:0] ? image_2921 : _GEN_12202; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12204 = 12'hb6a == _T_121[11:0] ? image_2922 : _GEN_12203; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12205 = 12'hb6b == _T_121[11:0] ? image_2923 : _GEN_12204; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12206 = 12'hb6c == _T_121[11:0] ? image_2924 : _GEN_12205; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12207 = 12'hb6d == _T_121[11:0] ? image_2925 : _GEN_12206; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12208 = 12'hb6e == _T_121[11:0] ? image_2926 : _GEN_12207; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12209 = 12'hb6f == _T_121[11:0] ? image_2927 : _GEN_12208; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12210 = 12'hb70 == _T_121[11:0] ? image_2928 : _GEN_12209; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12211 = 12'hb71 == _T_121[11:0] ? image_2929 : _GEN_12210; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12212 = 12'hb72 == _T_121[11:0] ? image_2930 : _GEN_12211; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12213 = 12'hb73 == _T_121[11:0] ? image_2931 : _GEN_12212; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12214 = 12'hb74 == _T_121[11:0] ? image_2932 : _GEN_12213; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12215 = 12'hb75 == _T_121[11:0] ? image_2933 : _GEN_12214; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12216 = 12'hb76 == _T_121[11:0] ? image_2934 : _GEN_12215; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12217 = 12'hb77 == _T_121[11:0] ? 4'h0 : _GEN_12216; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12218 = 12'hb78 == _T_121[11:0] ? 4'h0 : _GEN_12217; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12219 = 12'hb79 == _T_121[11:0] ? 4'h0 : _GEN_12218; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12220 = 12'hb7a == _T_121[11:0] ? 4'h0 : _GEN_12219; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12221 = 12'hb7b == _T_121[11:0] ? 4'h0 : _GEN_12220; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12222 = 12'hb7c == _T_121[11:0] ? 4'h0 : _GEN_12221; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12223 = 12'hb7d == _T_121[11:0] ? 4'h0 : _GEN_12222; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12224 = 12'hb7e == _T_121[11:0] ? 4'h0 : _GEN_12223; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12225 = 12'hb7f == _T_121[11:0] ? 4'h0 : _GEN_12224; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12226 = 12'hb80 == _T_121[11:0] ? 4'h0 : _GEN_12225; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12227 = 12'hb81 == _T_121[11:0] ? 4'h0 : _GEN_12226; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12228 = 12'hb82 == _T_121[11:0] ? 4'h0 : _GEN_12227; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12229 = 12'hb83 == _T_121[11:0] ? 4'h0 : _GEN_12228; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12230 = 12'hb84 == _T_121[11:0] ? 4'h0 : _GEN_12229; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12231 = 12'hb85 == _T_121[11:0] ? 4'h0 : _GEN_12230; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12232 = 12'hb86 == _T_121[11:0] ? 4'h0 : _GEN_12231; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12233 = 12'hb87 == _T_121[11:0] ? 4'h0 : _GEN_12232; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12234 = 12'hb88 == _T_121[11:0] ? 4'h0 : _GEN_12233; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12235 = 12'hb89 == _T_121[11:0] ? 4'h0 : _GEN_12234; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12236 = 12'hb8a == _T_121[11:0] ? 4'h0 : _GEN_12235; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12237 = 12'hb8b == _T_121[11:0] ? 4'h0 : _GEN_12236; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12238 = 12'hb8c == _T_121[11:0] ? 4'h0 : _GEN_12237; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12239 = 12'hb8d == _T_121[11:0] ? 4'h0 : _GEN_12238; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12240 = 12'hb8e == _T_121[11:0] ? 4'h0 : _GEN_12239; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12241 = 12'hb8f == _T_121[11:0] ? 4'h0 : _GEN_12240; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12242 = 12'hb90 == _T_121[11:0] ? 4'h0 : _GEN_12241; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12243 = 12'hb91 == _T_121[11:0] ? 4'h0 : _GEN_12242; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12244 = 12'hb92 == _T_121[11:0] ? 4'h0 : _GEN_12243; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12245 = 12'hb93 == _T_121[11:0] ? 4'h0 : _GEN_12244; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12246 = 12'hb94 == _T_121[11:0] ? 4'h0 : _GEN_12245; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12247 = 12'hb95 == _T_121[11:0] ? image_2965 : _GEN_12246; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12248 = 12'hb96 == _T_121[11:0] ? image_2966 : _GEN_12247; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12249 = 12'hb97 == _T_121[11:0] ? image_2967 : _GEN_12248; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12250 = 12'hb98 == _T_121[11:0] ? image_2968 : _GEN_12249; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12251 = 12'hb99 == _T_121[11:0] ? image_2969 : _GEN_12250; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12252 = 12'hb9a == _T_121[11:0] ? image_2970 : _GEN_12251; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12253 = 12'hb9b == _T_121[11:0] ? image_2971 : _GEN_12252; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12254 = 12'hb9c == _T_121[11:0] ? image_2972 : _GEN_12253; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12255 = 12'hb9d == _T_121[11:0] ? image_2973 : _GEN_12254; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12256 = 12'hb9e == _T_121[11:0] ? image_2974 : _GEN_12255; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12257 = 12'hb9f == _T_121[11:0] ? image_2975 : _GEN_12256; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12258 = 12'hba0 == _T_121[11:0] ? image_2976 : _GEN_12257; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12259 = 12'hba1 == _T_121[11:0] ? image_2977 : _GEN_12258; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12260 = 12'hba2 == _T_121[11:0] ? image_2978 : _GEN_12259; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12261 = 12'hba3 == _T_121[11:0] ? image_2979 : _GEN_12260; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12262 = 12'hba4 == _T_121[11:0] ? image_2980 : _GEN_12261; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12263 = 12'hba5 == _T_121[11:0] ? image_2981 : _GEN_12262; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12264 = 12'hba6 == _T_121[11:0] ? image_2982 : _GEN_12263; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12265 = 12'hba7 == _T_121[11:0] ? image_2983 : _GEN_12264; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12266 = 12'hba8 == _T_121[11:0] ? image_2984 : _GEN_12265; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12267 = 12'hba9 == _T_121[11:0] ? image_2985 : _GEN_12266; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12268 = 12'hbaa == _T_121[11:0] ? image_2986 : _GEN_12267; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12269 = 12'hbab == _T_121[11:0] ? image_2987 : _GEN_12268; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12270 = 12'hbac == _T_121[11:0] ? image_2988 : _GEN_12269; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12271 = 12'hbad == _T_121[11:0] ? image_2989 : _GEN_12270; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12272 = 12'hbae == _T_121[11:0] ? image_2990 : _GEN_12271; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12273 = 12'hbaf == _T_121[11:0] ? image_2991 : _GEN_12272; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12274 = 12'hbb0 == _T_121[11:0] ? image_2992 : _GEN_12273; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12275 = 12'hbb1 == _T_121[11:0] ? image_2993 : _GEN_12274; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12276 = 12'hbb2 == _T_121[11:0] ? image_2994 : _GEN_12275; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12277 = 12'hbb3 == _T_121[11:0] ? image_2995 : _GEN_12276; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12278 = 12'hbb4 == _T_121[11:0] ? image_2996 : _GEN_12277; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12279 = 12'hbb5 == _T_121[11:0] ? 4'h0 : _GEN_12278; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12280 = 12'hbb6 == _T_121[11:0] ? 4'h0 : _GEN_12279; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12281 = 12'hbb7 == _T_121[11:0] ? 4'h0 : _GEN_12280; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12282 = 12'hbb8 == _T_121[11:0] ? 4'h0 : _GEN_12281; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12283 = 12'hbb9 == _T_121[11:0] ? 4'h0 : _GEN_12282; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12284 = 12'hbba == _T_121[11:0] ? 4'h0 : _GEN_12283; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12285 = 12'hbbb == _T_121[11:0] ? 4'h0 : _GEN_12284; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12286 = 12'hbbc == _T_121[11:0] ? 4'h0 : _GEN_12285; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12287 = 12'hbbd == _T_121[11:0] ? 4'h0 : _GEN_12286; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12288 = 12'hbbe == _T_121[11:0] ? 4'h0 : _GEN_12287; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12289 = 12'hbbf == _T_121[11:0] ? 4'h0 : _GEN_12288; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12290 = 12'hbc0 == _T_121[11:0] ? 4'h0 : _GEN_12289; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12291 = 12'hbc1 == _T_121[11:0] ? 4'h0 : _GEN_12290; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12292 = 12'hbc2 == _T_121[11:0] ? 4'h0 : _GEN_12291; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12293 = 12'hbc3 == _T_121[11:0] ? 4'h0 : _GEN_12292; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12294 = 12'hbc4 == _T_121[11:0] ? 4'h0 : _GEN_12293; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12295 = 12'hbc5 == _T_121[11:0] ? 4'h0 : _GEN_12294; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12296 = 12'hbc6 == _T_121[11:0] ? 4'h0 : _GEN_12295; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12297 = 12'hbc7 == _T_121[11:0] ? 4'h0 : _GEN_12296; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12298 = 12'hbc8 == _T_121[11:0] ? 4'h0 : _GEN_12297; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12299 = 12'hbc9 == _T_121[11:0] ? 4'h0 : _GEN_12298; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12300 = 12'hbca == _T_121[11:0] ? 4'h0 : _GEN_12299; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12301 = 12'hbcb == _T_121[11:0] ? 4'h0 : _GEN_12300; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12302 = 12'hbcc == _T_121[11:0] ? 4'h0 : _GEN_12301; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12303 = 12'hbcd == _T_121[11:0] ? 4'h0 : _GEN_12302; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12304 = 12'hbce == _T_121[11:0] ? 4'h0 : _GEN_12303; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12305 = 12'hbcf == _T_121[11:0] ? 4'h0 : _GEN_12304; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12306 = 12'hbd0 == _T_121[11:0] ? 4'h0 : _GEN_12305; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12307 = 12'hbd1 == _T_121[11:0] ? 4'h0 : _GEN_12306; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12308 = 12'hbd2 == _T_121[11:0] ? 4'h0 : _GEN_12307; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12309 = 12'hbd3 == _T_121[11:0] ? 4'h0 : _GEN_12308; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12310 = 12'hbd4 == _T_121[11:0] ? 4'h0 : _GEN_12309; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12311 = 12'hbd5 == _T_121[11:0] ? 4'h0 : _GEN_12310; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12312 = 12'hbd6 == _T_121[11:0] ? 4'h0 : _GEN_12311; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12313 = 12'hbd7 == _T_121[11:0] ? 4'h0 : _GEN_12312; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12314 = 12'hbd8 == _T_121[11:0] ? 4'h0 : _GEN_12313; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12315 = 12'hbd9 == _T_121[11:0] ? 4'h0 : _GEN_12314; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12316 = 12'hbda == _T_121[11:0] ? 4'h0 : _GEN_12315; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12317 = 12'hbdb == _T_121[11:0] ? image_3035 : _GEN_12316; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12318 = 12'hbdc == _T_121[11:0] ? image_3036 : _GEN_12317; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12319 = 12'hbdd == _T_121[11:0] ? image_3037 : _GEN_12318; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12320 = 12'hbde == _T_121[11:0] ? image_3038 : _GEN_12319; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12321 = 12'hbdf == _T_121[11:0] ? image_3039 : _GEN_12320; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12322 = 12'hbe0 == _T_121[11:0] ? image_3040 : _GEN_12321; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12323 = 12'hbe1 == _T_121[11:0] ? image_3041 : _GEN_12322; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12324 = 12'hbe2 == _T_121[11:0] ? image_3042 : _GEN_12323; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12325 = 12'hbe3 == _T_121[11:0] ? image_3043 : _GEN_12324; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12326 = 12'hbe4 == _T_121[11:0] ? image_3044 : _GEN_12325; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12327 = 12'hbe5 == _T_121[11:0] ? image_3045 : _GEN_12326; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12328 = 12'hbe6 == _T_121[11:0] ? image_3046 : _GEN_12327; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12329 = 12'hbe7 == _T_121[11:0] ? image_3047 : _GEN_12328; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12330 = 12'hbe8 == _T_121[11:0] ? image_3048 : _GEN_12329; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12331 = 12'hbe9 == _T_121[11:0] ? image_3049 : _GEN_12330; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12332 = 12'hbea == _T_121[11:0] ? image_3050 : _GEN_12331; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12333 = 12'hbeb == _T_121[11:0] ? image_3051 : _GEN_12332; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12334 = 12'hbec == _T_121[11:0] ? image_3052 : _GEN_12333; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12335 = 12'hbed == _T_121[11:0] ? image_3053 : _GEN_12334; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12336 = 12'hbee == _T_121[11:0] ? image_3054 : _GEN_12335; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12337 = 12'hbef == _T_121[11:0] ? image_3055 : _GEN_12336; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12338 = 12'hbf0 == _T_121[11:0] ? image_3056 : _GEN_12337; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12339 = 12'hbf1 == _T_121[11:0] ? 4'h0 : _GEN_12338; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12340 = 12'hbf2 == _T_121[11:0] ? 4'h0 : _GEN_12339; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12341 = 12'hbf3 == _T_121[11:0] ? 4'h0 : _GEN_12340; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12342 = 12'hbf4 == _T_121[11:0] ? 4'h0 : _GEN_12341; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12343 = 12'hbf5 == _T_121[11:0] ? 4'h0 : _GEN_12342; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12344 = 12'hbf6 == _T_121[11:0] ? 4'h0 : _GEN_12343; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12345 = 12'hbf7 == _T_121[11:0] ? 4'h0 : _GEN_12344; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12346 = 12'hbf8 == _T_121[11:0] ? 4'h0 : _GEN_12345; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12347 = 12'hbf9 == _T_121[11:0] ? 4'h0 : _GEN_12346; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12348 = 12'hbfa == _T_121[11:0] ? 4'h0 : _GEN_12347; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12349 = 12'hbfb == _T_121[11:0] ? 4'h0 : _GEN_12348; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12350 = 12'hbfc == _T_121[11:0] ? 4'h0 : _GEN_12349; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12351 = 12'hbfd == _T_121[11:0] ? 4'h0 : _GEN_12350; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12352 = 12'hbfe == _T_121[11:0] ? 4'h0 : _GEN_12351; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12353 = 12'hbff == _T_121[11:0] ? 4'h0 : _GEN_12352; // @[Filter.scala 138:46]
  wire [31:0] _T_124 = pixelIndex + 32'h4; // @[Filter.scala 133:29]
  wire [31:0] _T_125 = _T_124 / 32'h40; // @[Filter.scala 133:36]
  wire [31:0] _T_127 = _T_125 + _GEN_24805; // @[Filter.scala 133:51]
  wire [31:0] _T_129 = _T_127 - 32'h1; // @[Filter.scala 133:67]
  wire [31:0] _GEN_4 = _T_124 % 32'h40; // @[Filter.scala 134:36]
  wire [6:0] _T_132 = _GEN_4[6:0]; // @[Filter.scala 134:36]
  wire [6:0] _T_134 = _T_132 + _GEN_24806; // @[Filter.scala 134:51]
  wire [6:0] _T_136 = _T_134 - 7'h1; // @[Filter.scala 134:67]
  wire  _T_138 = _T_129 >= 32'h40; // @[Filter.scala 135:27]
  wire  _T_142 = _T_136 >= 7'h30; // @[Filter.scala 135:59]
  wire  _T_143 = _T_138 | _T_142; // @[Filter.scala 135:54]
  wire [13:0] _T_144 = _T_136 * 7'h40; // @[Filter.scala 138:57]
  wire [31:0] _GEN_24819 = {{18'd0}, _T_144}; // @[Filter.scala 138:72]
  wire [31:0] _T_146 = _GEN_24819 + _T_129; // @[Filter.scala 138:72]
  wire [3:0] _GEN_12367 = 12'hc == _T_146[11:0] ? image_12 : 4'h0; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12368 = 12'hd == _T_146[11:0] ? 4'h0 : _GEN_12367; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12369 = 12'he == _T_146[11:0] ? image_14 : _GEN_12368; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12370 = 12'hf == _T_146[11:0] ? image_15 : _GEN_12369; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12371 = 12'h10 == _T_146[11:0] ? image_16 : _GEN_12370; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12372 = 12'h11 == _T_146[11:0] ? image_17 : _GEN_12371; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12373 = 12'h12 == _T_146[11:0] ? image_18 : _GEN_12372; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12374 = 12'h13 == _T_146[11:0] ? image_19 : _GEN_12373; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12375 = 12'h14 == _T_146[11:0] ? image_20 : _GEN_12374; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12376 = 12'h15 == _T_146[11:0] ? image_21 : _GEN_12375; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12377 = 12'h16 == _T_146[11:0] ? image_22 : _GEN_12376; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12378 = 12'h17 == _T_146[11:0] ? image_23 : _GEN_12377; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12379 = 12'h18 == _T_146[11:0] ? 4'h0 : _GEN_12378; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12380 = 12'h19 == _T_146[11:0] ? 4'h0 : _GEN_12379; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12381 = 12'h1a == _T_146[11:0] ? 4'h0 : _GEN_12380; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12382 = 12'h1b == _T_146[11:0] ? 4'h0 : _GEN_12381; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12383 = 12'h1c == _T_146[11:0] ? 4'h0 : _GEN_12382; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12384 = 12'h1d == _T_146[11:0] ? 4'h0 : _GEN_12383; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12385 = 12'h1e == _T_146[11:0] ? 4'h0 : _GEN_12384; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12386 = 12'h1f == _T_146[11:0] ? 4'h0 : _GEN_12385; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12387 = 12'h20 == _T_146[11:0] ? 4'h0 : _GEN_12386; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12388 = 12'h21 == _T_146[11:0] ? 4'h0 : _GEN_12387; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12389 = 12'h22 == _T_146[11:0] ? 4'h0 : _GEN_12388; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12390 = 12'h23 == _T_146[11:0] ? image_35 : _GEN_12389; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12391 = 12'h24 == _T_146[11:0] ? image_36 : _GEN_12390; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12392 = 12'h25 == _T_146[11:0] ? image_37 : _GEN_12391; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12393 = 12'h26 == _T_146[11:0] ? image_38 : _GEN_12392; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12394 = 12'h27 == _T_146[11:0] ? image_39 : _GEN_12393; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12395 = 12'h28 == _T_146[11:0] ? image_40 : _GEN_12394; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12396 = 12'h29 == _T_146[11:0] ? image_41 : _GEN_12395; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12397 = 12'h2a == _T_146[11:0] ? image_42 : _GEN_12396; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12398 = 12'h2b == _T_146[11:0] ? 4'h0 : _GEN_12397; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12399 = 12'h2c == _T_146[11:0] ? 4'h0 : _GEN_12398; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12400 = 12'h2d == _T_146[11:0] ? 4'h0 : _GEN_12399; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12401 = 12'h2e == _T_146[11:0] ? 4'h0 : _GEN_12400; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12402 = 12'h2f == _T_146[11:0] ? 4'h0 : _GEN_12401; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12403 = 12'h30 == _T_146[11:0] ? 4'h0 : _GEN_12402; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12404 = 12'h31 == _T_146[11:0] ? 4'h0 : _GEN_12403; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12405 = 12'h32 == _T_146[11:0] ? 4'h0 : _GEN_12404; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12406 = 12'h33 == _T_146[11:0] ? 4'h0 : _GEN_12405; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12407 = 12'h34 == _T_146[11:0] ? 4'h0 : _GEN_12406; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12408 = 12'h35 == _T_146[11:0] ? 4'h0 : _GEN_12407; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12409 = 12'h36 == _T_146[11:0] ? 4'h0 : _GEN_12408; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12410 = 12'h37 == _T_146[11:0] ? 4'h0 : _GEN_12409; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12411 = 12'h38 == _T_146[11:0] ? 4'h0 : _GEN_12410; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12412 = 12'h39 == _T_146[11:0] ? 4'h0 : _GEN_12411; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12413 = 12'h3a == _T_146[11:0] ? 4'h0 : _GEN_12412; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12414 = 12'h3b == _T_146[11:0] ? 4'h0 : _GEN_12413; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12415 = 12'h3c == _T_146[11:0] ? 4'h0 : _GEN_12414; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12416 = 12'h3d == _T_146[11:0] ? 4'h0 : _GEN_12415; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12417 = 12'h3e == _T_146[11:0] ? 4'h0 : _GEN_12416; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12418 = 12'h3f == _T_146[11:0] ? 4'h0 : _GEN_12417; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12419 = 12'h40 == _T_146[11:0] ? 4'h0 : _GEN_12418; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12420 = 12'h41 == _T_146[11:0] ? 4'h0 : _GEN_12419; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12421 = 12'h42 == _T_146[11:0] ? 4'h0 : _GEN_12420; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12422 = 12'h43 == _T_146[11:0] ? 4'h0 : _GEN_12421; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12423 = 12'h44 == _T_146[11:0] ? 4'h0 : _GEN_12422; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12424 = 12'h45 == _T_146[11:0] ? 4'h0 : _GEN_12423; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12425 = 12'h46 == _T_146[11:0] ? 4'h0 : _GEN_12424; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12426 = 12'h47 == _T_146[11:0] ? 4'h0 : _GEN_12425; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12427 = 12'h48 == _T_146[11:0] ? 4'h0 : _GEN_12426; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12428 = 12'h49 == _T_146[11:0] ? 4'h0 : _GEN_12427; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12429 = 12'h4a == _T_146[11:0] ? 4'h0 : _GEN_12428; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12430 = 12'h4b == _T_146[11:0] ? image_75 : _GEN_12429; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12431 = 12'h4c == _T_146[11:0] ? image_76 : _GEN_12430; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12432 = 12'h4d == _T_146[11:0] ? image_77 : _GEN_12431; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12433 = 12'h4e == _T_146[11:0] ? image_78 : _GEN_12432; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12434 = 12'h4f == _T_146[11:0] ? image_79 : _GEN_12433; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12435 = 12'h50 == _T_146[11:0] ? image_80 : _GEN_12434; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12436 = 12'h51 == _T_146[11:0] ? image_81 : _GEN_12435; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12437 = 12'h52 == _T_146[11:0] ? image_82 : _GEN_12436; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12438 = 12'h53 == _T_146[11:0] ? image_83 : _GEN_12437; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12439 = 12'h54 == _T_146[11:0] ? image_84 : _GEN_12438; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12440 = 12'h55 == _T_146[11:0] ? image_85 : _GEN_12439; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12441 = 12'h56 == _T_146[11:0] ? image_86 : _GEN_12440; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12442 = 12'h57 == _T_146[11:0] ? image_87 : _GEN_12441; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12443 = 12'h58 == _T_146[11:0] ? image_88 : _GEN_12442; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12444 = 12'h59 == _T_146[11:0] ? image_89 : _GEN_12443; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12445 = 12'h5a == _T_146[11:0] ? image_90 : _GEN_12444; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12446 = 12'h5b == _T_146[11:0] ? 4'h0 : _GEN_12445; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12447 = 12'h5c == _T_146[11:0] ? 4'h0 : _GEN_12446; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12448 = 12'h5d == _T_146[11:0] ? image_93 : _GEN_12447; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12449 = 12'h5e == _T_146[11:0] ? 4'h0 : _GEN_12448; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12450 = 12'h5f == _T_146[11:0] ? image_95 : _GEN_12449; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12451 = 12'h60 == _T_146[11:0] ? image_96 : _GEN_12450; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12452 = 12'h61 == _T_146[11:0] ? image_97 : _GEN_12451; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12453 = 12'h62 == _T_146[11:0] ? image_98 : _GEN_12452; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12454 = 12'h63 == _T_146[11:0] ? image_99 : _GEN_12453; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12455 = 12'h64 == _T_146[11:0] ? image_100 : _GEN_12454; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12456 = 12'h65 == _T_146[11:0] ? image_101 : _GEN_12455; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12457 = 12'h66 == _T_146[11:0] ? image_102 : _GEN_12456; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12458 = 12'h67 == _T_146[11:0] ? image_103 : _GEN_12457; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12459 = 12'h68 == _T_146[11:0] ? image_104 : _GEN_12458; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12460 = 12'h69 == _T_146[11:0] ? image_105 : _GEN_12459; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12461 = 12'h6a == _T_146[11:0] ? image_106 : _GEN_12460; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12462 = 12'h6b == _T_146[11:0] ? image_107 : _GEN_12461; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12463 = 12'h6c == _T_146[11:0] ? image_108 : _GEN_12462; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12464 = 12'h6d == _T_146[11:0] ? 4'h0 : _GEN_12463; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12465 = 12'h6e == _T_146[11:0] ? 4'h0 : _GEN_12464; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12466 = 12'h6f == _T_146[11:0] ? 4'h0 : _GEN_12465; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12467 = 12'h70 == _T_146[11:0] ? 4'h0 : _GEN_12466; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12468 = 12'h71 == _T_146[11:0] ? 4'h0 : _GEN_12467; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12469 = 12'h72 == _T_146[11:0] ? 4'h0 : _GEN_12468; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12470 = 12'h73 == _T_146[11:0] ? 4'h0 : _GEN_12469; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12471 = 12'h74 == _T_146[11:0] ? 4'h0 : _GEN_12470; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12472 = 12'h75 == _T_146[11:0] ? 4'h0 : _GEN_12471; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12473 = 12'h76 == _T_146[11:0] ? 4'h0 : _GEN_12472; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12474 = 12'h77 == _T_146[11:0] ? 4'h0 : _GEN_12473; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12475 = 12'h78 == _T_146[11:0] ? 4'h0 : _GEN_12474; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12476 = 12'h79 == _T_146[11:0] ? 4'h0 : _GEN_12475; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12477 = 12'h7a == _T_146[11:0] ? 4'h0 : _GEN_12476; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12478 = 12'h7b == _T_146[11:0] ? 4'h0 : _GEN_12477; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12479 = 12'h7c == _T_146[11:0] ? 4'h0 : _GEN_12478; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12480 = 12'h7d == _T_146[11:0] ? 4'h0 : _GEN_12479; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12481 = 12'h7e == _T_146[11:0] ? 4'h0 : _GEN_12480; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12482 = 12'h7f == _T_146[11:0] ? 4'h0 : _GEN_12481; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12483 = 12'h80 == _T_146[11:0] ? 4'h0 : _GEN_12482; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12484 = 12'h81 == _T_146[11:0] ? 4'h0 : _GEN_12483; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12485 = 12'h82 == _T_146[11:0] ? 4'h0 : _GEN_12484; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12486 = 12'h83 == _T_146[11:0] ? 4'h0 : _GEN_12485; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12487 = 12'h84 == _T_146[11:0] ? 4'h0 : _GEN_12486; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12488 = 12'h85 == _T_146[11:0] ? 4'h0 : _GEN_12487; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12489 = 12'h86 == _T_146[11:0] ? 4'h0 : _GEN_12488; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12490 = 12'h87 == _T_146[11:0] ? 4'h0 : _GEN_12489; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12491 = 12'h88 == _T_146[11:0] ? image_136 : _GEN_12490; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12492 = 12'h89 == _T_146[11:0] ? image_137 : _GEN_12491; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12493 = 12'h8a == _T_146[11:0] ? image_138 : _GEN_12492; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12494 = 12'h8b == _T_146[11:0] ? image_139 : _GEN_12493; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12495 = 12'h8c == _T_146[11:0] ? image_140 : _GEN_12494; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12496 = 12'h8d == _T_146[11:0] ? image_141 : _GEN_12495; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12497 = 12'h8e == _T_146[11:0] ? image_142 : _GEN_12496; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12498 = 12'h8f == _T_146[11:0] ? image_143 : _GEN_12497; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12499 = 12'h90 == _T_146[11:0] ? image_144 : _GEN_12498; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12500 = 12'h91 == _T_146[11:0] ? image_145 : _GEN_12499; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12501 = 12'h92 == _T_146[11:0] ? image_146 : _GEN_12500; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12502 = 12'h93 == _T_146[11:0] ? image_147 : _GEN_12501; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12503 = 12'h94 == _T_146[11:0] ? image_148 : _GEN_12502; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12504 = 12'h95 == _T_146[11:0] ? image_149 : _GEN_12503; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12505 = 12'h96 == _T_146[11:0] ? image_150 : _GEN_12504; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12506 = 12'h97 == _T_146[11:0] ? image_151 : _GEN_12505; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12507 = 12'h98 == _T_146[11:0] ? image_152 : _GEN_12506; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12508 = 12'h99 == _T_146[11:0] ? image_153 : _GEN_12507; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12509 = 12'h9a == _T_146[11:0] ? image_154 : _GEN_12508; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12510 = 12'h9b == _T_146[11:0] ? image_155 : _GEN_12509; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12511 = 12'h9c == _T_146[11:0] ? 4'h0 : _GEN_12510; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12512 = 12'h9d == _T_146[11:0] ? image_157 : _GEN_12511; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12513 = 12'h9e == _T_146[11:0] ? image_158 : _GEN_12512; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12514 = 12'h9f == _T_146[11:0] ? image_159 : _GEN_12513; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12515 = 12'ha0 == _T_146[11:0] ? image_160 : _GEN_12514; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12516 = 12'ha1 == _T_146[11:0] ? image_161 : _GEN_12515; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12517 = 12'ha2 == _T_146[11:0] ? image_162 : _GEN_12516; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12518 = 12'ha3 == _T_146[11:0] ? image_163 : _GEN_12517; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12519 = 12'ha4 == _T_146[11:0] ? image_164 : _GEN_12518; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12520 = 12'ha5 == _T_146[11:0] ? image_165 : _GEN_12519; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12521 = 12'ha6 == _T_146[11:0] ? image_166 : _GEN_12520; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12522 = 12'ha7 == _T_146[11:0] ? image_167 : _GEN_12521; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12523 = 12'ha8 == _T_146[11:0] ? image_168 : _GEN_12522; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12524 = 12'ha9 == _T_146[11:0] ? image_169 : _GEN_12523; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12525 = 12'haa == _T_146[11:0] ? image_170 : _GEN_12524; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12526 = 12'hab == _T_146[11:0] ? image_171 : _GEN_12525; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12527 = 12'hac == _T_146[11:0] ? image_172 : _GEN_12526; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12528 = 12'had == _T_146[11:0] ? image_173 : _GEN_12527; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12529 = 12'hae == _T_146[11:0] ? image_174 : _GEN_12528; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12530 = 12'haf == _T_146[11:0] ? image_175 : _GEN_12529; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12531 = 12'hb0 == _T_146[11:0] ? image_176 : _GEN_12530; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12532 = 12'hb1 == _T_146[11:0] ? image_177 : _GEN_12531; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12533 = 12'hb2 == _T_146[11:0] ? image_178 : _GEN_12532; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12534 = 12'hb3 == _T_146[11:0] ? image_179 : _GEN_12533; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12535 = 12'hb4 == _T_146[11:0] ? 4'h0 : _GEN_12534; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12536 = 12'hb5 == _T_146[11:0] ? 4'h0 : _GEN_12535; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12537 = 12'hb6 == _T_146[11:0] ? 4'h0 : _GEN_12536; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12538 = 12'hb7 == _T_146[11:0] ? 4'h0 : _GEN_12537; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12539 = 12'hb8 == _T_146[11:0] ? 4'h0 : _GEN_12538; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12540 = 12'hb9 == _T_146[11:0] ? 4'h0 : _GEN_12539; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12541 = 12'hba == _T_146[11:0] ? 4'h0 : _GEN_12540; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12542 = 12'hbb == _T_146[11:0] ? 4'h0 : _GEN_12541; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12543 = 12'hbc == _T_146[11:0] ? 4'h0 : _GEN_12542; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12544 = 12'hbd == _T_146[11:0] ? 4'h0 : _GEN_12543; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12545 = 12'hbe == _T_146[11:0] ? 4'h0 : _GEN_12544; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12546 = 12'hbf == _T_146[11:0] ? 4'h0 : _GEN_12545; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12547 = 12'hc0 == _T_146[11:0] ? 4'h0 : _GEN_12546; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12548 = 12'hc1 == _T_146[11:0] ? 4'h0 : _GEN_12547; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12549 = 12'hc2 == _T_146[11:0] ? 4'h0 : _GEN_12548; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12550 = 12'hc3 == _T_146[11:0] ? 4'h0 : _GEN_12549; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12551 = 12'hc4 == _T_146[11:0] ? 4'h0 : _GEN_12550; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12552 = 12'hc5 == _T_146[11:0] ? 4'h0 : _GEN_12551; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12553 = 12'hc6 == _T_146[11:0] ? 4'h0 : _GEN_12552; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12554 = 12'hc7 == _T_146[11:0] ? image_199 : _GEN_12553; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12555 = 12'hc8 == _T_146[11:0] ? image_200 : _GEN_12554; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12556 = 12'hc9 == _T_146[11:0] ? image_201 : _GEN_12555; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12557 = 12'hca == _T_146[11:0] ? image_202 : _GEN_12556; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12558 = 12'hcb == _T_146[11:0] ? image_203 : _GEN_12557; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12559 = 12'hcc == _T_146[11:0] ? image_204 : _GEN_12558; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12560 = 12'hcd == _T_146[11:0] ? image_205 : _GEN_12559; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12561 = 12'hce == _T_146[11:0] ? image_206 : _GEN_12560; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12562 = 12'hcf == _T_146[11:0] ? image_207 : _GEN_12561; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12563 = 12'hd0 == _T_146[11:0] ? image_208 : _GEN_12562; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12564 = 12'hd1 == _T_146[11:0] ? image_209 : _GEN_12563; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12565 = 12'hd2 == _T_146[11:0] ? image_210 : _GEN_12564; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12566 = 12'hd3 == _T_146[11:0] ? image_211 : _GEN_12565; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12567 = 12'hd4 == _T_146[11:0] ? image_212 : _GEN_12566; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12568 = 12'hd5 == _T_146[11:0] ? image_213 : _GEN_12567; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12569 = 12'hd6 == _T_146[11:0] ? image_214 : _GEN_12568; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12570 = 12'hd7 == _T_146[11:0] ? image_215 : _GEN_12569; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12571 = 12'hd8 == _T_146[11:0] ? image_216 : _GEN_12570; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12572 = 12'hd9 == _T_146[11:0] ? image_217 : _GEN_12571; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12573 = 12'hda == _T_146[11:0] ? image_218 : _GEN_12572; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12574 = 12'hdb == _T_146[11:0] ? image_219 : _GEN_12573; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12575 = 12'hdc == _T_146[11:0] ? image_220 : _GEN_12574; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12576 = 12'hdd == _T_146[11:0] ? image_221 : _GEN_12575; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12577 = 12'hde == _T_146[11:0] ? image_222 : _GEN_12576; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12578 = 12'hdf == _T_146[11:0] ? image_223 : _GEN_12577; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12579 = 12'he0 == _T_146[11:0] ? image_224 : _GEN_12578; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12580 = 12'he1 == _T_146[11:0] ? image_225 : _GEN_12579; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12581 = 12'he2 == _T_146[11:0] ? image_226 : _GEN_12580; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12582 = 12'he3 == _T_146[11:0] ? image_227 : _GEN_12581; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12583 = 12'he4 == _T_146[11:0] ? image_228 : _GEN_12582; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12584 = 12'he5 == _T_146[11:0] ? image_229 : _GEN_12583; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12585 = 12'he6 == _T_146[11:0] ? image_230 : _GEN_12584; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12586 = 12'he7 == _T_146[11:0] ? image_231 : _GEN_12585; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12587 = 12'he8 == _T_146[11:0] ? image_232 : _GEN_12586; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12588 = 12'he9 == _T_146[11:0] ? image_233 : _GEN_12587; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12589 = 12'hea == _T_146[11:0] ? image_234 : _GEN_12588; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12590 = 12'heb == _T_146[11:0] ? image_235 : _GEN_12589; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12591 = 12'hec == _T_146[11:0] ? image_236 : _GEN_12590; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12592 = 12'hed == _T_146[11:0] ? image_237 : _GEN_12591; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12593 = 12'hee == _T_146[11:0] ? image_238 : _GEN_12592; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12594 = 12'hef == _T_146[11:0] ? image_239 : _GEN_12593; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12595 = 12'hf0 == _T_146[11:0] ? image_240 : _GEN_12594; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12596 = 12'hf1 == _T_146[11:0] ? image_241 : _GEN_12595; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12597 = 12'hf2 == _T_146[11:0] ? image_242 : _GEN_12596; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12598 = 12'hf3 == _T_146[11:0] ? image_243 : _GEN_12597; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12599 = 12'hf4 == _T_146[11:0] ? image_244 : _GEN_12598; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12600 = 12'hf5 == _T_146[11:0] ? image_245 : _GEN_12599; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12601 = 12'hf6 == _T_146[11:0] ? image_246 : _GEN_12600; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12602 = 12'hf7 == _T_146[11:0] ? 4'h0 : _GEN_12601; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12603 = 12'hf8 == _T_146[11:0] ? 4'h0 : _GEN_12602; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12604 = 12'hf9 == _T_146[11:0] ? 4'h0 : _GEN_12603; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12605 = 12'hfa == _T_146[11:0] ? 4'h0 : _GEN_12604; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12606 = 12'hfb == _T_146[11:0] ? 4'h0 : _GEN_12605; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12607 = 12'hfc == _T_146[11:0] ? 4'h0 : _GEN_12606; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12608 = 12'hfd == _T_146[11:0] ? 4'h0 : _GEN_12607; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12609 = 12'hfe == _T_146[11:0] ? 4'h0 : _GEN_12608; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12610 = 12'hff == _T_146[11:0] ? 4'h0 : _GEN_12609; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12611 = 12'h100 == _T_146[11:0] ? 4'h0 : _GEN_12610; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12612 = 12'h101 == _T_146[11:0] ? 4'h0 : _GEN_12611; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12613 = 12'h102 == _T_146[11:0] ? 4'h0 : _GEN_12612; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12614 = 12'h103 == _T_146[11:0] ? 4'h0 : _GEN_12613; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12615 = 12'h104 == _T_146[11:0] ? 4'h0 : _GEN_12614; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12616 = 12'h105 == _T_146[11:0] ? 4'h0 : _GEN_12615; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12617 = 12'h106 == _T_146[11:0] ? image_262 : _GEN_12616; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12618 = 12'h107 == _T_146[11:0] ? image_263 : _GEN_12617; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12619 = 12'h108 == _T_146[11:0] ? image_264 : _GEN_12618; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12620 = 12'h109 == _T_146[11:0] ? image_265 : _GEN_12619; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12621 = 12'h10a == _T_146[11:0] ? image_266 : _GEN_12620; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12622 = 12'h10b == _T_146[11:0] ? image_267 : _GEN_12621; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12623 = 12'h10c == _T_146[11:0] ? image_268 : _GEN_12622; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12624 = 12'h10d == _T_146[11:0] ? image_269 : _GEN_12623; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12625 = 12'h10e == _T_146[11:0] ? image_270 : _GEN_12624; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12626 = 12'h10f == _T_146[11:0] ? image_271 : _GEN_12625; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12627 = 12'h110 == _T_146[11:0] ? image_272 : _GEN_12626; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12628 = 12'h111 == _T_146[11:0] ? image_273 : _GEN_12627; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12629 = 12'h112 == _T_146[11:0] ? image_274 : _GEN_12628; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12630 = 12'h113 == _T_146[11:0] ? image_275 : _GEN_12629; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12631 = 12'h114 == _T_146[11:0] ? image_276 : _GEN_12630; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12632 = 12'h115 == _T_146[11:0] ? image_277 : _GEN_12631; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12633 = 12'h116 == _T_146[11:0] ? image_278 : _GEN_12632; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12634 = 12'h117 == _T_146[11:0] ? image_279 : _GEN_12633; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12635 = 12'h118 == _T_146[11:0] ? image_280 : _GEN_12634; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12636 = 12'h119 == _T_146[11:0] ? image_281 : _GEN_12635; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12637 = 12'h11a == _T_146[11:0] ? image_282 : _GEN_12636; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12638 = 12'h11b == _T_146[11:0] ? image_283 : _GEN_12637; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12639 = 12'h11c == _T_146[11:0] ? image_284 : _GEN_12638; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12640 = 12'h11d == _T_146[11:0] ? image_285 : _GEN_12639; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12641 = 12'h11e == _T_146[11:0] ? image_286 : _GEN_12640; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12642 = 12'h11f == _T_146[11:0] ? image_287 : _GEN_12641; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12643 = 12'h120 == _T_146[11:0] ? image_288 : _GEN_12642; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12644 = 12'h121 == _T_146[11:0] ? image_289 : _GEN_12643; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12645 = 12'h122 == _T_146[11:0] ? image_290 : _GEN_12644; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12646 = 12'h123 == _T_146[11:0] ? image_291 : _GEN_12645; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12647 = 12'h124 == _T_146[11:0] ? image_292 : _GEN_12646; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12648 = 12'h125 == _T_146[11:0] ? image_293 : _GEN_12647; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12649 = 12'h126 == _T_146[11:0] ? image_294 : _GEN_12648; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12650 = 12'h127 == _T_146[11:0] ? image_295 : _GEN_12649; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12651 = 12'h128 == _T_146[11:0] ? image_296 : _GEN_12650; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12652 = 12'h129 == _T_146[11:0] ? image_297 : _GEN_12651; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12653 = 12'h12a == _T_146[11:0] ? image_298 : _GEN_12652; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12654 = 12'h12b == _T_146[11:0] ? image_299 : _GEN_12653; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12655 = 12'h12c == _T_146[11:0] ? image_300 : _GEN_12654; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12656 = 12'h12d == _T_146[11:0] ? image_301 : _GEN_12655; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12657 = 12'h12e == _T_146[11:0] ? image_302 : _GEN_12656; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12658 = 12'h12f == _T_146[11:0] ? image_303 : _GEN_12657; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12659 = 12'h130 == _T_146[11:0] ? image_304 : _GEN_12658; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12660 = 12'h131 == _T_146[11:0] ? image_305 : _GEN_12659; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12661 = 12'h132 == _T_146[11:0] ? image_306 : _GEN_12660; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12662 = 12'h133 == _T_146[11:0] ? image_307 : _GEN_12661; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12663 = 12'h134 == _T_146[11:0] ? image_308 : _GEN_12662; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12664 = 12'h135 == _T_146[11:0] ? image_309 : _GEN_12663; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12665 = 12'h136 == _T_146[11:0] ? image_310 : _GEN_12664; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12666 = 12'h137 == _T_146[11:0] ? image_311 : _GEN_12665; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12667 = 12'h138 == _T_146[11:0] ? image_312 : _GEN_12666; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12668 = 12'h139 == _T_146[11:0] ? image_313 : _GEN_12667; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12669 = 12'h13a == _T_146[11:0] ? image_314 : _GEN_12668; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12670 = 12'h13b == _T_146[11:0] ? image_315 : _GEN_12669; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12671 = 12'h13c == _T_146[11:0] ? 4'h0 : _GEN_12670; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12672 = 12'h13d == _T_146[11:0] ? 4'h0 : _GEN_12671; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12673 = 12'h13e == _T_146[11:0] ? 4'h0 : _GEN_12672; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12674 = 12'h13f == _T_146[11:0] ? 4'h0 : _GEN_12673; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12675 = 12'h140 == _T_146[11:0] ? 4'h0 : _GEN_12674; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12676 = 12'h141 == _T_146[11:0] ? 4'h0 : _GEN_12675; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12677 = 12'h142 == _T_146[11:0] ? 4'h0 : _GEN_12676; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12678 = 12'h143 == _T_146[11:0] ? 4'h0 : _GEN_12677; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12679 = 12'h144 == _T_146[11:0] ? 4'h0 : _GEN_12678; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12680 = 12'h145 == _T_146[11:0] ? image_325 : _GEN_12679; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12681 = 12'h146 == _T_146[11:0] ? image_326 : _GEN_12680; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12682 = 12'h147 == _T_146[11:0] ? image_327 : _GEN_12681; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12683 = 12'h148 == _T_146[11:0] ? image_328 : _GEN_12682; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12684 = 12'h149 == _T_146[11:0] ? image_329 : _GEN_12683; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12685 = 12'h14a == _T_146[11:0] ? image_330 : _GEN_12684; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12686 = 12'h14b == _T_146[11:0] ? image_331 : _GEN_12685; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12687 = 12'h14c == _T_146[11:0] ? image_332 : _GEN_12686; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12688 = 12'h14d == _T_146[11:0] ? image_333 : _GEN_12687; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12689 = 12'h14e == _T_146[11:0] ? image_334 : _GEN_12688; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12690 = 12'h14f == _T_146[11:0] ? image_335 : _GEN_12689; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12691 = 12'h150 == _T_146[11:0] ? image_336 : _GEN_12690; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12692 = 12'h151 == _T_146[11:0] ? image_337 : _GEN_12691; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12693 = 12'h152 == _T_146[11:0] ? image_338 : _GEN_12692; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12694 = 12'h153 == _T_146[11:0] ? image_339 : _GEN_12693; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12695 = 12'h154 == _T_146[11:0] ? image_340 : _GEN_12694; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12696 = 12'h155 == _T_146[11:0] ? image_341 : _GEN_12695; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12697 = 12'h156 == _T_146[11:0] ? image_342 : _GEN_12696; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12698 = 12'h157 == _T_146[11:0] ? image_343 : _GEN_12697; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12699 = 12'h158 == _T_146[11:0] ? image_344 : _GEN_12698; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12700 = 12'h159 == _T_146[11:0] ? image_345 : _GEN_12699; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12701 = 12'h15a == _T_146[11:0] ? image_346 : _GEN_12700; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12702 = 12'h15b == _T_146[11:0] ? image_347 : _GEN_12701; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12703 = 12'h15c == _T_146[11:0] ? image_348 : _GEN_12702; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12704 = 12'h15d == _T_146[11:0] ? image_349 : _GEN_12703; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12705 = 12'h15e == _T_146[11:0] ? image_350 : _GEN_12704; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12706 = 12'h15f == _T_146[11:0] ? image_351 : _GEN_12705; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12707 = 12'h160 == _T_146[11:0] ? image_352 : _GEN_12706; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12708 = 12'h161 == _T_146[11:0] ? image_353 : _GEN_12707; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12709 = 12'h162 == _T_146[11:0] ? image_354 : _GEN_12708; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12710 = 12'h163 == _T_146[11:0] ? image_355 : _GEN_12709; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12711 = 12'h164 == _T_146[11:0] ? image_356 : _GEN_12710; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12712 = 12'h165 == _T_146[11:0] ? image_357 : _GEN_12711; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12713 = 12'h166 == _T_146[11:0] ? image_358 : _GEN_12712; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12714 = 12'h167 == _T_146[11:0] ? image_359 : _GEN_12713; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12715 = 12'h168 == _T_146[11:0] ? image_360 : _GEN_12714; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12716 = 12'h169 == _T_146[11:0] ? image_361 : _GEN_12715; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12717 = 12'h16a == _T_146[11:0] ? image_362 : _GEN_12716; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12718 = 12'h16b == _T_146[11:0] ? image_363 : _GEN_12717; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12719 = 12'h16c == _T_146[11:0] ? image_364 : _GEN_12718; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12720 = 12'h16d == _T_146[11:0] ? image_365 : _GEN_12719; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12721 = 12'h16e == _T_146[11:0] ? image_366 : _GEN_12720; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12722 = 12'h16f == _T_146[11:0] ? image_367 : _GEN_12721; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12723 = 12'h170 == _T_146[11:0] ? image_368 : _GEN_12722; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12724 = 12'h171 == _T_146[11:0] ? image_369 : _GEN_12723; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12725 = 12'h172 == _T_146[11:0] ? image_370 : _GEN_12724; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12726 = 12'h173 == _T_146[11:0] ? image_371 : _GEN_12725; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12727 = 12'h174 == _T_146[11:0] ? image_372 : _GEN_12726; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12728 = 12'h175 == _T_146[11:0] ? image_373 : _GEN_12727; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12729 = 12'h176 == _T_146[11:0] ? image_374 : _GEN_12728; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12730 = 12'h177 == _T_146[11:0] ? image_375 : _GEN_12729; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12731 = 12'h178 == _T_146[11:0] ? image_376 : _GEN_12730; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12732 = 12'h179 == _T_146[11:0] ? image_377 : _GEN_12731; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12733 = 12'h17a == _T_146[11:0] ? image_378 : _GEN_12732; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12734 = 12'h17b == _T_146[11:0] ? image_379 : _GEN_12733; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12735 = 12'h17c == _T_146[11:0] ? 4'h0 : _GEN_12734; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12736 = 12'h17d == _T_146[11:0] ? 4'h0 : _GEN_12735; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12737 = 12'h17e == _T_146[11:0] ? 4'h0 : _GEN_12736; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12738 = 12'h17f == _T_146[11:0] ? 4'h0 : _GEN_12737; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12739 = 12'h180 == _T_146[11:0] ? 4'h0 : _GEN_12738; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12740 = 12'h181 == _T_146[11:0] ? 4'h0 : _GEN_12739; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12741 = 12'h182 == _T_146[11:0] ? 4'h0 : _GEN_12740; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12742 = 12'h183 == _T_146[11:0] ? 4'h0 : _GEN_12741; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12743 = 12'h184 == _T_146[11:0] ? image_388 : _GEN_12742; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12744 = 12'h185 == _T_146[11:0] ? image_389 : _GEN_12743; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12745 = 12'h186 == _T_146[11:0] ? image_390 : _GEN_12744; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12746 = 12'h187 == _T_146[11:0] ? image_391 : _GEN_12745; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12747 = 12'h188 == _T_146[11:0] ? image_392 : _GEN_12746; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12748 = 12'h189 == _T_146[11:0] ? image_393 : _GEN_12747; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12749 = 12'h18a == _T_146[11:0] ? image_394 : _GEN_12748; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12750 = 12'h18b == _T_146[11:0] ? image_395 : _GEN_12749; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12751 = 12'h18c == _T_146[11:0] ? image_396 : _GEN_12750; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12752 = 12'h18d == _T_146[11:0] ? image_397 : _GEN_12751; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12753 = 12'h18e == _T_146[11:0] ? image_398 : _GEN_12752; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12754 = 12'h18f == _T_146[11:0] ? image_399 : _GEN_12753; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12755 = 12'h190 == _T_146[11:0] ? image_400 : _GEN_12754; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12756 = 12'h191 == _T_146[11:0] ? image_401 : _GEN_12755; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12757 = 12'h192 == _T_146[11:0] ? image_402 : _GEN_12756; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12758 = 12'h193 == _T_146[11:0] ? image_403 : _GEN_12757; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12759 = 12'h194 == _T_146[11:0] ? image_404 : _GEN_12758; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12760 = 12'h195 == _T_146[11:0] ? image_405 : _GEN_12759; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12761 = 12'h196 == _T_146[11:0] ? image_406 : _GEN_12760; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12762 = 12'h197 == _T_146[11:0] ? image_407 : _GEN_12761; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12763 = 12'h198 == _T_146[11:0] ? image_408 : _GEN_12762; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12764 = 12'h199 == _T_146[11:0] ? image_409 : _GEN_12763; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12765 = 12'h19a == _T_146[11:0] ? image_410 : _GEN_12764; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12766 = 12'h19b == _T_146[11:0] ? image_411 : _GEN_12765; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12767 = 12'h19c == _T_146[11:0] ? image_412 : _GEN_12766; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12768 = 12'h19d == _T_146[11:0] ? image_413 : _GEN_12767; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12769 = 12'h19e == _T_146[11:0] ? image_414 : _GEN_12768; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12770 = 12'h19f == _T_146[11:0] ? image_415 : _GEN_12769; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12771 = 12'h1a0 == _T_146[11:0] ? image_416 : _GEN_12770; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12772 = 12'h1a1 == _T_146[11:0] ? image_417 : _GEN_12771; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12773 = 12'h1a2 == _T_146[11:0] ? image_418 : _GEN_12772; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12774 = 12'h1a3 == _T_146[11:0] ? image_419 : _GEN_12773; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12775 = 12'h1a4 == _T_146[11:0] ? image_420 : _GEN_12774; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12776 = 12'h1a5 == _T_146[11:0] ? image_421 : _GEN_12775; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12777 = 12'h1a6 == _T_146[11:0] ? image_422 : _GEN_12776; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12778 = 12'h1a7 == _T_146[11:0] ? image_423 : _GEN_12777; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12779 = 12'h1a8 == _T_146[11:0] ? image_424 : _GEN_12778; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12780 = 12'h1a9 == _T_146[11:0] ? image_425 : _GEN_12779; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12781 = 12'h1aa == _T_146[11:0] ? image_426 : _GEN_12780; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12782 = 12'h1ab == _T_146[11:0] ? image_427 : _GEN_12781; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12783 = 12'h1ac == _T_146[11:0] ? image_428 : _GEN_12782; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12784 = 12'h1ad == _T_146[11:0] ? image_429 : _GEN_12783; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12785 = 12'h1ae == _T_146[11:0] ? image_430 : _GEN_12784; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12786 = 12'h1af == _T_146[11:0] ? image_431 : _GEN_12785; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12787 = 12'h1b0 == _T_146[11:0] ? image_432 : _GEN_12786; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12788 = 12'h1b1 == _T_146[11:0] ? image_433 : _GEN_12787; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12789 = 12'h1b2 == _T_146[11:0] ? image_434 : _GEN_12788; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12790 = 12'h1b3 == _T_146[11:0] ? image_435 : _GEN_12789; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12791 = 12'h1b4 == _T_146[11:0] ? image_436 : _GEN_12790; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12792 = 12'h1b5 == _T_146[11:0] ? image_437 : _GEN_12791; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12793 = 12'h1b6 == _T_146[11:0] ? image_438 : _GEN_12792; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12794 = 12'h1b7 == _T_146[11:0] ? image_439 : _GEN_12793; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12795 = 12'h1b8 == _T_146[11:0] ? image_440 : _GEN_12794; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12796 = 12'h1b9 == _T_146[11:0] ? image_441 : _GEN_12795; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12797 = 12'h1ba == _T_146[11:0] ? image_442 : _GEN_12796; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12798 = 12'h1bb == _T_146[11:0] ? image_443 : _GEN_12797; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12799 = 12'h1bc == _T_146[11:0] ? image_444 : _GEN_12798; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12800 = 12'h1bd == _T_146[11:0] ? 4'h0 : _GEN_12799; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12801 = 12'h1be == _T_146[11:0] ? 4'h0 : _GEN_12800; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12802 = 12'h1bf == _T_146[11:0] ? 4'h0 : _GEN_12801; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12803 = 12'h1c0 == _T_146[11:0] ? 4'h0 : _GEN_12802; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12804 = 12'h1c1 == _T_146[11:0] ? 4'h0 : _GEN_12803; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12805 = 12'h1c2 == _T_146[11:0] ? 4'h0 : _GEN_12804; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12806 = 12'h1c3 == _T_146[11:0] ? image_451 : _GEN_12805; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12807 = 12'h1c4 == _T_146[11:0] ? image_452 : _GEN_12806; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12808 = 12'h1c5 == _T_146[11:0] ? image_453 : _GEN_12807; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12809 = 12'h1c6 == _T_146[11:0] ? image_454 : _GEN_12808; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12810 = 12'h1c7 == _T_146[11:0] ? image_455 : _GEN_12809; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12811 = 12'h1c8 == _T_146[11:0] ? image_456 : _GEN_12810; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12812 = 12'h1c9 == _T_146[11:0] ? image_457 : _GEN_12811; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12813 = 12'h1ca == _T_146[11:0] ? image_458 : _GEN_12812; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12814 = 12'h1cb == _T_146[11:0] ? image_459 : _GEN_12813; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12815 = 12'h1cc == _T_146[11:0] ? image_460 : _GEN_12814; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12816 = 12'h1cd == _T_146[11:0] ? image_461 : _GEN_12815; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12817 = 12'h1ce == _T_146[11:0] ? image_462 : _GEN_12816; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12818 = 12'h1cf == _T_146[11:0] ? image_463 : _GEN_12817; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12819 = 12'h1d0 == _T_146[11:0] ? image_464 : _GEN_12818; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12820 = 12'h1d1 == _T_146[11:0] ? image_465 : _GEN_12819; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12821 = 12'h1d2 == _T_146[11:0] ? image_466 : _GEN_12820; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12822 = 12'h1d3 == _T_146[11:0] ? image_467 : _GEN_12821; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12823 = 12'h1d4 == _T_146[11:0] ? image_468 : _GEN_12822; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12824 = 12'h1d5 == _T_146[11:0] ? image_469 : _GEN_12823; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12825 = 12'h1d6 == _T_146[11:0] ? image_470 : _GEN_12824; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12826 = 12'h1d7 == _T_146[11:0] ? image_471 : _GEN_12825; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12827 = 12'h1d8 == _T_146[11:0] ? image_472 : _GEN_12826; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12828 = 12'h1d9 == _T_146[11:0] ? image_473 : _GEN_12827; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12829 = 12'h1da == _T_146[11:0] ? image_474 : _GEN_12828; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12830 = 12'h1db == _T_146[11:0] ? image_475 : _GEN_12829; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12831 = 12'h1dc == _T_146[11:0] ? image_476 : _GEN_12830; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12832 = 12'h1dd == _T_146[11:0] ? image_477 : _GEN_12831; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12833 = 12'h1de == _T_146[11:0] ? image_478 : _GEN_12832; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12834 = 12'h1df == _T_146[11:0] ? image_479 : _GEN_12833; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12835 = 12'h1e0 == _T_146[11:0] ? image_480 : _GEN_12834; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12836 = 12'h1e1 == _T_146[11:0] ? image_481 : _GEN_12835; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12837 = 12'h1e2 == _T_146[11:0] ? image_482 : _GEN_12836; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12838 = 12'h1e3 == _T_146[11:0] ? image_483 : _GEN_12837; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12839 = 12'h1e4 == _T_146[11:0] ? image_484 : _GEN_12838; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12840 = 12'h1e5 == _T_146[11:0] ? image_485 : _GEN_12839; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12841 = 12'h1e6 == _T_146[11:0] ? image_486 : _GEN_12840; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12842 = 12'h1e7 == _T_146[11:0] ? image_487 : _GEN_12841; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12843 = 12'h1e8 == _T_146[11:0] ? image_488 : _GEN_12842; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12844 = 12'h1e9 == _T_146[11:0] ? image_489 : _GEN_12843; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12845 = 12'h1ea == _T_146[11:0] ? image_490 : _GEN_12844; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12846 = 12'h1eb == _T_146[11:0] ? image_491 : _GEN_12845; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12847 = 12'h1ec == _T_146[11:0] ? image_492 : _GEN_12846; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12848 = 12'h1ed == _T_146[11:0] ? image_493 : _GEN_12847; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12849 = 12'h1ee == _T_146[11:0] ? image_494 : _GEN_12848; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12850 = 12'h1ef == _T_146[11:0] ? image_495 : _GEN_12849; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12851 = 12'h1f0 == _T_146[11:0] ? image_496 : _GEN_12850; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12852 = 12'h1f1 == _T_146[11:0] ? image_497 : _GEN_12851; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12853 = 12'h1f2 == _T_146[11:0] ? image_498 : _GEN_12852; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12854 = 12'h1f3 == _T_146[11:0] ? image_499 : _GEN_12853; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12855 = 12'h1f4 == _T_146[11:0] ? image_500 : _GEN_12854; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12856 = 12'h1f5 == _T_146[11:0] ? image_501 : _GEN_12855; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12857 = 12'h1f6 == _T_146[11:0] ? image_502 : _GEN_12856; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12858 = 12'h1f7 == _T_146[11:0] ? image_503 : _GEN_12857; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12859 = 12'h1f8 == _T_146[11:0] ? image_504 : _GEN_12858; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12860 = 12'h1f9 == _T_146[11:0] ? image_505 : _GEN_12859; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12861 = 12'h1fa == _T_146[11:0] ? image_506 : _GEN_12860; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12862 = 12'h1fb == _T_146[11:0] ? image_507 : _GEN_12861; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12863 = 12'h1fc == _T_146[11:0] ? image_508 : _GEN_12862; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12864 = 12'h1fd == _T_146[11:0] ? image_509 : _GEN_12863; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12865 = 12'h1fe == _T_146[11:0] ? 4'h0 : _GEN_12864; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12866 = 12'h1ff == _T_146[11:0] ? 4'h0 : _GEN_12865; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12867 = 12'h200 == _T_146[11:0] ? 4'h0 : _GEN_12866; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12868 = 12'h201 == _T_146[11:0] ? 4'h0 : _GEN_12867; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12869 = 12'h202 == _T_146[11:0] ? 4'h0 : _GEN_12868; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12870 = 12'h203 == _T_146[11:0] ? image_515 : _GEN_12869; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12871 = 12'h204 == _T_146[11:0] ? image_516 : _GEN_12870; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12872 = 12'h205 == _T_146[11:0] ? image_517 : _GEN_12871; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12873 = 12'h206 == _T_146[11:0] ? image_518 : _GEN_12872; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12874 = 12'h207 == _T_146[11:0] ? image_519 : _GEN_12873; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12875 = 12'h208 == _T_146[11:0] ? image_520 : _GEN_12874; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12876 = 12'h209 == _T_146[11:0] ? image_521 : _GEN_12875; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12877 = 12'h20a == _T_146[11:0] ? image_522 : _GEN_12876; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12878 = 12'h20b == _T_146[11:0] ? image_523 : _GEN_12877; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12879 = 12'h20c == _T_146[11:0] ? image_524 : _GEN_12878; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12880 = 12'h20d == _T_146[11:0] ? image_525 : _GEN_12879; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12881 = 12'h20e == _T_146[11:0] ? image_526 : _GEN_12880; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12882 = 12'h20f == _T_146[11:0] ? image_527 : _GEN_12881; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12883 = 12'h210 == _T_146[11:0] ? image_528 : _GEN_12882; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12884 = 12'h211 == _T_146[11:0] ? image_529 : _GEN_12883; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12885 = 12'h212 == _T_146[11:0] ? image_530 : _GEN_12884; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12886 = 12'h213 == _T_146[11:0] ? image_531 : _GEN_12885; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12887 = 12'h214 == _T_146[11:0] ? image_532 : _GEN_12886; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12888 = 12'h215 == _T_146[11:0] ? image_533 : _GEN_12887; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12889 = 12'h216 == _T_146[11:0] ? image_534 : _GEN_12888; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12890 = 12'h217 == _T_146[11:0] ? image_535 : _GEN_12889; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12891 = 12'h218 == _T_146[11:0] ? image_536 : _GEN_12890; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12892 = 12'h219 == _T_146[11:0] ? image_537 : _GEN_12891; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12893 = 12'h21a == _T_146[11:0] ? image_538 : _GEN_12892; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12894 = 12'h21b == _T_146[11:0] ? image_539 : _GEN_12893; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12895 = 12'h21c == _T_146[11:0] ? image_540 : _GEN_12894; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12896 = 12'h21d == _T_146[11:0] ? image_541 : _GEN_12895; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12897 = 12'h21e == _T_146[11:0] ? image_542 : _GEN_12896; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12898 = 12'h21f == _T_146[11:0] ? image_543 : _GEN_12897; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12899 = 12'h220 == _T_146[11:0] ? image_544 : _GEN_12898; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12900 = 12'h221 == _T_146[11:0] ? image_545 : _GEN_12899; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12901 = 12'h222 == _T_146[11:0] ? image_546 : _GEN_12900; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12902 = 12'h223 == _T_146[11:0] ? image_547 : _GEN_12901; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12903 = 12'h224 == _T_146[11:0] ? image_548 : _GEN_12902; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12904 = 12'h225 == _T_146[11:0] ? image_549 : _GEN_12903; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12905 = 12'h226 == _T_146[11:0] ? image_550 : _GEN_12904; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12906 = 12'h227 == _T_146[11:0] ? image_551 : _GEN_12905; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12907 = 12'h228 == _T_146[11:0] ? image_552 : _GEN_12906; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12908 = 12'h229 == _T_146[11:0] ? image_553 : _GEN_12907; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12909 = 12'h22a == _T_146[11:0] ? image_554 : _GEN_12908; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12910 = 12'h22b == _T_146[11:0] ? image_555 : _GEN_12909; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12911 = 12'h22c == _T_146[11:0] ? image_556 : _GEN_12910; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12912 = 12'h22d == _T_146[11:0] ? image_557 : _GEN_12911; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12913 = 12'h22e == _T_146[11:0] ? image_558 : _GEN_12912; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12914 = 12'h22f == _T_146[11:0] ? image_559 : _GEN_12913; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12915 = 12'h230 == _T_146[11:0] ? image_560 : _GEN_12914; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12916 = 12'h231 == _T_146[11:0] ? image_561 : _GEN_12915; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12917 = 12'h232 == _T_146[11:0] ? image_562 : _GEN_12916; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12918 = 12'h233 == _T_146[11:0] ? image_563 : _GEN_12917; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12919 = 12'h234 == _T_146[11:0] ? image_564 : _GEN_12918; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12920 = 12'h235 == _T_146[11:0] ? image_565 : _GEN_12919; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12921 = 12'h236 == _T_146[11:0] ? image_566 : _GEN_12920; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12922 = 12'h237 == _T_146[11:0] ? 4'h0 : _GEN_12921; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12923 = 12'h238 == _T_146[11:0] ? 4'h0 : _GEN_12922; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12924 = 12'h239 == _T_146[11:0] ? 4'h0 : _GEN_12923; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12925 = 12'h23a == _T_146[11:0] ? 4'h0 : _GEN_12924; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12926 = 12'h23b == _T_146[11:0] ? image_571 : _GEN_12925; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12927 = 12'h23c == _T_146[11:0] ? image_572 : _GEN_12926; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12928 = 12'h23d == _T_146[11:0] ? image_573 : _GEN_12927; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12929 = 12'h23e == _T_146[11:0] ? image_574 : _GEN_12928; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12930 = 12'h23f == _T_146[11:0] ? 4'h0 : _GEN_12929; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12931 = 12'h240 == _T_146[11:0] ? 4'h0 : _GEN_12930; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12932 = 12'h241 == _T_146[11:0] ? 4'h0 : _GEN_12931; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12933 = 12'h242 == _T_146[11:0] ? image_578 : _GEN_12932; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12934 = 12'h243 == _T_146[11:0] ? image_579 : _GEN_12933; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12935 = 12'h244 == _T_146[11:0] ? image_580 : _GEN_12934; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12936 = 12'h245 == _T_146[11:0] ? image_581 : _GEN_12935; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12937 = 12'h246 == _T_146[11:0] ? image_582 : _GEN_12936; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12938 = 12'h247 == _T_146[11:0] ? image_583 : _GEN_12937; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12939 = 12'h248 == _T_146[11:0] ? image_584 : _GEN_12938; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12940 = 12'h249 == _T_146[11:0] ? image_585 : _GEN_12939; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12941 = 12'h24a == _T_146[11:0] ? image_586 : _GEN_12940; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12942 = 12'h24b == _T_146[11:0] ? image_587 : _GEN_12941; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12943 = 12'h24c == _T_146[11:0] ? image_588 : _GEN_12942; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12944 = 12'h24d == _T_146[11:0] ? image_589 : _GEN_12943; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12945 = 12'h24e == _T_146[11:0] ? image_590 : _GEN_12944; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12946 = 12'h24f == _T_146[11:0] ? image_591 : _GEN_12945; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12947 = 12'h250 == _T_146[11:0] ? image_592 : _GEN_12946; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12948 = 12'h251 == _T_146[11:0] ? image_593 : _GEN_12947; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12949 = 12'h252 == _T_146[11:0] ? image_594 : _GEN_12948; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12950 = 12'h253 == _T_146[11:0] ? image_595 : _GEN_12949; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12951 = 12'h254 == _T_146[11:0] ? image_596 : _GEN_12950; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12952 = 12'h255 == _T_146[11:0] ? image_597 : _GEN_12951; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12953 = 12'h256 == _T_146[11:0] ? image_598 : _GEN_12952; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12954 = 12'h257 == _T_146[11:0] ? image_599 : _GEN_12953; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12955 = 12'h258 == _T_146[11:0] ? image_600 : _GEN_12954; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12956 = 12'h259 == _T_146[11:0] ? image_601 : _GEN_12955; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12957 = 12'h25a == _T_146[11:0] ? image_602 : _GEN_12956; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12958 = 12'h25b == _T_146[11:0] ? image_603 : _GEN_12957; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12959 = 12'h25c == _T_146[11:0] ? image_604 : _GEN_12958; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12960 = 12'h25d == _T_146[11:0] ? image_605 : _GEN_12959; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12961 = 12'h25e == _T_146[11:0] ? image_606 : _GEN_12960; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12962 = 12'h25f == _T_146[11:0] ? image_607 : _GEN_12961; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12963 = 12'h260 == _T_146[11:0] ? 4'h0 : _GEN_12962; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12964 = 12'h261 == _T_146[11:0] ? 4'h0 : _GEN_12963; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12965 = 12'h262 == _T_146[11:0] ? 4'h0 : _GEN_12964; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12966 = 12'h263 == _T_146[11:0] ? 4'h0 : _GEN_12965; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12967 = 12'h264 == _T_146[11:0] ? 4'h0 : _GEN_12966; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12968 = 12'h265 == _T_146[11:0] ? 4'h0 : _GEN_12967; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12969 = 12'h266 == _T_146[11:0] ? image_614 : _GEN_12968; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12970 = 12'h267 == _T_146[11:0] ? image_615 : _GEN_12969; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12971 = 12'h268 == _T_146[11:0] ? image_616 : _GEN_12970; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12972 = 12'h269 == _T_146[11:0] ? image_617 : _GEN_12971; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12973 = 12'h26a == _T_146[11:0] ? image_618 : _GEN_12972; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12974 = 12'h26b == _T_146[11:0] ? image_619 : _GEN_12973; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12975 = 12'h26c == _T_146[11:0] ? image_620 : _GEN_12974; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12976 = 12'h26d == _T_146[11:0] ? image_621 : _GEN_12975; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12977 = 12'h26e == _T_146[11:0] ? image_622 : _GEN_12976; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12978 = 12'h26f == _T_146[11:0] ? image_623 : _GEN_12977; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12979 = 12'h270 == _T_146[11:0] ? image_624 : _GEN_12978; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12980 = 12'h271 == _T_146[11:0] ? image_625 : _GEN_12979; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12981 = 12'h272 == _T_146[11:0] ? image_626 : _GEN_12980; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12982 = 12'h273 == _T_146[11:0] ? image_627 : _GEN_12981; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12983 = 12'h274 == _T_146[11:0] ? image_628 : _GEN_12982; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12984 = 12'h275 == _T_146[11:0] ? 4'h0 : _GEN_12983; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12985 = 12'h276 == _T_146[11:0] ? 4'h0 : _GEN_12984; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12986 = 12'h277 == _T_146[11:0] ? 4'h0 : _GEN_12985; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12987 = 12'h278 == _T_146[11:0] ? 4'h0 : _GEN_12986; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12988 = 12'h279 == _T_146[11:0] ? 4'h0 : _GEN_12987; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12989 = 12'h27a == _T_146[11:0] ? 4'h0 : _GEN_12988; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12990 = 12'h27b == _T_146[11:0] ? 4'h0 : _GEN_12989; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12991 = 12'h27c == _T_146[11:0] ? image_636 : _GEN_12990; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12992 = 12'h27d == _T_146[11:0] ? image_637 : _GEN_12991; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12993 = 12'h27e == _T_146[11:0] ? image_638 : _GEN_12992; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12994 = 12'h27f == _T_146[11:0] ? image_639 : _GEN_12993; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12995 = 12'h280 == _T_146[11:0] ? 4'h0 : _GEN_12994; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12996 = 12'h281 == _T_146[11:0] ? 4'h0 : _GEN_12995; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12997 = 12'h282 == _T_146[11:0] ? image_642 : _GEN_12996; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12998 = 12'h283 == _T_146[11:0] ? image_643 : _GEN_12997; // @[Filter.scala 138:46]
  wire [3:0] _GEN_12999 = 12'h284 == _T_146[11:0] ? image_644 : _GEN_12998; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13000 = 12'h285 == _T_146[11:0] ? image_645 : _GEN_12999; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13001 = 12'h286 == _T_146[11:0] ? image_646 : _GEN_13000; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13002 = 12'h287 == _T_146[11:0] ? image_647 : _GEN_13001; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13003 = 12'h288 == _T_146[11:0] ? image_648 : _GEN_13002; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13004 = 12'h289 == _T_146[11:0] ? image_649 : _GEN_13003; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13005 = 12'h28a == _T_146[11:0] ? image_650 : _GEN_13004; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13006 = 12'h28b == _T_146[11:0] ? image_651 : _GEN_13005; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13007 = 12'h28c == _T_146[11:0] ? image_652 : _GEN_13006; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13008 = 12'h28d == _T_146[11:0] ? image_653 : _GEN_13007; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13009 = 12'h28e == _T_146[11:0] ? image_654 : _GEN_13008; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13010 = 12'h28f == _T_146[11:0] ? image_655 : _GEN_13009; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13011 = 12'h290 == _T_146[11:0] ? image_656 : _GEN_13010; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13012 = 12'h291 == _T_146[11:0] ? image_657 : _GEN_13011; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13013 = 12'h292 == _T_146[11:0] ? image_658 : _GEN_13012; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13014 = 12'h293 == _T_146[11:0] ? image_659 : _GEN_13013; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13015 = 12'h294 == _T_146[11:0] ? image_660 : _GEN_13014; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13016 = 12'h295 == _T_146[11:0] ? image_661 : _GEN_13015; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13017 = 12'h296 == _T_146[11:0] ? image_662 : _GEN_13016; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13018 = 12'h297 == _T_146[11:0] ? image_663 : _GEN_13017; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13019 = 12'h298 == _T_146[11:0] ? image_664 : _GEN_13018; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13020 = 12'h299 == _T_146[11:0] ? image_665 : _GEN_13019; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13021 = 12'h29a == _T_146[11:0] ? image_666 : _GEN_13020; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13022 = 12'h29b == _T_146[11:0] ? image_667 : _GEN_13021; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13023 = 12'h29c == _T_146[11:0] ? image_668 : _GEN_13022; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13024 = 12'h29d == _T_146[11:0] ? image_669 : _GEN_13023; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13025 = 12'h29e == _T_146[11:0] ? image_670 : _GEN_13024; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13026 = 12'h29f == _T_146[11:0] ? 4'h0 : _GEN_13025; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13027 = 12'h2a0 == _T_146[11:0] ? 4'h0 : _GEN_13026; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13028 = 12'h2a1 == _T_146[11:0] ? 4'h0 : _GEN_13027; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13029 = 12'h2a2 == _T_146[11:0] ? 4'h0 : _GEN_13028; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13030 = 12'h2a3 == _T_146[11:0] ? 4'h0 : _GEN_13029; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13031 = 12'h2a4 == _T_146[11:0] ? 4'h0 : _GEN_13030; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13032 = 12'h2a5 == _T_146[11:0] ? 4'h0 : _GEN_13031; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13033 = 12'h2a6 == _T_146[11:0] ? 4'h0 : _GEN_13032; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13034 = 12'h2a7 == _T_146[11:0] ? image_679 : _GEN_13033; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13035 = 12'h2a8 == _T_146[11:0] ? image_680 : _GEN_13034; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13036 = 12'h2a9 == _T_146[11:0] ? image_681 : _GEN_13035; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13037 = 12'h2aa == _T_146[11:0] ? image_682 : _GEN_13036; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13038 = 12'h2ab == _T_146[11:0] ? image_683 : _GEN_13037; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13039 = 12'h2ac == _T_146[11:0] ? image_684 : _GEN_13038; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13040 = 12'h2ad == _T_146[11:0] ? image_685 : _GEN_13039; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13041 = 12'h2ae == _T_146[11:0] ? image_686 : _GEN_13040; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13042 = 12'h2af == _T_146[11:0] ? image_687 : _GEN_13041; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13043 = 12'h2b0 == _T_146[11:0] ? image_688 : _GEN_13042; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13044 = 12'h2b1 == _T_146[11:0] ? image_689 : _GEN_13043; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13045 = 12'h2b2 == _T_146[11:0] ? image_690 : _GEN_13044; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13046 = 12'h2b3 == _T_146[11:0] ? image_691 : _GEN_13045; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13047 = 12'h2b4 == _T_146[11:0] ? image_692 : _GEN_13046; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13048 = 12'h2b5 == _T_146[11:0] ? image_693 : _GEN_13047; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13049 = 12'h2b6 == _T_146[11:0] ? image_694 : _GEN_13048; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13050 = 12'h2b7 == _T_146[11:0] ? image_695 : _GEN_13049; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13051 = 12'h2b8 == _T_146[11:0] ? image_696 : _GEN_13050; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13052 = 12'h2b9 == _T_146[11:0] ? image_697 : _GEN_13051; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13053 = 12'h2ba == _T_146[11:0] ? image_698 : _GEN_13052; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13054 = 12'h2bb == _T_146[11:0] ? 4'h0 : _GEN_13053; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13055 = 12'h2bc == _T_146[11:0] ? 4'h0 : _GEN_13054; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13056 = 12'h2bd == _T_146[11:0] ? image_701 : _GEN_13055; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13057 = 12'h2be == _T_146[11:0] ? image_702 : _GEN_13056; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13058 = 12'h2bf == _T_146[11:0] ? image_703 : _GEN_13057; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13059 = 12'h2c0 == _T_146[11:0] ? 4'h0 : _GEN_13058; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13060 = 12'h2c1 == _T_146[11:0] ? image_705 : _GEN_13059; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13061 = 12'h2c2 == _T_146[11:0] ? image_706 : _GEN_13060; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13062 = 12'h2c3 == _T_146[11:0] ? image_707 : _GEN_13061; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13063 = 12'h2c4 == _T_146[11:0] ? image_708 : _GEN_13062; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13064 = 12'h2c5 == _T_146[11:0] ? image_709 : _GEN_13063; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13065 = 12'h2c6 == _T_146[11:0] ? image_710 : _GEN_13064; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13066 = 12'h2c7 == _T_146[11:0] ? image_711 : _GEN_13065; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13067 = 12'h2c8 == _T_146[11:0] ? image_712 : _GEN_13066; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13068 = 12'h2c9 == _T_146[11:0] ? image_713 : _GEN_13067; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13069 = 12'h2ca == _T_146[11:0] ? image_714 : _GEN_13068; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13070 = 12'h2cb == _T_146[11:0] ? image_715 : _GEN_13069; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13071 = 12'h2cc == _T_146[11:0] ? image_716 : _GEN_13070; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13072 = 12'h2cd == _T_146[11:0] ? image_717 : _GEN_13071; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13073 = 12'h2ce == _T_146[11:0] ? image_718 : _GEN_13072; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13074 = 12'h2cf == _T_146[11:0] ? image_719 : _GEN_13073; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13075 = 12'h2d0 == _T_146[11:0] ? image_720 : _GEN_13074; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13076 = 12'h2d1 == _T_146[11:0] ? image_721 : _GEN_13075; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13077 = 12'h2d2 == _T_146[11:0] ? image_722 : _GEN_13076; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13078 = 12'h2d3 == _T_146[11:0] ? image_723 : _GEN_13077; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13079 = 12'h2d4 == _T_146[11:0] ? image_724 : _GEN_13078; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13080 = 12'h2d5 == _T_146[11:0] ? image_725 : _GEN_13079; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13081 = 12'h2d6 == _T_146[11:0] ? image_726 : _GEN_13080; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13082 = 12'h2d7 == _T_146[11:0] ? image_727 : _GEN_13081; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13083 = 12'h2d8 == _T_146[11:0] ? image_728 : _GEN_13082; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13084 = 12'h2d9 == _T_146[11:0] ? image_729 : _GEN_13083; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13085 = 12'h2da == _T_146[11:0] ? image_730 : _GEN_13084; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13086 = 12'h2db == _T_146[11:0] ? image_731 : _GEN_13085; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13087 = 12'h2dc == _T_146[11:0] ? image_732 : _GEN_13086; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13088 = 12'h2dd == _T_146[11:0] ? image_733 : _GEN_13087; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13089 = 12'h2de == _T_146[11:0] ? image_734 : _GEN_13088; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13090 = 12'h2df == _T_146[11:0] ? 4'h0 : _GEN_13089; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13091 = 12'h2e0 == _T_146[11:0] ? image_736 : _GEN_13090; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13092 = 12'h2e1 == _T_146[11:0] ? image_737 : _GEN_13091; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13093 = 12'h2e2 == _T_146[11:0] ? 4'h0 : _GEN_13092; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13094 = 12'h2e3 == _T_146[11:0] ? image_739 : _GEN_13093; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13095 = 12'h2e4 == _T_146[11:0] ? image_740 : _GEN_13094; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13096 = 12'h2e5 == _T_146[11:0] ? image_741 : _GEN_13095; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13097 = 12'h2e6 == _T_146[11:0] ? 4'h0 : _GEN_13096; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13098 = 12'h2e7 == _T_146[11:0] ? 4'h0 : _GEN_13097; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13099 = 12'h2e8 == _T_146[11:0] ? image_744 : _GEN_13098; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13100 = 12'h2e9 == _T_146[11:0] ? image_745 : _GEN_13099; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13101 = 12'h2ea == _T_146[11:0] ? image_746 : _GEN_13100; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13102 = 12'h2eb == _T_146[11:0] ? image_747 : _GEN_13101; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13103 = 12'h2ec == _T_146[11:0] ? image_748 : _GEN_13102; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13104 = 12'h2ed == _T_146[11:0] ? image_749 : _GEN_13103; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13105 = 12'h2ee == _T_146[11:0] ? image_750 : _GEN_13104; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13106 = 12'h2ef == _T_146[11:0] ? image_751 : _GEN_13105; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13107 = 12'h2f0 == _T_146[11:0] ? image_752 : _GEN_13106; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13108 = 12'h2f1 == _T_146[11:0] ? image_753 : _GEN_13107; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13109 = 12'h2f2 == _T_146[11:0] ? image_754 : _GEN_13108; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13110 = 12'h2f3 == _T_146[11:0] ? image_755 : _GEN_13109; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13111 = 12'h2f4 == _T_146[11:0] ? image_756 : _GEN_13110; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13112 = 12'h2f5 == _T_146[11:0] ? 4'h0 : _GEN_13111; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13113 = 12'h2f6 == _T_146[11:0] ? image_758 : _GEN_13112; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13114 = 12'h2f7 == _T_146[11:0] ? 4'h0 : _GEN_13113; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13115 = 12'h2f8 == _T_146[11:0] ? image_760 : _GEN_13114; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13116 = 12'h2f9 == _T_146[11:0] ? image_761 : _GEN_13115; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13117 = 12'h2fa == _T_146[11:0] ? image_762 : _GEN_13116; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13118 = 12'h2fb == _T_146[11:0] ? image_763 : _GEN_13117; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13119 = 12'h2fc == _T_146[11:0] ? 4'h0 : _GEN_13118; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13120 = 12'h2fd == _T_146[11:0] ? image_765 : _GEN_13119; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13121 = 12'h2fe == _T_146[11:0] ? image_766 : _GEN_13120; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13122 = 12'h2ff == _T_146[11:0] ? image_767 : _GEN_13121; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13123 = 12'h300 == _T_146[11:0] ? image_768 : _GEN_13122; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13124 = 12'h301 == _T_146[11:0] ? image_769 : _GEN_13123; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13125 = 12'h302 == _T_146[11:0] ? image_770 : _GEN_13124; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13126 = 12'h303 == _T_146[11:0] ? image_771 : _GEN_13125; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13127 = 12'h304 == _T_146[11:0] ? image_772 : _GEN_13126; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13128 = 12'h305 == _T_146[11:0] ? image_773 : _GEN_13127; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13129 = 12'h306 == _T_146[11:0] ? image_774 : _GEN_13128; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13130 = 12'h307 == _T_146[11:0] ? image_775 : _GEN_13129; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13131 = 12'h308 == _T_146[11:0] ? image_776 : _GEN_13130; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13132 = 12'h309 == _T_146[11:0] ? image_777 : _GEN_13131; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13133 = 12'h30a == _T_146[11:0] ? image_778 : _GEN_13132; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13134 = 12'h30b == _T_146[11:0] ? image_779 : _GEN_13133; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13135 = 12'h30c == _T_146[11:0] ? image_780 : _GEN_13134; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13136 = 12'h30d == _T_146[11:0] ? image_781 : _GEN_13135; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13137 = 12'h30e == _T_146[11:0] ? image_782 : _GEN_13136; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13138 = 12'h30f == _T_146[11:0] ? image_783 : _GEN_13137; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13139 = 12'h310 == _T_146[11:0] ? image_784 : _GEN_13138; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13140 = 12'h311 == _T_146[11:0] ? image_785 : _GEN_13139; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13141 = 12'h312 == _T_146[11:0] ? image_786 : _GEN_13140; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13142 = 12'h313 == _T_146[11:0] ? image_787 : _GEN_13141; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13143 = 12'h314 == _T_146[11:0] ? image_788 : _GEN_13142; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13144 = 12'h315 == _T_146[11:0] ? image_789 : _GEN_13143; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13145 = 12'h316 == _T_146[11:0] ? image_790 : _GEN_13144; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13146 = 12'h317 == _T_146[11:0] ? image_791 : _GEN_13145; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13147 = 12'h318 == _T_146[11:0] ? image_792 : _GEN_13146; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13148 = 12'h319 == _T_146[11:0] ? image_793 : _GEN_13147; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13149 = 12'h31a == _T_146[11:0] ? image_794 : _GEN_13148; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13150 = 12'h31b == _T_146[11:0] ? image_795 : _GEN_13149; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13151 = 12'h31c == _T_146[11:0] ? image_796 : _GEN_13150; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13152 = 12'h31d == _T_146[11:0] ? image_797 : _GEN_13151; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13153 = 12'h31e == _T_146[11:0] ? 4'h0 : _GEN_13152; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13154 = 12'h31f == _T_146[11:0] ? 4'h0 : _GEN_13153; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13155 = 12'h320 == _T_146[11:0] ? image_800 : _GEN_13154; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13156 = 12'h321 == _T_146[11:0] ? image_801 : _GEN_13155; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13157 = 12'h322 == _T_146[11:0] ? image_802 : _GEN_13156; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13158 = 12'h323 == _T_146[11:0] ? image_803 : _GEN_13157; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13159 = 12'h324 == _T_146[11:0] ? image_804 : _GEN_13158; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13160 = 12'h325 == _T_146[11:0] ? image_805 : _GEN_13159; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13161 = 12'h326 == _T_146[11:0] ? image_806 : _GEN_13160; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13162 = 12'h327 == _T_146[11:0] ? 4'h0 : _GEN_13161; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13163 = 12'h328 == _T_146[11:0] ? image_808 : _GEN_13162; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13164 = 12'h329 == _T_146[11:0] ? image_809 : _GEN_13163; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13165 = 12'h32a == _T_146[11:0] ? image_810 : _GEN_13164; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13166 = 12'h32b == _T_146[11:0] ? image_811 : _GEN_13165; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13167 = 12'h32c == _T_146[11:0] ? image_812 : _GEN_13166; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13168 = 12'h32d == _T_146[11:0] ? image_813 : _GEN_13167; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13169 = 12'h32e == _T_146[11:0] ? image_814 : _GEN_13168; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13170 = 12'h32f == _T_146[11:0] ? image_815 : _GEN_13169; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13171 = 12'h330 == _T_146[11:0] ? image_816 : _GEN_13170; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13172 = 12'h331 == _T_146[11:0] ? image_817 : _GEN_13171; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13173 = 12'h332 == _T_146[11:0] ? image_818 : _GEN_13172; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13174 = 12'h333 == _T_146[11:0] ? image_819 : _GEN_13173; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13175 = 12'h334 == _T_146[11:0] ? image_820 : _GEN_13174; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13176 = 12'h335 == _T_146[11:0] ? 4'h0 : _GEN_13175; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13177 = 12'h336 == _T_146[11:0] ? image_822 : _GEN_13176; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13178 = 12'h337 == _T_146[11:0] ? image_823 : _GEN_13177; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13179 = 12'h338 == _T_146[11:0] ? image_824 : _GEN_13178; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13180 = 12'h339 == _T_146[11:0] ? image_825 : _GEN_13179; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13181 = 12'h33a == _T_146[11:0] ? image_826 : _GEN_13180; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13182 = 12'h33b == _T_146[11:0] ? 4'h0 : _GEN_13181; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13183 = 12'h33c == _T_146[11:0] ? image_828 : _GEN_13182; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13184 = 12'h33d == _T_146[11:0] ? image_829 : _GEN_13183; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13185 = 12'h33e == _T_146[11:0] ? image_830 : _GEN_13184; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13186 = 12'h33f == _T_146[11:0] ? image_831 : _GEN_13185; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13187 = 12'h340 == _T_146[11:0] ? 4'h0 : _GEN_13186; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13188 = 12'h341 == _T_146[11:0] ? image_833 : _GEN_13187; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13189 = 12'h342 == _T_146[11:0] ? image_834 : _GEN_13188; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13190 = 12'h343 == _T_146[11:0] ? image_835 : _GEN_13189; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13191 = 12'h344 == _T_146[11:0] ? image_836 : _GEN_13190; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13192 = 12'h345 == _T_146[11:0] ? image_837 : _GEN_13191; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13193 = 12'h346 == _T_146[11:0] ? image_838 : _GEN_13192; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13194 = 12'h347 == _T_146[11:0] ? image_839 : _GEN_13193; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13195 = 12'h348 == _T_146[11:0] ? image_840 : _GEN_13194; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13196 = 12'h349 == _T_146[11:0] ? image_841 : _GEN_13195; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13197 = 12'h34a == _T_146[11:0] ? image_842 : _GEN_13196; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13198 = 12'h34b == _T_146[11:0] ? image_843 : _GEN_13197; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13199 = 12'h34c == _T_146[11:0] ? image_844 : _GEN_13198; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13200 = 12'h34d == _T_146[11:0] ? image_845 : _GEN_13199; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13201 = 12'h34e == _T_146[11:0] ? image_846 : _GEN_13200; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13202 = 12'h34f == _T_146[11:0] ? image_847 : _GEN_13201; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13203 = 12'h350 == _T_146[11:0] ? image_848 : _GEN_13202; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13204 = 12'h351 == _T_146[11:0] ? image_849 : _GEN_13203; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13205 = 12'h352 == _T_146[11:0] ? image_850 : _GEN_13204; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13206 = 12'h353 == _T_146[11:0] ? image_851 : _GEN_13205; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13207 = 12'h354 == _T_146[11:0] ? image_852 : _GEN_13206; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13208 = 12'h355 == _T_146[11:0] ? image_853 : _GEN_13207; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13209 = 12'h356 == _T_146[11:0] ? image_854 : _GEN_13208; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13210 = 12'h357 == _T_146[11:0] ? image_855 : _GEN_13209; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13211 = 12'h358 == _T_146[11:0] ? image_856 : _GEN_13210; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13212 = 12'h359 == _T_146[11:0] ? image_857 : _GEN_13211; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13213 = 12'h35a == _T_146[11:0] ? image_858 : _GEN_13212; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13214 = 12'h35b == _T_146[11:0] ? image_859 : _GEN_13213; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13215 = 12'h35c == _T_146[11:0] ? image_860 : _GEN_13214; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13216 = 12'h35d == _T_146[11:0] ? image_861 : _GEN_13215; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13217 = 12'h35e == _T_146[11:0] ? image_862 : _GEN_13216; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13218 = 12'h35f == _T_146[11:0] ? 4'h0 : _GEN_13217; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13219 = 12'h360 == _T_146[11:0] ? 4'h0 : _GEN_13218; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13220 = 12'h361 == _T_146[11:0] ? image_865 : _GEN_13219; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13221 = 12'h362 == _T_146[11:0] ? image_866 : _GEN_13220; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13222 = 12'h363 == _T_146[11:0] ? image_867 : _GEN_13221; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13223 = 12'h364 == _T_146[11:0] ? image_868 : _GEN_13222; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13224 = 12'h365 == _T_146[11:0] ? image_869 : _GEN_13223; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13225 = 12'h366 == _T_146[11:0] ? 4'h0 : _GEN_13224; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13226 = 12'h367 == _T_146[11:0] ? 4'h0 : _GEN_13225; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13227 = 12'h368 == _T_146[11:0] ? image_872 : _GEN_13226; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13228 = 12'h369 == _T_146[11:0] ? image_873 : _GEN_13227; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13229 = 12'h36a == _T_146[11:0] ? image_874 : _GEN_13228; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13230 = 12'h36b == _T_146[11:0] ? image_875 : _GEN_13229; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13231 = 12'h36c == _T_146[11:0] ? image_876 : _GEN_13230; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13232 = 12'h36d == _T_146[11:0] ? image_877 : _GEN_13231; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13233 = 12'h36e == _T_146[11:0] ? image_878 : _GEN_13232; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13234 = 12'h36f == _T_146[11:0] ? image_879 : _GEN_13233; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13235 = 12'h370 == _T_146[11:0] ? image_880 : _GEN_13234; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13236 = 12'h371 == _T_146[11:0] ? image_881 : _GEN_13235; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13237 = 12'h372 == _T_146[11:0] ? image_882 : _GEN_13236; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13238 = 12'h373 == _T_146[11:0] ? image_883 : _GEN_13237; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13239 = 12'h374 == _T_146[11:0] ? image_884 : _GEN_13238; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13240 = 12'h375 == _T_146[11:0] ? image_885 : _GEN_13239; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13241 = 12'h376 == _T_146[11:0] ? 4'h0 : _GEN_13240; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13242 = 12'h377 == _T_146[11:0] ? 4'h0 : _GEN_13241; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13243 = 12'h378 == _T_146[11:0] ? 4'h0 : _GEN_13242; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13244 = 12'h379 == _T_146[11:0] ? 4'h0 : _GEN_13243; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13245 = 12'h37a == _T_146[11:0] ? 4'h0 : _GEN_13244; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13246 = 12'h37b == _T_146[11:0] ? image_891 : _GEN_13245; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13247 = 12'h37c == _T_146[11:0] ? image_892 : _GEN_13246; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13248 = 12'h37d == _T_146[11:0] ? image_893 : _GEN_13247; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13249 = 12'h37e == _T_146[11:0] ? image_894 : _GEN_13248; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13250 = 12'h37f == _T_146[11:0] ? image_895 : _GEN_13249; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13251 = 12'h380 == _T_146[11:0] ? 4'h0 : _GEN_13250; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13252 = 12'h381 == _T_146[11:0] ? image_897 : _GEN_13251; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13253 = 12'h382 == _T_146[11:0] ? image_898 : _GEN_13252; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13254 = 12'h383 == _T_146[11:0] ? image_899 : _GEN_13253; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13255 = 12'h384 == _T_146[11:0] ? image_900 : _GEN_13254; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13256 = 12'h385 == _T_146[11:0] ? image_901 : _GEN_13255; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13257 = 12'h386 == _T_146[11:0] ? image_902 : _GEN_13256; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13258 = 12'h387 == _T_146[11:0] ? image_903 : _GEN_13257; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13259 = 12'h388 == _T_146[11:0] ? image_904 : _GEN_13258; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13260 = 12'h389 == _T_146[11:0] ? image_905 : _GEN_13259; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13261 = 12'h38a == _T_146[11:0] ? image_906 : _GEN_13260; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13262 = 12'h38b == _T_146[11:0] ? image_907 : _GEN_13261; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13263 = 12'h38c == _T_146[11:0] ? image_908 : _GEN_13262; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13264 = 12'h38d == _T_146[11:0] ? image_909 : _GEN_13263; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13265 = 12'h38e == _T_146[11:0] ? image_910 : _GEN_13264; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13266 = 12'h38f == _T_146[11:0] ? image_911 : _GEN_13265; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13267 = 12'h390 == _T_146[11:0] ? image_912 : _GEN_13266; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13268 = 12'h391 == _T_146[11:0] ? image_913 : _GEN_13267; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13269 = 12'h392 == _T_146[11:0] ? image_914 : _GEN_13268; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13270 = 12'h393 == _T_146[11:0] ? image_915 : _GEN_13269; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13271 = 12'h394 == _T_146[11:0] ? image_916 : _GEN_13270; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13272 = 12'h395 == _T_146[11:0] ? image_917 : _GEN_13271; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13273 = 12'h396 == _T_146[11:0] ? image_918 : _GEN_13272; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13274 = 12'h397 == _T_146[11:0] ? image_919 : _GEN_13273; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13275 = 12'h398 == _T_146[11:0] ? image_920 : _GEN_13274; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13276 = 12'h399 == _T_146[11:0] ? image_921 : _GEN_13275; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13277 = 12'h39a == _T_146[11:0] ? image_922 : _GEN_13276; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13278 = 12'h39b == _T_146[11:0] ? image_923 : _GEN_13277; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13279 = 12'h39c == _T_146[11:0] ? image_924 : _GEN_13278; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13280 = 12'h39d == _T_146[11:0] ? image_925 : _GEN_13279; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13281 = 12'h39e == _T_146[11:0] ? image_926 : _GEN_13280; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13282 = 12'h39f == _T_146[11:0] ? image_927 : _GEN_13281; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13283 = 12'h3a0 == _T_146[11:0] ? 4'h0 : _GEN_13282; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13284 = 12'h3a1 == _T_146[11:0] ? image_929 : _GEN_13283; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13285 = 12'h3a2 == _T_146[11:0] ? image_930 : _GEN_13284; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13286 = 12'h3a3 == _T_146[11:0] ? 4'h0 : _GEN_13285; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13287 = 12'h3a4 == _T_146[11:0] ? 4'h0 : _GEN_13286; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13288 = 12'h3a5 == _T_146[11:0] ? 4'h0 : _GEN_13287; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13289 = 12'h3a6 == _T_146[11:0] ? 4'h0 : _GEN_13288; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13290 = 12'h3a7 == _T_146[11:0] ? image_935 : _GEN_13289; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13291 = 12'h3a8 == _T_146[11:0] ? image_936 : _GEN_13290; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13292 = 12'h3a9 == _T_146[11:0] ? image_937 : _GEN_13291; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13293 = 12'h3aa == _T_146[11:0] ? image_938 : _GEN_13292; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13294 = 12'h3ab == _T_146[11:0] ? image_939 : _GEN_13293; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13295 = 12'h3ac == _T_146[11:0] ? image_940 : _GEN_13294; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13296 = 12'h3ad == _T_146[11:0] ? image_941 : _GEN_13295; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13297 = 12'h3ae == _T_146[11:0] ? image_942 : _GEN_13296; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13298 = 12'h3af == _T_146[11:0] ? image_943 : _GEN_13297; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13299 = 12'h3b0 == _T_146[11:0] ? image_944 : _GEN_13298; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13300 = 12'h3b1 == _T_146[11:0] ? image_945 : _GEN_13299; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13301 = 12'h3b2 == _T_146[11:0] ? image_946 : _GEN_13300; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13302 = 12'h3b3 == _T_146[11:0] ? image_947 : _GEN_13301; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13303 = 12'h3b4 == _T_146[11:0] ? image_948 : _GEN_13302; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13304 = 12'h3b5 == _T_146[11:0] ? image_949 : _GEN_13303; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13305 = 12'h3b6 == _T_146[11:0] ? image_950 : _GEN_13304; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13306 = 12'h3b7 == _T_146[11:0] ? image_951 : _GEN_13305; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13307 = 12'h3b8 == _T_146[11:0] ? image_952 : _GEN_13306; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13308 = 12'h3b9 == _T_146[11:0] ? image_953 : _GEN_13307; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13309 = 12'h3ba == _T_146[11:0] ? image_954 : _GEN_13308; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13310 = 12'h3bb == _T_146[11:0] ? image_955 : _GEN_13309; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13311 = 12'h3bc == _T_146[11:0] ? image_956 : _GEN_13310; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13312 = 12'h3bd == _T_146[11:0] ? image_957 : _GEN_13311; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13313 = 12'h3be == _T_146[11:0] ? image_958 : _GEN_13312; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13314 = 12'h3bf == _T_146[11:0] ? image_959 : _GEN_13313; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13315 = 12'h3c0 == _T_146[11:0] ? 4'h0 : _GEN_13314; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13316 = 12'h3c1 == _T_146[11:0] ? image_961 : _GEN_13315; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13317 = 12'h3c2 == _T_146[11:0] ? image_962 : _GEN_13316; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13318 = 12'h3c3 == _T_146[11:0] ? image_963 : _GEN_13317; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13319 = 12'h3c4 == _T_146[11:0] ? image_964 : _GEN_13318; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13320 = 12'h3c5 == _T_146[11:0] ? image_965 : _GEN_13319; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13321 = 12'h3c6 == _T_146[11:0] ? image_966 : _GEN_13320; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13322 = 12'h3c7 == _T_146[11:0] ? image_967 : _GEN_13321; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13323 = 12'h3c8 == _T_146[11:0] ? image_968 : _GEN_13322; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13324 = 12'h3c9 == _T_146[11:0] ? image_969 : _GEN_13323; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13325 = 12'h3ca == _T_146[11:0] ? image_970 : _GEN_13324; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13326 = 12'h3cb == _T_146[11:0] ? image_971 : _GEN_13325; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13327 = 12'h3cc == _T_146[11:0] ? image_972 : _GEN_13326; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13328 = 12'h3cd == _T_146[11:0] ? image_973 : _GEN_13327; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13329 = 12'h3ce == _T_146[11:0] ? image_974 : _GEN_13328; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13330 = 12'h3cf == _T_146[11:0] ? image_975 : _GEN_13329; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13331 = 12'h3d0 == _T_146[11:0] ? image_976 : _GEN_13330; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13332 = 12'h3d1 == _T_146[11:0] ? image_977 : _GEN_13331; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13333 = 12'h3d2 == _T_146[11:0] ? image_978 : _GEN_13332; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13334 = 12'h3d3 == _T_146[11:0] ? image_979 : _GEN_13333; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13335 = 12'h3d4 == _T_146[11:0] ? image_980 : _GEN_13334; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13336 = 12'h3d5 == _T_146[11:0] ? image_981 : _GEN_13335; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13337 = 12'h3d6 == _T_146[11:0] ? image_982 : _GEN_13336; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13338 = 12'h3d7 == _T_146[11:0] ? image_983 : _GEN_13337; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13339 = 12'h3d8 == _T_146[11:0] ? image_984 : _GEN_13338; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13340 = 12'h3d9 == _T_146[11:0] ? image_985 : _GEN_13339; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13341 = 12'h3da == _T_146[11:0] ? image_986 : _GEN_13340; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13342 = 12'h3db == _T_146[11:0] ? image_987 : _GEN_13341; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13343 = 12'h3dc == _T_146[11:0] ? image_988 : _GEN_13342; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13344 = 12'h3dd == _T_146[11:0] ? image_989 : _GEN_13343; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13345 = 12'h3de == _T_146[11:0] ? image_990 : _GEN_13344; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13346 = 12'h3df == _T_146[11:0] ? image_991 : _GEN_13345; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13347 = 12'h3e0 == _T_146[11:0] ? image_992 : _GEN_13346; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13348 = 12'h3e1 == _T_146[11:0] ? 4'h0 : _GEN_13347; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13349 = 12'h3e2 == _T_146[11:0] ? 4'h0 : _GEN_13348; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13350 = 12'h3e3 == _T_146[11:0] ? 4'h0 : _GEN_13349; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13351 = 12'h3e4 == _T_146[11:0] ? 4'h0 : _GEN_13350; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13352 = 12'h3e5 == _T_146[11:0] ? image_997 : _GEN_13351; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13353 = 12'h3e6 == _T_146[11:0] ? image_998 : _GEN_13352; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13354 = 12'h3e7 == _T_146[11:0] ? image_999 : _GEN_13353; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13355 = 12'h3e8 == _T_146[11:0] ? image_1000 : _GEN_13354; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13356 = 12'h3e9 == _T_146[11:0] ? image_1001 : _GEN_13355; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13357 = 12'h3ea == _T_146[11:0] ? image_1002 : _GEN_13356; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13358 = 12'h3eb == _T_146[11:0] ? image_1003 : _GEN_13357; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13359 = 12'h3ec == _T_146[11:0] ? image_1004 : _GEN_13358; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13360 = 12'h3ed == _T_146[11:0] ? image_1005 : _GEN_13359; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13361 = 12'h3ee == _T_146[11:0] ? image_1006 : _GEN_13360; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13362 = 12'h3ef == _T_146[11:0] ? image_1007 : _GEN_13361; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13363 = 12'h3f0 == _T_146[11:0] ? image_1008 : _GEN_13362; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13364 = 12'h3f1 == _T_146[11:0] ? image_1009 : _GEN_13363; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13365 = 12'h3f2 == _T_146[11:0] ? image_1010 : _GEN_13364; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13366 = 12'h3f3 == _T_146[11:0] ? image_1011 : _GEN_13365; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13367 = 12'h3f4 == _T_146[11:0] ? image_1012 : _GEN_13366; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13368 = 12'h3f5 == _T_146[11:0] ? image_1013 : _GEN_13367; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13369 = 12'h3f6 == _T_146[11:0] ? image_1014 : _GEN_13368; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13370 = 12'h3f7 == _T_146[11:0] ? image_1015 : _GEN_13369; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13371 = 12'h3f8 == _T_146[11:0] ? image_1016 : _GEN_13370; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13372 = 12'h3f9 == _T_146[11:0] ? image_1017 : _GEN_13371; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13373 = 12'h3fa == _T_146[11:0] ? image_1018 : _GEN_13372; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13374 = 12'h3fb == _T_146[11:0] ? image_1019 : _GEN_13373; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13375 = 12'h3fc == _T_146[11:0] ? image_1020 : _GEN_13374; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13376 = 12'h3fd == _T_146[11:0] ? 4'h0 : _GEN_13375; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13377 = 12'h3fe == _T_146[11:0] ? 4'h0 : _GEN_13376; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13378 = 12'h3ff == _T_146[11:0] ? 4'h0 : _GEN_13377; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13379 = 12'h400 == _T_146[11:0] ? image_1024 : _GEN_13378; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13380 = 12'h401 == _T_146[11:0] ? image_1025 : _GEN_13379; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13381 = 12'h402 == _T_146[11:0] ? image_1026 : _GEN_13380; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13382 = 12'h403 == _T_146[11:0] ? image_1027 : _GEN_13381; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13383 = 12'h404 == _T_146[11:0] ? image_1028 : _GEN_13382; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13384 = 12'h405 == _T_146[11:0] ? image_1029 : _GEN_13383; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13385 = 12'h406 == _T_146[11:0] ? image_1030 : _GEN_13384; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13386 = 12'h407 == _T_146[11:0] ? image_1031 : _GEN_13385; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13387 = 12'h408 == _T_146[11:0] ? image_1032 : _GEN_13386; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13388 = 12'h409 == _T_146[11:0] ? image_1033 : _GEN_13387; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13389 = 12'h40a == _T_146[11:0] ? image_1034 : _GEN_13388; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13390 = 12'h40b == _T_146[11:0] ? image_1035 : _GEN_13389; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13391 = 12'h40c == _T_146[11:0] ? image_1036 : _GEN_13390; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13392 = 12'h40d == _T_146[11:0] ? image_1037 : _GEN_13391; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13393 = 12'h40e == _T_146[11:0] ? image_1038 : _GEN_13392; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13394 = 12'h40f == _T_146[11:0] ? image_1039 : _GEN_13393; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13395 = 12'h410 == _T_146[11:0] ? image_1040 : _GEN_13394; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13396 = 12'h411 == _T_146[11:0] ? image_1041 : _GEN_13395; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13397 = 12'h412 == _T_146[11:0] ? image_1042 : _GEN_13396; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13398 = 12'h413 == _T_146[11:0] ? image_1043 : _GEN_13397; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13399 = 12'h414 == _T_146[11:0] ? image_1044 : _GEN_13398; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13400 = 12'h415 == _T_146[11:0] ? image_1045 : _GEN_13399; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13401 = 12'h416 == _T_146[11:0] ? image_1046 : _GEN_13400; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13402 = 12'h417 == _T_146[11:0] ? image_1047 : _GEN_13401; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13403 = 12'h418 == _T_146[11:0] ? image_1048 : _GEN_13402; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13404 = 12'h419 == _T_146[11:0] ? image_1049 : _GEN_13403; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13405 = 12'h41a == _T_146[11:0] ? image_1050 : _GEN_13404; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13406 = 12'h41b == _T_146[11:0] ? image_1051 : _GEN_13405; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13407 = 12'h41c == _T_146[11:0] ? image_1052 : _GEN_13406; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13408 = 12'h41d == _T_146[11:0] ? image_1053 : _GEN_13407; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13409 = 12'h41e == _T_146[11:0] ? image_1054 : _GEN_13408; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13410 = 12'h41f == _T_146[11:0] ? image_1055 : _GEN_13409; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13411 = 12'h420 == _T_146[11:0] ? image_1056 : _GEN_13410; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13412 = 12'h421 == _T_146[11:0] ? image_1057 : _GEN_13411; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13413 = 12'h422 == _T_146[11:0] ? image_1058 : _GEN_13412; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13414 = 12'h423 == _T_146[11:0] ? image_1059 : _GEN_13413; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13415 = 12'h424 == _T_146[11:0] ? image_1060 : _GEN_13414; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13416 = 12'h425 == _T_146[11:0] ? image_1061 : _GEN_13415; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13417 = 12'h426 == _T_146[11:0] ? image_1062 : _GEN_13416; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13418 = 12'h427 == _T_146[11:0] ? image_1063 : _GEN_13417; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13419 = 12'h428 == _T_146[11:0] ? image_1064 : _GEN_13418; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13420 = 12'h429 == _T_146[11:0] ? image_1065 : _GEN_13419; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13421 = 12'h42a == _T_146[11:0] ? image_1066 : _GEN_13420; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13422 = 12'h42b == _T_146[11:0] ? image_1067 : _GEN_13421; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13423 = 12'h42c == _T_146[11:0] ? image_1068 : _GEN_13422; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13424 = 12'h42d == _T_146[11:0] ? image_1069 : _GEN_13423; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13425 = 12'h42e == _T_146[11:0] ? image_1070 : _GEN_13424; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13426 = 12'h42f == _T_146[11:0] ? image_1071 : _GEN_13425; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13427 = 12'h430 == _T_146[11:0] ? image_1072 : _GEN_13426; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13428 = 12'h431 == _T_146[11:0] ? image_1073 : _GEN_13427; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13429 = 12'h432 == _T_146[11:0] ? image_1074 : _GEN_13428; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13430 = 12'h433 == _T_146[11:0] ? image_1075 : _GEN_13429; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13431 = 12'h434 == _T_146[11:0] ? image_1076 : _GEN_13430; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13432 = 12'h435 == _T_146[11:0] ? image_1077 : _GEN_13431; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13433 = 12'h436 == _T_146[11:0] ? image_1078 : _GEN_13432; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13434 = 12'h437 == _T_146[11:0] ? image_1079 : _GEN_13433; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13435 = 12'h438 == _T_146[11:0] ? image_1080 : _GEN_13434; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13436 = 12'h439 == _T_146[11:0] ? image_1081 : _GEN_13435; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13437 = 12'h43a == _T_146[11:0] ? image_1082 : _GEN_13436; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13438 = 12'h43b == _T_146[11:0] ? image_1083 : _GEN_13437; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13439 = 12'h43c == _T_146[11:0] ? image_1084 : _GEN_13438; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13440 = 12'h43d == _T_146[11:0] ? image_1085 : _GEN_13439; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13441 = 12'h43e == _T_146[11:0] ? 4'h0 : _GEN_13440; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13442 = 12'h43f == _T_146[11:0] ? 4'h0 : _GEN_13441; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13443 = 12'h440 == _T_146[11:0] ? image_1088 : _GEN_13442; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13444 = 12'h441 == _T_146[11:0] ? image_1089 : _GEN_13443; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13445 = 12'h442 == _T_146[11:0] ? image_1090 : _GEN_13444; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13446 = 12'h443 == _T_146[11:0] ? image_1091 : _GEN_13445; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13447 = 12'h444 == _T_146[11:0] ? image_1092 : _GEN_13446; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13448 = 12'h445 == _T_146[11:0] ? image_1093 : _GEN_13447; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13449 = 12'h446 == _T_146[11:0] ? image_1094 : _GEN_13448; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13450 = 12'h447 == _T_146[11:0] ? image_1095 : _GEN_13449; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13451 = 12'h448 == _T_146[11:0] ? image_1096 : _GEN_13450; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13452 = 12'h449 == _T_146[11:0] ? image_1097 : _GEN_13451; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13453 = 12'h44a == _T_146[11:0] ? image_1098 : _GEN_13452; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13454 = 12'h44b == _T_146[11:0] ? image_1099 : _GEN_13453; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13455 = 12'h44c == _T_146[11:0] ? image_1100 : _GEN_13454; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13456 = 12'h44d == _T_146[11:0] ? image_1101 : _GEN_13455; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13457 = 12'h44e == _T_146[11:0] ? image_1102 : _GEN_13456; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13458 = 12'h44f == _T_146[11:0] ? image_1103 : _GEN_13457; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13459 = 12'h450 == _T_146[11:0] ? image_1104 : _GEN_13458; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13460 = 12'h451 == _T_146[11:0] ? image_1105 : _GEN_13459; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13461 = 12'h452 == _T_146[11:0] ? image_1106 : _GEN_13460; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13462 = 12'h453 == _T_146[11:0] ? image_1107 : _GEN_13461; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13463 = 12'h454 == _T_146[11:0] ? image_1108 : _GEN_13462; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13464 = 12'h455 == _T_146[11:0] ? image_1109 : _GEN_13463; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13465 = 12'h456 == _T_146[11:0] ? image_1110 : _GEN_13464; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13466 = 12'h457 == _T_146[11:0] ? image_1111 : _GEN_13465; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13467 = 12'h458 == _T_146[11:0] ? image_1112 : _GEN_13466; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13468 = 12'h459 == _T_146[11:0] ? image_1113 : _GEN_13467; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13469 = 12'h45a == _T_146[11:0] ? image_1114 : _GEN_13468; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13470 = 12'h45b == _T_146[11:0] ? image_1115 : _GEN_13469; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13471 = 12'h45c == _T_146[11:0] ? image_1116 : _GEN_13470; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13472 = 12'h45d == _T_146[11:0] ? image_1117 : _GEN_13471; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13473 = 12'h45e == _T_146[11:0] ? image_1118 : _GEN_13472; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13474 = 12'h45f == _T_146[11:0] ? image_1119 : _GEN_13473; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13475 = 12'h460 == _T_146[11:0] ? image_1120 : _GEN_13474; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13476 = 12'h461 == _T_146[11:0] ? image_1121 : _GEN_13475; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13477 = 12'h462 == _T_146[11:0] ? image_1122 : _GEN_13476; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13478 = 12'h463 == _T_146[11:0] ? image_1123 : _GEN_13477; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13479 = 12'h464 == _T_146[11:0] ? image_1124 : _GEN_13478; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13480 = 12'h465 == _T_146[11:0] ? image_1125 : _GEN_13479; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13481 = 12'h466 == _T_146[11:0] ? image_1126 : _GEN_13480; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13482 = 12'h467 == _T_146[11:0] ? image_1127 : _GEN_13481; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13483 = 12'h468 == _T_146[11:0] ? image_1128 : _GEN_13482; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13484 = 12'h469 == _T_146[11:0] ? image_1129 : _GEN_13483; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13485 = 12'h46a == _T_146[11:0] ? image_1130 : _GEN_13484; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13486 = 12'h46b == _T_146[11:0] ? image_1131 : _GEN_13485; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13487 = 12'h46c == _T_146[11:0] ? image_1132 : _GEN_13486; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13488 = 12'h46d == _T_146[11:0] ? image_1133 : _GEN_13487; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13489 = 12'h46e == _T_146[11:0] ? image_1134 : _GEN_13488; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13490 = 12'h46f == _T_146[11:0] ? image_1135 : _GEN_13489; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13491 = 12'h470 == _T_146[11:0] ? image_1136 : _GEN_13490; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13492 = 12'h471 == _T_146[11:0] ? image_1137 : _GEN_13491; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13493 = 12'h472 == _T_146[11:0] ? image_1138 : _GEN_13492; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13494 = 12'h473 == _T_146[11:0] ? image_1139 : _GEN_13493; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13495 = 12'h474 == _T_146[11:0] ? image_1140 : _GEN_13494; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13496 = 12'h475 == _T_146[11:0] ? image_1141 : _GEN_13495; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13497 = 12'h476 == _T_146[11:0] ? image_1142 : _GEN_13496; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13498 = 12'h477 == _T_146[11:0] ? image_1143 : _GEN_13497; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13499 = 12'h478 == _T_146[11:0] ? image_1144 : _GEN_13498; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13500 = 12'h479 == _T_146[11:0] ? image_1145 : _GEN_13499; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13501 = 12'h47a == _T_146[11:0] ? image_1146 : _GEN_13500; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13502 = 12'h47b == _T_146[11:0] ? image_1147 : _GEN_13501; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13503 = 12'h47c == _T_146[11:0] ? image_1148 : _GEN_13502; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13504 = 12'h47d == _T_146[11:0] ? 4'h0 : _GEN_13503; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13505 = 12'h47e == _T_146[11:0] ? 4'h0 : _GEN_13504; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13506 = 12'h47f == _T_146[11:0] ? 4'h0 : _GEN_13505; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13507 = 12'h480 == _T_146[11:0] ? image_1152 : _GEN_13506; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13508 = 12'h481 == _T_146[11:0] ? image_1153 : _GEN_13507; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13509 = 12'h482 == _T_146[11:0] ? image_1154 : _GEN_13508; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13510 = 12'h483 == _T_146[11:0] ? image_1155 : _GEN_13509; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13511 = 12'h484 == _T_146[11:0] ? image_1156 : _GEN_13510; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13512 = 12'h485 == _T_146[11:0] ? image_1157 : _GEN_13511; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13513 = 12'h486 == _T_146[11:0] ? image_1158 : _GEN_13512; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13514 = 12'h487 == _T_146[11:0] ? image_1159 : _GEN_13513; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13515 = 12'h488 == _T_146[11:0] ? image_1160 : _GEN_13514; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13516 = 12'h489 == _T_146[11:0] ? image_1161 : _GEN_13515; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13517 = 12'h48a == _T_146[11:0] ? image_1162 : _GEN_13516; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13518 = 12'h48b == _T_146[11:0] ? image_1163 : _GEN_13517; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13519 = 12'h48c == _T_146[11:0] ? image_1164 : _GEN_13518; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13520 = 12'h48d == _T_146[11:0] ? image_1165 : _GEN_13519; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13521 = 12'h48e == _T_146[11:0] ? image_1166 : _GEN_13520; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13522 = 12'h48f == _T_146[11:0] ? image_1167 : _GEN_13521; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13523 = 12'h490 == _T_146[11:0] ? image_1168 : _GEN_13522; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13524 = 12'h491 == _T_146[11:0] ? image_1169 : _GEN_13523; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13525 = 12'h492 == _T_146[11:0] ? image_1170 : _GEN_13524; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13526 = 12'h493 == _T_146[11:0] ? image_1171 : _GEN_13525; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13527 = 12'h494 == _T_146[11:0] ? image_1172 : _GEN_13526; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13528 = 12'h495 == _T_146[11:0] ? image_1173 : _GEN_13527; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13529 = 12'h496 == _T_146[11:0] ? image_1174 : _GEN_13528; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13530 = 12'h497 == _T_146[11:0] ? image_1175 : _GEN_13529; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13531 = 12'h498 == _T_146[11:0] ? image_1176 : _GEN_13530; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13532 = 12'h499 == _T_146[11:0] ? image_1177 : _GEN_13531; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13533 = 12'h49a == _T_146[11:0] ? image_1178 : _GEN_13532; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13534 = 12'h49b == _T_146[11:0] ? image_1179 : _GEN_13533; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13535 = 12'h49c == _T_146[11:0] ? image_1180 : _GEN_13534; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13536 = 12'h49d == _T_146[11:0] ? image_1181 : _GEN_13535; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13537 = 12'h49e == _T_146[11:0] ? image_1182 : _GEN_13536; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13538 = 12'h49f == _T_146[11:0] ? image_1183 : _GEN_13537; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13539 = 12'h4a0 == _T_146[11:0] ? image_1184 : _GEN_13538; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13540 = 12'h4a1 == _T_146[11:0] ? image_1185 : _GEN_13539; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13541 = 12'h4a2 == _T_146[11:0] ? image_1186 : _GEN_13540; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13542 = 12'h4a3 == _T_146[11:0] ? image_1187 : _GEN_13541; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13543 = 12'h4a4 == _T_146[11:0] ? image_1188 : _GEN_13542; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13544 = 12'h4a5 == _T_146[11:0] ? image_1189 : _GEN_13543; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13545 = 12'h4a6 == _T_146[11:0] ? image_1190 : _GEN_13544; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13546 = 12'h4a7 == _T_146[11:0] ? image_1191 : _GEN_13545; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13547 = 12'h4a8 == _T_146[11:0] ? image_1192 : _GEN_13546; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13548 = 12'h4a9 == _T_146[11:0] ? image_1193 : _GEN_13547; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13549 = 12'h4aa == _T_146[11:0] ? image_1194 : _GEN_13548; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13550 = 12'h4ab == _T_146[11:0] ? image_1195 : _GEN_13549; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13551 = 12'h4ac == _T_146[11:0] ? image_1196 : _GEN_13550; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13552 = 12'h4ad == _T_146[11:0] ? image_1197 : _GEN_13551; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13553 = 12'h4ae == _T_146[11:0] ? image_1198 : _GEN_13552; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13554 = 12'h4af == _T_146[11:0] ? image_1199 : _GEN_13553; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13555 = 12'h4b0 == _T_146[11:0] ? image_1200 : _GEN_13554; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13556 = 12'h4b1 == _T_146[11:0] ? image_1201 : _GEN_13555; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13557 = 12'h4b2 == _T_146[11:0] ? image_1202 : _GEN_13556; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13558 = 12'h4b3 == _T_146[11:0] ? image_1203 : _GEN_13557; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13559 = 12'h4b4 == _T_146[11:0] ? image_1204 : _GEN_13558; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13560 = 12'h4b5 == _T_146[11:0] ? image_1205 : _GEN_13559; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13561 = 12'h4b6 == _T_146[11:0] ? image_1206 : _GEN_13560; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13562 = 12'h4b7 == _T_146[11:0] ? image_1207 : _GEN_13561; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13563 = 12'h4b8 == _T_146[11:0] ? image_1208 : _GEN_13562; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13564 = 12'h4b9 == _T_146[11:0] ? 4'h0 : _GEN_13563; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13565 = 12'h4ba == _T_146[11:0] ? 4'h0 : _GEN_13564; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13566 = 12'h4bb == _T_146[11:0] ? 4'h0 : _GEN_13565; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13567 = 12'h4bc == _T_146[11:0] ? 4'h0 : _GEN_13566; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13568 = 12'h4bd == _T_146[11:0] ? 4'h0 : _GEN_13567; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13569 = 12'h4be == _T_146[11:0] ? 4'h0 : _GEN_13568; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13570 = 12'h4bf == _T_146[11:0] ? 4'h0 : _GEN_13569; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13571 = 12'h4c0 == _T_146[11:0] ? image_1216 : _GEN_13570; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13572 = 12'h4c1 == _T_146[11:0] ? image_1217 : _GEN_13571; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13573 = 12'h4c2 == _T_146[11:0] ? image_1218 : _GEN_13572; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13574 = 12'h4c3 == _T_146[11:0] ? image_1219 : _GEN_13573; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13575 = 12'h4c4 == _T_146[11:0] ? image_1220 : _GEN_13574; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13576 = 12'h4c5 == _T_146[11:0] ? image_1221 : _GEN_13575; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13577 = 12'h4c6 == _T_146[11:0] ? image_1222 : _GEN_13576; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13578 = 12'h4c7 == _T_146[11:0] ? image_1223 : _GEN_13577; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13579 = 12'h4c8 == _T_146[11:0] ? image_1224 : _GEN_13578; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13580 = 12'h4c9 == _T_146[11:0] ? image_1225 : _GEN_13579; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13581 = 12'h4ca == _T_146[11:0] ? image_1226 : _GEN_13580; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13582 = 12'h4cb == _T_146[11:0] ? image_1227 : _GEN_13581; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13583 = 12'h4cc == _T_146[11:0] ? image_1228 : _GEN_13582; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13584 = 12'h4cd == _T_146[11:0] ? image_1229 : _GEN_13583; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13585 = 12'h4ce == _T_146[11:0] ? image_1230 : _GEN_13584; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13586 = 12'h4cf == _T_146[11:0] ? image_1231 : _GEN_13585; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13587 = 12'h4d0 == _T_146[11:0] ? image_1232 : _GEN_13586; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13588 = 12'h4d1 == _T_146[11:0] ? image_1233 : _GEN_13587; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13589 = 12'h4d2 == _T_146[11:0] ? image_1234 : _GEN_13588; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13590 = 12'h4d3 == _T_146[11:0] ? image_1235 : _GEN_13589; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13591 = 12'h4d4 == _T_146[11:0] ? image_1236 : _GEN_13590; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13592 = 12'h4d5 == _T_146[11:0] ? image_1237 : _GEN_13591; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13593 = 12'h4d6 == _T_146[11:0] ? image_1238 : _GEN_13592; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13594 = 12'h4d7 == _T_146[11:0] ? image_1239 : _GEN_13593; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13595 = 12'h4d8 == _T_146[11:0] ? image_1240 : _GEN_13594; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13596 = 12'h4d9 == _T_146[11:0] ? image_1241 : _GEN_13595; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13597 = 12'h4da == _T_146[11:0] ? image_1242 : _GEN_13596; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13598 = 12'h4db == _T_146[11:0] ? image_1243 : _GEN_13597; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13599 = 12'h4dc == _T_146[11:0] ? image_1244 : _GEN_13598; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13600 = 12'h4dd == _T_146[11:0] ? image_1245 : _GEN_13599; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13601 = 12'h4de == _T_146[11:0] ? image_1246 : _GEN_13600; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13602 = 12'h4df == _T_146[11:0] ? image_1247 : _GEN_13601; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13603 = 12'h4e0 == _T_146[11:0] ? image_1248 : _GEN_13602; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13604 = 12'h4e1 == _T_146[11:0] ? image_1249 : _GEN_13603; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13605 = 12'h4e2 == _T_146[11:0] ? image_1250 : _GEN_13604; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13606 = 12'h4e3 == _T_146[11:0] ? image_1251 : _GEN_13605; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13607 = 12'h4e4 == _T_146[11:0] ? image_1252 : _GEN_13606; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13608 = 12'h4e5 == _T_146[11:0] ? image_1253 : _GEN_13607; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13609 = 12'h4e6 == _T_146[11:0] ? image_1254 : _GEN_13608; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13610 = 12'h4e7 == _T_146[11:0] ? image_1255 : _GEN_13609; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13611 = 12'h4e8 == _T_146[11:0] ? image_1256 : _GEN_13610; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13612 = 12'h4e9 == _T_146[11:0] ? image_1257 : _GEN_13611; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13613 = 12'h4ea == _T_146[11:0] ? image_1258 : _GEN_13612; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13614 = 12'h4eb == _T_146[11:0] ? image_1259 : _GEN_13613; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13615 = 12'h4ec == _T_146[11:0] ? image_1260 : _GEN_13614; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13616 = 12'h4ed == _T_146[11:0] ? image_1261 : _GEN_13615; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13617 = 12'h4ee == _T_146[11:0] ? image_1262 : _GEN_13616; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13618 = 12'h4ef == _T_146[11:0] ? image_1263 : _GEN_13617; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13619 = 12'h4f0 == _T_146[11:0] ? image_1264 : _GEN_13618; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13620 = 12'h4f1 == _T_146[11:0] ? image_1265 : _GEN_13619; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13621 = 12'h4f2 == _T_146[11:0] ? image_1266 : _GEN_13620; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13622 = 12'h4f3 == _T_146[11:0] ? image_1267 : _GEN_13621; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13623 = 12'h4f4 == _T_146[11:0] ? image_1268 : _GEN_13622; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13624 = 12'h4f5 == _T_146[11:0] ? image_1269 : _GEN_13623; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13625 = 12'h4f6 == _T_146[11:0] ? image_1270 : _GEN_13624; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13626 = 12'h4f7 == _T_146[11:0] ? image_1271 : _GEN_13625; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13627 = 12'h4f8 == _T_146[11:0] ? image_1272 : _GEN_13626; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13628 = 12'h4f9 == _T_146[11:0] ? image_1273 : _GEN_13627; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13629 = 12'h4fa == _T_146[11:0] ? image_1274 : _GEN_13628; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13630 = 12'h4fb == _T_146[11:0] ? image_1275 : _GEN_13629; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13631 = 12'h4fc == _T_146[11:0] ? 4'h0 : _GEN_13630; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13632 = 12'h4fd == _T_146[11:0] ? 4'h0 : _GEN_13631; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13633 = 12'h4fe == _T_146[11:0] ? 4'h0 : _GEN_13632; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13634 = 12'h4ff == _T_146[11:0] ? 4'h0 : _GEN_13633; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13635 = 12'h500 == _T_146[11:0] ? image_1280 : _GEN_13634; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13636 = 12'h501 == _T_146[11:0] ? image_1281 : _GEN_13635; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13637 = 12'h502 == _T_146[11:0] ? image_1282 : _GEN_13636; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13638 = 12'h503 == _T_146[11:0] ? image_1283 : _GEN_13637; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13639 = 12'h504 == _T_146[11:0] ? image_1284 : _GEN_13638; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13640 = 12'h505 == _T_146[11:0] ? image_1285 : _GEN_13639; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13641 = 12'h506 == _T_146[11:0] ? image_1286 : _GEN_13640; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13642 = 12'h507 == _T_146[11:0] ? image_1287 : _GEN_13641; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13643 = 12'h508 == _T_146[11:0] ? image_1288 : _GEN_13642; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13644 = 12'h509 == _T_146[11:0] ? image_1289 : _GEN_13643; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13645 = 12'h50a == _T_146[11:0] ? image_1290 : _GEN_13644; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13646 = 12'h50b == _T_146[11:0] ? image_1291 : _GEN_13645; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13647 = 12'h50c == _T_146[11:0] ? image_1292 : _GEN_13646; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13648 = 12'h50d == _T_146[11:0] ? image_1293 : _GEN_13647; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13649 = 12'h50e == _T_146[11:0] ? image_1294 : _GEN_13648; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13650 = 12'h50f == _T_146[11:0] ? image_1295 : _GEN_13649; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13651 = 12'h510 == _T_146[11:0] ? image_1296 : _GEN_13650; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13652 = 12'h511 == _T_146[11:0] ? image_1297 : _GEN_13651; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13653 = 12'h512 == _T_146[11:0] ? image_1298 : _GEN_13652; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13654 = 12'h513 == _T_146[11:0] ? image_1299 : _GEN_13653; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13655 = 12'h514 == _T_146[11:0] ? image_1300 : _GEN_13654; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13656 = 12'h515 == _T_146[11:0] ? image_1301 : _GEN_13655; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13657 = 12'h516 == _T_146[11:0] ? image_1302 : _GEN_13656; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13658 = 12'h517 == _T_146[11:0] ? image_1303 : _GEN_13657; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13659 = 12'h518 == _T_146[11:0] ? image_1304 : _GEN_13658; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13660 = 12'h519 == _T_146[11:0] ? image_1305 : _GEN_13659; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13661 = 12'h51a == _T_146[11:0] ? image_1306 : _GEN_13660; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13662 = 12'h51b == _T_146[11:0] ? image_1307 : _GEN_13661; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13663 = 12'h51c == _T_146[11:0] ? image_1308 : _GEN_13662; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13664 = 12'h51d == _T_146[11:0] ? image_1309 : _GEN_13663; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13665 = 12'h51e == _T_146[11:0] ? image_1310 : _GEN_13664; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13666 = 12'h51f == _T_146[11:0] ? image_1311 : _GEN_13665; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13667 = 12'h520 == _T_146[11:0] ? image_1312 : _GEN_13666; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13668 = 12'h521 == _T_146[11:0] ? image_1313 : _GEN_13667; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13669 = 12'h522 == _T_146[11:0] ? image_1314 : _GEN_13668; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13670 = 12'h523 == _T_146[11:0] ? image_1315 : _GEN_13669; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13671 = 12'h524 == _T_146[11:0] ? image_1316 : _GEN_13670; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13672 = 12'h525 == _T_146[11:0] ? image_1317 : _GEN_13671; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13673 = 12'h526 == _T_146[11:0] ? image_1318 : _GEN_13672; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13674 = 12'h527 == _T_146[11:0] ? image_1319 : _GEN_13673; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13675 = 12'h528 == _T_146[11:0] ? image_1320 : _GEN_13674; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13676 = 12'h529 == _T_146[11:0] ? image_1321 : _GEN_13675; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13677 = 12'h52a == _T_146[11:0] ? image_1322 : _GEN_13676; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13678 = 12'h52b == _T_146[11:0] ? image_1323 : _GEN_13677; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13679 = 12'h52c == _T_146[11:0] ? image_1324 : _GEN_13678; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13680 = 12'h52d == _T_146[11:0] ? image_1325 : _GEN_13679; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13681 = 12'h52e == _T_146[11:0] ? image_1326 : _GEN_13680; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13682 = 12'h52f == _T_146[11:0] ? image_1327 : _GEN_13681; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13683 = 12'h530 == _T_146[11:0] ? image_1328 : _GEN_13682; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13684 = 12'h531 == _T_146[11:0] ? image_1329 : _GEN_13683; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13685 = 12'h532 == _T_146[11:0] ? image_1330 : _GEN_13684; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13686 = 12'h533 == _T_146[11:0] ? image_1331 : _GEN_13685; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13687 = 12'h534 == _T_146[11:0] ? image_1332 : _GEN_13686; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13688 = 12'h535 == _T_146[11:0] ? image_1333 : _GEN_13687; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13689 = 12'h536 == _T_146[11:0] ? image_1334 : _GEN_13688; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13690 = 12'h537 == _T_146[11:0] ? image_1335 : _GEN_13689; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13691 = 12'h538 == _T_146[11:0] ? image_1336 : _GEN_13690; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13692 = 12'h539 == _T_146[11:0] ? image_1337 : _GEN_13691; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13693 = 12'h53a == _T_146[11:0] ? image_1338 : _GEN_13692; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13694 = 12'h53b == _T_146[11:0] ? image_1339 : _GEN_13693; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13695 = 12'h53c == _T_146[11:0] ? image_1340 : _GEN_13694; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13696 = 12'h53d == _T_146[11:0] ? image_1341 : _GEN_13695; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13697 = 12'h53e == _T_146[11:0] ? 4'h0 : _GEN_13696; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13698 = 12'h53f == _T_146[11:0] ? 4'h0 : _GEN_13697; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13699 = 12'h540 == _T_146[11:0] ? image_1344 : _GEN_13698; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13700 = 12'h541 == _T_146[11:0] ? image_1345 : _GEN_13699; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13701 = 12'h542 == _T_146[11:0] ? image_1346 : _GEN_13700; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13702 = 12'h543 == _T_146[11:0] ? image_1347 : _GEN_13701; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13703 = 12'h544 == _T_146[11:0] ? image_1348 : _GEN_13702; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13704 = 12'h545 == _T_146[11:0] ? image_1349 : _GEN_13703; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13705 = 12'h546 == _T_146[11:0] ? image_1350 : _GEN_13704; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13706 = 12'h547 == _T_146[11:0] ? image_1351 : _GEN_13705; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13707 = 12'h548 == _T_146[11:0] ? image_1352 : _GEN_13706; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13708 = 12'h549 == _T_146[11:0] ? image_1353 : _GEN_13707; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13709 = 12'h54a == _T_146[11:0] ? image_1354 : _GEN_13708; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13710 = 12'h54b == _T_146[11:0] ? image_1355 : _GEN_13709; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13711 = 12'h54c == _T_146[11:0] ? image_1356 : _GEN_13710; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13712 = 12'h54d == _T_146[11:0] ? image_1357 : _GEN_13711; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13713 = 12'h54e == _T_146[11:0] ? image_1358 : _GEN_13712; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13714 = 12'h54f == _T_146[11:0] ? image_1359 : _GEN_13713; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13715 = 12'h550 == _T_146[11:0] ? image_1360 : _GEN_13714; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13716 = 12'h551 == _T_146[11:0] ? image_1361 : _GEN_13715; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13717 = 12'h552 == _T_146[11:0] ? image_1362 : _GEN_13716; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13718 = 12'h553 == _T_146[11:0] ? image_1363 : _GEN_13717; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13719 = 12'h554 == _T_146[11:0] ? image_1364 : _GEN_13718; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13720 = 12'h555 == _T_146[11:0] ? image_1365 : _GEN_13719; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13721 = 12'h556 == _T_146[11:0] ? image_1366 : _GEN_13720; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13722 = 12'h557 == _T_146[11:0] ? image_1367 : _GEN_13721; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13723 = 12'h558 == _T_146[11:0] ? image_1368 : _GEN_13722; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13724 = 12'h559 == _T_146[11:0] ? image_1369 : _GEN_13723; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13725 = 12'h55a == _T_146[11:0] ? image_1370 : _GEN_13724; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13726 = 12'h55b == _T_146[11:0] ? image_1371 : _GEN_13725; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13727 = 12'h55c == _T_146[11:0] ? image_1372 : _GEN_13726; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13728 = 12'h55d == _T_146[11:0] ? image_1373 : _GEN_13727; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13729 = 12'h55e == _T_146[11:0] ? image_1374 : _GEN_13728; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13730 = 12'h55f == _T_146[11:0] ? image_1375 : _GEN_13729; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13731 = 12'h560 == _T_146[11:0] ? image_1376 : _GEN_13730; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13732 = 12'h561 == _T_146[11:0] ? image_1377 : _GEN_13731; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13733 = 12'h562 == _T_146[11:0] ? image_1378 : _GEN_13732; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13734 = 12'h563 == _T_146[11:0] ? image_1379 : _GEN_13733; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13735 = 12'h564 == _T_146[11:0] ? image_1380 : _GEN_13734; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13736 = 12'h565 == _T_146[11:0] ? image_1381 : _GEN_13735; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13737 = 12'h566 == _T_146[11:0] ? image_1382 : _GEN_13736; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13738 = 12'h567 == _T_146[11:0] ? image_1383 : _GEN_13737; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13739 = 12'h568 == _T_146[11:0] ? image_1384 : _GEN_13738; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13740 = 12'h569 == _T_146[11:0] ? image_1385 : _GEN_13739; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13741 = 12'h56a == _T_146[11:0] ? image_1386 : _GEN_13740; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13742 = 12'h56b == _T_146[11:0] ? image_1387 : _GEN_13741; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13743 = 12'h56c == _T_146[11:0] ? image_1388 : _GEN_13742; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13744 = 12'h56d == _T_146[11:0] ? image_1389 : _GEN_13743; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13745 = 12'h56e == _T_146[11:0] ? image_1390 : _GEN_13744; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13746 = 12'h56f == _T_146[11:0] ? image_1391 : _GEN_13745; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13747 = 12'h570 == _T_146[11:0] ? image_1392 : _GEN_13746; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13748 = 12'h571 == _T_146[11:0] ? image_1393 : _GEN_13747; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13749 = 12'h572 == _T_146[11:0] ? image_1394 : _GEN_13748; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13750 = 12'h573 == _T_146[11:0] ? image_1395 : _GEN_13749; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13751 = 12'h574 == _T_146[11:0] ? image_1396 : _GEN_13750; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13752 = 12'h575 == _T_146[11:0] ? image_1397 : _GEN_13751; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13753 = 12'h576 == _T_146[11:0] ? image_1398 : _GEN_13752; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13754 = 12'h577 == _T_146[11:0] ? image_1399 : _GEN_13753; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13755 = 12'h578 == _T_146[11:0] ? image_1400 : _GEN_13754; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13756 = 12'h579 == _T_146[11:0] ? image_1401 : _GEN_13755; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13757 = 12'h57a == _T_146[11:0] ? image_1402 : _GEN_13756; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13758 = 12'h57b == _T_146[11:0] ? image_1403 : _GEN_13757; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13759 = 12'h57c == _T_146[11:0] ? image_1404 : _GEN_13758; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13760 = 12'h57d == _T_146[11:0] ? image_1405 : _GEN_13759; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13761 = 12'h57e == _T_146[11:0] ? 4'h0 : _GEN_13760; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13762 = 12'h57f == _T_146[11:0] ? 4'h0 : _GEN_13761; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13763 = 12'h580 == _T_146[11:0] ? image_1408 : _GEN_13762; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13764 = 12'h581 == _T_146[11:0] ? image_1409 : _GEN_13763; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13765 = 12'h582 == _T_146[11:0] ? image_1410 : _GEN_13764; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13766 = 12'h583 == _T_146[11:0] ? image_1411 : _GEN_13765; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13767 = 12'h584 == _T_146[11:0] ? image_1412 : _GEN_13766; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13768 = 12'h585 == _T_146[11:0] ? image_1413 : _GEN_13767; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13769 = 12'h586 == _T_146[11:0] ? image_1414 : _GEN_13768; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13770 = 12'h587 == _T_146[11:0] ? image_1415 : _GEN_13769; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13771 = 12'h588 == _T_146[11:0] ? image_1416 : _GEN_13770; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13772 = 12'h589 == _T_146[11:0] ? image_1417 : _GEN_13771; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13773 = 12'h58a == _T_146[11:0] ? image_1418 : _GEN_13772; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13774 = 12'h58b == _T_146[11:0] ? image_1419 : _GEN_13773; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13775 = 12'h58c == _T_146[11:0] ? image_1420 : _GEN_13774; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13776 = 12'h58d == _T_146[11:0] ? image_1421 : _GEN_13775; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13777 = 12'h58e == _T_146[11:0] ? image_1422 : _GEN_13776; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13778 = 12'h58f == _T_146[11:0] ? image_1423 : _GEN_13777; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13779 = 12'h590 == _T_146[11:0] ? image_1424 : _GEN_13778; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13780 = 12'h591 == _T_146[11:0] ? image_1425 : _GEN_13779; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13781 = 12'h592 == _T_146[11:0] ? image_1426 : _GEN_13780; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13782 = 12'h593 == _T_146[11:0] ? image_1427 : _GEN_13781; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13783 = 12'h594 == _T_146[11:0] ? image_1428 : _GEN_13782; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13784 = 12'h595 == _T_146[11:0] ? image_1429 : _GEN_13783; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13785 = 12'h596 == _T_146[11:0] ? image_1430 : _GEN_13784; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13786 = 12'h597 == _T_146[11:0] ? image_1431 : _GEN_13785; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13787 = 12'h598 == _T_146[11:0] ? image_1432 : _GEN_13786; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13788 = 12'h599 == _T_146[11:0] ? image_1433 : _GEN_13787; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13789 = 12'h59a == _T_146[11:0] ? image_1434 : _GEN_13788; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13790 = 12'h59b == _T_146[11:0] ? image_1435 : _GEN_13789; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13791 = 12'h59c == _T_146[11:0] ? image_1436 : _GEN_13790; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13792 = 12'h59d == _T_146[11:0] ? image_1437 : _GEN_13791; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13793 = 12'h59e == _T_146[11:0] ? image_1438 : _GEN_13792; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13794 = 12'h59f == _T_146[11:0] ? image_1439 : _GEN_13793; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13795 = 12'h5a0 == _T_146[11:0] ? image_1440 : _GEN_13794; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13796 = 12'h5a1 == _T_146[11:0] ? image_1441 : _GEN_13795; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13797 = 12'h5a2 == _T_146[11:0] ? image_1442 : _GEN_13796; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13798 = 12'h5a3 == _T_146[11:0] ? image_1443 : _GEN_13797; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13799 = 12'h5a4 == _T_146[11:0] ? image_1444 : _GEN_13798; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13800 = 12'h5a5 == _T_146[11:0] ? image_1445 : _GEN_13799; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13801 = 12'h5a6 == _T_146[11:0] ? image_1446 : _GEN_13800; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13802 = 12'h5a7 == _T_146[11:0] ? image_1447 : _GEN_13801; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13803 = 12'h5a8 == _T_146[11:0] ? image_1448 : _GEN_13802; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13804 = 12'h5a9 == _T_146[11:0] ? image_1449 : _GEN_13803; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13805 = 12'h5aa == _T_146[11:0] ? image_1450 : _GEN_13804; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13806 = 12'h5ab == _T_146[11:0] ? image_1451 : _GEN_13805; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13807 = 12'h5ac == _T_146[11:0] ? image_1452 : _GEN_13806; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13808 = 12'h5ad == _T_146[11:0] ? image_1453 : _GEN_13807; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13809 = 12'h5ae == _T_146[11:0] ? image_1454 : _GEN_13808; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13810 = 12'h5af == _T_146[11:0] ? image_1455 : _GEN_13809; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13811 = 12'h5b0 == _T_146[11:0] ? image_1456 : _GEN_13810; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13812 = 12'h5b1 == _T_146[11:0] ? image_1457 : _GEN_13811; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13813 = 12'h5b2 == _T_146[11:0] ? image_1458 : _GEN_13812; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13814 = 12'h5b3 == _T_146[11:0] ? image_1459 : _GEN_13813; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13815 = 12'h5b4 == _T_146[11:0] ? image_1460 : _GEN_13814; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13816 = 12'h5b5 == _T_146[11:0] ? image_1461 : _GEN_13815; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13817 = 12'h5b6 == _T_146[11:0] ? image_1462 : _GEN_13816; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13818 = 12'h5b7 == _T_146[11:0] ? image_1463 : _GEN_13817; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13819 = 12'h5b8 == _T_146[11:0] ? image_1464 : _GEN_13818; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13820 = 12'h5b9 == _T_146[11:0] ? image_1465 : _GEN_13819; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13821 = 12'h5ba == _T_146[11:0] ? image_1466 : _GEN_13820; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13822 = 12'h5bb == _T_146[11:0] ? image_1467 : _GEN_13821; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13823 = 12'h5bc == _T_146[11:0] ? image_1468 : _GEN_13822; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13824 = 12'h5bd == _T_146[11:0] ? image_1469 : _GEN_13823; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13825 = 12'h5be == _T_146[11:0] ? 4'h0 : _GEN_13824; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13826 = 12'h5bf == _T_146[11:0] ? 4'h0 : _GEN_13825; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13827 = 12'h5c0 == _T_146[11:0] ? image_1472 : _GEN_13826; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13828 = 12'h5c1 == _T_146[11:0] ? image_1473 : _GEN_13827; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13829 = 12'h5c2 == _T_146[11:0] ? image_1474 : _GEN_13828; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13830 = 12'h5c3 == _T_146[11:0] ? image_1475 : _GEN_13829; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13831 = 12'h5c4 == _T_146[11:0] ? image_1476 : _GEN_13830; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13832 = 12'h5c5 == _T_146[11:0] ? image_1477 : _GEN_13831; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13833 = 12'h5c6 == _T_146[11:0] ? image_1478 : _GEN_13832; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13834 = 12'h5c7 == _T_146[11:0] ? image_1479 : _GEN_13833; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13835 = 12'h5c8 == _T_146[11:0] ? image_1480 : _GEN_13834; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13836 = 12'h5c9 == _T_146[11:0] ? image_1481 : _GEN_13835; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13837 = 12'h5ca == _T_146[11:0] ? image_1482 : _GEN_13836; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13838 = 12'h5cb == _T_146[11:0] ? image_1483 : _GEN_13837; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13839 = 12'h5cc == _T_146[11:0] ? image_1484 : _GEN_13838; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13840 = 12'h5cd == _T_146[11:0] ? image_1485 : _GEN_13839; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13841 = 12'h5ce == _T_146[11:0] ? image_1486 : _GEN_13840; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13842 = 12'h5cf == _T_146[11:0] ? image_1487 : _GEN_13841; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13843 = 12'h5d0 == _T_146[11:0] ? image_1488 : _GEN_13842; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13844 = 12'h5d1 == _T_146[11:0] ? image_1489 : _GEN_13843; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13845 = 12'h5d2 == _T_146[11:0] ? image_1490 : _GEN_13844; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13846 = 12'h5d3 == _T_146[11:0] ? image_1491 : _GEN_13845; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13847 = 12'h5d4 == _T_146[11:0] ? image_1492 : _GEN_13846; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13848 = 12'h5d5 == _T_146[11:0] ? image_1493 : _GEN_13847; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13849 = 12'h5d6 == _T_146[11:0] ? image_1494 : _GEN_13848; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13850 = 12'h5d7 == _T_146[11:0] ? image_1495 : _GEN_13849; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13851 = 12'h5d8 == _T_146[11:0] ? image_1496 : _GEN_13850; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13852 = 12'h5d9 == _T_146[11:0] ? image_1497 : _GEN_13851; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13853 = 12'h5da == _T_146[11:0] ? image_1498 : _GEN_13852; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13854 = 12'h5db == _T_146[11:0] ? image_1499 : _GEN_13853; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13855 = 12'h5dc == _T_146[11:0] ? image_1500 : _GEN_13854; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13856 = 12'h5dd == _T_146[11:0] ? image_1501 : _GEN_13855; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13857 = 12'h5de == _T_146[11:0] ? image_1502 : _GEN_13856; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13858 = 12'h5df == _T_146[11:0] ? image_1503 : _GEN_13857; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13859 = 12'h5e0 == _T_146[11:0] ? image_1504 : _GEN_13858; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13860 = 12'h5e1 == _T_146[11:0] ? image_1505 : _GEN_13859; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13861 = 12'h5e2 == _T_146[11:0] ? image_1506 : _GEN_13860; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13862 = 12'h5e3 == _T_146[11:0] ? image_1507 : _GEN_13861; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13863 = 12'h5e4 == _T_146[11:0] ? image_1508 : _GEN_13862; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13864 = 12'h5e5 == _T_146[11:0] ? image_1509 : _GEN_13863; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13865 = 12'h5e6 == _T_146[11:0] ? image_1510 : _GEN_13864; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13866 = 12'h5e7 == _T_146[11:0] ? image_1511 : _GEN_13865; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13867 = 12'h5e8 == _T_146[11:0] ? image_1512 : _GEN_13866; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13868 = 12'h5e9 == _T_146[11:0] ? image_1513 : _GEN_13867; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13869 = 12'h5ea == _T_146[11:0] ? image_1514 : _GEN_13868; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13870 = 12'h5eb == _T_146[11:0] ? image_1515 : _GEN_13869; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13871 = 12'h5ec == _T_146[11:0] ? image_1516 : _GEN_13870; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13872 = 12'h5ed == _T_146[11:0] ? image_1517 : _GEN_13871; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13873 = 12'h5ee == _T_146[11:0] ? image_1518 : _GEN_13872; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13874 = 12'h5ef == _T_146[11:0] ? image_1519 : _GEN_13873; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13875 = 12'h5f0 == _T_146[11:0] ? image_1520 : _GEN_13874; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13876 = 12'h5f1 == _T_146[11:0] ? image_1521 : _GEN_13875; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13877 = 12'h5f2 == _T_146[11:0] ? image_1522 : _GEN_13876; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13878 = 12'h5f3 == _T_146[11:0] ? image_1523 : _GEN_13877; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13879 = 12'h5f4 == _T_146[11:0] ? image_1524 : _GEN_13878; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13880 = 12'h5f5 == _T_146[11:0] ? image_1525 : _GEN_13879; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13881 = 12'h5f6 == _T_146[11:0] ? image_1526 : _GEN_13880; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13882 = 12'h5f7 == _T_146[11:0] ? image_1527 : _GEN_13881; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13883 = 12'h5f8 == _T_146[11:0] ? image_1528 : _GEN_13882; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13884 = 12'h5f9 == _T_146[11:0] ? image_1529 : _GEN_13883; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13885 = 12'h5fa == _T_146[11:0] ? image_1530 : _GEN_13884; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13886 = 12'h5fb == _T_146[11:0] ? image_1531 : _GEN_13885; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13887 = 12'h5fc == _T_146[11:0] ? image_1532 : _GEN_13886; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13888 = 12'h5fd == _T_146[11:0] ? image_1533 : _GEN_13887; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13889 = 12'h5fe == _T_146[11:0] ? 4'h0 : _GEN_13888; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13890 = 12'h5ff == _T_146[11:0] ? 4'h0 : _GEN_13889; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13891 = 12'h600 == _T_146[11:0] ? image_1536 : _GEN_13890; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13892 = 12'h601 == _T_146[11:0] ? image_1537 : _GEN_13891; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13893 = 12'h602 == _T_146[11:0] ? image_1538 : _GEN_13892; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13894 = 12'h603 == _T_146[11:0] ? image_1539 : _GEN_13893; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13895 = 12'h604 == _T_146[11:0] ? image_1540 : _GEN_13894; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13896 = 12'h605 == _T_146[11:0] ? image_1541 : _GEN_13895; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13897 = 12'h606 == _T_146[11:0] ? image_1542 : _GEN_13896; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13898 = 12'h607 == _T_146[11:0] ? image_1543 : _GEN_13897; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13899 = 12'h608 == _T_146[11:0] ? image_1544 : _GEN_13898; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13900 = 12'h609 == _T_146[11:0] ? image_1545 : _GEN_13899; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13901 = 12'h60a == _T_146[11:0] ? image_1546 : _GEN_13900; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13902 = 12'h60b == _T_146[11:0] ? image_1547 : _GEN_13901; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13903 = 12'h60c == _T_146[11:0] ? image_1548 : _GEN_13902; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13904 = 12'h60d == _T_146[11:0] ? image_1549 : _GEN_13903; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13905 = 12'h60e == _T_146[11:0] ? image_1550 : _GEN_13904; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13906 = 12'h60f == _T_146[11:0] ? image_1551 : _GEN_13905; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13907 = 12'h610 == _T_146[11:0] ? image_1552 : _GEN_13906; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13908 = 12'h611 == _T_146[11:0] ? image_1553 : _GEN_13907; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13909 = 12'h612 == _T_146[11:0] ? image_1554 : _GEN_13908; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13910 = 12'h613 == _T_146[11:0] ? image_1555 : _GEN_13909; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13911 = 12'h614 == _T_146[11:0] ? image_1556 : _GEN_13910; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13912 = 12'h615 == _T_146[11:0] ? image_1557 : _GEN_13911; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13913 = 12'h616 == _T_146[11:0] ? image_1558 : _GEN_13912; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13914 = 12'h617 == _T_146[11:0] ? image_1559 : _GEN_13913; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13915 = 12'h618 == _T_146[11:0] ? image_1560 : _GEN_13914; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13916 = 12'h619 == _T_146[11:0] ? image_1561 : _GEN_13915; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13917 = 12'h61a == _T_146[11:0] ? image_1562 : _GEN_13916; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13918 = 12'h61b == _T_146[11:0] ? image_1563 : _GEN_13917; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13919 = 12'h61c == _T_146[11:0] ? image_1564 : _GEN_13918; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13920 = 12'h61d == _T_146[11:0] ? image_1565 : _GEN_13919; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13921 = 12'h61e == _T_146[11:0] ? image_1566 : _GEN_13920; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13922 = 12'h61f == _T_146[11:0] ? image_1567 : _GEN_13921; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13923 = 12'h620 == _T_146[11:0] ? image_1568 : _GEN_13922; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13924 = 12'h621 == _T_146[11:0] ? image_1569 : _GEN_13923; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13925 = 12'h622 == _T_146[11:0] ? image_1570 : _GEN_13924; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13926 = 12'h623 == _T_146[11:0] ? image_1571 : _GEN_13925; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13927 = 12'h624 == _T_146[11:0] ? image_1572 : _GEN_13926; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13928 = 12'h625 == _T_146[11:0] ? image_1573 : _GEN_13927; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13929 = 12'h626 == _T_146[11:0] ? image_1574 : _GEN_13928; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13930 = 12'h627 == _T_146[11:0] ? image_1575 : _GEN_13929; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13931 = 12'h628 == _T_146[11:0] ? image_1576 : _GEN_13930; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13932 = 12'h629 == _T_146[11:0] ? image_1577 : _GEN_13931; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13933 = 12'h62a == _T_146[11:0] ? image_1578 : _GEN_13932; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13934 = 12'h62b == _T_146[11:0] ? image_1579 : _GEN_13933; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13935 = 12'h62c == _T_146[11:0] ? image_1580 : _GEN_13934; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13936 = 12'h62d == _T_146[11:0] ? image_1581 : _GEN_13935; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13937 = 12'h62e == _T_146[11:0] ? image_1582 : _GEN_13936; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13938 = 12'h62f == _T_146[11:0] ? image_1583 : _GEN_13937; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13939 = 12'h630 == _T_146[11:0] ? image_1584 : _GEN_13938; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13940 = 12'h631 == _T_146[11:0] ? image_1585 : _GEN_13939; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13941 = 12'h632 == _T_146[11:0] ? image_1586 : _GEN_13940; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13942 = 12'h633 == _T_146[11:0] ? image_1587 : _GEN_13941; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13943 = 12'h634 == _T_146[11:0] ? image_1588 : _GEN_13942; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13944 = 12'h635 == _T_146[11:0] ? image_1589 : _GEN_13943; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13945 = 12'h636 == _T_146[11:0] ? image_1590 : _GEN_13944; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13946 = 12'h637 == _T_146[11:0] ? image_1591 : _GEN_13945; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13947 = 12'h638 == _T_146[11:0] ? image_1592 : _GEN_13946; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13948 = 12'h639 == _T_146[11:0] ? image_1593 : _GEN_13947; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13949 = 12'h63a == _T_146[11:0] ? image_1594 : _GEN_13948; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13950 = 12'h63b == _T_146[11:0] ? image_1595 : _GEN_13949; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13951 = 12'h63c == _T_146[11:0] ? image_1596 : _GEN_13950; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13952 = 12'h63d == _T_146[11:0] ? image_1597 : _GEN_13951; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13953 = 12'h63e == _T_146[11:0] ? 4'h0 : _GEN_13952; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13954 = 12'h63f == _T_146[11:0] ? 4'h0 : _GEN_13953; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13955 = 12'h640 == _T_146[11:0] ? image_1600 : _GEN_13954; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13956 = 12'h641 == _T_146[11:0] ? image_1601 : _GEN_13955; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13957 = 12'h642 == _T_146[11:0] ? image_1602 : _GEN_13956; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13958 = 12'h643 == _T_146[11:0] ? image_1603 : _GEN_13957; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13959 = 12'h644 == _T_146[11:0] ? image_1604 : _GEN_13958; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13960 = 12'h645 == _T_146[11:0] ? image_1605 : _GEN_13959; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13961 = 12'h646 == _T_146[11:0] ? image_1606 : _GEN_13960; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13962 = 12'h647 == _T_146[11:0] ? image_1607 : _GEN_13961; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13963 = 12'h648 == _T_146[11:0] ? image_1608 : _GEN_13962; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13964 = 12'h649 == _T_146[11:0] ? image_1609 : _GEN_13963; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13965 = 12'h64a == _T_146[11:0] ? image_1610 : _GEN_13964; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13966 = 12'h64b == _T_146[11:0] ? image_1611 : _GEN_13965; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13967 = 12'h64c == _T_146[11:0] ? image_1612 : _GEN_13966; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13968 = 12'h64d == _T_146[11:0] ? image_1613 : _GEN_13967; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13969 = 12'h64e == _T_146[11:0] ? image_1614 : _GEN_13968; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13970 = 12'h64f == _T_146[11:0] ? image_1615 : _GEN_13969; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13971 = 12'h650 == _T_146[11:0] ? image_1616 : _GEN_13970; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13972 = 12'h651 == _T_146[11:0] ? image_1617 : _GEN_13971; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13973 = 12'h652 == _T_146[11:0] ? image_1618 : _GEN_13972; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13974 = 12'h653 == _T_146[11:0] ? image_1619 : _GEN_13973; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13975 = 12'h654 == _T_146[11:0] ? image_1620 : _GEN_13974; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13976 = 12'h655 == _T_146[11:0] ? image_1621 : _GEN_13975; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13977 = 12'h656 == _T_146[11:0] ? image_1622 : _GEN_13976; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13978 = 12'h657 == _T_146[11:0] ? image_1623 : _GEN_13977; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13979 = 12'h658 == _T_146[11:0] ? image_1624 : _GEN_13978; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13980 = 12'h659 == _T_146[11:0] ? image_1625 : _GEN_13979; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13981 = 12'h65a == _T_146[11:0] ? image_1626 : _GEN_13980; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13982 = 12'h65b == _T_146[11:0] ? image_1627 : _GEN_13981; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13983 = 12'h65c == _T_146[11:0] ? image_1628 : _GEN_13982; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13984 = 12'h65d == _T_146[11:0] ? image_1629 : _GEN_13983; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13985 = 12'h65e == _T_146[11:0] ? image_1630 : _GEN_13984; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13986 = 12'h65f == _T_146[11:0] ? image_1631 : _GEN_13985; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13987 = 12'h660 == _T_146[11:0] ? image_1632 : _GEN_13986; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13988 = 12'h661 == _T_146[11:0] ? image_1633 : _GEN_13987; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13989 = 12'h662 == _T_146[11:0] ? image_1634 : _GEN_13988; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13990 = 12'h663 == _T_146[11:0] ? image_1635 : _GEN_13989; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13991 = 12'h664 == _T_146[11:0] ? image_1636 : _GEN_13990; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13992 = 12'h665 == _T_146[11:0] ? image_1637 : _GEN_13991; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13993 = 12'h666 == _T_146[11:0] ? image_1638 : _GEN_13992; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13994 = 12'h667 == _T_146[11:0] ? image_1639 : _GEN_13993; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13995 = 12'h668 == _T_146[11:0] ? image_1640 : _GEN_13994; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13996 = 12'h669 == _T_146[11:0] ? image_1641 : _GEN_13995; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13997 = 12'h66a == _T_146[11:0] ? image_1642 : _GEN_13996; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13998 = 12'h66b == _T_146[11:0] ? image_1643 : _GEN_13997; // @[Filter.scala 138:46]
  wire [3:0] _GEN_13999 = 12'h66c == _T_146[11:0] ? image_1644 : _GEN_13998; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14000 = 12'h66d == _T_146[11:0] ? image_1645 : _GEN_13999; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14001 = 12'h66e == _T_146[11:0] ? image_1646 : _GEN_14000; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14002 = 12'h66f == _T_146[11:0] ? image_1647 : _GEN_14001; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14003 = 12'h670 == _T_146[11:0] ? image_1648 : _GEN_14002; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14004 = 12'h671 == _T_146[11:0] ? image_1649 : _GEN_14003; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14005 = 12'h672 == _T_146[11:0] ? image_1650 : _GEN_14004; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14006 = 12'h673 == _T_146[11:0] ? image_1651 : _GEN_14005; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14007 = 12'h674 == _T_146[11:0] ? image_1652 : _GEN_14006; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14008 = 12'h675 == _T_146[11:0] ? image_1653 : _GEN_14007; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14009 = 12'h676 == _T_146[11:0] ? image_1654 : _GEN_14008; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14010 = 12'h677 == _T_146[11:0] ? image_1655 : _GEN_14009; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14011 = 12'h678 == _T_146[11:0] ? image_1656 : _GEN_14010; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14012 = 12'h679 == _T_146[11:0] ? image_1657 : _GEN_14011; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14013 = 12'h67a == _T_146[11:0] ? image_1658 : _GEN_14012; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14014 = 12'h67b == _T_146[11:0] ? image_1659 : _GEN_14013; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14015 = 12'h67c == _T_146[11:0] ? image_1660 : _GEN_14014; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14016 = 12'h67d == _T_146[11:0] ? 4'h0 : _GEN_14015; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14017 = 12'h67e == _T_146[11:0] ? 4'h0 : _GEN_14016; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14018 = 12'h67f == _T_146[11:0] ? 4'h0 : _GEN_14017; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14019 = 12'h680 == _T_146[11:0] ? image_1664 : _GEN_14018; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14020 = 12'h681 == _T_146[11:0] ? image_1665 : _GEN_14019; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14021 = 12'h682 == _T_146[11:0] ? image_1666 : _GEN_14020; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14022 = 12'h683 == _T_146[11:0] ? image_1667 : _GEN_14021; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14023 = 12'h684 == _T_146[11:0] ? image_1668 : _GEN_14022; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14024 = 12'h685 == _T_146[11:0] ? image_1669 : _GEN_14023; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14025 = 12'h686 == _T_146[11:0] ? image_1670 : _GEN_14024; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14026 = 12'h687 == _T_146[11:0] ? image_1671 : _GEN_14025; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14027 = 12'h688 == _T_146[11:0] ? image_1672 : _GEN_14026; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14028 = 12'h689 == _T_146[11:0] ? image_1673 : _GEN_14027; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14029 = 12'h68a == _T_146[11:0] ? image_1674 : _GEN_14028; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14030 = 12'h68b == _T_146[11:0] ? image_1675 : _GEN_14029; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14031 = 12'h68c == _T_146[11:0] ? image_1676 : _GEN_14030; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14032 = 12'h68d == _T_146[11:0] ? image_1677 : _GEN_14031; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14033 = 12'h68e == _T_146[11:0] ? image_1678 : _GEN_14032; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14034 = 12'h68f == _T_146[11:0] ? image_1679 : _GEN_14033; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14035 = 12'h690 == _T_146[11:0] ? image_1680 : _GEN_14034; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14036 = 12'h691 == _T_146[11:0] ? image_1681 : _GEN_14035; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14037 = 12'h692 == _T_146[11:0] ? image_1682 : _GEN_14036; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14038 = 12'h693 == _T_146[11:0] ? image_1683 : _GEN_14037; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14039 = 12'h694 == _T_146[11:0] ? image_1684 : _GEN_14038; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14040 = 12'h695 == _T_146[11:0] ? image_1685 : _GEN_14039; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14041 = 12'h696 == _T_146[11:0] ? image_1686 : _GEN_14040; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14042 = 12'h697 == _T_146[11:0] ? image_1687 : _GEN_14041; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14043 = 12'h698 == _T_146[11:0] ? image_1688 : _GEN_14042; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14044 = 12'h699 == _T_146[11:0] ? image_1689 : _GEN_14043; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14045 = 12'h69a == _T_146[11:0] ? image_1690 : _GEN_14044; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14046 = 12'h69b == _T_146[11:0] ? image_1691 : _GEN_14045; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14047 = 12'h69c == _T_146[11:0] ? image_1692 : _GEN_14046; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14048 = 12'h69d == _T_146[11:0] ? image_1693 : _GEN_14047; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14049 = 12'h69e == _T_146[11:0] ? image_1694 : _GEN_14048; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14050 = 12'h69f == _T_146[11:0] ? image_1695 : _GEN_14049; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14051 = 12'h6a0 == _T_146[11:0] ? image_1696 : _GEN_14050; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14052 = 12'h6a1 == _T_146[11:0] ? image_1697 : _GEN_14051; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14053 = 12'h6a2 == _T_146[11:0] ? image_1698 : _GEN_14052; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14054 = 12'h6a3 == _T_146[11:0] ? image_1699 : _GEN_14053; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14055 = 12'h6a4 == _T_146[11:0] ? image_1700 : _GEN_14054; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14056 = 12'h6a5 == _T_146[11:0] ? image_1701 : _GEN_14055; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14057 = 12'h6a6 == _T_146[11:0] ? image_1702 : _GEN_14056; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14058 = 12'h6a7 == _T_146[11:0] ? image_1703 : _GEN_14057; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14059 = 12'h6a8 == _T_146[11:0] ? image_1704 : _GEN_14058; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14060 = 12'h6a9 == _T_146[11:0] ? image_1705 : _GEN_14059; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14061 = 12'h6aa == _T_146[11:0] ? image_1706 : _GEN_14060; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14062 = 12'h6ab == _T_146[11:0] ? image_1707 : _GEN_14061; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14063 = 12'h6ac == _T_146[11:0] ? image_1708 : _GEN_14062; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14064 = 12'h6ad == _T_146[11:0] ? image_1709 : _GEN_14063; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14065 = 12'h6ae == _T_146[11:0] ? image_1710 : _GEN_14064; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14066 = 12'h6af == _T_146[11:0] ? image_1711 : _GEN_14065; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14067 = 12'h6b0 == _T_146[11:0] ? image_1712 : _GEN_14066; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14068 = 12'h6b1 == _T_146[11:0] ? image_1713 : _GEN_14067; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14069 = 12'h6b2 == _T_146[11:0] ? image_1714 : _GEN_14068; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14070 = 12'h6b3 == _T_146[11:0] ? image_1715 : _GEN_14069; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14071 = 12'h6b4 == _T_146[11:0] ? image_1716 : _GEN_14070; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14072 = 12'h6b5 == _T_146[11:0] ? image_1717 : _GEN_14071; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14073 = 12'h6b6 == _T_146[11:0] ? image_1718 : _GEN_14072; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14074 = 12'h6b7 == _T_146[11:0] ? image_1719 : _GEN_14073; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14075 = 12'h6b8 == _T_146[11:0] ? image_1720 : _GEN_14074; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14076 = 12'h6b9 == _T_146[11:0] ? image_1721 : _GEN_14075; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14077 = 12'h6ba == _T_146[11:0] ? image_1722 : _GEN_14076; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14078 = 12'h6bb == _T_146[11:0] ? image_1723 : _GEN_14077; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14079 = 12'h6bc == _T_146[11:0] ? 4'h0 : _GEN_14078; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14080 = 12'h6bd == _T_146[11:0] ? 4'h0 : _GEN_14079; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14081 = 12'h6be == _T_146[11:0] ? 4'h0 : _GEN_14080; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14082 = 12'h6bf == _T_146[11:0] ? 4'h0 : _GEN_14081; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14083 = 12'h6c0 == _T_146[11:0] ? image_1728 : _GEN_14082; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14084 = 12'h6c1 == _T_146[11:0] ? image_1729 : _GEN_14083; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14085 = 12'h6c2 == _T_146[11:0] ? image_1730 : _GEN_14084; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14086 = 12'h6c3 == _T_146[11:0] ? image_1731 : _GEN_14085; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14087 = 12'h6c4 == _T_146[11:0] ? image_1732 : _GEN_14086; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14088 = 12'h6c5 == _T_146[11:0] ? image_1733 : _GEN_14087; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14089 = 12'h6c6 == _T_146[11:0] ? image_1734 : _GEN_14088; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14090 = 12'h6c7 == _T_146[11:0] ? image_1735 : _GEN_14089; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14091 = 12'h6c8 == _T_146[11:0] ? image_1736 : _GEN_14090; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14092 = 12'h6c9 == _T_146[11:0] ? image_1737 : _GEN_14091; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14093 = 12'h6ca == _T_146[11:0] ? image_1738 : _GEN_14092; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14094 = 12'h6cb == _T_146[11:0] ? image_1739 : _GEN_14093; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14095 = 12'h6cc == _T_146[11:0] ? image_1740 : _GEN_14094; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14096 = 12'h6cd == _T_146[11:0] ? image_1741 : _GEN_14095; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14097 = 12'h6ce == _T_146[11:0] ? image_1742 : _GEN_14096; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14098 = 12'h6cf == _T_146[11:0] ? image_1743 : _GEN_14097; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14099 = 12'h6d0 == _T_146[11:0] ? image_1744 : _GEN_14098; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14100 = 12'h6d1 == _T_146[11:0] ? image_1745 : _GEN_14099; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14101 = 12'h6d2 == _T_146[11:0] ? image_1746 : _GEN_14100; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14102 = 12'h6d3 == _T_146[11:0] ? image_1747 : _GEN_14101; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14103 = 12'h6d4 == _T_146[11:0] ? image_1748 : _GEN_14102; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14104 = 12'h6d5 == _T_146[11:0] ? image_1749 : _GEN_14103; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14105 = 12'h6d6 == _T_146[11:0] ? image_1750 : _GEN_14104; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14106 = 12'h6d7 == _T_146[11:0] ? image_1751 : _GEN_14105; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14107 = 12'h6d8 == _T_146[11:0] ? image_1752 : _GEN_14106; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14108 = 12'h6d9 == _T_146[11:0] ? image_1753 : _GEN_14107; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14109 = 12'h6da == _T_146[11:0] ? image_1754 : _GEN_14108; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14110 = 12'h6db == _T_146[11:0] ? image_1755 : _GEN_14109; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14111 = 12'h6dc == _T_146[11:0] ? image_1756 : _GEN_14110; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14112 = 12'h6dd == _T_146[11:0] ? image_1757 : _GEN_14111; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14113 = 12'h6de == _T_146[11:0] ? image_1758 : _GEN_14112; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14114 = 12'h6df == _T_146[11:0] ? image_1759 : _GEN_14113; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14115 = 12'h6e0 == _T_146[11:0] ? image_1760 : _GEN_14114; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14116 = 12'h6e1 == _T_146[11:0] ? image_1761 : _GEN_14115; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14117 = 12'h6e2 == _T_146[11:0] ? image_1762 : _GEN_14116; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14118 = 12'h6e3 == _T_146[11:0] ? image_1763 : _GEN_14117; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14119 = 12'h6e4 == _T_146[11:0] ? image_1764 : _GEN_14118; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14120 = 12'h6e5 == _T_146[11:0] ? image_1765 : _GEN_14119; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14121 = 12'h6e6 == _T_146[11:0] ? image_1766 : _GEN_14120; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14122 = 12'h6e7 == _T_146[11:0] ? image_1767 : _GEN_14121; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14123 = 12'h6e8 == _T_146[11:0] ? image_1768 : _GEN_14122; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14124 = 12'h6e9 == _T_146[11:0] ? image_1769 : _GEN_14123; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14125 = 12'h6ea == _T_146[11:0] ? image_1770 : _GEN_14124; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14126 = 12'h6eb == _T_146[11:0] ? image_1771 : _GEN_14125; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14127 = 12'h6ec == _T_146[11:0] ? image_1772 : _GEN_14126; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14128 = 12'h6ed == _T_146[11:0] ? image_1773 : _GEN_14127; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14129 = 12'h6ee == _T_146[11:0] ? image_1774 : _GEN_14128; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14130 = 12'h6ef == _T_146[11:0] ? image_1775 : _GEN_14129; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14131 = 12'h6f0 == _T_146[11:0] ? image_1776 : _GEN_14130; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14132 = 12'h6f1 == _T_146[11:0] ? image_1777 : _GEN_14131; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14133 = 12'h6f2 == _T_146[11:0] ? image_1778 : _GEN_14132; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14134 = 12'h6f3 == _T_146[11:0] ? image_1779 : _GEN_14133; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14135 = 12'h6f4 == _T_146[11:0] ? image_1780 : _GEN_14134; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14136 = 12'h6f5 == _T_146[11:0] ? image_1781 : _GEN_14135; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14137 = 12'h6f6 == _T_146[11:0] ? image_1782 : _GEN_14136; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14138 = 12'h6f7 == _T_146[11:0] ? image_1783 : _GEN_14137; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14139 = 12'h6f8 == _T_146[11:0] ? image_1784 : _GEN_14138; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14140 = 12'h6f9 == _T_146[11:0] ? image_1785 : _GEN_14139; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14141 = 12'h6fa == _T_146[11:0] ? image_1786 : _GEN_14140; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14142 = 12'h6fb == _T_146[11:0] ? 4'h0 : _GEN_14141; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14143 = 12'h6fc == _T_146[11:0] ? 4'h0 : _GEN_14142; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14144 = 12'h6fd == _T_146[11:0] ? 4'h0 : _GEN_14143; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14145 = 12'h6fe == _T_146[11:0] ? 4'h0 : _GEN_14144; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14146 = 12'h6ff == _T_146[11:0] ? 4'h0 : _GEN_14145; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14147 = 12'h700 == _T_146[11:0] ? 4'h0 : _GEN_14146; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14148 = 12'h701 == _T_146[11:0] ? image_1793 : _GEN_14147; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14149 = 12'h702 == _T_146[11:0] ? image_1794 : _GEN_14148; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14150 = 12'h703 == _T_146[11:0] ? image_1795 : _GEN_14149; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14151 = 12'h704 == _T_146[11:0] ? image_1796 : _GEN_14150; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14152 = 12'h705 == _T_146[11:0] ? image_1797 : _GEN_14151; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14153 = 12'h706 == _T_146[11:0] ? image_1798 : _GEN_14152; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14154 = 12'h707 == _T_146[11:0] ? image_1799 : _GEN_14153; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14155 = 12'h708 == _T_146[11:0] ? image_1800 : _GEN_14154; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14156 = 12'h709 == _T_146[11:0] ? image_1801 : _GEN_14155; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14157 = 12'h70a == _T_146[11:0] ? image_1802 : _GEN_14156; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14158 = 12'h70b == _T_146[11:0] ? image_1803 : _GEN_14157; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14159 = 12'h70c == _T_146[11:0] ? image_1804 : _GEN_14158; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14160 = 12'h70d == _T_146[11:0] ? image_1805 : _GEN_14159; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14161 = 12'h70e == _T_146[11:0] ? image_1806 : _GEN_14160; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14162 = 12'h70f == _T_146[11:0] ? image_1807 : _GEN_14161; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14163 = 12'h710 == _T_146[11:0] ? image_1808 : _GEN_14162; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14164 = 12'h711 == _T_146[11:0] ? image_1809 : _GEN_14163; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14165 = 12'h712 == _T_146[11:0] ? image_1810 : _GEN_14164; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14166 = 12'h713 == _T_146[11:0] ? image_1811 : _GEN_14165; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14167 = 12'h714 == _T_146[11:0] ? image_1812 : _GEN_14166; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14168 = 12'h715 == _T_146[11:0] ? image_1813 : _GEN_14167; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14169 = 12'h716 == _T_146[11:0] ? image_1814 : _GEN_14168; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14170 = 12'h717 == _T_146[11:0] ? image_1815 : _GEN_14169; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14171 = 12'h718 == _T_146[11:0] ? image_1816 : _GEN_14170; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14172 = 12'h719 == _T_146[11:0] ? image_1817 : _GEN_14171; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14173 = 12'h71a == _T_146[11:0] ? image_1818 : _GEN_14172; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14174 = 12'h71b == _T_146[11:0] ? image_1819 : _GEN_14173; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14175 = 12'h71c == _T_146[11:0] ? image_1820 : _GEN_14174; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14176 = 12'h71d == _T_146[11:0] ? image_1821 : _GEN_14175; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14177 = 12'h71e == _T_146[11:0] ? image_1822 : _GEN_14176; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14178 = 12'h71f == _T_146[11:0] ? image_1823 : _GEN_14177; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14179 = 12'h720 == _T_146[11:0] ? image_1824 : _GEN_14178; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14180 = 12'h721 == _T_146[11:0] ? image_1825 : _GEN_14179; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14181 = 12'h722 == _T_146[11:0] ? image_1826 : _GEN_14180; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14182 = 12'h723 == _T_146[11:0] ? image_1827 : _GEN_14181; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14183 = 12'h724 == _T_146[11:0] ? image_1828 : _GEN_14182; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14184 = 12'h725 == _T_146[11:0] ? image_1829 : _GEN_14183; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14185 = 12'h726 == _T_146[11:0] ? image_1830 : _GEN_14184; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14186 = 12'h727 == _T_146[11:0] ? image_1831 : _GEN_14185; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14187 = 12'h728 == _T_146[11:0] ? image_1832 : _GEN_14186; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14188 = 12'h729 == _T_146[11:0] ? image_1833 : _GEN_14187; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14189 = 12'h72a == _T_146[11:0] ? image_1834 : _GEN_14188; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14190 = 12'h72b == _T_146[11:0] ? image_1835 : _GEN_14189; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14191 = 12'h72c == _T_146[11:0] ? image_1836 : _GEN_14190; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14192 = 12'h72d == _T_146[11:0] ? image_1837 : _GEN_14191; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14193 = 12'h72e == _T_146[11:0] ? image_1838 : _GEN_14192; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14194 = 12'h72f == _T_146[11:0] ? image_1839 : _GEN_14193; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14195 = 12'h730 == _T_146[11:0] ? image_1840 : _GEN_14194; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14196 = 12'h731 == _T_146[11:0] ? image_1841 : _GEN_14195; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14197 = 12'h732 == _T_146[11:0] ? image_1842 : _GEN_14196; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14198 = 12'h733 == _T_146[11:0] ? image_1843 : _GEN_14197; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14199 = 12'h734 == _T_146[11:0] ? image_1844 : _GEN_14198; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14200 = 12'h735 == _T_146[11:0] ? image_1845 : _GEN_14199; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14201 = 12'h736 == _T_146[11:0] ? image_1846 : _GEN_14200; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14202 = 12'h737 == _T_146[11:0] ? image_1847 : _GEN_14201; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14203 = 12'h738 == _T_146[11:0] ? image_1848 : _GEN_14202; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14204 = 12'h739 == _T_146[11:0] ? image_1849 : _GEN_14203; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14205 = 12'h73a == _T_146[11:0] ? 4'h0 : _GEN_14204; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14206 = 12'h73b == _T_146[11:0] ? 4'h0 : _GEN_14205; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14207 = 12'h73c == _T_146[11:0] ? 4'h0 : _GEN_14206; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14208 = 12'h73d == _T_146[11:0] ? 4'h0 : _GEN_14207; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14209 = 12'h73e == _T_146[11:0] ? 4'h0 : _GEN_14208; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14210 = 12'h73f == _T_146[11:0] ? 4'h0 : _GEN_14209; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14211 = 12'h740 == _T_146[11:0] ? 4'h0 : _GEN_14210; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14212 = 12'h741 == _T_146[11:0] ? image_1857 : _GEN_14211; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14213 = 12'h742 == _T_146[11:0] ? image_1858 : _GEN_14212; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14214 = 12'h743 == _T_146[11:0] ? image_1859 : _GEN_14213; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14215 = 12'h744 == _T_146[11:0] ? image_1860 : _GEN_14214; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14216 = 12'h745 == _T_146[11:0] ? image_1861 : _GEN_14215; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14217 = 12'h746 == _T_146[11:0] ? image_1862 : _GEN_14216; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14218 = 12'h747 == _T_146[11:0] ? image_1863 : _GEN_14217; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14219 = 12'h748 == _T_146[11:0] ? image_1864 : _GEN_14218; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14220 = 12'h749 == _T_146[11:0] ? image_1865 : _GEN_14219; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14221 = 12'h74a == _T_146[11:0] ? image_1866 : _GEN_14220; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14222 = 12'h74b == _T_146[11:0] ? image_1867 : _GEN_14221; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14223 = 12'h74c == _T_146[11:0] ? image_1868 : _GEN_14222; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14224 = 12'h74d == _T_146[11:0] ? image_1869 : _GEN_14223; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14225 = 12'h74e == _T_146[11:0] ? image_1870 : _GEN_14224; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14226 = 12'h74f == _T_146[11:0] ? image_1871 : _GEN_14225; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14227 = 12'h750 == _T_146[11:0] ? image_1872 : _GEN_14226; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14228 = 12'h751 == _T_146[11:0] ? image_1873 : _GEN_14227; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14229 = 12'h752 == _T_146[11:0] ? image_1874 : _GEN_14228; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14230 = 12'h753 == _T_146[11:0] ? image_1875 : _GEN_14229; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14231 = 12'h754 == _T_146[11:0] ? image_1876 : _GEN_14230; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14232 = 12'h755 == _T_146[11:0] ? image_1877 : _GEN_14231; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14233 = 12'h756 == _T_146[11:0] ? image_1878 : _GEN_14232; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14234 = 12'h757 == _T_146[11:0] ? image_1879 : _GEN_14233; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14235 = 12'h758 == _T_146[11:0] ? image_1880 : _GEN_14234; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14236 = 12'h759 == _T_146[11:0] ? image_1881 : _GEN_14235; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14237 = 12'h75a == _T_146[11:0] ? image_1882 : _GEN_14236; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14238 = 12'h75b == _T_146[11:0] ? image_1883 : _GEN_14237; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14239 = 12'h75c == _T_146[11:0] ? image_1884 : _GEN_14238; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14240 = 12'h75d == _T_146[11:0] ? image_1885 : _GEN_14239; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14241 = 12'h75e == _T_146[11:0] ? image_1886 : _GEN_14240; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14242 = 12'h75f == _T_146[11:0] ? image_1887 : _GEN_14241; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14243 = 12'h760 == _T_146[11:0] ? image_1888 : _GEN_14242; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14244 = 12'h761 == _T_146[11:0] ? image_1889 : _GEN_14243; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14245 = 12'h762 == _T_146[11:0] ? image_1890 : _GEN_14244; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14246 = 12'h763 == _T_146[11:0] ? image_1891 : _GEN_14245; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14247 = 12'h764 == _T_146[11:0] ? image_1892 : _GEN_14246; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14248 = 12'h765 == _T_146[11:0] ? image_1893 : _GEN_14247; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14249 = 12'h766 == _T_146[11:0] ? image_1894 : _GEN_14248; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14250 = 12'h767 == _T_146[11:0] ? image_1895 : _GEN_14249; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14251 = 12'h768 == _T_146[11:0] ? image_1896 : _GEN_14250; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14252 = 12'h769 == _T_146[11:0] ? image_1897 : _GEN_14251; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14253 = 12'h76a == _T_146[11:0] ? image_1898 : _GEN_14252; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14254 = 12'h76b == _T_146[11:0] ? image_1899 : _GEN_14253; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14255 = 12'h76c == _T_146[11:0] ? image_1900 : _GEN_14254; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14256 = 12'h76d == _T_146[11:0] ? image_1901 : _GEN_14255; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14257 = 12'h76e == _T_146[11:0] ? image_1902 : _GEN_14256; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14258 = 12'h76f == _T_146[11:0] ? image_1903 : _GEN_14257; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14259 = 12'h770 == _T_146[11:0] ? image_1904 : _GEN_14258; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14260 = 12'h771 == _T_146[11:0] ? image_1905 : _GEN_14259; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14261 = 12'h772 == _T_146[11:0] ? image_1906 : _GEN_14260; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14262 = 12'h773 == _T_146[11:0] ? image_1907 : _GEN_14261; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14263 = 12'h774 == _T_146[11:0] ? image_1908 : _GEN_14262; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14264 = 12'h775 == _T_146[11:0] ? image_1909 : _GEN_14263; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14265 = 12'h776 == _T_146[11:0] ? image_1910 : _GEN_14264; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14266 = 12'h777 == _T_146[11:0] ? image_1911 : _GEN_14265; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14267 = 12'h778 == _T_146[11:0] ? image_1912 : _GEN_14266; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14268 = 12'h779 == _T_146[11:0] ? image_1913 : _GEN_14267; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14269 = 12'h77a == _T_146[11:0] ? 4'h0 : _GEN_14268; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14270 = 12'h77b == _T_146[11:0] ? 4'h0 : _GEN_14269; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14271 = 12'h77c == _T_146[11:0] ? 4'h0 : _GEN_14270; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14272 = 12'h77d == _T_146[11:0] ? 4'h0 : _GEN_14271; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14273 = 12'h77e == _T_146[11:0] ? 4'h0 : _GEN_14272; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14274 = 12'h77f == _T_146[11:0] ? 4'h0 : _GEN_14273; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14275 = 12'h780 == _T_146[11:0] ? 4'h0 : _GEN_14274; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14276 = 12'h781 == _T_146[11:0] ? image_1921 : _GEN_14275; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14277 = 12'h782 == _T_146[11:0] ? image_1922 : _GEN_14276; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14278 = 12'h783 == _T_146[11:0] ? image_1923 : _GEN_14277; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14279 = 12'h784 == _T_146[11:0] ? image_1924 : _GEN_14278; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14280 = 12'h785 == _T_146[11:0] ? image_1925 : _GEN_14279; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14281 = 12'h786 == _T_146[11:0] ? image_1926 : _GEN_14280; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14282 = 12'h787 == _T_146[11:0] ? image_1927 : _GEN_14281; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14283 = 12'h788 == _T_146[11:0] ? image_1928 : _GEN_14282; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14284 = 12'h789 == _T_146[11:0] ? image_1929 : _GEN_14283; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14285 = 12'h78a == _T_146[11:0] ? image_1930 : _GEN_14284; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14286 = 12'h78b == _T_146[11:0] ? image_1931 : _GEN_14285; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14287 = 12'h78c == _T_146[11:0] ? image_1932 : _GEN_14286; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14288 = 12'h78d == _T_146[11:0] ? image_1933 : _GEN_14287; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14289 = 12'h78e == _T_146[11:0] ? image_1934 : _GEN_14288; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14290 = 12'h78f == _T_146[11:0] ? image_1935 : _GEN_14289; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14291 = 12'h790 == _T_146[11:0] ? image_1936 : _GEN_14290; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14292 = 12'h791 == _T_146[11:0] ? image_1937 : _GEN_14291; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14293 = 12'h792 == _T_146[11:0] ? image_1938 : _GEN_14292; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14294 = 12'h793 == _T_146[11:0] ? image_1939 : _GEN_14293; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14295 = 12'h794 == _T_146[11:0] ? image_1940 : _GEN_14294; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14296 = 12'h795 == _T_146[11:0] ? image_1941 : _GEN_14295; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14297 = 12'h796 == _T_146[11:0] ? image_1942 : _GEN_14296; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14298 = 12'h797 == _T_146[11:0] ? image_1943 : _GEN_14297; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14299 = 12'h798 == _T_146[11:0] ? image_1944 : _GEN_14298; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14300 = 12'h799 == _T_146[11:0] ? image_1945 : _GEN_14299; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14301 = 12'h79a == _T_146[11:0] ? image_1946 : _GEN_14300; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14302 = 12'h79b == _T_146[11:0] ? image_1947 : _GEN_14301; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14303 = 12'h79c == _T_146[11:0] ? image_1948 : _GEN_14302; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14304 = 12'h79d == _T_146[11:0] ? image_1949 : _GEN_14303; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14305 = 12'h79e == _T_146[11:0] ? image_1950 : _GEN_14304; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14306 = 12'h79f == _T_146[11:0] ? image_1951 : _GEN_14305; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14307 = 12'h7a0 == _T_146[11:0] ? image_1952 : _GEN_14306; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14308 = 12'h7a1 == _T_146[11:0] ? image_1953 : _GEN_14307; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14309 = 12'h7a2 == _T_146[11:0] ? image_1954 : _GEN_14308; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14310 = 12'h7a3 == _T_146[11:0] ? image_1955 : _GEN_14309; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14311 = 12'h7a4 == _T_146[11:0] ? image_1956 : _GEN_14310; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14312 = 12'h7a5 == _T_146[11:0] ? image_1957 : _GEN_14311; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14313 = 12'h7a6 == _T_146[11:0] ? image_1958 : _GEN_14312; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14314 = 12'h7a7 == _T_146[11:0] ? image_1959 : _GEN_14313; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14315 = 12'h7a8 == _T_146[11:0] ? image_1960 : _GEN_14314; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14316 = 12'h7a9 == _T_146[11:0] ? image_1961 : _GEN_14315; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14317 = 12'h7aa == _T_146[11:0] ? image_1962 : _GEN_14316; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14318 = 12'h7ab == _T_146[11:0] ? image_1963 : _GEN_14317; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14319 = 12'h7ac == _T_146[11:0] ? image_1964 : _GEN_14318; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14320 = 12'h7ad == _T_146[11:0] ? image_1965 : _GEN_14319; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14321 = 12'h7ae == _T_146[11:0] ? image_1966 : _GEN_14320; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14322 = 12'h7af == _T_146[11:0] ? image_1967 : _GEN_14321; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14323 = 12'h7b0 == _T_146[11:0] ? image_1968 : _GEN_14322; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14324 = 12'h7b1 == _T_146[11:0] ? image_1969 : _GEN_14323; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14325 = 12'h7b2 == _T_146[11:0] ? image_1970 : _GEN_14324; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14326 = 12'h7b3 == _T_146[11:0] ? image_1971 : _GEN_14325; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14327 = 12'h7b4 == _T_146[11:0] ? image_1972 : _GEN_14326; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14328 = 12'h7b5 == _T_146[11:0] ? image_1973 : _GEN_14327; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14329 = 12'h7b6 == _T_146[11:0] ? image_1974 : _GEN_14328; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14330 = 12'h7b7 == _T_146[11:0] ? image_1975 : _GEN_14329; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14331 = 12'h7b8 == _T_146[11:0] ? image_1976 : _GEN_14330; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14332 = 12'h7b9 == _T_146[11:0] ? image_1977 : _GEN_14331; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14333 = 12'h7ba == _T_146[11:0] ? 4'h0 : _GEN_14332; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14334 = 12'h7bb == _T_146[11:0] ? 4'h0 : _GEN_14333; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14335 = 12'h7bc == _T_146[11:0] ? 4'h0 : _GEN_14334; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14336 = 12'h7bd == _T_146[11:0] ? 4'h0 : _GEN_14335; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14337 = 12'h7be == _T_146[11:0] ? 4'h0 : _GEN_14336; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14338 = 12'h7bf == _T_146[11:0] ? 4'h0 : _GEN_14337; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14339 = 12'h7c0 == _T_146[11:0] ? 4'h0 : _GEN_14338; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14340 = 12'h7c1 == _T_146[11:0] ? image_1985 : _GEN_14339; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14341 = 12'h7c2 == _T_146[11:0] ? image_1986 : _GEN_14340; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14342 = 12'h7c3 == _T_146[11:0] ? image_1987 : _GEN_14341; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14343 = 12'h7c4 == _T_146[11:0] ? image_1988 : _GEN_14342; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14344 = 12'h7c5 == _T_146[11:0] ? image_1989 : _GEN_14343; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14345 = 12'h7c6 == _T_146[11:0] ? image_1990 : _GEN_14344; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14346 = 12'h7c7 == _T_146[11:0] ? image_1991 : _GEN_14345; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14347 = 12'h7c8 == _T_146[11:0] ? image_1992 : _GEN_14346; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14348 = 12'h7c9 == _T_146[11:0] ? image_1993 : _GEN_14347; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14349 = 12'h7ca == _T_146[11:0] ? image_1994 : _GEN_14348; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14350 = 12'h7cb == _T_146[11:0] ? image_1995 : _GEN_14349; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14351 = 12'h7cc == _T_146[11:0] ? image_1996 : _GEN_14350; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14352 = 12'h7cd == _T_146[11:0] ? image_1997 : _GEN_14351; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14353 = 12'h7ce == _T_146[11:0] ? image_1998 : _GEN_14352; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14354 = 12'h7cf == _T_146[11:0] ? image_1999 : _GEN_14353; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14355 = 12'h7d0 == _T_146[11:0] ? image_2000 : _GEN_14354; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14356 = 12'h7d1 == _T_146[11:0] ? image_2001 : _GEN_14355; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14357 = 12'h7d2 == _T_146[11:0] ? image_2002 : _GEN_14356; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14358 = 12'h7d3 == _T_146[11:0] ? image_2003 : _GEN_14357; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14359 = 12'h7d4 == _T_146[11:0] ? image_2004 : _GEN_14358; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14360 = 12'h7d5 == _T_146[11:0] ? image_2005 : _GEN_14359; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14361 = 12'h7d6 == _T_146[11:0] ? image_2006 : _GEN_14360; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14362 = 12'h7d7 == _T_146[11:0] ? image_2007 : _GEN_14361; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14363 = 12'h7d8 == _T_146[11:0] ? image_2008 : _GEN_14362; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14364 = 12'h7d9 == _T_146[11:0] ? image_2009 : _GEN_14363; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14365 = 12'h7da == _T_146[11:0] ? image_2010 : _GEN_14364; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14366 = 12'h7db == _T_146[11:0] ? image_2011 : _GEN_14365; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14367 = 12'h7dc == _T_146[11:0] ? image_2012 : _GEN_14366; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14368 = 12'h7dd == _T_146[11:0] ? image_2013 : _GEN_14367; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14369 = 12'h7de == _T_146[11:0] ? image_2014 : _GEN_14368; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14370 = 12'h7df == _T_146[11:0] ? image_2015 : _GEN_14369; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14371 = 12'h7e0 == _T_146[11:0] ? image_2016 : _GEN_14370; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14372 = 12'h7e1 == _T_146[11:0] ? image_2017 : _GEN_14371; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14373 = 12'h7e2 == _T_146[11:0] ? image_2018 : _GEN_14372; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14374 = 12'h7e3 == _T_146[11:0] ? image_2019 : _GEN_14373; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14375 = 12'h7e4 == _T_146[11:0] ? image_2020 : _GEN_14374; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14376 = 12'h7e5 == _T_146[11:0] ? image_2021 : _GEN_14375; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14377 = 12'h7e6 == _T_146[11:0] ? image_2022 : _GEN_14376; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14378 = 12'h7e7 == _T_146[11:0] ? image_2023 : _GEN_14377; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14379 = 12'h7e8 == _T_146[11:0] ? image_2024 : _GEN_14378; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14380 = 12'h7e9 == _T_146[11:0] ? image_2025 : _GEN_14379; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14381 = 12'h7ea == _T_146[11:0] ? image_2026 : _GEN_14380; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14382 = 12'h7eb == _T_146[11:0] ? image_2027 : _GEN_14381; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14383 = 12'h7ec == _T_146[11:0] ? image_2028 : _GEN_14382; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14384 = 12'h7ed == _T_146[11:0] ? image_2029 : _GEN_14383; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14385 = 12'h7ee == _T_146[11:0] ? image_2030 : _GEN_14384; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14386 = 12'h7ef == _T_146[11:0] ? image_2031 : _GEN_14385; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14387 = 12'h7f0 == _T_146[11:0] ? image_2032 : _GEN_14386; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14388 = 12'h7f1 == _T_146[11:0] ? image_2033 : _GEN_14387; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14389 = 12'h7f2 == _T_146[11:0] ? image_2034 : _GEN_14388; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14390 = 12'h7f3 == _T_146[11:0] ? image_2035 : _GEN_14389; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14391 = 12'h7f4 == _T_146[11:0] ? image_2036 : _GEN_14390; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14392 = 12'h7f5 == _T_146[11:0] ? image_2037 : _GEN_14391; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14393 = 12'h7f6 == _T_146[11:0] ? image_2038 : _GEN_14392; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14394 = 12'h7f7 == _T_146[11:0] ? image_2039 : _GEN_14393; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14395 = 12'h7f8 == _T_146[11:0] ? image_2040 : _GEN_14394; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14396 = 12'h7f9 == _T_146[11:0] ? image_2041 : _GEN_14395; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14397 = 12'h7fa == _T_146[11:0] ? 4'h0 : _GEN_14396; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14398 = 12'h7fb == _T_146[11:0] ? 4'h0 : _GEN_14397; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14399 = 12'h7fc == _T_146[11:0] ? 4'h0 : _GEN_14398; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14400 = 12'h7fd == _T_146[11:0] ? 4'h0 : _GEN_14399; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14401 = 12'h7fe == _T_146[11:0] ? 4'h0 : _GEN_14400; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14402 = 12'h7ff == _T_146[11:0] ? 4'h0 : _GEN_14401; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14403 = 12'h800 == _T_146[11:0] ? 4'h0 : _GEN_14402; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14404 = 12'h801 == _T_146[11:0] ? image_2049 : _GEN_14403; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14405 = 12'h802 == _T_146[11:0] ? image_2050 : _GEN_14404; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14406 = 12'h803 == _T_146[11:0] ? image_2051 : _GEN_14405; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14407 = 12'h804 == _T_146[11:0] ? image_2052 : _GEN_14406; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14408 = 12'h805 == _T_146[11:0] ? image_2053 : _GEN_14407; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14409 = 12'h806 == _T_146[11:0] ? image_2054 : _GEN_14408; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14410 = 12'h807 == _T_146[11:0] ? image_2055 : _GEN_14409; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14411 = 12'h808 == _T_146[11:0] ? image_2056 : _GEN_14410; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14412 = 12'h809 == _T_146[11:0] ? image_2057 : _GEN_14411; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14413 = 12'h80a == _T_146[11:0] ? image_2058 : _GEN_14412; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14414 = 12'h80b == _T_146[11:0] ? image_2059 : _GEN_14413; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14415 = 12'h80c == _T_146[11:0] ? image_2060 : _GEN_14414; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14416 = 12'h80d == _T_146[11:0] ? image_2061 : _GEN_14415; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14417 = 12'h80e == _T_146[11:0] ? image_2062 : _GEN_14416; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14418 = 12'h80f == _T_146[11:0] ? image_2063 : _GEN_14417; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14419 = 12'h810 == _T_146[11:0] ? image_2064 : _GEN_14418; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14420 = 12'h811 == _T_146[11:0] ? image_2065 : _GEN_14419; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14421 = 12'h812 == _T_146[11:0] ? image_2066 : _GEN_14420; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14422 = 12'h813 == _T_146[11:0] ? image_2067 : _GEN_14421; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14423 = 12'h814 == _T_146[11:0] ? image_2068 : _GEN_14422; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14424 = 12'h815 == _T_146[11:0] ? image_2069 : _GEN_14423; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14425 = 12'h816 == _T_146[11:0] ? image_2070 : _GEN_14424; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14426 = 12'h817 == _T_146[11:0] ? image_2071 : _GEN_14425; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14427 = 12'h818 == _T_146[11:0] ? image_2072 : _GEN_14426; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14428 = 12'h819 == _T_146[11:0] ? image_2073 : _GEN_14427; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14429 = 12'h81a == _T_146[11:0] ? image_2074 : _GEN_14428; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14430 = 12'h81b == _T_146[11:0] ? image_2075 : _GEN_14429; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14431 = 12'h81c == _T_146[11:0] ? image_2076 : _GEN_14430; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14432 = 12'h81d == _T_146[11:0] ? image_2077 : _GEN_14431; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14433 = 12'h81e == _T_146[11:0] ? image_2078 : _GEN_14432; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14434 = 12'h81f == _T_146[11:0] ? image_2079 : _GEN_14433; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14435 = 12'h820 == _T_146[11:0] ? image_2080 : _GEN_14434; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14436 = 12'h821 == _T_146[11:0] ? image_2081 : _GEN_14435; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14437 = 12'h822 == _T_146[11:0] ? image_2082 : _GEN_14436; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14438 = 12'h823 == _T_146[11:0] ? image_2083 : _GEN_14437; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14439 = 12'h824 == _T_146[11:0] ? image_2084 : _GEN_14438; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14440 = 12'h825 == _T_146[11:0] ? image_2085 : _GEN_14439; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14441 = 12'h826 == _T_146[11:0] ? image_2086 : _GEN_14440; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14442 = 12'h827 == _T_146[11:0] ? image_2087 : _GEN_14441; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14443 = 12'h828 == _T_146[11:0] ? image_2088 : _GEN_14442; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14444 = 12'h829 == _T_146[11:0] ? image_2089 : _GEN_14443; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14445 = 12'h82a == _T_146[11:0] ? image_2090 : _GEN_14444; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14446 = 12'h82b == _T_146[11:0] ? image_2091 : _GEN_14445; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14447 = 12'h82c == _T_146[11:0] ? image_2092 : _GEN_14446; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14448 = 12'h82d == _T_146[11:0] ? image_2093 : _GEN_14447; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14449 = 12'h82e == _T_146[11:0] ? image_2094 : _GEN_14448; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14450 = 12'h82f == _T_146[11:0] ? image_2095 : _GEN_14449; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14451 = 12'h830 == _T_146[11:0] ? image_2096 : _GEN_14450; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14452 = 12'h831 == _T_146[11:0] ? image_2097 : _GEN_14451; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14453 = 12'h832 == _T_146[11:0] ? image_2098 : _GEN_14452; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14454 = 12'h833 == _T_146[11:0] ? image_2099 : _GEN_14453; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14455 = 12'h834 == _T_146[11:0] ? image_2100 : _GEN_14454; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14456 = 12'h835 == _T_146[11:0] ? image_2101 : _GEN_14455; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14457 = 12'h836 == _T_146[11:0] ? image_2102 : _GEN_14456; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14458 = 12'h837 == _T_146[11:0] ? image_2103 : _GEN_14457; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14459 = 12'h838 == _T_146[11:0] ? image_2104 : _GEN_14458; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14460 = 12'h839 == _T_146[11:0] ? image_2105 : _GEN_14459; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14461 = 12'h83a == _T_146[11:0] ? image_2106 : _GEN_14460; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14462 = 12'h83b == _T_146[11:0] ? 4'h0 : _GEN_14461; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14463 = 12'h83c == _T_146[11:0] ? 4'h0 : _GEN_14462; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14464 = 12'h83d == _T_146[11:0] ? 4'h0 : _GEN_14463; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14465 = 12'h83e == _T_146[11:0] ? 4'h0 : _GEN_14464; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14466 = 12'h83f == _T_146[11:0] ? 4'h0 : _GEN_14465; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14467 = 12'h840 == _T_146[11:0] ? 4'h0 : _GEN_14466; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14468 = 12'h841 == _T_146[11:0] ? 4'h0 : _GEN_14467; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14469 = 12'h842 == _T_146[11:0] ? image_2114 : _GEN_14468; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14470 = 12'h843 == _T_146[11:0] ? image_2115 : _GEN_14469; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14471 = 12'h844 == _T_146[11:0] ? image_2116 : _GEN_14470; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14472 = 12'h845 == _T_146[11:0] ? image_2117 : _GEN_14471; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14473 = 12'h846 == _T_146[11:0] ? image_2118 : _GEN_14472; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14474 = 12'h847 == _T_146[11:0] ? image_2119 : _GEN_14473; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14475 = 12'h848 == _T_146[11:0] ? image_2120 : _GEN_14474; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14476 = 12'h849 == _T_146[11:0] ? image_2121 : _GEN_14475; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14477 = 12'h84a == _T_146[11:0] ? image_2122 : _GEN_14476; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14478 = 12'h84b == _T_146[11:0] ? image_2123 : _GEN_14477; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14479 = 12'h84c == _T_146[11:0] ? image_2124 : _GEN_14478; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14480 = 12'h84d == _T_146[11:0] ? image_2125 : _GEN_14479; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14481 = 12'h84e == _T_146[11:0] ? image_2126 : _GEN_14480; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14482 = 12'h84f == _T_146[11:0] ? image_2127 : _GEN_14481; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14483 = 12'h850 == _T_146[11:0] ? image_2128 : _GEN_14482; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14484 = 12'h851 == _T_146[11:0] ? image_2129 : _GEN_14483; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14485 = 12'h852 == _T_146[11:0] ? image_2130 : _GEN_14484; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14486 = 12'h853 == _T_146[11:0] ? image_2131 : _GEN_14485; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14487 = 12'h854 == _T_146[11:0] ? image_2132 : _GEN_14486; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14488 = 12'h855 == _T_146[11:0] ? image_2133 : _GEN_14487; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14489 = 12'h856 == _T_146[11:0] ? image_2134 : _GEN_14488; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14490 = 12'h857 == _T_146[11:0] ? image_2135 : _GEN_14489; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14491 = 12'h858 == _T_146[11:0] ? image_2136 : _GEN_14490; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14492 = 12'h859 == _T_146[11:0] ? image_2137 : _GEN_14491; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14493 = 12'h85a == _T_146[11:0] ? image_2138 : _GEN_14492; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14494 = 12'h85b == _T_146[11:0] ? image_2139 : _GEN_14493; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14495 = 12'h85c == _T_146[11:0] ? image_2140 : _GEN_14494; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14496 = 12'h85d == _T_146[11:0] ? image_2141 : _GEN_14495; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14497 = 12'h85e == _T_146[11:0] ? image_2142 : _GEN_14496; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14498 = 12'h85f == _T_146[11:0] ? image_2143 : _GEN_14497; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14499 = 12'h860 == _T_146[11:0] ? image_2144 : _GEN_14498; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14500 = 12'h861 == _T_146[11:0] ? image_2145 : _GEN_14499; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14501 = 12'h862 == _T_146[11:0] ? image_2146 : _GEN_14500; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14502 = 12'h863 == _T_146[11:0] ? image_2147 : _GEN_14501; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14503 = 12'h864 == _T_146[11:0] ? image_2148 : _GEN_14502; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14504 = 12'h865 == _T_146[11:0] ? image_2149 : _GEN_14503; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14505 = 12'h866 == _T_146[11:0] ? image_2150 : _GEN_14504; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14506 = 12'h867 == _T_146[11:0] ? image_2151 : _GEN_14505; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14507 = 12'h868 == _T_146[11:0] ? image_2152 : _GEN_14506; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14508 = 12'h869 == _T_146[11:0] ? image_2153 : _GEN_14507; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14509 = 12'h86a == _T_146[11:0] ? image_2154 : _GEN_14508; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14510 = 12'h86b == _T_146[11:0] ? image_2155 : _GEN_14509; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14511 = 12'h86c == _T_146[11:0] ? image_2156 : _GEN_14510; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14512 = 12'h86d == _T_146[11:0] ? image_2157 : _GEN_14511; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14513 = 12'h86e == _T_146[11:0] ? image_2158 : _GEN_14512; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14514 = 12'h86f == _T_146[11:0] ? image_2159 : _GEN_14513; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14515 = 12'h870 == _T_146[11:0] ? image_2160 : _GEN_14514; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14516 = 12'h871 == _T_146[11:0] ? image_2161 : _GEN_14515; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14517 = 12'h872 == _T_146[11:0] ? image_2162 : _GEN_14516; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14518 = 12'h873 == _T_146[11:0] ? image_2163 : _GEN_14517; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14519 = 12'h874 == _T_146[11:0] ? image_2164 : _GEN_14518; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14520 = 12'h875 == _T_146[11:0] ? image_2165 : _GEN_14519; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14521 = 12'h876 == _T_146[11:0] ? image_2166 : _GEN_14520; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14522 = 12'h877 == _T_146[11:0] ? image_2167 : _GEN_14521; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14523 = 12'h878 == _T_146[11:0] ? image_2168 : _GEN_14522; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14524 = 12'h879 == _T_146[11:0] ? image_2169 : _GEN_14523; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14525 = 12'h87a == _T_146[11:0] ? image_2170 : _GEN_14524; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14526 = 12'h87b == _T_146[11:0] ? 4'h0 : _GEN_14525; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14527 = 12'h87c == _T_146[11:0] ? 4'h0 : _GEN_14526; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14528 = 12'h87d == _T_146[11:0] ? 4'h0 : _GEN_14527; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14529 = 12'h87e == _T_146[11:0] ? 4'h0 : _GEN_14528; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14530 = 12'h87f == _T_146[11:0] ? 4'h0 : _GEN_14529; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14531 = 12'h880 == _T_146[11:0] ? 4'h0 : _GEN_14530; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14532 = 12'h881 == _T_146[11:0] ? image_2177 : _GEN_14531; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14533 = 12'h882 == _T_146[11:0] ? image_2178 : _GEN_14532; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14534 = 12'h883 == _T_146[11:0] ? image_2179 : _GEN_14533; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14535 = 12'h884 == _T_146[11:0] ? image_2180 : _GEN_14534; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14536 = 12'h885 == _T_146[11:0] ? image_2181 : _GEN_14535; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14537 = 12'h886 == _T_146[11:0] ? image_2182 : _GEN_14536; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14538 = 12'h887 == _T_146[11:0] ? image_2183 : _GEN_14537; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14539 = 12'h888 == _T_146[11:0] ? image_2184 : _GEN_14538; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14540 = 12'h889 == _T_146[11:0] ? image_2185 : _GEN_14539; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14541 = 12'h88a == _T_146[11:0] ? image_2186 : _GEN_14540; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14542 = 12'h88b == _T_146[11:0] ? image_2187 : _GEN_14541; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14543 = 12'h88c == _T_146[11:0] ? image_2188 : _GEN_14542; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14544 = 12'h88d == _T_146[11:0] ? image_2189 : _GEN_14543; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14545 = 12'h88e == _T_146[11:0] ? image_2190 : _GEN_14544; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14546 = 12'h88f == _T_146[11:0] ? image_2191 : _GEN_14545; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14547 = 12'h890 == _T_146[11:0] ? image_2192 : _GEN_14546; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14548 = 12'h891 == _T_146[11:0] ? image_2193 : _GEN_14547; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14549 = 12'h892 == _T_146[11:0] ? image_2194 : _GEN_14548; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14550 = 12'h893 == _T_146[11:0] ? image_2195 : _GEN_14549; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14551 = 12'h894 == _T_146[11:0] ? image_2196 : _GEN_14550; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14552 = 12'h895 == _T_146[11:0] ? image_2197 : _GEN_14551; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14553 = 12'h896 == _T_146[11:0] ? image_2198 : _GEN_14552; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14554 = 12'h897 == _T_146[11:0] ? image_2199 : _GEN_14553; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14555 = 12'h898 == _T_146[11:0] ? image_2200 : _GEN_14554; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14556 = 12'h899 == _T_146[11:0] ? image_2201 : _GEN_14555; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14557 = 12'h89a == _T_146[11:0] ? image_2202 : _GEN_14556; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14558 = 12'h89b == _T_146[11:0] ? image_2203 : _GEN_14557; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14559 = 12'h89c == _T_146[11:0] ? image_2204 : _GEN_14558; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14560 = 12'h89d == _T_146[11:0] ? image_2205 : _GEN_14559; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14561 = 12'h89e == _T_146[11:0] ? image_2206 : _GEN_14560; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14562 = 12'h89f == _T_146[11:0] ? image_2207 : _GEN_14561; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14563 = 12'h8a0 == _T_146[11:0] ? image_2208 : _GEN_14562; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14564 = 12'h8a1 == _T_146[11:0] ? image_2209 : _GEN_14563; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14565 = 12'h8a2 == _T_146[11:0] ? image_2210 : _GEN_14564; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14566 = 12'h8a3 == _T_146[11:0] ? image_2211 : _GEN_14565; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14567 = 12'h8a4 == _T_146[11:0] ? image_2212 : _GEN_14566; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14568 = 12'h8a5 == _T_146[11:0] ? image_2213 : _GEN_14567; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14569 = 12'h8a6 == _T_146[11:0] ? image_2214 : _GEN_14568; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14570 = 12'h8a7 == _T_146[11:0] ? image_2215 : _GEN_14569; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14571 = 12'h8a8 == _T_146[11:0] ? image_2216 : _GEN_14570; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14572 = 12'h8a9 == _T_146[11:0] ? image_2217 : _GEN_14571; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14573 = 12'h8aa == _T_146[11:0] ? image_2218 : _GEN_14572; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14574 = 12'h8ab == _T_146[11:0] ? image_2219 : _GEN_14573; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14575 = 12'h8ac == _T_146[11:0] ? image_2220 : _GEN_14574; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14576 = 12'h8ad == _T_146[11:0] ? image_2221 : _GEN_14575; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14577 = 12'h8ae == _T_146[11:0] ? image_2222 : _GEN_14576; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14578 = 12'h8af == _T_146[11:0] ? image_2223 : _GEN_14577; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14579 = 12'h8b0 == _T_146[11:0] ? image_2224 : _GEN_14578; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14580 = 12'h8b1 == _T_146[11:0] ? image_2225 : _GEN_14579; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14581 = 12'h8b2 == _T_146[11:0] ? image_2226 : _GEN_14580; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14582 = 12'h8b3 == _T_146[11:0] ? image_2227 : _GEN_14581; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14583 = 12'h8b4 == _T_146[11:0] ? image_2228 : _GEN_14582; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14584 = 12'h8b5 == _T_146[11:0] ? image_2229 : _GEN_14583; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14585 = 12'h8b6 == _T_146[11:0] ? image_2230 : _GEN_14584; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14586 = 12'h8b7 == _T_146[11:0] ? image_2231 : _GEN_14585; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14587 = 12'h8b8 == _T_146[11:0] ? image_2232 : _GEN_14586; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14588 = 12'h8b9 == _T_146[11:0] ? image_2233 : _GEN_14587; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14589 = 12'h8ba == _T_146[11:0] ? image_2234 : _GEN_14588; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14590 = 12'h8bb == _T_146[11:0] ? 4'h0 : _GEN_14589; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14591 = 12'h8bc == _T_146[11:0] ? 4'h0 : _GEN_14590; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14592 = 12'h8bd == _T_146[11:0] ? 4'h0 : _GEN_14591; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14593 = 12'h8be == _T_146[11:0] ? 4'h0 : _GEN_14592; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14594 = 12'h8bf == _T_146[11:0] ? 4'h0 : _GEN_14593; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14595 = 12'h8c0 == _T_146[11:0] ? 4'h0 : _GEN_14594; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14596 = 12'h8c1 == _T_146[11:0] ? 4'h0 : _GEN_14595; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14597 = 12'h8c2 == _T_146[11:0] ? 4'h0 : _GEN_14596; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14598 = 12'h8c3 == _T_146[11:0] ? image_2243 : _GEN_14597; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14599 = 12'h8c4 == _T_146[11:0] ? image_2244 : _GEN_14598; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14600 = 12'h8c5 == _T_146[11:0] ? image_2245 : _GEN_14599; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14601 = 12'h8c6 == _T_146[11:0] ? image_2246 : _GEN_14600; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14602 = 12'h8c7 == _T_146[11:0] ? image_2247 : _GEN_14601; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14603 = 12'h8c8 == _T_146[11:0] ? image_2248 : _GEN_14602; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14604 = 12'h8c9 == _T_146[11:0] ? image_2249 : _GEN_14603; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14605 = 12'h8ca == _T_146[11:0] ? image_2250 : _GEN_14604; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14606 = 12'h8cb == _T_146[11:0] ? image_2251 : _GEN_14605; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14607 = 12'h8cc == _T_146[11:0] ? image_2252 : _GEN_14606; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14608 = 12'h8cd == _T_146[11:0] ? image_2253 : _GEN_14607; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14609 = 12'h8ce == _T_146[11:0] ? image_2254 : _GEN_14608; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14610 = 12'h8cf == _T_146[11:0] ? image_2255 : _GEN_14609; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14611 = 12'h8d0 == _T_146[11:0] ? image_2256 : _GEN_14610; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14612 = 12'h8d1 == _T_146[11:0] ? image_2257 : _GEN_14611; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14613 = 12'h8d2 == _T_146[11:0] ? image_2258 : _GEN_14612; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14614 = 12'h8d3 == _T_146[11:0] ? image_2259 : _GEN_14613; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14615 = 12'h8d4 == _T_146[11:0] ? image_2260 : _GEN_14614; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14616 = 12'h8d5 == _T_146[11:0] ? image_2261 : _GEN_14615; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14617 = 12'h8d6 == _T_146[11:0] ? image_2262 : _GEN_14616; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14618 = 12'h8d7 == _T_146[11:0] ? image_2263 : _GEN_14617; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14619 = 12'h8d8 == _T_146[11:0] ? image_2264 : _GEN_14618; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14620 = 12'h8d9 == _T_146[11:0] ? image_2265 : _GEN_14619; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14621 = 12'h8da == _T_146[11:0] ? image_2266 : _GEN_14620; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14622 = 12'h8db == _T_146[11:0] ? image_2267 : _GEN_14621; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14623 = 12'h8dc == _T_146[11:0] ? image_2268 : _GEN_14622; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14624 = 12'h8dd == _T_146[11:0] ? image_2269 : _GEN_14623; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14625 = 12'h8de == _T_146[11:0] ? image_2270 : _GEN_14624; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14626 = 12'h8df == _T_146[11:0] ? image_2271 : _GEN_14625; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14627 = 12'h8e0 == _T_146[11:0] ? image_2272 : _GEN_14626; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14628 = 12'h8e1 == _T_146[11:0] ? image_2273 : _GEN_14627; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14629 = 12'h8e2 == _T_146[11:0] ? image_2274 : _GEN_14628; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14630 = 12'h8e3 == _T_146[11:0] ? image_2275 : _GEN_14629; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14631 = 12'h8e4 == _T_146[11:0] ? image_2276 : _GEN_14630; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14632 = 12'h8e5 == _T_146[11:0] ? image_2277 : _GEN_14631; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14633 = 12'h8e6 == _T_146[11:0] ? image_2278 : _GEN_14632; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14634 = 12'h8e7 == _T_146[11:0] ? image_2279 : _GEN_14633; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14635 = 12'h8e8 == _T_146[11:0] ? image_2280 : _GEN_14634; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14636 = 12'h8e9 == _T_146[11:0] ? image_2281 : _GEN_14635; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14637 = 12'h8ea == _T_146[11:0] ? image_2282 : _GEN_14636; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14638 = 12'h8eb == _T_146[11:0] ? image_2283 : _GEN_14637; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14639 = 12'h8ec == _T_146[11:0] ? image_2284 : _GEN_14638; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14640 = 12'h8ed == _T_146[11:0] ? image_2285 : _GEN_14639; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14641 = 12'h8ee == _T_146[11:0] ? image_2286 : _GEN_14640; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14642 = 12'h8ef == _T_146[11:0] ? image_2287 : _GEN_14641; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14643 = 12'h8f0 == _T_146[11:0] ? image_2288 : _GEN_14642; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14644 = 12'h8f1 == _T_146[11:0] ? image_2289 : _GEN_14643; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14645 = 12'h8f2 == _T_146[11:0] ? image_2290 : _GEN_14644; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14646 = 12'h8f3 == _T_146[11:0] ? image_2291 : _GEN_14645; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14647 = 12'h8f4 == _T_146[11:0] ? image_2292 : _GEN_14646; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14648 = 12'h8f5 == _T_146[11:0] ? image_2293 : _GEN_14647; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14649 = 12'h8f6 == _T_146[11:0] ? image_2294 : _GEN_14648; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14650 = 12'h8f7 == _T_146[11:0] ? image_2295 : _GEN_14649; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14651 = 12'h8f8 == _T_146[11:0] ? image_2296 : _GEN_14650; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14652 = 12'h8f9 == _T_146[11:0] ? image_2297 : _GEN_14651; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14653 = 12'h8fa == _T_146[11:0] ? image_2298 : _GEN_14652; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14654 = 12'h8fb == _T_146[11:0] ? 4'h0 : _GEN_14653; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14655 = 12'h8fc == _T_146[11:0] ? 4'h0 : _GEN_14654; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14656 = 12'h8fd == _T_146[11:0] ? 4'h0 : _GEN_14655; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14657 = 12'h8fe == _T_146[11:0] ? 4'h0 : _GEN_14656; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14658 = 12'h8ff == _T_146[11:0] ? 4'h0 : _GEN_14657; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14659 = 12'h900 == _T_146[11:0] ? 4'h0 : _GEN_14658; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14660 = 12'h901 == _T_146[11:0] ? 4'h0 : _GEN_14659; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14661 = 12'h902 == _T_146[11:0] ? 4'h0 : _GEN_14660; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14662 = 12'h903 == _T_146[11:0] ? image_2307 : _GEN_14661; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14663 = 12'h904 == _T_146[11:0] ? image_2308 : _GEN_14662; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14664 = 12'h905 == _T_146[11:0] ? image_2309 : _GEN_14663; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14665 = 12'h906 == _T_146[11:0] ? image_2310 : _GEN_14664; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14666 = 12'h907 == _T_146[11:0] ? image_2311 : _GEN_14665; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14667 = 12'h908 == _T_146[11:0] ? image_2312 : _GEN_14666; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14668 = 12'h909 == _T_146[11:0] ? image_2313 : _GEN_14667; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14669 = 12'h90a == _T_146[11:0] ? image_2314 : _GEN_14668; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14670 = 12'h90b == _T_146[11:0] ? image_2315 : _GEN_14669; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14671 = 12'h90c == _T_146[11:0] ? image_2316 : _GEN_14670; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14672 = 12'h90d == _T_146[11:0] ? image_2317 : _GEN_14671; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14673 = 12'h90e == _T_146[11:0] ? image_2318 : _GEN_14672; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14674 = 12'h90f == _T_146[11:0] ? image_2319 : _GEN_14673; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14675 = 12'h910 == _T_146[11:0] ? image_2320 : _GEN_14674; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14676 = 12'h911 == _T_146[11:0] ? image_2321 : _GEN_14675; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14677 = 12'h912 == _T_146[11:0] ? image_2322 : _GEN_14676; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14678 = 12'h913 == _T_146[11:0] ? image_2323 : _GEN_14677; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14679 = 12'h914 == _T_146[11:0] ? image_2324 : _GEN_14678; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14680 = 12'h915 == _T_146[11:0] ? image_2325 : _GEN_14679; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14681 = 12'h916 == _T_146[11:0] ? image_2326 : _GEN_14680; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14682 = 12'h917 == _T_146[11:0] ? image_2327 : _GEN_14681; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14683 = 12'h918 == _T_146[11:0] ? image_2328 : _GEN_14682; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14684 = 12'h919 == _T_146[11:0] ? image_2329 : _GEN_14683; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14685 = 12'h91a == _T_146[11:0] ? image_2330 : _GEN_14684; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14686 = 12'h91b == _T_146[11:0] ? image_2331 : _GEN_14685; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14687 = 12'h91c == _T_146[11:0] ? image_2332 : _GEN_14686; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14688 = 12'h91d == _T_146[11:0] ? image_2333 : _GEN_14687; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14689 = 12'h91e == _T_146[11:0] ? image_2334 : _GEN_14688; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14690 = 12'h91f == _T_146[11:0] ? image_2335 : _GEN_14689; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14691 = 12'h920 == _T_146[11:0] ? image_2336 : _GEN_14690; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14692 = 12'h921 == _T_146[11:0] ? image_2337 : _GEN_14691; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14693 = 12'h922 == _T_146[11:0] ? image_2338 : _GEN_14692; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14694 = 12'h923 == _T_146[11:0] ? image_2339 : _GEN_14693; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14695 = 12'h924 == _T_146[11:0] ? image_2340 : _GEN_14694; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14696 = 12'h925 == _T_146[11:0] ? image_2341 : _GEN_14695; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14697 = 12'h926 == _T_146[11:0] ? image_2342 : _GEN_14696; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14698 = 12'h927 == _T_146[11:0] ? image_2343 : _GEN_14697; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14699 = 12'h928 == _T_146[11:0] ? image_2344 : _GEN_14698; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14700 = 12'h929 == _T_146[11:0] ? image_2345 : _GEN_14699; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14701 = 12'h92a == _T_146[11:0] ? image_2346 : _GEN_14700; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14702 = 12'h92b == _T_146[11:0] ? image_2347 : _GEN_14701; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14703 = 12'h92c == _T_146[11:0] ? image_2348 : _GEN_14702; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14704 = 12'h92d == _T_146[11:0] ? image_2349 : _GEN_14703; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14705 = 12'h92e == _T_146[11:0] ? image_2350 : _GEN_14704; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14706 = 12'h92f == _T_146[11:0] ? image_2351 : _GEN_14705; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14707 = 12'h930 == _T_146[11:0] ? image_2352 : _GEN_14706; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14708 = 12'h931 == _T_146[11:0] ? image_2353 : _GEN_14707; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14709 = 12'h932 == _T_146[11:0] ? image_2354 : _GEN_14708; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14710 = 12'h933 == _T_146[11:0] ? image_2355 : _GEN_14709; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14711 = 12'h934 == _T_146[11:0] ? image_2356 : _GEN_14710; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14712 = 12'h935 == _T_146[11:0] ? image_2357 : _GEN_14711; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14713 = 12'h936 == _T_146[11:0] ? image_2358 : _GEN_14712; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14714 = 12'h937 == _T_146[11:0] ? image_2359 : _GEN_14713; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14715 = 12'h938 == _T_146[11:0] ? image_2360 : _GEN_14714; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14716 = 12'h939 == _T_146[11:0] ? image_2361 : _GEN_14715; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14717 = 12'h93a == _T_146[11:0] ? image_2362 : _GEN_14716; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14718 = 12'h93b == _T_146[11:0] ? 4'h0 : _GEN_14717; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14719 = 12'h93c == _T_146[11:0] ? 4'h0 : _GEN_14718; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14720 = 12'h93d == _T_146[11:0] ? 4'h0 : _GEN_14719; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14721 = 12'h93e == _T_146[11:0] ? 4'h0 : _GEN_14720; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14722 = 12'h93f == _T_146[11:0] ? 4'h0 : _GEN_14721; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14723 = 12'h940 == _T_146[11:0] ? 4'h0 : _GEN_14722; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14724 = 12'h941 == _T_146[11:0] ? 4'h0 : _GEN_14723; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14725 = 12'h942 == _T_146[11:0] ? 4'h0 : _GEN_14724; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14726 = 12'h943 == _T_146[11:0] ? 4'h0 : _GEN_14725; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14727 = 12'h944 == _T_146[11:0] ? image_2372 : _GEN_14726; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14728 = 12'h945 == _T_146[11:0] ? image_2373 : _GEN_14727; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14729 = 12'h946 == _T_146[11:0] ? image_2374 : _GEN_14728; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14730 = 12'h947 == _T_146[11:0] ? image_2375 : _GEN_14729; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14731 = 12'h948 == _T_146[11:0] ? image_2376 : _GEN_14730; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14732 = 12'h949 == _T_146[11:0] ? image_2377 : _GEN_14731; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14733 = 12'h94a == _T_146[11:0] ? image_2378 : _GEN_14732; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14734 = 12'h94b == _T_146[11:0] ? image_2379 : _GEN_14733; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14735 = 12'h94c == _T_146[11:0] ? image_2380 : _GEN_14734; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14736 = 12'h94d == _T_146[11:0] ? image_2381 : _GEN_14735; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14737 = 12'h94e == _T_146[11:0] ? image_2382 : _GEN_14736; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14738 = 12'h94f == _T_146[11:0] ? image_2383 : _GEN_14737; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14739 = 12'h950 == _T_146[11:0] ? image_2384 : _GEN_14738; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14740 = 12'h951 == _T_146[11:0] ? image_2385 : _GEN_14739; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14741 = 12'h952 == _T_146[11:0] ? image_2386 : _GEN_14740; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14742 = 12'h953 == _T_146[11:0] ? image_2387 : _GEN_14741; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14743 = 12'h954 == _T_146[11:0] ? image_2388 : _GEN_14742; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14744 = 12'h955 == _T_146[11:0] ? image_2389 : _GEN_14743; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14745 = 12'h956 == _T_146[11:0] ? image_2390 : _GEN_14744; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14746 = 12'h957 == _T_146[11:0] ? image_2391 : _GEN_14745; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14747 = 12'h958 == _T_146[11:0] ? image_2392 : _GEN_14746; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14748 = 12'h959 == _T_146[11:0] ? image_2393 : _GEN_14747; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14749 = 12'h95a == _T_146[11:0] ? image_2394 : _GEN_14748; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14750 = 12'h95b == _T_146[11:0] ? image_2395 : _GEN_14749; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14751 = 12'h95c == _T_146[11:0] ? image_2396 : _GEN_14750; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14752 = 12'h95d == _T_146[11:0] ? image_2397 : _GEN_14751; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14753 = 12'h95e == _T_146[11:0] ? image_2398 : _GEN_14752; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14754 = 12'h95f == _T_146[11:0] ? image_2399 : _GEN_14753; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14755 = 12'h960 == _T_146[11:0] ? image_2400 : _GEN_14754; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14756 = 12'h961 == _T_146[11:0] ? image_2401 : _GEN_14755; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14757 = 12'h962 == _T_146[11:0] ? image_2402 : _GEN_14756; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14758 = 12'h963 == _T_146[11:0] ? image_2403 : _GEN_14757; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14759 = 12'h964 == _T_146[11:0] ? image_2404 : _GEN_14758; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14760 = 12'h965 == _T_146[11:0] ? image_2405 : _GEN_14759; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14761 = 12'h966 == _T_146[11:0] ? image_2406 : _GEN_14760; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14762 = 12'h967 == _T_146[11:0] ? image_2407 : _GEN_14761; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14763 = 12'h968 == _T_146[11:0] ? image_2408 : _GEN_14762; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14764 = 12'h969 == _T_146[11:0] ? image_2409 : _GEN_14763; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14765 = 12'h96a == _T_146[11:0] ? image_2410 : _GEN_14764; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14766 = 12'h96b == _T_146[11:0] ? image_2411 : _GEN_14765; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14767 = 12'h96c == _T_146[11:0] ? image_2412 : _GEN_14766; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14768 = 12'h96d == _T_146[11:0] ? image_2413 : _GEN_14767; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14769 = 12'h96e == _T_146[11:0] ? image_2414 : _GEN_14768; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14770 = 12'h96f == _T_146[11:0] ? image_2415 : _GEN_14769; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14771 = 12'h970 == _T_146[11:0] ? image_2416 : _GEN_14770; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14772 = 12'h971 == _T_146[11:0] ? image_2417 : _GEN_14771; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14773 = 12'h972 == _T_146[11:0] ? image_2418 : _GEN_14772; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14774 = 12'h973 == _T_146[11:0] ? image_2419 : _GEN_14773; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14775 = 12'h974 == _T_146[11:0] ? image_2420 : _GEN_14774; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14776 = 12'h975 == _T_146[11:0] ? image_2421 : _GEN_14775; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14777 = 12'h976 == _T_146[11:0] ? image_2422 : _GEN_14776; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14778 = 12'h977 == _T_146[11:0] ? image_2423 : _GEN_14777; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14779 = 12'h978 == _T_146[11:0] ? image_2424 : _GEN_14778; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14780 = 12'h979 == _T_146[11:0] ? image_2425 : _GEN_14779; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14781 = 12'h97a == _T_146[11:0] ? image_2426 : _GEN_14780; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14782 = 12'h97b == _T_146[11:0] ? 4'h0 : _GEN_14781; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14783 = 12'h97c == _T_146[11:0] ? 4'h0 : _GEN_14782; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14784 = 12'h97d == _T_146[11:0] ? 4'h0 : _GEN_14783; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14785 = 12'h97e == _T_146[11:0] ? 4'h0 : _GEN_14784; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14786 = 12'h97f == _T_146[11:0] ? 4'h0 : _GEN_14785; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14787 = 12'h980 == _T_146[11:0] ? 4'h0 : _GEN_14786; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14788 = 12'h981 == _T_146[11:0] ? 4'h0 : _GEN_14787; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14789 = 12'h982 == _T_146[11:0] ? 4'h0 : _GEN_14788; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14790 = 12'h983 == _T_146[11:0] ? 4'h0 : _GEN_14789; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14791 = 12'h984 == _T_146[11:0] ? 4'h0 : _GEN_14790; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14792 = 12'h985 == _T_146[11:0] ? image_2437 : _GEN_14791; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14793 = 12'h986 == _T_146[11:0] ? image_2438 : _GEN_14792; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14794 = 12'h987 == _T_146[11:0] ? image_2439 : _GEN_14793; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14795 = 12'h988 == _T_146[11:0] ? image_2440 : _GEN_14794; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14796 = 12'h989 == _T_146[11:0] ? image_2441 : _GEN_14795; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14797 = 12'h98a == _T_146[11:0] ? image_2442 : _GEN_14796; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14798 = 12'h98b == _T_146[11:0] ? image_2443 : _GEN_14797; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14799 = 12'h98c == _T_146[11:0] ? image_2444 : _GEN_14798; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14800 = 12'h98d == _T_146[11:0] ? image_2445 : _GEN_14799; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14801 = 12'h98e == _T_146[11:0] ? image_2446 : _GEN_14800; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14802 = 12'h98f == _T_146[11:0] ? image_2447 : _GEN_14801; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14803 = 12'h990 == _T_146[11:0] ? image_2448 : _GEN_14802; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14804 = 12'h991 == _T_146[11:0] ? image_2449 : _GEN_14803; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14805 = 12'h992 == _T_146[11:0] ? image_2450 : _GEN_14804; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14806 = 12'h993 == _T_146[11:0] ? image_2451 : _GEN_14805; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14807 = 12'h994 == _T_146[11:0] ? image_2452 : _GEN_14806; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14808 = 12'h995 == _T_146[11:0] ? image_2453 : _GEN_14807; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14809 = 12'h996 == _T_146[11:0] ? image_2454 : _GEN_14808; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14810 = 12'h997 == _T_146[11:0] ? image_2455 : _GEN_14809; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14811 = 12'h998 == _T_146[11:0] ? image_2456 : _GEN_14810; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14812 = 12'h999 == _T_146[11:0] ? image_2457 : _GEN_14811; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14813 = 12'h99a == _T_146[11:0] ? image_2458 : _GEN_14812; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14814 = 12'h99b == _T_146[11:0] ? image_2459 : _GEN_14813; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14815 = 12'h99c == _T_146[11:0] ? image_2460 : _GEN_14814; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14816 = 12'h99d == _T_146[11:0] ? image_2461 : _GEN_14815; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14817 = 12'h99e == _T_146[11:0] ? image_2462 : _GEN_14816; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14818 = 12'h99f == _T_146[11:0] ? image_2463 : _GEN_14817; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14819 = 12'h9a0 == _T_146[11:0] ? image_2464 : _GEN_14818; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14820 = 12'h9a1 == _T_146[11:0] ? image_2465 : _GEN_14819; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14821 = 12'h9a2 == _T_146[11:0] ? image_2466 : _GEN_14820; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14822 = 12'h9a3 == _T_146[11:0] ? image_2467 : _GEN_14821; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14823 = 12'h9a4 == _T_146[11:0] ? image_2468 : _GEN_14822; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14824 = 12'h9a5 == _T_146[11:0] ? image_2469 : _GEN_14823; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14825 = 12'h9a6 == _T_146[11:0] ? image_2470 : _GEN_14824; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14826 = 12'h9a7 == _T_146[11:0] ? image_2471 : _GEN_14825; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14827 = 12'h9a8 == _T_146[11:0] ? image_2472 : _GEN_14826; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14828 = 12'h9a9 == _T_146[11:0] ? image_2473 : _GEN_14827; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14829 = 12'h9aa == _T_146[11:0] ? image_2474 : _GEN_14828; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14830 = 12'h9ab == _T_146[11:0] ? image_2475 : _GEN_14829; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14831 = 12'h9ac == _T_146[11:0] ? image_2476 : _GEN_14830; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14832 = 12'h9ad == _T_146[11:0] ? image_2477 : _GEN_14831; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14833 = 12'h9ae == _T_146[11:0] ? image_2478 : _GEN_14832; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14834 = 12'h9af == _T_146[11:0] ? image_2479 : _GEN_14833; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14835 = 12'h9b0 == _T_146[11:0] ? image_2480 : _GEN_14834; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14836 = 12'h9b1 == _T_146[11:0] ? image_2481 : _GEN_14835; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14837 = 12'h9b2 == _T_146[11:0] ? image_2482 : _GEN_14836; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14838 = 12'h9b3 == _T_146[11:0] ? image_2483 : _GEN_14837; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14839 = 12'h9b4 == _T_146[11:0] ? image_2484 : _GEN_14838; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14840 = 12'h9b5 == _T_146[11:0] ? image_2485 : _GEN_14839; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14841 = 12'h9b6 == _T_146[11:0] ? image_2486 : _GEN_14840; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14842 = 12'h9b7 == _T_146[11:0] ? image_2487 : _GEN_14841; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14843 = 12'h9b8 == _T_146[11:0] ? image_2488 : _GEN_14842; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14844 = 12'h9b9 == _T_146[11:0] ? image_2489 : _GEN_14843; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14845 = 12'h9ba == _T_146[11:0] ? image_2490 : _GEN_14844; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14846 = 12'h9bb == _T_146[11:0] ? 4'h0 : _GEN_14845; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14847 = 12'h9bc == _T_146[11:0] ? 4'h0 : _GEN_14846; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14848 = 12'h9bd == _T_146[11:0] ? 4'h0 : _GEN_14847; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14849 = 12'h9be == _T_146[11:0] ? 4'h0 : _GEN_14848; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14850 = 12'h9bf == _T_146[11:0] ? 4'h0 : _GEN_14849; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14851 = 12'h9c0 == _T_146[11:0] ? 4'h0 : _GEN_14850; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14852 = 12'h9c1 == _T_146[11:0] ? 4'h0 : _GEN_14851; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14853 = 12'h9c2 == _T_146[11:0] ? 4'h0 : _GEN_14852; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14854 = 12'h9c3 == _T_146[11:0] ? 4'h0 : _GEN_14853; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14855 = 12'h9c4 == _T_146[11:0] ? 4'h0 : _GEN_14854; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14856 = 12'h9c5 == _T_146[11:0] ? 4'h0 : _GEN_14855; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14857 = 12'h9c6 == _T_146[11:0] ? image_2502 : _GEN_14856; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14858 = 12'h9c7 == _T_146[11:0] ? image_2503 : _GEN_14857; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14859 = 12'h9c8 == _T_146[11:0] ? image_2504 : _GEN_14858; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14860 = 12'h9c9 == _T_146[11:0] ? image_2505 : _GEN_14859; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14861 = 12'h9ca == _T_146[11:0] ? image_2506 : _GEN_14860; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14862 = 12'h9cb == _T_146[11:0] ? image_2507 : _GEN_14861; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14863 = 12'h9cc == _T_146[11:0] ? image_2508 : _GEN_14862; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14864 = 12'h9cd == _T_146[11:0] ? image_2509 : _GEN_14863; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14865 = 12'h9ce == _T_146[11:0] ? image_2510 : _GEN_14864; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14866 = 12'h9cf == _T_146[11:0] ? image_2511 : _GEN_14865; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14867 = 12'h9d0 == _T_146[11:0] ? image_2512 : _GEN_14866; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14868 = 12'h9d1 == _T_146[11:0] ? image_2513 : _GEN_14867; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14869 = 12'h9d2 == _T_146[11:0] ? image_2514 : _GEN_14868; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14870 = 12'h9d3 == _T_146[11:0] ? image_2515 : _GEN_14869; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14871 = 12'h9d4 == _T_146[11:0] ? image_2516 : _GEN_14870; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14872 = 12'h9d5 == _T_146[11:0] ? image_2517 : _GEN_14871; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14873 = 12'h9d6 == _T_146[11:0] ? image_2518 : _GEN_14872; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14874 = 12'h9d7 == _T_146[11:0] ? image_2519 : _GEN_14873; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14875 = 12'h9d8 == _T_146[11:0] ? image_2520 : _GEN_14874; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14876 = 12'h9d9 == _T_146[11:0] ? image_2521 : _GEN_14875; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14877 = 12'h9da == _T_146[11:0] ? image_2522 : _GEN_14876; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14878 = 12'h9db == _T_146[11:0] ? image_2523 : _GEN_14877; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14879 = 12'h9dc == _T_146[11:0] ? image_2524 : _GEN_14878; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14880 = 12'h9dd == _T_146[11:0] ? image_2525 : _GEN_14879; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14881 = 12'h9de == _T_146[11:0] ? image_2526 : _GEN_14880; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14882 = 12'h9df == _T_146[11:0] ? image_2527 : _GEN_14881; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14883 = 12'h9e0 == _T_146[11:0] ? image_2528 : _GEN_14882; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14884 = 12'h9e1 == _T_146[11:0] ? image_2529 : _GEN_14883; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14885 = 12'h9e2 == _T_146[11:0] ? image_2530 : _GEN_14884; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14886 = 12'h9e3 == _T_146[11:0] ? image_2531 : _GEN_14885; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14887 = 12'h9e4 == _T_146[11:0] ? image_2532 : _GEN_14886; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14888 = 12'h9e5 == _T_146[11:0] ? image_2533 : _GEN_14887; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14889 = 12'h9e6 == _T_146[11:0] ? image_2534 : _GEN_14888; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14890 = 12'h9e7 == _T_146[11:0] ? image_2535 : _GEN_14889; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14891 = 12'h9e8 == _T_146[11:0] ? image_2536 : _GEN_14890; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14892 = 12'h9e9 == _T_146[11:0] ? image_2537 : _GEN_14891; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14893 = 12'h9ea == _T_146[11:0] ? image_2538 : _GEN_14892; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14894 = 12'h9eb == _T_146[11:0] ? image_2539 : _GEN_14893; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14895 = 12'h9ec == _T_146[11:0] ? image_2540 : _GEN_14894; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14896 = 12'h9ed == _T_146[11:0] ? image_2541 : _GEN_14895; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14897 = 12'h9ee == _T_146[11:0] ? image_2542 : _GEN_14896; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14898 = 12'h9ef == _T_146[11:0] ? image_2543 : _GEN_14897; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14899 = 12'h9f0 == _T_146[11:0] ? image_2544 : _GEN_14898; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14900 = 12'h9f1 == _T_146[11:0] ? image_2545 : _GEN_14899; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14901 = 12'h9f2 == _T_146[11:0] ? image_2546 : _GEN_14900; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14902 = 12'h9f3 == _T_146[11:0] ? image_2547 : _GEN_14901; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14903 = 12'h9f4 == _T_146[11:0] ? image_2548 : _GEN_14902; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14904 = 12'h9f5 == _T_146[11:0] ? image_2549 : _GEN_14903; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14905 = 12'h9f6 == _T_146[11:0] ? image_2550 : _GEN_14904; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14906 = 12'h9f7 == _T_146[11:0] ? image_2551 : _GEN_14905; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14907 = 12'h9f8 == _T_146[11:0] ? image_2552 : _GEN_14906; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14908 = 12'h9f9 == _T_146[11:0] ? image_2553 : _GEN_14907; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14909 = 12'h9fa == _T_146[11:0] ? image_2554 : _GEN_14908; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14910 = 12'h9fb == _T_146[11:0] ? 4'h0 : _GEN_14909; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14911 = 12'h9fc == _T_146[11:0] ? 4'h0 : _GEN_14910; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14912 = 12'h9fd == _T_146[11:0] ? 4'h0 : _GEN_14911; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14913 = 12'h9fe == _T_146[11:0] ? 4'h0 : _GEN_14912; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14914 = 12'h9ff == _T_146[11:0] ? 4'h0 : _GEN_14913; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14915 = 12'ha00 == _T_146[11:0] ? 4'h0 : _GEN_14914; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14916 = 12'ha01 == _T_146[11:0] ? 4'h0 : _GEN_14915; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14917 = 12'ha02 == _T_146[11:0] ? 4'h0 : _GEN_14916; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14918 = 12'ha03 == _T_146[11:0] ? 4'h0 : _GEN_14917; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14919 = 12'ha04 == _T_146[11:0] ? 4'h0 : _GEN_14918; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14920 = 12'ha05 == _T_146[11:0] ? 4'h0 : _GEN_14919; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14921 = 12'ha06 == _T_146[11:0] ? 4'h0 : _GEN_14920; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14922 = 12'ha07 == _T_146[11:0] ? image_2567 : _GEN_14921; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14923 = 12'ha08 == _T_146[11:0] ? image_2568 : _GEN_14922; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14924 = 12'ha09 == _T_146[11:0] ? image_2569 : _GEN_14923; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14925 = 12'ha0a == _T_146[11:0] ? image_2570 : _GEN_14924; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14926 = 12'ha0b == _T_146[11:0] ? image_2571 : _GEN_14925; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14927 = 12'ha0c == _T_146[11:0] ? image_2572 : _GEN_14926; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14928 = 12'ha0d == _T_146[11:0] ? image_2573 : _GEN_14927; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14929 = 12'ha0e == _T_146[11:0] ? image_2574 : _GEN_14928; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14930 = 12'ha0f == _T_146[11:0] ? image_2575 : _GEN_14929; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14931 = 12'ha10 == _T_146[11:0] ? image_2576 : _GEN_14930; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14932 = 12'ha11 == _T_146[11:0] ? image_2577 : _GEN_14931; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14933 = 12'ha12 == _T_146[11:0] ? image_2578 : _GEN_14932; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14934 = 12'ha13 == _T_146[11:0] ? image_2579 : _GEN_14933; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14935 = 12'ha14 == _T_146[11:0] ? image_2580 : _GEN_14934; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14936 = 12'ha15 == _T_146[11:0] ? image_2581 : _GEN_14935; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14937 = 12'ha16 == _T_146[11:0] ? image_2582 : _GEN_14936; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14938 = 12'ha17 == _T_146[11:0] ? image_2583 : _GEN_14937; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14939 = 12'ha18 == _T_146[11:0] ? image_2584 : _GEN_14938; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14940 = 12'ha19 == _T_146[11:0] ? image_2585 : _GEN_14939; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14941 = 12'ha1a == _T_146[11:0] ? image_2586 : _GEN_14940; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14942 = 12'ha1b == _T_146[11:0] ? image_2587 : _GEN_14941; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14943 = 12'ha1c == _T_146[11:0] ? image_2588 : _GEN_14942; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14944 = 12'ha1d == _T_146[11:0] ? image_2589 : _GEN_14943; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14945 = 12'ha1e == _T_146[11:0] ? image_2590 : _GEN_14944; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14946 = 12'ha1f == _T_146[11:0] ? image_2591 : _GEN_14945; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14947 = 12'ha20 == _T_146[11:0] ? image_2592 : _GEN_14946; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14948 = 12'ha21 == _T_146[11:0] ? image_2593 : _GEN_14947; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14949 = 12'ha22 == _T_146[11:0] ? image_2594 : _GEN_14948; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14950 = 12'ha23 == _T_146[11:0] ? image_2595 : _GEN_14949; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14951 = 12'ha24 == _T_146[11:0] ? image_2596 : _GEN_14950; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14952 = 12'ha25 == _T_146[11:0] ? image_2597 : _GEN_14951; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14953 = 12'ha26 == _T_146[11:0] ? image_2598 : _GEN_14952; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14954 = 12'ha27 == _T_146[11:0] ? image_2599 : _GEN_14953; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14955 = 12'ha28 == _T_146[11:0] ? image_2600 : _GEN_14954; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14956 = 12'ha29 == _T_146[11:0] ? image_2601 : _GEN_14955; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14957 = 12'ha2a == _T_146[11:0] ? image_2602 : _GEN_14956; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14958 = 12'ha2b == _T_146[11:0] ? image_2603 : _GEN_14957; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14959 = 12'ha2c == _T_146[11:0] ? image_2604 : _GEN_14958; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14960 = 12'ha2d == _T_146[11:0] ? image_2605 : _GEN_14959; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14961 = 12'ha2e == _T_146[11:0] ? image_2606 : _GEN_14960; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14962 = 12'ha2f == _T_146[11:0] ? image_2607 : _GEN_14961; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14963 = 12'ha30 == _T_146[11:0] ? image_2608 : _GEN_14962; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14964 = 12'ha31 == _T_146[11:0] ? image_2609 : _GEN_14963; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14965 = 12'ha32 == _T_146[11:0] ? image_2610 : _GEN_14964; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14966 = 12'ha33 == _T_146[11:0] ? image_2611 : _GEN_14965; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14967 = 12'ha34 == _T_146[11:0] ? image_2612 : _GEN_14966; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14968 = 12'ha35 == _T_146[11:0] ? image_2613 : _GEN_14967; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14969 = 12'ha36 == _T_146[11:0] ? image_2614 : _GEN_14968; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14970 = 12'ha37 == _T_146[11:0] ? image_2615 : _GEN_14969; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14971 = 12'ha38 == _T_146[11:0] ? image_2616 : _GEN_14970; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14972 = 12'ha39 == _T_146[11:0] ? image_2617 : _GEN_14971; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14973 = 12'ha3a == _T_146[11:0] ? image_2618 : _GEN_14972; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14974 = 12'ha3b == _T_146[11:0] ? 4'h0 : _GEN_14973; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14975 = 12'ha3c == _T_146[11:0] ? 4'h0 : _GEN_14974; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14976 = 12'ha3d == _T_146[11:0] ? 4'h0 : _GEN_14975; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14977 = 12'ha3e == _T_146[11:0] ? 4'h0 : _GEN_14976; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14978 = 12'ha3f == _T_146[11:0] ? 4'h0 : _GEN_14977; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14979 = 12'ha40 == _T_146[11:0] ? 4'h0 : _GEN_14978; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14980 = 12'ha41 == _T_146[11:0] ? 4'h0 : _GEN_14979; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14981 = 12'ha42 == _T_146[11:0] ? 4'h0 : _GEN_14980; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14982 = 12'ha43 == _T_146[11:0] ? 4'h0 : _GEN_14981; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14983 = 12'ha44 == _T_146[11:0] ? 4'h0 : _GEN_14982; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14984 = 12'ha45 == _T_146[11:0] ? 4'h0 : _GEN_14983; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14985 = 12'ha46 == _T_146[11:0] ? 4'h0 : _GEN_14984; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14986 = 12'ha47 == _T_146[11:0] ? 4'h0 : _GEN_14985; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14987 = 12'ha48 == _T_146[11:0] ? image_2632 : _GEN_14986; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14988 = 12'ha49 == _T_146[11:0] ? image_2633 : _GEN_14987; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14989 = 12'ha4a == _T_146[11:0] ? image_2634 : _GEN_14988; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14990 = 12'ha4b == _T_146[11:0] ? image_2635 : _GEN_14989; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14991 = 12'ha4c == _T_146[11:0] ? image_2636 : _GEN_14990; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14992 = 12'ha4d == _T_146[11:0] ? image_2637 : _GEN_14991; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14993 = 12'ha4e == _T_146[11:0] ? image_2638 : _GEN_14992; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14994 = 12'ha4f == _T_146[11:0] ? image_2639 : _GEN_14993; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14995 = 12'ha50 == _T_146[11:0] ? image_2640 : _GEN_14994; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14996 = 12'ha51 == _T_146[11:0] ? image_2641 : _GEN_14995; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14997 = 12'ha52 == _T_146[11:0] ? image_2642 : _GEN_14996; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14998 = 12'ha53 == _T_146[11:0] ? image_2643 : _GEN_14997; // @[Filter.scala 138:46]
  wire [3:0] _GEN_14999 = 12'ha54 == _T_146[11:0] ? image_2644 : _GEN_14998; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15000 = 12'ha55 == _T_146[11:0] ? image_2645 : _GEN_14999; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15001 = 12'ha56 == _T_146[11:0] ? image_2646 : _GEN_15000; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15002 = 12'ha57 == _T_146[11:0] ? image_2647 : _GEN_15001; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15003 = 12'ha58 == _T_146[11:0] ? image_2648 : _GEN_15002; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15004 = 12'ha59 == _T_146[11:0] ? image_2649 : _GEN_15003; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15005 = 12'ha5a == _T_146[11:0] ? image_2650 : _GEN_15004; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15006 = 12'ha5b == _T_146[11:0] ? image_2651 : _GEN_15005; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15007 = 12'ha5c == _T_146[11:0] ? image_2652 : _GEN_15006; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15008 = 12'ha5d == _T_146[11:0] ? image_2653 : _GEN_15007; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15009 = 12'ha5e == _T_146[11:0] ? image_2654 : _GEN_15008; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15010 = 12'ha5f == _T_146[11:0] ? image_2655 : _GEN_15009; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15011 = 12'ha60 == _T_146[11:0] ? image_2656 : _GEN_15010; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15012 = 12'ha61 == _T_146[11:0] ? image_2657 : _GEN_15011; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15013 = 12'ha62 == _T_146[11:0] ? image_2658 : _GEN_15012; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15014 = 12'ha63 == _T_146[11:0] ? image_2659 : _GEN_15013; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15015 = 12'ha64 == _T_146[11:0] ? image_2660 : _GEN_15014; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15016 = 12'ha65 == _T_146[11:0] ? image_2661 : _GEN_15015; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15017 = 12'ha66 == _T_146[11:0] ? image_2662 : _GEN_15016; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15018 = 12'ha67 == _T_146[11:0] ? image_2663 : _GEN_15017; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15019 = 12'ha68 == _T_146[11:0] ? image_2664 : _GEN_15018; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15020 = 12'ha69 == _T_146[11:0] ? image_2665 : _GEN_15019; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15021 = 12'ha6a == _T_146[11:0] ? image_2666 : _GEN_15020; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15022 = 12'ha6b == _T_146[11:0] ? image_2667 : _GEN_15021; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15023 = 12'ha6c == _T_146[11:0] ? image_2668 : _GEN_15022; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15024 = 12'ha6d == _T_146[11:0] ? image_2669 : _GEN_15023; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15025 = 12'ha6e == _T_146[11:0] ? image_2670 : _GEN_15024; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15026 = 12'ha6f == _T_146[11:0] ? image_2671 : _GEN_15025; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15027 = 12'ha70 == _T_146[11:0] ? image_2672 : _GEN_15026; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15028 = 12'ha71 == _T_146[11:0] ? image_2673 : _GEN_15027; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15029 = 12'ha72 == _T_146[11:0] ? image_2674 : _GEN_15028; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15030 = 12'ha73 == _T_146[11:0] ? image_2675 : _GEN_15029; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15031 = 12'ha74 == _T_146[11:0] ? image_2676 : _GEN_15030; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15032 = 12'ha75 == _T_146[11:0] ? image_2677 : _GEN_15031; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15033 = 12'ha76 == _T_146[11:0] ? image_2678 : _GEN_15032; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15034 = 12'ha77 == _T_146[11:0] ? image_2679 : _GEN_15033; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15035 = 12'ha78 == _T_146[11:0] ? image_2680 : _GEN_15034; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15036 = 12'ha79 == _T_146[11:0] ? image_2681 : _GEN_15035; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15037 = 12'ha7a == _T_146[11:0] ? image_2682 : _GEN_15036; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15038 = 12'ha7b == _T_146[11:0] ? 4'h0 : _GEN_15037; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15039 = 12'ha7c == _T_146[11:0] ? 4'h0 : _GEN_15038; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15040 = 12'ha7d == _T_146[11:0] ? 4'h0 : _GEN_15039; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15041 = 12'ha7e == _T_146[11:0] ? 4'h0 : _GEN_15040; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15042 = 12'ha7f == _T_146[11:0] ? 4'h0 : _GEN_15041; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15043 = 12'ha80 == _T_146[11:0] ? 4'h0 : _GEN_15042; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15044 = 12'ha81 == _T_146[11:0] ? 4'h0 : _GEN_15043; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15045 = 12'ha82 == _T_146[11:0] ? 4'h0 : _GEN_15044; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15046 = 12'ha83 == _T_146[11:0] ? 4'h0 : _GEN_15045; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15047 = 12'ha84 == _T_146[11:0] ? 4'h0 : _GEN_15046; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15048 = 12'ha85 == _T_146[11:0] ? 4'h0 : _GEN_15047; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15049 = 12'ha86 == _T_146[11:0] ? 4'h0 : _GEN_15048; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15050 = 12'ha87 == _T_146[11:0] ? 4'h0 : _GEN_15049; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15051 = 12'ha88 == _T_146[11:0] ? 4'h0 : _GEN_15050; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15052 = 12'ha89 == _T_146[11:0] ? image_2697 : _GEN_15051; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15053 = 12'ha8a == _T_146[11:0] ? image_2698 : _GEN_15052; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15054 = 12'ha8b == _T_146[11:0] ? image_2699 : _GEN_15053; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15055 = 12'ha8c == _T_146[11:0] ? image_2700 : _GEN_15054; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15056 = 12'ha8d == _T_146[11:0] ? image_2701 : _GEN_15055; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15057 = 12'ha8e == _T_146[11:0] ? image_2702 : _GEN_15056; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15058 = 12'ha8f == _T_146[11:0] ? image_2703 : _GEN_15057; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15059 = 12'ha90 == _T_146[11:0] ? image_2704 : _GEN_15058; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15060 = 12'ha91 == _T_146[11:0] ? image_2705 : _GEN_15059; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15061 = 12'ha92 == _T_146[11:0] ? image_2706 : _GEN_15060; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15062 = 12'ha93 == _T_146[11:0] ? image_2707 : _GEN_15061; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15063 = 12'ha94 == _T_146[11:0] ? image_2708 : _GEN_15062; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15064 = 12'ha95 == _T_146[11:0] ? image_2709 : _GEN_15063; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15065 = 12'ha96 == _T_146[11:0] ? image_2710 : _GEN_15064; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15066 = 12'ha97 == _T_146[11:0] ? image_2711 : _GEN_15065; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15067 = 12'ha98 == _T_146[11:0] ? image_2712 : _GEN_15066; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15068 = 12'ha99 == _T_146[11:0] ? image_2713 : _GEN_15067; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15069 = 12'ha9a == _T_146[11:0] ? image_2714 : _GEN_15068; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15070 = 12'ha9b == _T_146[11:0] ? image_2715 : _GEN_15069; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15071 = 12'ha9c == _T_146[11:0] ? image_2716 : _GEN_15070; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15072 = 12'ha9d == _T_146[11:0] ? image_2717 : _GEN_15071; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15073 = 12'ha9e == _T_146[11:0] ? image_2718 : _GEN_15072; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15074 = 12'ha9f == _T_146[11:0] ? image_2719 : _GEN_15073; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15075 = 12'haa0 == _T_146[11:0] ? image_2720 : _GEN_15074; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15076 = 12'haa1 == _T_146[11:0] ? image_2721 : _GEN_15075; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15077 = 12'haa2 == _T_146[11:0] ? image_2722 : _GEN_15076; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15078 = 12'haa3 == _T_146[11:0] ? image_2723 : _GEN_15077; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15079 = 12'haa4 == _T_146[11:0] ? image_2724 : _GEN_15078; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15080 = 12'haa5 == _T_146[11:0] ? image_2725 : _GEN_15079; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15081 = 12'haa6 == _T_146[11:0] ? image_2726 : _GEN_15080; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15082 = 12'haa7 == _T_146[11:0] ? image_2727 : _GEN_15081; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15083 = 12'haa8 == _T_146[11:0] ? image_2728 : _GEN_15082; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15084 = 12'haa9 == _T_146[11:0] ? image_2729 : _GEN_15083; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15085 = 12'haaa == _T_146[11:0] ? image_2730 : _GEN_15084; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15086 = 12'haab == _T_146[11:0] ? image_2731 : _GEN_15085; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15087 = 12'haac == _T_146[11:0] ? image_2732 : _GEN_15086; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15088 = 12'haad == _T_146[11:0] ? image_2733 : _GEN_15087; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15089 = 12'haae == _T_146[11:0] ? image_2734 : _GEN_15088; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15090 = 12'haaf == _T_146[11:0] ? image_2735 : _GEN_15089; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15091 = 12'hab0 == _T_146[11:0] ? image_2736 : _GEN_15090; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15092 = 12'hab1 == _T_146[11:0] ? image_2737 : _GEN_15091; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15093 = 12'hab2 == _T_146[11:0] ? image_2738 : _GEN_15092; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15094 = 12'hab3 == _T_146[11:0] ? image_2739 : _GEN_15093; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15095 = 12'hab4 == _T_146[11:0] ? image_2740 : _GEN_15094; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15096 = 12'hab5 == _T_146[11:0] ? image_2741 : _GEN_15095; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15097 = 12'hab6 == _T_146[11:0] ? image_2742 : _GEN_15096; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15098 = 12'hab7 == _T_146[11:0] ? image_2743 : _GEN_15097; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15099 = 12'hab8 == _T_146[11:0] ? image_2744 : _GEN_15098; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15100 = 12'hab9 == _T_146[11:0] ? image_2745 : _GEN_15099; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15101 = 12'haba == _T_146[11:0] ? 4'h0 : _GEN_15100; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15102 = 12'habb == _T_146[11:0] ? 4'h0 : _GEN_15101; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15103 = 12'habc == _T_146[11:0] ? 4'h0 : _GEN_15102; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15104 = 12'habd == _T_146[11:0] ? 4'h0 : _GEN_15103; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15105 = 12'habe == _T_146[11:0] ? 4'h0 : _GEN_15104; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15106 = 12'habf == _T_146[11:0] ? 4'h0 : _GEN_15105; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15107 = 12'hac0 == _T_146[11:0] ? 4'h0 : _GEN_15106; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15108 = 12'hac1 == _T_146[11:0] ? 4'h0 : _GEN_15107; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15109 = 12'hac2 == _T_146[11:0] ? 4'h0 : _GEN_15108; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15110 = 12'hac3 == _T_146[11:0] ? 4'h0 : _GEN_15109; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15111 = 12'hac4 == _T_146[11:0] ? 4'h0 : _GEN_15110; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15112 = 12'hac5 == _T_146[11:0] ? 4'h0 : _GEN_15111; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15113 = 12'hac6 == _T_146[11:0] ? 4'h0 : _GEN_15112; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15114 = 12'hac7 == _T_146[11:0] ? 4'h0 : _GEN_15113; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15115 = 12'hac8 == _T_146[11:0] ? 4'h0 : _GEN_15114; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15116 = 12'hac9 == _T_146[11:0] ? 4'h0 : _GEN_15115; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15117 = 12'haca == _T_146[11:0] ? 4'h0 : _GEN_15116; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15118 = 12'hacb == _T_146[11:0] ? image_2763 : _GEN_15117; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15119 = 12'hacc == _T_146[11:0] ? image_2764 : _GEN_15118; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15120 = 12'hacd == _T_146[11:0] ? image_2765 : _GEN_15119; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15121 = 12'hace == _T_146[11:0] ? image_2766 : _GEN_15120; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15122 = 12'hacf == _T_146[11:0] ? image_2767 : _GEN_15121; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15123 = 12'had0 == _T_146[11:0] ? image_2768 : _GEN_15122; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15124 = 12'had1 == _T_146[11:0] ? image_2769 : _GEN_15123; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15125 = 12'had2 == _T_146[11:0] ? image_2770 : _GEN_15124; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15126 = 12'had3 == _T_146[11:0] ? image_2771 : _GEN_15125; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15127 = 12'had4 == _T_146[11:0] ? image_2772 : _GEN_15126; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15128 = 12'had5 == _T_146[11:0] ? image_2773 : _GEN_15127; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15129 = 12'had6 == _T_146[11:0] ? image_2774 : _GEN_15128; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15130 = 12'had7 == _T_146[11:0] ? image_2775 : _GEN_15129; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15131 = 12'had8 == _T_146[11:0] ? image_2776 : _GEN_15130; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15132 = 12'had9 == _T_146[11:0] ? image_2777 : _GEN_15131; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15133 = 12'hada == _T_146[11:0] ? image_2778 : _GEN_15132; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15134 = 12'hadb == _T_146[11:0] ? image_2779 : _GEN_15133; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15135 = 12'hadc == _T_146[11:0] ? image_2780 : _GEN_15134; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15136 = 12'hadd == _T_146[11:0] ? image_2781 : _GEN_15135; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15137 = 12'hade == _T_146[11:0] ? image_2782 : _GEN_15136; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15138 = 12'hadf == _T_146[11:0] ? image_2783 : _GEN_15137; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15139 = 12'hae0 == _T_146[11:0] ? image_2784 : _GEN_15138; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15140 = 12'hae1 == _T_146[11:0] ? image_2785 : _GEN_15139; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15141 = 12'hae2 == _T_146[11:0] ? image_2786 : _GEN_15140; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15142 = 12'hae3 == _T_146[11:0] ? image_2787 : _GEN_15141; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15143 = 12'hae4 == _T_146[11:0] ? image_2788 : _GEN_15142; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15144 = 12'hae5 == _T_146[11:0] ? image_2789 : _GEN_15143; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15145 = 12'hae6 == _T_146[11:0] ? image_2790 : _GEN_15144; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15146 = 12'hae7 == _T_146[11:0] ? image_2791 : _GEN_15145; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15147 = 12'hae8 == _T_146[11:0] ? image_2792 : _GEN_15146; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15148 = 12'hae9 == _T_146[11:0] ? image_2793 : _GEN_15147; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15149 = 12'haea == _T_146[11:0] ? image_2794 : _GEN_15148; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15150 = 12'haeb == _T_146[11:0] ? image_2795 : _GEN_15149; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15151 = 12'haec == _T_146[11:0] ? image_2796 : _GEN_15150; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15152 = 12'haed == _T_146[11:0] ? image_2797 : _GEN_15151; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15153 = 12'haee == _T_146[11:0] ? image_2798 : _GEN_15152; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15154 = 12'haef == _T_146[11:0] ? image_2799 : _GEN_15153; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15155 = 12'haf0 == _T_146[11:0] ? image_2800 : _GEN_15154; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15156 = 12'haf1 == _T_146[11:0] ? image_2801 : _GEN_15155; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15157 = 12'haf2 == _T_146[11:0] ? image_2802 : _GEN_15156; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15158 = 12'haf3 == _T_146[11:0] ? image_2803 : _GEN_15157; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15159 = 12'haf4 == _T_146[11:0] ? image_2804 : _GEN_15158; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15160 = 12'haf5 == _T_146[11:0] ? image_2805 : _GEN_15159; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15161 = 12'haf6 == _T_146[11:0] ? image_2806 : _GEN_15160; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15162 = 12'haf7 == _T_146[11:0] ? image_2807 : _GEN_15161; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15163 = 12'haf8 == _T_146[11:0] ? image_2808 : _GEN_15162; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15164 = 12'haf9 == _T_146[11:0] ? 4'h0 : _GEN_15163; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15165 = 12'hafa == _T_146[11:0] ? 4'h0 : _GEN_15164; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15166 = 12'hafb == _T_146[11:0] ? 4'h0 : _GEN_15165; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15167 = 12'hafc == _T_146[11:0] ? 4'h0 : _GEN_15166; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15168 = 12'hafd == _T_146[11:0] ? 4'h0 : _GEN_15167; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15169 = 12'hafe == _T_146[11:0] ? 4'h0 : _GEN_15168; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15170 = 12'haff == _T_146[11:0] ? 4'h0 : _GEN_15169; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15171 = 12'hb00 == _T_146[11:0] ? 4'h0 : _GEN_15170; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15172 = 12'hb01 == _T_146[11:0] ? 4'h0 : _GEN_15171; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15173 = 12'hb02 == _T_146[11:0] ? 4'h0 : _GEN_15172; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15174 = 12'hb03 == _T_146[11:0] ? 4'h0 : _GEN_15173; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15175 = 12'hb04 == _T_146[11:0] ? 4'h0 : _GEN_15174; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15176 = 12'hb05 == _T_146[11:0] ? 4'h0 : _GEN_15175; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15177 = 12'hb06 == _T_146[11:0] ? 4'h0 : _GEN_15176; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15178 = 12'hb07 == _T_146[11:0] ? 4'h0 : _GEN_15177; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15179 = 12'hb08 == _T_146[11:0] ? 4'h0 : _GEN_15178; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15180 = 12'hb09 == _T_146[11:0] ? 4'h0 : _GEN_15179; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15181 = 12'hb0a == _T_146[11:0] ? 4'h0 : _GEN_15180; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15182 = 12'hb0b == _T_146[11:0] ? 4'h0 : _GEN_15181; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15183 = 12'hb0c == _T_146[11:0] ? image_2828 : _GEN_15182; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15184 = 12'hb0d == _T_146[11:0] ? image_2829 : _GEN_15183; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15185 = 12'hb0e == _T_146[11:0] ? image_2830 : _GEN_15184; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15186 = 12'hb0f == _T_146[11:0] ? image_2831 : _GEN_15185; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15187 = 12'hb10 == _T_146[11:0] ? image_2832 : _GEN_15186; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15188 = 12'hb11 == _T_146[11:0] ? image_2833 : _GEN_15187; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15189 = 12'hb12 == _T_146[11:0] ? image_2834 : _GEN_15188; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15190 = 12'hb13 == _T_146[11:0] ? image_2835 : _GEN_15189; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15191 = 12'hb14 == _T_146[11:0] ? image_2836 : _GEN_15190; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15192 = 12'hb15 == _T_146[11:0] ? image_2837 : _GEN_15191; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15193 = 12'hb16 == _T_146[11:0] ? image_2838 : _GEN_15192; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15194 = 12'hb17 == _T_146[11:0] ? image_2839 : _GEN_15193; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15195 = 12'hb18 == _T_146[11:0] ? image_2840 : _GEN_15194; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15196 = 12'hb19 == _T_146[11:0] ? image_2841 : _GEN_15195; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15197 = 12'hb1a == _T_146[11:0] ? image_2842 : _GEN_15196; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15198 = 12'hb1b == _T_146[11:0] ? image_2843 : _GEN_15197; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15199 = 12'hb1c == _T_146[11:0] ? image_2844 : _GEN_15198; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15200 = 12'hb1d == _T_146[11:0] ? image_2845 : _GEN_15199; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15201 = 12'hb1e == _T_146[11:0] ? image_2846 : _GEN_15200; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15202 = 12'hb1f == _T_146[11:0] ? image_2847 : _GEN_15201; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15203 = 12'hb20 == _T_146[11:0] ? image_2848 : _GEN_15202; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15204 = 12'hb21 == _T_146[11:0] ? image_2849 : _GEN_15203; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15205 = 12'hb22 == _T_146[11:0] ? image_2850 : _GEN_15204; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15206 = 12'hb23 == _T_146[11:0] ? image_2851 : _GEN_15205; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15207 = 12'hb24 == _T_146[11:0] ? image_2852 : _GEN_15206; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15208 = 12'hb25 == _T_146[11:0] ? image_2853 : _GEN_15207; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15209 = 12'hb26 == _T_146[11:0] ? image_2854 : _GEN_15208; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15210 = 12'hb27 == _T_146[11:0] ? image_2855 : _GEN_15209; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15211 = 12'hb28 == _T_146[11:0] ? image_2856 : _GEN_15210; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15212 = 12'hb29 == _T_146[11:0] ? image_2857 : _GEN_15211; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15213 = 12'hb2a == _T_146[11:0] ? image_2858 : _GEN_15212; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15214 = 12'hb2b == _T_146[11:0] ? image_2859 : _GEN_15213; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15215 = 12'hb2c == _T_146[11:0] ? image_2860 : _GEN_15214; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15216 = 12'hb2d == _T_146[11:0] ? image_2861 : _GEN_15215; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15217 = 12'hb2e == _T_146[11:0] ? image_2862 : _GEN_15216; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15218 = 12'hb2f == _T_146[11:0] ? image_2863 : _GEN_15217; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15219 = 12'hb30 == _T_146[11:0] ? image_2864 : _GEN_15218; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15220 = 12'hb31 == _T_146[11:0] ? image_2865 : _GEN_15219; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15221 = 12'hb32 == _T_146[11:0] ? image_2866 : _GEN_15220; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15222 = 12'hb33 == _T_146[11:0] ? image_2867 : _GEN_15221; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15223 = 12'hb34 == _T_146[11:0] ? image_2868 : _GEN_15222; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15224 = 12'hb35 == _T_146[11:0] ? image_2869 : _GEN_15223; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15225 = 12'hb36 == _T_146[11:0] ? image_2870 : _GEN_15224; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15226 = 12'hb37 == _T_146[11:0] ? image_2871 : _GEN_15225; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15227 = 12'hb38 == _T_146[11:0] ? 4'h0 : _GEN_15226; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15228 = 12'hb39 == _T_146[11:0] ? 4'h0 : _GEN_15227; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15229 = 12'hb3a == _T_146[11:0] ? 4'h0 : _GEN_15228; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15230 = 12'hb3b == _T_146[11:0] ? 4'h0 : _GEN_15229; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15231 = 12'hb3c == _T_146[11:0] ? 4'h0 : _GEN_15230; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15232 = 12'hb3d == _T_146[11:0] ? 4'h0 : _GEN_15231; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15233 = 12'hb3e == _T_146[11:0] ? 4'h0 : _GEN_15232; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15234 = 12'hb3f == _T_146[11:0] ? 4'h0 : _GEN_15233; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15235 = 12'hb40 == _T_146[11:0] ? 4'h0 : _GEN_15234; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15236 = 12'hb41 == _T_146[11:0] ? 4'h0 : _GEN_15235; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15237 = 12'hb42 == _T_146[11:0] ? 4'h0 : _GEN_15236; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15238 = 12'hb43 == _T_146[11:0] ? 4'h0 : _GEN_15237; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15239 = 12'hb44 == _T_146[11:0] ? 4'h0 : _GEN_15238; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15240 = 12'hb45 == _T_146[11:0] ? 4'h0 : _GEN_15239; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15241 = 12'hb46 == _T_146[11:0] ? 4'h0 : _GEN_15240; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15242 = 12'hb47 == _T_146[11:0] ? 4'h0 : _GEN_15241; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15243 = 12'hb48 == _T_146[11:0] ? 4'h0 : _GEN_15242; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15244 = 12'hb49 == _T_146[11:0] ? 4'h0 : _GEN_15243; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15245 = 12'hb4a == _T_146[11:0] ? 4'h0 : _GEN_15244; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15246 = 12'hb4b == _T_146[11:0] ? 4'h0 : _GEN_15245; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15247 = 12'hb4c == _T_146[11:0] ? 4'h0 : _GEN_15246; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15248 = 12'hb4d == _T_146[11:0] ? 4'h0 : _GEN_15247; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15249 = 12'hb4e == _T_146[11:0] ? 4'h0 : _GEN_15248; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15250 = 12'hb4f == _T_146[11:0] ? image_2895 : _GEN_15249; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15251 = 12'hb50 == _T_146[11:0] ? image_2896 : _GEN_15250; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15252 = 12'hb51 == _T_146[11:0] ? image_2897 : _GEN_15251; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15253 = 12'hb52 == _T_146[11:0] ? image_2898 : _GEN_15252; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15254 = 12'hb53 == _T_146[11:0] ? image_2899 : _GEN_15253; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15255 = 12'hb54 == _T_146[11:0] ? image_2900 : _GEN_15254; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15256 = 12'hb55 == _T_146[11:0] ? image_2901 : _GEN_15255; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15257 = 12'hb56 == _T_146[11:0] ? image_2902 : _GEN_15256; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15258 = 12'hb57 == _T_146[11:0] ? image_2903 : _GEN_15257; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15259 = 12'hb58 == _T_146[11:0] ? image_2904 : _GEN_15258; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15260 = 12'hb59 == _T_146[11:0] ? image_2905 : _GEN_15259; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15261 = 12'hb5a == _T_146[11:0] ? image_2906 : _GEN_15260; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15262 = 12'hb5b == _T_146[11:0] ? image_2907 : _GEN_15261; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15263 = 12'hb5c == _T_146[11:0] ? image_2908 : _GEN_15262; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15264 = 12'hb5d == _T_146[11:0] ? image_2909 : _GEN_15263; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15265 = 12'hb5e == _T_146[11:0] ? image_2910 : _GEN_15264; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15266 = 12'hb5f == _T_146[11:0] ? image_2911 : _GEN_15265; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15267 = 12'hb60 == _T_146[11:0] ? image_2912 : _GEN_15266; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15268 = 12'hb61 == _T_146[11:0] ? image_2913 : _GEN_15267; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15269 = 12'hb62 == _T_146[11:0] ? image_2914 : _GEN_15268; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15270 = 12'hb63 == _T_146[11:0] ? image_2915 : _GEN_15269; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15271 = 12'hb64 == _T_146[11:0] ? image_2916 : _GEN_15270; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15272 = 12'hb65 == _T_146[11:0] ? image_2917 : _GEN_15271; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15273 = 12'hb66 == _T_146[11:0] ? image_2918 : _GEN_15272; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15274 = 12'hb67 == _T_146[11:0] ? image_2919 : _GEN_15273; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15275 = 12'hb68 == _T_146[11:0] ? image_2920 : _GEN_15274; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15276 = 12'hb69 == _T_146[11:0] ? image_2921 : _GEN_15275; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15277 = 12'hb6a == _T_146[11:0] ? image_2922 : _GEN_15276; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15278 = 12'hb6b == _T_146[11:0] ? image_2923 : _GEN_15277; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15279 = 12'hb6c == _T_146[11:0] ? image_2924 : _GEN_15278; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15280 = 12'hb6d == _T_146[11:0] ? image_2925 : _GEN_15279; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15281 = 12'hb6e == _T_146[11:0] ? image_2926 : _GEN_15280; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15282 = 12'hb6f == _T_146[11:0] ? image_2927 : _GEN_15281; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15283 = 12'hb70 == _T_146[11:0] ? image_2928 : _GEN_15282; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15284 = 12'hb71 == _T_146[11:0] ? image_2929 : _GEN_15283; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15285 = 12'hb72 == _T_146[11:0] ? image_2930 : _GEN_15284; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15286 = 12'hb73 == _T_146[11:0] ? image_2931 : _GEN_15285; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15287 = 12'hb74 == _T_146[11:0] ? image_2932 : _GEN_15286; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15288 = 12'hb75 == _T_146[11:0] ? image_2933 : _GEN_15287; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15289 = 12'hb76 == _T_146[11:0] ? image_2934 : _GEN_15288; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15290 = 12'hb77 == _T_146[11:0] ? 4'h0 : _GEN_15289; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15291 = 12'hb78 == _T_146[11:0] ? 4'h0 : _GEN_15290; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15292 = 12'hb79 == _T_146[11:0] ? 4'h0 : _GEN_15291; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15293 = 12'hb7a == _T_146[11:0] ? 4'h0 : _GEN_15292; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15294 = 12'hb7b == _T_146[11:0] ? 4'h0 : _GEN_15293; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15295 = 12'hb7c == _T_146[11:0] ? 4'h0 : _GEN_15294; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15296 = 12'hb7d == _T_146[11:0] ? 4'h0 : _GEN_15295; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15297 = 12'hb7e == _T_146[11:0] ? 4'h0 : _GEN_15296; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15298 = 12'hb7f == _T_146[11:0] ? 4'h0 : _GEN_15297; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15299 = 12'hb80 == _T_146[11:0] ? 4'h0 : _GEN_15298; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15300 = 12'hb81 == _T_146[11:0] ? 4'h0 : _GEN_15299; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15301 = 12'hb82 == _T_146[11:0] ? 4'h0 : _GEN_15300; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15302 = 12'hb83 == _T_146[11:0] ? 4'h0 : _GEN_15301; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15303 = 12'hb84 == _T_146[11:0] ? 4'h0 : _GEN_15302; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15304 = 12'hb85 == _T_146[11:0] ? 4'h0 : _GEN_15303; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15305 = 12'hb86 == _T_146[11:0] ? 4'h0 : _GEN_15304; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15306 = 12'hb87 == _T_146[11:0] ? 4'h0 : _GEN_15305; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15307 = 12'hb88 == _T_146[11:0] ? 4'h0 : _GEN_15306; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15308 = 12'hb89 == _T_146[11:0] ? 4'h0 : _GEN_15307; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15309 = 12'hb8a == _T_146[11:0] ? 4'h0 : _GEN_15308; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15310 = 12'hb8b == _T_146[11:0] ? 4'h0 : _GEN_15309; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15311 = 12'hb8c == _T_146[11:0] ? 4'h0 : _GEN_15310; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15312 = 12'hb8d == _T_146[11:0] ? 4'h0 : _GEN_15311; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15313 = 12'hb8e == _T_146[11:0] ? 4'h0 : _GEN_15312; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15314 = 12'hb8f == _T_146[11:0] ? 4'h0 : _GEN_15313; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15315 = 12'hb90 == _T_146[11:0] ? 4'h0 : _GEN_15314; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15316 = 12'hb91 == _T_146[11:0] ? 4'h0 : _GEN_15315; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15317 = 12'hb92 == _T_146[11:0] ? 4'h0 : _GEN_15316; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15318 = 12'hb93 == _T_146[11:0] ? 4'h0 : _GEN_15317; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15319 = 12'hb94 == _T_146[11:0] ? 4'h0 : _GEN_15318; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15320 = 12'hb95 == _T_146[11:0] ? image_2965 : _GEN_15319; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15321 = 12'hb96 == _T_146[11:0] ? image_2966 : _GEN_15320; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15322 = 12'hb97 == _T_146[11:0] ? image_2967 : _GEN_15321; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15323 = 12'hb98 == _T_146[11:0] ? image_2968 : _GEN_15322; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15324 = 12'hb99 == _T_146[11:0] ? image_2969 : _GEN_15323; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15325 = 12'hb9a == _T_146[11:0] ? image_2970 : _GEN_15324; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15326 = 12'hb9b == _T_146[11:0] ? image_2971 : _GEN_15325; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15327 = 12'hb9c == _T_146[11:0] ? image_2972 : _GEN_15326; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15328 = 12'hb9d == _T_146[11:0] ? image_2973 : _GEN_15327; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15329 = 12'hb9e == _T_146[11:0] ? image_2974 : _GEN_15328; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15330 = 12'hb9f == _T_146[11:0] ? image_2975 : _GEN_15329; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15331 = 12'hba0 == _T_146[11:0] ? image_2976 : _GEN_15330; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15332 = 12'hba1 == _T_146[11:0] ? image_2977 : _GEN_15331; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15333 = 12'hba2 == _T_146[11:0] ? image_2978 : _GEN_15332; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15334 = 12'hba3 == _T_146[11:0] ? image_2979 : _GEN_15333; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15335 = 12'hba4 == _T_146[11:0] ? image_2980 : _GEN_15334; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15336 = 12'hba5 == _T_146[11:0] ? image_2981 : _GEN_15335; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15337 = 12'hba6 == _T_146[11:0] ? image_2982 : _GEN_15336; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15338 = 12'hba7 == _T_146[11:0] ? image_2983 : _GEN_15337; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15339 = 12'hba8 == _T_146[11:0] ? image_2984 : _GEN_15338; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15340 = 12'hba9 == _T_146[11:0] ? image_2985 : _GEN_15339; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15341 = 12'hbaa == _T_146[11:0] ? image_2986 : _GEN_15340; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15342 = 12'hbab == _T_146[11:0] ? image_2987 : _GEN_15341; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15343 = 12'hbac == _T_146[11:0] ? image_2988 : _GEN_15342; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15344 = 12'hbad == _T_146[11:0] ? image_2989 : _GEN_15343; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15345 = 12'hbae == _T_146[11:0] ? image_2990 : _GEN_15344; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15346 = 12'hbaf == _T_146[11:0] ? image_2991 : _GEN_15345; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15347 = 12'hbb0 == _T_146[11:0] ? image_2992 : _GEN_15346; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15348 = 12'hbb1 == _T_146[11:0] ? image_2993 : _GEN_15347; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15349 = 12'hbb2 == _T_146[11:0] ? image_2994 : _GEN_15348; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15350 = 12'hbb3 == _T_146[11:0] ? image_2995 : _GEN_15349; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15351 = 12'hbb4 == _T_146[11:0] ? image_2996 : _GEN_15350; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15352 = 12'hbb5 == _T_146[11:0] ? 4'h0 : _GEN_15351; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15353 = 12'hbb6 == _T_146[11:0] ? 4'h0 : _GEN_15352; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15354 = 12'hbb7 == _T_146[11:0] ? 4'h0 : _GEN_15353; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15355 = 12'hbb8 == _T_146[11:0] ? 4'h0 : _GEN_15354; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15356 = 12'hbb9 == _T_146[11:0] ? 4'h0 : _GEN_15355; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15357 = 12'hbba == _T_146[11:0] ? 4'h0 : _GEN_15356; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15358 = 12'hbbb == _T_146[11:0] ? 4'h0 : _GEN_15357; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15359 = 12'hbbc == _T_146[11:0] ? 4'h0 : _GEN_15358; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15360 = 12'hbbd == _T_146[11:0] ? 4'h0 : _GEN_15359; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15361 = 12'hbbe == _T_146[11:0] ? 4'h0 : _GEN_15360; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15362 = 12'hbbf == _T_146[11:0] ? 4'h0 : _GEN_15361; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15363 = 12'hbc0 == _T_146[11:0] ? 4'h0 : _GEN_15362; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15364 = 12'hbc1 == _T_146[11:0] ? 4'h0 : _GEN_15363; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15365 = 12'hbc2 == _T_146[11:0] ? 4'h0 : _GEN_15364; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15366 = 12'hbc3 == _T_146[11:0] ? 4'h0 : _GEN_15365; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15367 = 12'hbc4 == _T_146[11:0] ? 4'h0 : _GEN_15366; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15368 = 12'hbc5 == _T_146[11:0] ? 4'h0 : _GEN_15367; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15369 = 12'hbc6 == _T_146[11:0] ? 4'h0 : _GEN_15368; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15370 = 12'hbc7 == _T_146[11:0] ? 4'h0 : _GEN_15369; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15371 = 12'hbc8 == _T_146[11:0] ? 4'h0 : _GEN_15370; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15372 = 12'hbc9 == _T_146[11:0] ? 4'h0 : _GEN_15371; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15373 = 12'hbca == _T_146[11:0] ? 4'h0 : _GEN_15372; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15374 = 12'hbcb == _T_146[11:0] ? 4'h0 : _GEN_15373; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15375 = 12'hbcc == _T_146[11:0] ? 4'h0 : _GEN_15374; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15376 = 12'hbcd == _T_146[11:0] ? 4'h0 : _GEN_15375; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15377 = 12'hbce == _T_146[11:0] ? 4'h0 : _GEN_15376; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15378 = 12'hbcf == _T_146[11:0] ? 4'h0 : _GEN_15377; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15379 = 12'hbd0 == _T_146[11:0] ? 4'h0 : _GEN_15378; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15380 = 12'hbd1 == _T_146[11:0] ? 4'h0 : _GEN_15379; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15381 = 12'hbd2 == _T_146[11:0] ? 4'h0 : _GEN_15380; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15382 = 12'hbd3 == _T_146[11:0] ? 4'h0 : _GEN_15381; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15383 = 12'hbd4 == _T_146[11:0] ? 4'h0 : _GEN_15382; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15384 = 12'hbd5 == _T_146[11:0] ? 4'h0 : _GEN_15383; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15385 = 12'hbd6 == _T_146[11:0] ? 4'h0 : _GEN_15384; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15386 = 12'hbd7 == _T_146[11:0] ? 4'h0 : _GEN_15385; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15387 = 12'hbd8 == _T_146[11:0] ? 4'h0 : _GEN_15386; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15388 = 12'hbd9 == _T_146[11:0] ? 4'h0 : _GEN_15387; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15389 = 12'hbda == _T_146[11:0] ? 4'h0 : _GEN_15388; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15390 = 12'hbdb == _T_146[11:0] ? image_3035 : _GEN_15389; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15391 = 12'hbdc == _T_146[11:0] ? image_3036 : _GEN_15390; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15392 = 12'hbdd == _T_146[11:0] ? image_3037 : _GEN_15391; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15393 = 12'hbde == _T_146[11:0] ? image_3038 : _GEN_15392; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15394 = 12'hbdf == _T_146[11:0] ? image_3039 : _GEN_15393; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15395 = 12'hbe0 == _T_146[11:0] ? image_3040 : _GEN_15394; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15396 = 12'hbe1 == _T_146[11:0] ? image_3041 : _GEN_15395; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15397 = 12'hbe2 == _T_146[11:0] ? image_3042 : _GEN_15396; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15398 = 12'hbe3 == _T_146[11:0] ? image_3043 : _GEN_15397; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15399 = 12'hbe4 == _T_146[11:0] ? image_3044 : _GEN_15398; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15400 = 12'hbe5 == _T_146[11:0] ? image_3045 : _GEN_15399; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15401 = 12'hbe6 == _T_146[11:0] ? image_3046 : _GEN_15400; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15402 = 12'hbe7 == _T_146[11:0] ? image_3047 : _GEN_15401; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15403 = 12'hbe8 == _T_146[11:0] ? image_3048 : _GEN_15402; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15404 = 12'hbe9 == _T_146[11:0] ? image_3049 : _GEN_15403; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15405 = 12'hbea == _T_146[11:0] ? image_3050 : _GEN_15404; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15406 = 12'hbeb == _T_146[11:0] ? image_3051 : _GEN_15405; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15407 = 12'hbec == _T_146[11:0] ? image_3052 : _GEN_15406; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15408 = 12'hbed == _T_146[11:0] ? image_3053 : _GEN_15407; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15409 = 12'hbee == _T_146[11:0] ? image_3054 : _GEN_15408; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15410 = 12'hbef == _T_146[11:0] ? image_3055 : _GEN_15409; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15411 = 12'hbf0 == _T_146[11:0] ? image_3056 : _GEN_15410; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15412 = 12'hbf1 == _T_146[11:0] ? 4'h0 : _GEN_15411; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15413 = 12'hbf2 == _T_146[11:0] ? 4'h0 : _GEN_15412; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15414 = 12'hbf3 == _T_146[11:0] ? 4'h0 : _GEN_15413; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15415 = 12'hbf4 == _T_146[11:0] ? 4'h0 : _GEN_15414; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15416 = 12'hbf5 == _T_146[11:0] ? 4'h0 : _GEN_15415; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15417 = 12'hbf6 == _T_146[11:0] ? 4'h0 : _GEN_15416; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15418 = 12'hbf7 == _T_146[11:0] ? 4'h0 : _GEN_15417; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15419 = 12'hbf8 == _T_146[11:0] ? 4'h0 : _GEN_15418; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15420 = 12'hbf9 == _T_146[11:0] ? 4'h0 : _GEN_15419; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15421 = 12'hbfa == _T_146[11:0] ? 4'h0 : _GEN_15420; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15422 = 12'hbfb == _T_146[11:0] ? 4'h0 : _GEN_15421; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15423 = 12'hbfc == _T_146[11:0] ? 4'h0 : _GEN_15422; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15424 = 12'hbfd == _T_146[11:0] ? 4'h0 : _GEN_15423; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15425 = 12'hbfe == _T_146[11:0] ? 4'h0 : _GEN_15424; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15426 = 12'hbff == _T_146[11:0] ? 4'h0 : _GEN_15425; // @[Filter.scala 138:46]
  wire [31:0] _T_149 = pixelIndex + 32'h5; // @[Filter.scala 133:29]
  wire [31:0] _T_150 = _T_149 / 32'h40; // @[Filter.scala 133:36]
  wire [31:0] _T_152 = _T_150 + _GEN_24805; // @[Filter.scala 133:51]
  wire [31:0] _T_154 = _T_152 - 32'h1; // @[Filter.scala 133:67]
  wire [31:0] _GEN_5 = _T_149 % 32'h40; // @[Filter.scala 134:36]
  wire [6:0] _T_157 = _GEN_5[6:0]; // @[Filter.scala 134:36]
  wire [6:0] _T_159 = _T_157 + _GEN_24806; // @[Filter.scala 134:51]
  wire [6:0] _T_161 = _T_159 - 7'h1; // @[Filter.scala 134:67]
  wire  _T_163 = _T_154 >= 32'h40; // @[Filter.scala 135:27]
  wire  _T_167 = _T_161 >= 7'h30; // @[Filter.scala 135:59]
  wire  _T_168 = _T_163 | _T_167; // @[Filter.scala 135:54]
  wire [13:0] _T_169 = _T_161 * 7'h40; // @[Filter.scala 138:57]
  wire [31:0] _GEN_24822 = {{18'd0}, _T_169}; // @[Filter.scala 138:72]
  wire [31:0] _T_171 = _GEN_24822 + _T_154; // @[Filter.scala 138:72]
  wire [3:0] _GEN_15440 = 12'hc == _T_171[11:0] ? image_12 : 4'h0; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15441 = 12'hd == _T_171[11:0] ? 4'h0 : _GEN_15440; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15442 = 12'he == _T_171[11:0] ? image_14 : _GEN_15441; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15443 = 12'hf == _T_171[11:0] ? image_15 : _GEN_15442; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15444 = 12'h10 == _T_171[11:0] ? image_16 : _GEN_15443; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15445 = 12'h11 == _T_171[11:0] ? image_17 : _GEN_15444; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15446 = 12'h12 == _T_171[11:0] ? image_18 : _GEN_15445; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15447 = 12'h13 == _T_171[11:0] ? image_19 : _GEN_15446; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15448 = 12'h14 == _T_171[11:0] ? image_20 : _GEN_15447; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15449 = 12'h15 == _T_171[11:0] ? image_21 : _GEN_15448; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15450 = 12'h16 == _T_171[11:0] ? image_22 : _GEN_15449; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15451 = 12'h17 == _T_171[11:0] ? image_23 : _GEN_15450; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15452 = 12'h18 == _T_171[11:0] ? 4'h0 : _GEN_15451; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15453 = 12'h19 == _T_171[11:0] ? 4'h0 : _GEN_15452; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15454 = 12'h1a == _T_171[11:0] ? 4'h0 : _GEN_15453; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15455 = 12'h1b == _T_171[11:0] ? 4'h0 : _GEN_15454; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15456 = 12'h1c == _T_171[11:0] ? 4'h0 : _GEN_15455; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15457 = 12'h1d == _T_171[11:0] ? 4'h0 : _GEN_15456; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15458 = 12'h1e == _T_171[11:0] ? 4'h0 : _GEN_15457; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15459 = 12'h1f == _T_171[11:0] ? 4'h0 : _GEN_15458; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15460 = 12'h20 == _T_171[11:0] ? 4'h0 : _GEN_15459; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15461 = 12'h21 == _T_171[11:0] ? 4'h0 : _GEN_15460; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15462 = 12'h22 == _T_171[11:0] ? 4'h0 : _GEN_15461; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15463 = 12'h23 == _T_171[11:0] ? image_35 : _GEN_15462; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15464 = 12'h24 == _T_171[11:0] ? image_36 : _GEN_15463; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15465 = 12'h25 == _T_171[11:0] ? image_37 : _GEN_15464; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15466 = 12'h26 == _T_171[11:0] ? image_38 : _GEN_15465; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15467 = 12'h27 == _T_171[11:0] ? image_39 : _GEN_15466; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15468 = 12'h28 == _T_171[11:0] ? image_40 : _GEN_15467; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15469 = 12'h29 == _T_171[11:0] ? image_41 : _GEN_15468; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15470 = 12'h2a == _T_171[11:0] ? image_42 : _GEN_15469; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15471 = 12'h2b == _T_171[11:0] ? 4'h0 : _GEN_15470; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15472 = 12'h2c == _T_171[11:0] ? 4'h0 : _GEN_15471; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15473 = 12'h2d == _T_171[11:0] ? 4'h0 : _GEN_15472; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15474 = 12'h2e == _T_171[11:0] ? 4'h0 : _GEN_15473; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15475 = 12'h2f == _T_171[11:0] ? 4'h0 : _GEN_15474; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15476 = 12'h30 == _T_171[11:0] ? 4'h0 : _GEN_15475; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15477 = 12'h31 == _T_171[11:0] ? 4'h0 : _GEN_15476; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15478 = 12'h32 == _T_171[11:0] ? 4'h0 : _GEN_15477; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15479 = 12'h33 == _T_171[11:0] ? 4'h0 : _GEN_15478; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15480 = 12'h34 == _T_171[11:0] ? 4'h0 : _GEN_15479; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15481 = 12'h35 == _T_171[11:0] ? 4'h0 : _GEN_15480; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15482 = 12'h36 == _T_171[11:0] ? 4'h0 : _GEN_15481; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15483 = 12'h37 == _T_171[11:0] ? 4'h0 : _GEN_15482; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15484 = 12'h38 == _T_171[11:0] ? 4'h0 : _GEN_15483; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15485 = 12'h39 == _T_171[11:0] ? 4'h0 : _GEN_15484; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15486 = 12'h3a == _T_171[11:0] ? 4'h0 : _GEN_15485; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15487 = 12'h3b == _T_171[11:0] ? 4'h0 : _GEN_15486; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15488 = 12'h3c == _T_171[11:0] ? 4'h0 : _GEN_15487; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15489 = 12'h3d == _T_171[11:0] ? 4'h0 : _GEN_15488; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15490 = 12'h3e == _T_171[11:0] ? 4'h0 : _GEN_15489; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15491 = 12'h3f == _T_171[11:0] ? 4'h0 : _GEN_15490; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15492 = 12'h40 == _T_171[11:0] ? 4'h0 : _GEN_15491; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15493 = 12'h41 == _T_171[11:0] ? 4'h0 : _GEN_15492; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15494 = 12'h42 == _T_171[11:0] ? 4'h0 : _GEN_15493; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15495 = 12'h43 == _T_171[11:0] ? 4'h0 : _GEN_15494; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15496 = 12'h44 == _T_171[11:0] ? 4'h0 : _GEN_15495; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15497 = 12'h45 == _T_171[11:0] ? 4'h0 : _GEN_15496; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15498 = 12'h46 == _T_171[11:0] ? 4'h0 : _GEN_15497; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15499 = 12'h47 == _T_171[11:0] ? 4'h0 : _GEN_15498; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15500 = 12'h48 == _T_171[11:0] ? 4'h0 : _GEN_15499; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15501 = 12'h49 == _T_171[11:0] ? 4'h0 : _GEN_15500; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15502 = 12'h4a == _T_171[11:0] ? 4'h0 : _GEN_15501; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15503 = 12'h4b == _T_171[11:0] ? image_75 : _GEN_15502; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15504 = 12'h4c == _T_171[11:0] ? image_76 : _GEN_15503; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15505 = 12'h4d == _T_171[11:0] ? image_77 : _GEN_15504; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15506 = 12'h4e == _T_171[11:0] ? image_78 : _GEN_15505; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15507 = 12'h4f == _T_171[11:0] ? image_79 : _GEN_15506; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15508 = 12'h50 == _T_171[11:0] ? image_80 : _GEN_15507; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15509 = 12'h51 == _T_171[11:0] ? image_81 : _GEN_15508; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15510 = 12'h52 == _T_171[11:0] ? image_82 : _GEN_15509; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15511 = 12'h53 == _T_171[11:0] ? image_83 : _GEN_15510; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15512 = 12'h54 == _T_171[11:0] ? image_84 : _GEN_15511; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15513 = 12'h55 == _T_171[11:0] ? image_85 : _GEN_15512; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15514 = 12'h56 == _T_171[11:0] ? image_86 : _GEN_15513; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15515 = 12'h57 == _T_171[11:0] ? image_87 : _GEN_15514; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15516 = 12'h58 == _T_171[11:0] ? image_88 : _GEN_15515; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15517 = 12'h59 == _T_171[11:0] ? image_89 : _GEN_15516; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15518 = 12'h5a == _T_171[11:0] ? image_90 : _GEN_15517; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15519 = 12'h5b == _T_171[11:0] ? 4'h0 : _GEN_15518; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15520 = 12'h5c == _T_171[11:0] ? 4'h0 : _GEN_15519; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15521 = 12'h5d == _T_171[11:0] ? image_93 : _GEN_15520; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15522 = 12'h5e == _T_171[11:0] ? 4'h0 : _GEN_15521; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15523 = 12'h5f == _T_171[11:0] ? image_95 : _GEN_15522; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15524 = 12'h60 == _T_171[11:0] ? image_96 : _GEN_15523; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15525 = 12'h61 == _T_171[11:0] ? image_97 : _GEN_15524; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15526 = 12'h62 == _T_171[11:0] ? image_98 : _GEN_15525; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15527 = 12'h63 == _T_171[11:0] ? image_99 : _GEN_15526; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15528 = 12'h64 == _T_171[11:0] ? image_100 : _GEN_15527; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15529 = 12'h65 == _T_171[11:0] ? image_101 : _GEN_15528; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15530 = 12'h66 == _T_171[11:0] ? image_102 : _GEN_15529; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15531 = 12'h67 == _T_171[11:0] ? image_103 : _GEN_15530; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15532 = 12'h68 == _T_171[11:0] ? image_104 : _GEN_15531; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15533 = 12'h69 == _T_171[11:0] ? image_105 : _GEN_15532; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15534 = 12'h6a == _T_171[11:0] ? image_106 : _GEN_15533; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15535 = 12'h6b == _T_171[11:0] ? image_107 : _GEN_15534; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15536 = 12'h6c == _T_171[11:0] ? image_108 : _GEN_15535; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15537 = 12'h6d == _T_171[11:0] ? 4'h0 : _GEN_15536; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15538 = 12'h6e == _T_171[11:0] ? 4'h0 : _GEN_15537; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15539 = 12'h6f == _T_171[11:0] ? 4'h0 : _GEN_15538; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15540 = 12'h70 == _T_171[11:0] ? 4'h0 : _GEN_15539; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15541 = 12'h71 == _T_171[11:0] ? 4'h0 : _GEN_15540; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15542 = 12'h72 == _T_171[11:0] ? 4'h0 : _GEN_15541; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15543 = 12'h73 == _T_171[11:0] ? 4'h0 : _GEN_15542; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15544 = 12'h74 == _T_171[11:0] ? 4'h0 : _GEN_15543; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15545 = 12'h75 == _T_171[11:0] ? 4'h0 : _GEN_15544; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15546 = 12'h76 == _T_171[11:0] ? 4'h0 : _GEN_15545; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15547 = 12'h77 == _T_171[11:0] ? 4'h0 : _GEN_15546; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15548 = 12'h78 == _T_171[11:0] ? 4'h0 : _GEN_15547; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15549 = 12'h79 == _T_171[11:0] ? 4'h0 : _GEN_15548; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15550 = 12'h7a == _T_171[11:0] ? 4'h0 : _GEN_15549; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15551 = 12'h7b == _T_171[11:0] ? 4'h0 : _GEN_15550; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15552 = 12'h7c == _T_171[11:0] ? 4'h0 : _GEN_15551; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15553 = 12'h7d == _T_171[11:0] ? 4'h0 : _GEN_15552; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15554 = 12'h7e == _T_171[11:0] ? 4'h0 : _GEN_15553; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15555 = 12'h7f == _T_171[11:0] ? 4'h0 : _GEN_15554; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15556 = 12'h80 == _T_171[11:0] ? 4'h0 : _GEN_15555; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15557 = 12'h81 == _T_171[11:0] ? 4'h0 : _GEN_15556; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15558 = 12'h82 == _T_171[11:0] ? 4'h0 : _GEN_15557; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15559 = 12'h83 == _T_171[11:0] ? 4'h0 : _GEN_15558; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15560 = 12'h84 == _T_171[11:0] ? 4'h0 : _GEN_15559; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15561 = 12'h85 == _T_171[11:0] ? 4'h0 : _GEN_15560; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15562 = 12'h86 == _T_171[11:0] ? 4'h0 : _GEN_15561; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15563 = 12'h87 == _T_171[11:0] ? 4'h0 : _GEN_15562; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15564 = 12'h88 == _T_171[11:0] ? image_136 : _GEN_15563; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15565 = 12'h89 == _T_171[11:0] ? image_137 : _GEN_15564; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15566 = 12'h8a == _T_171[11:0] ? image_138 : _GEN_15565; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15567 = 12'h8b == _T_171[11:0] ? image_139 : _GEN_15566; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15568 = 12'h8c == _T_171[11:0] ? image_140 : _GEN_15567; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15569 = 12'h8d == _T_171[11:0] ? image_141 : _GEN_15568; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15570 = 12'h8e == _T_171[11:0] ? image_142 : _GEN_15569; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15571 = 12'h8f == _T_171[11:0] ? image_143 : _GEN_15570; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15572 = 12'h90 == _T_171[11:0] ? image_144 : _GEN_15571; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15573 = 12'h91 == _T_171[11:0] ? image_145 : _GEN_15572; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15574 = 12'h92 == _T_171[11:0] ? image_146 : _GEN_15573; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15575 = 12'h93 == _T_171[11:0] ? image_147 : _GEN_15574; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15576 = 12'h94 == _T_171[11:0] ? image_148 : _GEN_15575; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15577 = 12'h95 == _T_171[11:0] ? image_149 : _GEN_15576; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15578 = 12'h96 == _T_171[11:0] ? image_150 : _GEN_15577; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15579 = 12'h97 == _T_171[11:0] ? image_151 : _GEN_15578; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15580 = 12'h98 == _T_171[11:0] ? image_152 : _GEN_15579; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15581 = 12'h99 == _T_171[11:0] ? image_153 : _GEN_15580; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15582 = 12'h9a == _T_171[11:0] ? image_154 : _GEN_15581; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15583 = 12'h9b == _T_171[11:0] ? image_155 : _GEN_15582; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15584 = 12'h9c == _T_171[11:0] ? 4'h0 : _GEN_15583; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15585 = 12'h9d == _T_171[11:0] ? image_157 : _GEN_15584; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15586 = 12'h9e == _T_171[11:0] ? image_158 : _GEN_15585; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15587 = 12'h9f == _T_171[11:0] ? image_159 : _GEN_15586; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15588 = 12'ha0 == _T_171[11:0] ? image_160 : _GEN_15587; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15589 = 12'ha1 == _T_171[11:0] ? image_161 : _GEN_15588; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15590 = 12'ha2 == _T_171[11:0] ? image_162 : _GEN_15589; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15591 = 12'ha3 == _T_171[11:0] ? image_163 : _GEN_15590; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15592 = 12'ha4 == _T_171[11:0] ? image_164 : _GEN_15591; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15593 = 12'ha5 == _T_171[11:0] ? image_165 : _GEN_15592; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15594 = 12'ha6 == _T_171[11:0] ? image_166 : _GEN_15593; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15595 = 12'ha7 == _T_171[11:0] ? image_167 : _GEN_15594; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15596 = 12'ha8 == _T_171[11:0] ? image_168 : _GEN_15595; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15597 = 12'ha9 == _T_171[11:0] ? image_169 : _GEN_15596; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15598 = 12'haa == _T_171[11:0] ? image_170 : _GEN_15597; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15599 = 12'hab == _T_171[11:0] ? image_171 : _GEN_15598; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15600 = 12'hac == _T_171[11:0] ? image_172 : _GEN_15599; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15601 = 12'had == _T_171[11:0] ? image_173 : _GEN_15600; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15602 = 12'hae == _T_171[11:0] ? image_174 : _GEN_15601; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15603 = 12'haf == _T_171[11:0] ? image_175 : _GEN_15602; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15604 = 12'hb0 == _T_171[11:0] ? image_176 : _GEN_15603; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15605 = 12'hb1 == _T_171[11:0] ? image_177 : _GEN_15604; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15606 = 12'hb2 == _T_171[11:0] ? image_178 : _GEN_15605; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15607 = 12'hb3 == _T_171[11:0] ? image_179 : _GEN_15606; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15608 = 12'hb4 == _T_171[11:0] ? 4'h0 : _GEN_15607; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15609 = 12'hb5 == _T_171[11:0] ? 4'h0 : _GEN_15608; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15610 = 12'hb6 == _T_171[11:0] ? 4'h0 : _GEN_15609; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15611 = 12'hb7 == _T_171[11:0] ? 4'h0 : _GEN_15610; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15612 = 12'hb8 == _T_171[11:0] ? 4'h0 : _GEN_15611; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15613 = 12'hb9 == _T_171[11:0] ? 4'h0 : _GEN_15612; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15614 = 12'hba == _T_171[11:0] ? 4'h0 : _GEN_15613; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15615 = 12'hbb == _T_171[11:0] ? 4'h0 : _GEN_15614; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15616 = 12'hbc == _T_171[11:0] ? 4'h0 : _GEN_15615; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15617 = 12'hbd == _T_171[11:0] ? 4'h0 : _GEN_15616; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15618 = 12'hbe == _T_171[11:0] ? 4'h0 : _GEN_15617; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15619 = 12'hbf == _T_171[11:0] ? 4'h0 : _GEN_15618; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15620 = 12'hc0 == _T_171[11:0] ? 4'h0 : _GEN_15619; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15621 = 12'hc1 == _T_171[11:0] ? 4'h0 : _GEN_15620; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15622 = 12'hc2 == _T_171[11:0] ? 4'h0 : _GEN_15621; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15623 = 12'hc3 == _T_171[11:0] ? 4'h0 : _GEN_15622; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15624 = 12'hc4 == _T_171[11:0] ? 4'h0 : _GEN_15623; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15625 = 12'hc5 == _T_171[11:0] ? 4'h0 : _GEN_15624; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15626 = 12'hc6 == _T_171[11:0] ? 4'h0 : _GEN_15625; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15627 = 12'hc7 == _T_171[11:0] ? image_199 : _GEN_15626; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15628 = 12'hc8 == _T_171[11:0] ? image_200 : _GEN_15627; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15629 = 12'hc9 == _T_171[11:0] ? image_201 : _GEN_15628; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15630 = 12'hca == _T_171[11:0] ? image_202 : _GEN_15629; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15631 = 12'hcb == _T_171[11:0] ? image_203 : _GEN_15630; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15632 = 12'hcc == _T_171[11:0] ? image_204 : _GEN_15631; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15633 = 12'hcd == _T_171[11:0] ? image_205 : _GEN_15632; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15634 = 12'hce == _T_171[11:0] ? image_206 : _GEN_15633; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15635 = 12'hcf == _T_171[11:0] ? image_207 : _GEN_15634; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15636 = 12'hd0 == _T_171[11:0] ? image_208 : _GEN_15635; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15637 = 12'hd1 == _T_171[11:0] ? image_209 : _GEN_15636; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15638 = 12'hd2 == _T_171[11:0] ? image_210 : _GEN_15637; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15639 = 12'hd3 == _T_171[11:0] ? image_211 : _GEN_15638; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15640 = 12'hd4 == _T_171[11:0] ? image_212 : _GEN_15639; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15641 = 12'hd5 == _T_171[11:0] ? image_213 : _GEN_15640; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15642 = 12'hd6 == _T_171[11:0] ? image_214 : _GEN_15641; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15643 = 12'hd7 == _T_171[11:0] ? image_215 : _GEN_15642; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15644 = 12'hd8 == _T_171[11:0] ? image_216 : _GEN_15643; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15645 = 12'hd9 == _T_171[11:0] ? image_217 : _GEN_15644; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15646 = 12'hda == _T_171[11:0] ? image_218 : _GEN_15645; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15647 = 12'hdb == _T_171[11:0] ? image_219 : _GEN_15646; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15648 = 12'hdc == _T_171[11:0] ? image_220 : _GEN_15647; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15649 = 12'hdd == _T_171[11:0] ? image_221 : _GEN_15648; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15650 = 12'hde == _T_171[11:0] ? image_222 : _GEN_15649; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15651 = 12'hdf == _T_171[11:0] ? image_223 : _GEN_15650; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15652 = 12'he0 == _T_171[11:0] ? image_224 : _GEN_15651; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15653 = 12'he1 == _T_171[11:0] ? image_225 : _GEN_15652; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15654 = 12'he2 == _T_171[11:0] ? image_226 : _GEN_15653; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15655 = 12'he3 == _T_171[11:0] ? image_227 : _GEN_15654; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15656 = 12'he4 == _T_171[11:0] ? image_228 : _GEN_15655; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15657 = 12'he5 == _T_171[11:0] ? image_229 : _GEN_15656; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15658 = 12'he6 == _T_171[11:0] ? image_230 : _GEN_15657; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15659 = 12'he7 == _T_171[11:0] ? image_231 : _GEN_15658; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15660 = 12'he8 == _T_171[11:0] ? image_232 : _GEN_15659; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15661 = 12'he9 == _T_171[11:0] ? image_233 : _GEN_15660; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15662 = 12'hea == _T_171[11:0] ? image_234 : _GEN_15661; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15663 = 12'heb == _T_171[11:0] ? image_235 : _GEN_15662; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15664 = 12'hec == _T_171[11:0] ? image_236 : _GEN_15663; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15665 = 12'hed == _T_171[11:0] ? image_237 : _GEN_15664; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15666 = 12'hee == _T_171[11:0] ? image_238 : _GEN_15665; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15667 = 12'hef == _T_171[11:0] ? image_239 : _GEN_15666; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15668 = 12'hf0 == _T_171[11:0] ? image_240 : _GEN_15667; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15669 = 12'hf1 == _T_171[11:0] ? image_241 : _GEN_15668; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15670 = 12'hf2 == _T_171[11:0] ? image_242 : _GEN_15669; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15671 = 12'hf3 == _T_171[11:0] ? image_243 : _GEN_15670; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15672 = 12'hf4 == _T_171[11:0] ? image_244 : _GEN_15671; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15673 = 12'hf5 == _T_171[11:0] ? image_245 : _GEN_15672; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15674 = 12'hf6 == _T_171[11:0] ? image_246 : _GEN_15673; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15675 = 12'hf7 == _T_171[11:0] ? 4'h0 : _GEN_15674; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15676 = 12'hf8 == _T_171[11:0] ? 4'h0 : _GEN_15675; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15677 = 12'hf9 == _T_171[11:0] ? 4'h0 : _GEN_15676; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15678 = 12'hfa == _T_171[11:0] ? 4'h0 : _GEN_15677; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15679 = 12'hfb == _T_171[11:0] ? 4'h0 : _GEN_15678; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15680 = 12'hfc == _T_171[11:0] ? 4'h0 : _GEN_15679; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15681 = 12'hfd == _T_171[11:0] ? 4'h0 : _GEN_15680; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15682 = 12'hfe == _T_171[11:0] ? 4'h0 : _GEN_15681; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15683 = 12'hff == _T_171[11:0] ? 4'h0 : _GEN_15682; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15684 = 12'h100 == _T_171[11:0] ? 4'h0 : _GEN_15683; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15685 = 12'h101 == _T_171[11:0] ? 4'h0 : _GEN_15684; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15686 = 12'h102 == _T_171[11:0] ? 4'h0 : _GEN_15685; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15687 = 12'h103 == _T_171[11:0] ? 4'h0 : _GEN_15686; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15688 = 12'h104 == _T_171[11:0] ? 4'h0 : _GEN_15687; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15689 = 12'h105 == _T_171[11:0] ? 4'h0 : _GEN_15688; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15690 = 12'h106 == _T_171[11:0] ? image_262 : _GEN_15689; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15691 = 12'h107 == _T_171[11:0] ? image_263 : _GEN_15690; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15692 = 12'h108 == _T_171[11:0] ? image_264 : _GEN_15691; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15693 = 12'h109 == _T_171[11:0] ? image_265 : _GEN_15692; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15694 = 12'h10a == _T_171[11:0] ? image_266 : _GEN_15693; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15695 = 12'h10b == _T_171[11:0] ? image_267 : _GEN_15694; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15696 = 12'h10c == _T_171[11:0] ? image_268 : _GEN_15695; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15697 = 12'h10d == _T_171[11:0] ? image_269 : _GEN_15696; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15698 = 12'h10e == _T_171[11:0] ? image_270 : _GEN_15697; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15699 = 12'h10f == _T_171[11:0] ? image_271 : _GEN_15698; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15700 = 12'h110 == _T_171[11:0] ? image_272 : _GEN_15699; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15701 = 12'h111 == _T_171[11:0] ? image_273 : _GEN_15700; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15702 = 12'h112 == _T_171[11:0] ? image_274 : _GEN_15701; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15703 = 12'h113 == _T_171[11:0] ? image_275 : _GEN_15702; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15704 = 12'h114 == _T_171[11:0] ? image_276 : _GEN_15703; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15705 = 12'h115 == _T_171[11:0] ? image_277 : _GEN_15704; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15706 = 12'h116 == _T_171[11:0] ? image_278 : _GEN_15705; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15707 = 12'h117 == _T_171[11:0] ? image_279 : _GEN_15706; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15708 = 12'h118 == _T_171[11:0] ? image_280 : _GEN_15707; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15709 = 12'h119 == _T_171[11:0] ? image_281 : _GEN_15708; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15710 = 12'h11a == _T_171[11:0] ? image_282 : _GEN_15709; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15711 = 12'h11b == _T_171[11:0] ? image_283 : _GEN_15710; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15712 = 12'h11c == _T_171[11:0] ? image_284 : _GEN_15711; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15713 = 12'h11d == _T_171[11:0] ? image_285 : _GEN_15712; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15714 = 12'h11e == _T_171[11:0] ? image_286 : _GEN_15713; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15715 = 12'h11f == _T_171[11:0] ? image_287 : _GEN_15714; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15716 = 12'h120 == _T_171[11:0] ? image_288 : _GEN_15715; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15717 = 12'h121 == _T_171[11:0] ? image_289 : _GEN_15716; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15718 = 12'h122 == _T_171[11:0] ? image_290 : _GEN_15717; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15719 = 12'h123 == _T_171[11:0] ? image_291 : _GEN_15718; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15720 = 12'h124 == _T_171[11:0] ? image_292 : _GEN_15719; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15721 = 12'h125 == _T_171[11:0] ? image_293 : _GEN_15720; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15722 = 12'h126 == _T_171[11:0] ? image_294 : _GEN_15721; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15723 = 12'h127 == _T_171[11:0] ? image_295 : _GEN_15722; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15724 = 12'h128 == _T_171[11:0] ? image_296 : _GEN_15723; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15725 = 12'h129 == _T_171[11:0] ? image_297 : _GEN_15724; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15726 = 12'h12a == _T_171[11:0] ? image_298 : _GEN_15725; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15727 = 12'h12b == _T_171[11:0] ? image_299 : _GEN_15726; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15728 = 12'h12c == _T_171[11:0] ? image_300 : _GEN_15727; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15729 = 12'h12d == _T_171[11:0] ? image_301 : _GEN_15728; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15730 = 12'h12e == _T_171[11:0] ? image_302 : _GEN_15729; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15731 = 12'h12f == _T_171[11:0] ? image_303 : _GEN_15730; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15732 = 12'h130 == _T_171[11:0] ? image_304 : _GEN_15731; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15733 = 12'h131 == _T_171[11:0] ? image_305 : _GEN_15732; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15734 = 12'h132 == _T_171[11:0] ? image_306 : _GEN_15733; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15735 = 12'h133 == _T_171[11:0] ? image_307 : _GEN_15734; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15736 = 12'h134 == _T_171[11:0] ? image_308 : _GEN_15735; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15737 = 12'h135 == _T_171[11:0] ? image_309 : _GEN_15736; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15738 = 12'h136 == _T_171[11:0] ? image_310 : _GEN_15737; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15739 = 12'h137 == _T_171[11:0] ? image_311 : _GEN_15738; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15740 = 12'h138 == _T_171[11:0] ? image_312 : _GEN_15739; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15741 = 12'h139 == _T_171[11:0] ? image_313 : _GEN_15740; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15742 = 12'h13a == _T_171[11:0] ? image_314 : _GEN_15741; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15743 = 12'h13b == _T_171[11:0] ? image_315 : _GEN_15742; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15744 = 12'h13c == _T_171[11:0] ? 4'h0 : _GEN_15743; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15745 = 12'h13d == _T_171[11:0] ? 4'h0 : _GEN_15744; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15746 = 12'h13e == _T_171[11:0] ? 4'h0 : _GEN_15745; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15747 = 12'h13f == _T_171[11:0] ? 4'h0 : _GEN_15746; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15748 = 12'h140 == _T_171[11:0] ? 4'h0 : _GEN_15747; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15749 = 12'h141 == _T_171[11:0] ? 4'h0 : _GEN_15748; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15750 = 12'h142 == _T_171[11:0] ? 4'h0 : _GEN_15749; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15751 = 12'h143 == _T_171[11:0] ? 4'h0 : _GEN_15750; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15752 = 12'h144 == _T_171[11:0] ? 4'h0 : _GEN_15751; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15753 = 12'h145 == _T_171[11:0] ? image_325 : _GEN_15752; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15754 = 12'h146 == _T_171[11:0] ? image_326 : _GEN_15753; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15755 = 12'h147 == _T_171[11:0] ? image_327 : _GEN_15754; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15756 = 12'h148 == _T_171[11:0] ? image_328 : _GEN_15755; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15757 = 12'h149 == _T_171[11:0] ? image_329 : _GEN_15756; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15758 = 12'h14a == _T_171[11:0] ? image_330 : _GEN_15757; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15759 = 12'h14b == _T_171[11:0] ? image_331 : _GEN_15758; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15760 = 12'h14c == _T_171[11:0] ? image_332 : _GEN_15759; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15761 = 12'h14d == _T_171[11:0] ? image_333 : _GEN_15760; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15762 = 12'h14e == _T_171[11:0] ? image_334 : _GEN_15761; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15763 = 12'h14f == _T_171[11:0] ? image_335 : _GEN_15762; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15764 = 12'h150 == _T_171[11:0] ? image_336 : _GEN_15763; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15765 = 12'h151 == _T_171[11:0] ? image_337 : _GEN_15764; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15766 = 12'h152 == _T_171[11:0] ? image_338 : _GEN_15765; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15767 = 12'h153 == _T_171[11:0] ? image_339 : _GEN_15766; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15768 = 12'h154 == _T_171[11:0] ? image_340 : _GEN_15767; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15769 = 12'h155 == _T_171[11:0] ? image_341 : _GEN_15768; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15770 = 12'h156 == _T_171[11:0] ? image_342 : _GEN_15769; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15771 = 12'h157 == _T_171[11:0] ? image_343 : _GEN_15770; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15772 = 12'h158 == _T_171[11:0] ? image_344 : _GEN_15771; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15773 = 12'h159 == _T_171[11:0] ? image_345 : _GEN_15772; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15774 = 12'h15a == _T_171[11:0] ? image_346 : _GEN_15773; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15775 = 12'h15b == _T_171[11:0] ? image_347 : _GEN_15774; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15776 = 12'h15c == _T_171[11:0] ? image_348 : _GEN_15775; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15777 = 12'h15d == _T_171[11:0] ? image_349 : _GEN_15776; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15778 = 12'h15e == _T_171[11:0] ? image_350 : _GEN_15777; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15779 = 12'h15f == _T_171[11:0] ? image_351 : _GEN_15778; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15780 = 12'h160 == _T_171[11:0] ? image_352 : _GEN_15779; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15781 = 12'h161 == _T_171[11:0] ? image_353 : _GEN_15780; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15782 = 12'h162 == _T_171[11:0] ? image_354 : _GEN_15781; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15783 = 12'h163 == _T_171[11:0] ? image_355 : _GEN_15782; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15784 = 12'h164 == _T_171[11:0] ? image_356 : _GEN_15783; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15785 = 12'h165 == _T_171[11:0] ? image_357 : _GEN_15784; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15786 = 12'h166 == _T_171[11:0] ? image_358 : _GEN_15785; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15787 = 12'h167 == _T_171[11:0] ? image_359 : _GEN_15786; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15788 = 12'h168 == _T_171[11:0] ? image_360 : _GEN_15787; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15789 = 12'h169 == _T_171[11:0] ? image_361 : _GEN_15788; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15790 = 12'h16a == _T_171[11:0] ? image_362 : _GEN_15789; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15791 = 12'h16b == _T_171[11:0] ? image_363 : _GEN_15790; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15792 = 12'h16c == _T_171[11:0] ? image_364 : _GEN_15791; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15793 = 12'h16d == _T_171[11:0] ? image_365 : _GEN_15792; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15794 = 12'h16e == _T_171[11:0] ? image_366 : _GEN_15793; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15795 = 12'h16f == _T_171[11:0] ? image_367 : _GEN_15794; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15796 = 12'h170 == _T_171[11:0] ? image_368 : _GEN_15795; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15797 = 12'h171 == _T_171[11:0] ? image_369 : _GEN_15796; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15798 = 12'h172 == _T_171[11:0] ? image_370 : _GEN_15797; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15799 = 12'h173 == _T_171[11:0] ? image_371 : _GEN_15798; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15800 = 12'h174 == _T_171[11:0] ? image_372 : _GEN_15799; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15801 = 12'h175 == _T_171[11:0] ? image_373 : _GEN_15800; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15802 = 12'h176 == _T_171[11:0] ? image_374 : _GEN_15801; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15803 = 12'h177 == _T_171[11:0] ? image_375 : _GEN_15802; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15804 = 12'h178 == _T_171[11:0] ? image_376 : _GEN_15803; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15805 = 12'h179 == _T_171[11:0] ? image_377 : _GEN_15804; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15806 = 12'h17a == _T_171[11:0] ? image_378 : _GEN_15805; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15807 = 12'h17b == _T_171[11:0] ? image_379 : _GEN_15806; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15808 = 12'h17c == _T_171[11:0] ? 4'h0 : _GEN_15807; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15809 = 12'h17d == _T_171[11:0] ? 4'h0 : _GEN_15808; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15810 = 12'h17e == _T_171[11:0] ? 4'h0 : _GEN_15809; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15811 = 12'h17f == _T_171[11:0] ? 4'h0 : _GEN_15810; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15812 = 12'h180 == _T_171[11:0] ? 4'h0 : _GEN_15811; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15813 = 12'h181 == _T_171[11:0] ? 4'h0 : _GEN_15812; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15814 = 12'h182 == _T_171[11:0] ? 4'h0 : _GEN_15813; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15815 = 12'h183 == _T_171[11:0] ? 4'h0 : _GEN_15814; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15816 = 12'h184 == _T_171[11:0] ? image_388 : _GEN_15815; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15817 = 12'h185 == _T_171[11:0] ? image_389 : _GEN_15816; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15818 = 12'h186 == _T_171[11:0] ? image_390 : _GEN_15817; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15819 = 12'h187 == _T_171[11:0] ? image_391 : _GEN_15818; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15820 = 12'h188 == _T_171[11:0] ? image_392 : _GEN_15819; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15821 = 12'h189 == _T_171[11:0] ? image_393 : _GEN_15820; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15822 = 12'h18a == _T_171[11:0] ? image_394 : _GEN_15821; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15823 = 12'h18b == _T_171[11:0] ? image_395 : _GEN_15822; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15824 = 12'h18c == _T_171[11:0] ? image_396 : _GEN_15823; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15825 = 12'h18d == _T_171[11:0] ? image_397 : _GEN_15824; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15826 = 12'h18e == _T_171[11:0] ? image_398 : _GEN_15825; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15827 = 12'h18f == _T_171[11:0] ? image_399 : _GEN_15826; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15828 = 12'h190 == _T_171[11:0] ? image_400 : _GEN_15827; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15829 = 12'h191 == _T_171[11:0] ? image_401 : _GEN_15828; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15830 = 12'h192 == _T_171[11:0] ? image_402 : _GEN_15829; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15831 = 12'h193 == _T_171[11:0] ? image_403 : _GEN_15830; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15832 = 12'h194 == _T_171[11:0] ? image_404 : _GEN_15831; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15833 = 12'h195 == _T_171[11:0] ? image_405 : _GEN_15832; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15834 = 12'h196 == _T_171[11:0] ? image_406 : _GEN_15833; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15835 = 12'h197 == _T_171[11:0] ? image_407 : _GEN_15834; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15836 = 12'h198 == _T_171[11:0] ? image_408 : _GEN_15835; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15837 = 12'h199 == _T_171[11:0] ? image_409 : _GEN_15836; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15838 = 12'h19a == _T_171[11:0] ? image_410 : _GEN_15837; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15839 = 12'h19b == _T_171[11:0] ? image_411 : _GEN_15838; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15840 = 12'h19c == _T_171[11:0] ? image_412 : _GEN_15839; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15841 = 12'h19d == _T_171[11:0] ? image_413 : _GEN_15840; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15842 = 12'h19e == _T_171[11:0] ? image_414 : _GEN_15841; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15843 = 12'h19f == _T_171[11:0] ? image_415 : _GEN_15842; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15844 = 12'h1a0 == _T_171[11:0] ? image_416 : _GEN_15843; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15845 = 12'h1a1 == _T_171[11:0] ? image_417 : _GEN_15844; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15846 = 12'h1a2 == _T_171[11:0] ? image_418 : _GEN_15845; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15847 = 12'h1a3 == _T_171[11:0] ? image_419 : _GEN_15846; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15848 = 12'h1a4 == _T_171[11:0] ? image_420 : _GEN_15847; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15849 = 12'h1a5 == _T_171[11:0] ? image_421 : _GEN_15848; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15850 = 12'h1a6 == _T_171[11:0] ? image_422 : _GEN_15849; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15851 = 12'h1a7 == _T_171[11:0] ? image_423 : _GEN_15850; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15852 = 12'h1a8 == _T_171[11:0] ? image_424 : _GEN_15851; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15853 = 12'h1a9 == _T_171[11:0] ? image_425 : _GEN_15852; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15854 = 12'h1aa == _T_171[11:0] ? image_426 : _GEN_15853; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15855 = 12'h1ab == _T_171[11:0] ? image_427 : _GEN_15854; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15856 = 12'h1ac == _T_171[11:0] ? image_428 : _GEN_15855; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15857 = 12'h1ad == _T_171[11:0] ? image_429 : _GEN_15856; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15858 = 12'h1ae == _T_171[11:0] ? image_430 : _GEN_15857; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15859 = 12'h1af == _T_171[11:0] ? image_431 : _GEN_15858; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15860 = 12'h1b0 == _T_171[11:0] ? image_432 : _GEN_15859; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15861 = 12'h1b1 == _T_171[11:0] ? image_433 : _GEN_15860; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15862 = 12'h1b2 == _T_171[11:0] ? image_434 : _GEN_15861; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15863 = 12'h1b3 == _T_171[11:0] ? image_435 : _GEN_15862; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15864 = 12'h1b4 == _T_171[11:0] ? image_436 : _GEN_15863; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15865 = 12'h1b5 == _T_171[11:0] ? image_437 : _GEN_15864; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15866 = 12'h1b6 == _T_171[11:0] ? image_438 : _GEN_15865; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15867 = 12'h1b7 == _T_171[11:0] ? image_439 : _GEN_15866; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15868 = 12'h1b8 == _T_171[11:0] ? image_440 : _GEN_15867; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15869 = 12'h1b9 == _T_171[11:0] ? image_441 : _GEN_15868; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15870 = 12'h1ba == _T_171[11:0] ? image_442 : _GEN_15869; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15871 = 12'h1bb == _T_171[11:0] ? image_443 : _GEN_15870; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15872 = 12'h1bc == _T_171[11:0] ? image_444 : _GEN_15871; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15873 = 12'h1bd == _T_171[11:0] ? 4'h0 : _GEN_15872; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15874 = 12'h1be == _T_171[11:0] ? 4'h0 : _GEN_15873; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15875 = 12'h1bf == _T_171[11:0] ? 4'h0 : _GEN_15874; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15876 = 12'h1c0 == _T_171[11:0] ? 4'h0 : _GEN_15875; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15877 = 12'h1c1 == _T_171[11:0] ? 4'h0 : _GEN_15876; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15878 = 12'h1c2 == _T_171[11:0] ? 4'h0 : _GEN_15877; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15879 = 12'h1c3 == _T_171[11:0] ? image_451 : _GEN_15878; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15880 = 12'h1c4 == _T_171[11:0] ? image_452 : _GEN_15879; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15881 = 12'h1c5 == _T_171[11:0] ? image_453 : _GEN_15880; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15882 = 12'h1c6 == _T_171[11:0] ? image_454 : _GEN_15881; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15883 = 12'h1c7 == _T_171[11:0] ? image_455 : _GEN_15882; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15884 = 12'h1c8 == _T_171[11:0] ? image_456 : _GEN_15883; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15885 = 12'h1c9 == _T_171[11:0] ? image_457 : _GEN_15884; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15886 = 12'h1ca == _T_171[11:0] ? image_458 : _GEN_15885; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15887 = 12'h1cb == _T_171[11:0] ? image_459 : _GEN_15886; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15888 = 12'h1cc == _T_171[11:0] ? image_460 : _GEN_15887; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15889 = 12'h1cd == _T_171[11:0] ? image_461 : _GEN_15888; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15890 = 12'h1ce == _T_171[11:0] ? image_462 : _GEN_15889; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15891 = 12'h1cf == _T_171[11:0] ? image_463 : _GEN_15890; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15892 = 12'h1d0 == _T_171[11:0] ? image_464 : _GEN_15891; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15893 = 12'h1d1 == _T_171[11:0] ? image_465 : _GEN_15892; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15894 = 12'h1d2 == _T_171[11:0] ? image_466 : _GEN_15893; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15895 = 12'h1d3 == _T_171[11:0] ? image_467 : _GEN_15894; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15896 = 12'h1d4 == _T_171[11:0] ? image_468 : _GEN_15895; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15897 = 12'h1d5 == _T_171[11:0] ? image_469 : _GEN_15896; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15898 = 12'h1d6 == _T_171[11:0] ? image_470 : _GEN_15897; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15899 = 12'h1d7 == _T_171[11:0] ? image_471 : _GEN_15898; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15900 = 12'h1d8 == _T_171[11:0] ? image_472 : _GEN_15899; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15901 = 12'h1d9 == _T_171[11:0] ? image_473 : _GEN_15900; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15902 = 12'h1da == _T_171[11:0] ? image_474 : _GEN_15901; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15903 = 12'h1db == _T_171[11:0] ? image_475 : _GEN_15902; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15904 = 12'h1dc == _T_171[11:0] ? image_476 : _GEN_15903; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15905 = 12'h1dd == _T_171[11:0] ? image_477 : _GEN_15904; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15906 = 12'h1de == _T_171[11:0] ? image_478 : _GEN_15905; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15907 = 12'h1df == _T_171[11:0] ? image_479 : _GEN_15906; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15908 = 12'h1e0 == _T_171[11:0] ? image_480 : _GEN_15907; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15909 = 12'h1e1 == _T_171[11:0] ? image_481 : _GEN_15908; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15910 = 12'h1e2 == _T_171[11:0] ? image_482 : _GEN_15909; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15911 = 12'h1e3 == _T_171[11:0] ? image_483 : _GEN_15910; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15912 = 12'h1e4 == _T_171[11:0] ? image_484 : _GEN_15911; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15913 = 12'h1e5 == _T_171[11:0] ? image_485 : _GEN_15912; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15914 = 12'h1e6 == _T_171[11:0] ? image_486 : _GEN_15913; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15915 = 12'h1e7 == _T_171[11:0] ? image_487 : _GEN_15914; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15916 = 12'h1e8 == _T_171[11:0] ? image_488 : _GEN_15915; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15917 = 12'h1e9 == _T_171[11:0] ? image_489 : _GEN_15916; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15918 = 12'h1ea == _T_171[11:0] ? image_490 : _GEN_15917; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15919 = 12'h1eb == _T_171[11:0] ? image_491 : _GEN_15918; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15920 = 12'h1ec == _T_171[11:0] ? image_492 : _GEN_15919; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15921 = 12'h1ed == _T_171[11:0] ? image_493 : _GEN_15920; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15922 = 12'h1ee == _T_171[11:0] ? image_494 : _GEN_15921; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15923 = 12'h1ef == _T_171[11:0] ? image_495 : _GEN_15922; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15924 = 12'h1f0 == _T_171[11:0] ? image_496 : _GEN_15923; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15925 = 12'h1f1 == _T_171[11:0] ? image_497 : _GEN_15924; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15926 = 12'h1f2 == _T_171[11:0] ? image_498 : _GEN_15925; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15927 = 12'h1f3 == _T_171[11:0] ? image_499 : _GEN_15926; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15928 = 12'h1f4 == _T_171[11:0] ? image_500 : _GEN_15927; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15929 = 12'h1f5 == _T_171[11:0] ? image_501 : _GEN_15928; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15930 = 12'h1f6 == _T_171[11:0] ? image_502 : _GEN_15929; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15931 = 12'h1f7 == _T_171[11:0] ? image_503 : _GEN_15930; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15932 = 12'h1f8 == _T_171[11:0] ? image_504 : _GEN_15931; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15933 = 12'h1f9 == _T_171[11:0] ? image_505 : _GEN_15932; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15934 = 12'h1fa == _T_171[11:0] ? image_506 : _GEN_15933; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15935 = 12'h1fb == _T_171[11:0] ? image_507 : _GEN_15934; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15936 = 12'h1fc == _T_171[11:0] ? image_508 : _GEN_15935; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15937 = 12'h1fd == _T_171[11:0] ? image_509 : _GEN_15936; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15938 = 12'h1fe == _T_171[11:0] ? 4'h0 : _GEN_15937; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15939 = 12'h1ff == _T_171[11:0] ? 4'h0 : _GEN_15938; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15940 = 12'h200 == _T_171[11:0] ? 4'h0 : _GEN_15939; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15941 = 12'h201 == _T_171[11:0] ? 4'h0 : _GEN_15940; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15942 = 12'h202 == _T_171[11:0] ? 4'h0 : _GEN_15941; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15943 = 12'h203 == _T_171[11:0] ? image_515 : _GEN_15942; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15944 = 12'h204 == _T_171[11:0] ? image_516 : _GEN_15943; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15945 = 12'h205 == _T_171[11:0] ? image_517 : _GEN_15944; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15946 = 12'h206 == _T_171[11:0] ? image_518 : _GEN_15945; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15947 = 12'h207 == _T_171[11:0] ? image_519 : _GEN_15946; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15948 = 12'h208 == _T_171[11:0] ? image_520 : _GEN_15947; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15949 = 12'h209 == _T_171[11:0] ? image_521 : _GEN_15948; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15950 = 12'h20a == _T_171[11:0] ? image_522 : _GEN_15949; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15951 = 12'h20b == _T_171[11:0] ? image_523 : _GEN_15950; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15952 = 12'h20c == _T_171[11:0] ? image_524 : _GEN_15951; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15953 = 12'h20d == _T_171[11:0] ? image_525 : _GEN_15952; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15954 = 12'h20e == _T_171[11:0] ? image_526 : _GEN_15953; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15955 = 12'h20f == _T_171[11:0] ? image_527 : _GEN_15954; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15956 = 12'h210 == _T_171[11:0] ? image_528 : _GEN_15955; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15957 = 12'h211 == _T_171[11:0] ? image_529 : _GEN_15956; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15958 = 12'h212 == _T_171[11:0] ? image_530 : _GEN_15957; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15959 = 12'h213 == _T_171[11:0] ? image_531 : _GEN_15958; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15960 = 12'h214 == _T_171[11:0] ? image_532 : _GEN_15959; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15961 = 12'h215 == _T_171[11:0] ? image_533 : _GEN_15960; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15962 = 12'h216 == _T_171[11:0] ? image_534 : _GEN_15961; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15963 = 12'h217 == _T_171[11:0] ? image_535 : _GEN_15962; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15964 = 12'h218 == _T_171[11:0] ? image_536 : _GEN_15963; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15965 = 12'h219 == _T_171[11:0] ? image_537 : _GEN_15964; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15966 = 12'h21a == _T_171[11:0] ? image_538 : _GEN_15965; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15967 = 12'h21b == _T_171[11:0] ? image_539 : _GEN_15966; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15968 = 12'h21c == _T_171[11:0] ? image_540 : _GEN_15967; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15969 = 12'h21d == _T_171[11:0] ? image_541 : _GEN_15968; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15970 = 12'h21e == _T_171[11:0] ? image_542 : _GEN_15969; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15971 = 12'h21f == _T_171[11:0] ? image_543 : _GEN_15970; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15972 = 12'h220 == _T_171[11:0] ? image_544 : _GEN_15971; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15973 = 12'h221 == _T_171[11:0] ? image_545 : _GEN_15972; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15974 = 12'h222 == _T_171[11:0] ? image_546 : _GEN_15973; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15975 = 12'h223 == _T_171[11:0] ? image_547 : _GEN_15974; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15976 = 12'h224 == _T_171[11:0] ? image_548 : _GEN_15975; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15977 = 12'h225 == _T_171[11:0] ? image_549 : _GEN_15976; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15978 = 12'h226 == _T_171[11:0] ? image_550 : _GEN_15977; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15979 = 12'h227 == _T_171[11:0] ? image_551 : _GEN_15978; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15980 = 12'h228 == _T_171[11:0] ? image_552 : _GEN_15979; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15981 = 12'h229 == _T_171[11:0] ? image_553 : _GEN_15980; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15982 = 12'h22a == _T_171[11:0] ? image_554 : _GEN_15981; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15983 = 12'h22b == _T_171[11:0] ? image_555 : _GEN_15982; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15984 = 12'h22c == _T_171[11:0] ? image_556 : _GEN_15983; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15985 = 12'h22d == _T_171[11:0] ? image_557 : _GEN_15984; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15986 = 12'h22e == _T_171[11:0] ? image_558 : _GEN_15985; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15987 = 12'h22f == _T_171[11:0] ? image_559 : _GEN_15986; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15988 = 12'h230 == _T_171[11:0] ? image_560 : _GEN_15987; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15989 = 12'h231 == _T_171[11:0] ? image_561 : _GEN_15988; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15990 = 12'h232 == _T_171[11:0] ? image_562 : _GEN_15989; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15991 = 12'h233 == _T_171[11:0] ? image_563 : _GEN_15990; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15992 = 12'h234 == _T_171[11:0] ? image_564 : _GEN_15991; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15993 = 12'h235 == _T_171[11:0] ? image_565 : _GEN_15992; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15994 = 12'h236 == _T_171[11:0] ? image_566 : _GEN_15993; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15995 = 12'h237 == _T_171[11:0] ? 4'h0 : _GEN_15994; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15996 = 12'h238 == _T_171[11:0] ? 4'h0 : _GEN_15995; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15997 = 12'h239 == _T_171[11:0] ? 4'h0 : _GEN_15996; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15998 = 12'h23a == _T_171[11:0] ? 4'h0 : _GEN_15997; // @[Filter.scala 138:46]
  wire [3:0] _GEN_15999 = 12'h23b == _T_171[11:0] ? image_571 : _GEN_15998; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16000 = 12'h23c == _T_171[11:0] ? image_572 : _GEN_15999; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16001 = 12'h23d == _T_171[11:0] ? image_573 : _GEN_16000; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16002 = 12'h23e == _T_171[11:0] ? image_574 : _GEN_16001; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16003 = 12'h23f == _T_171[11:0] ? 4'h0 : _GEN_16002; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16004 = 12'h240 == _T_171[11:0] ? 4'h0 : _GEN_16003; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16005 = 12'h241 == _T_171[11:0] ? 4'h0 : _GEN_16004; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16006 = 12'h242 == _T_171[11:0] ? image_578 : _GEN_16005; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16007 = 12'h243 == _T_171[11:0] ? image_579 : _GEN_16006; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16008 = 12'h244 == _T_171[11:0] ? image_580 : _GEN_16007; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16009 = 12'h245 == _T_171[11:0] ? image_581 : _GEN_16008; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16010 = 12'h246 == _T_171[11:0] ? image_582 : _GEN_16009; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16011 = 12'h247 == _T_171[11:0] ? image_583 : _GEN_16010; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16012 = 12'h248 == _T_171[11:0] ? image_584 : _GEN_16011; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16013 = 12'h249 == _T_171[11:0] ? image_585 : _GEN_16012; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16014 = 12'h24a == _T_171[11:0] ? image_586 : _GEN_16013; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16015 = 12'h24b == _T_171[11:0] ? image_587 : _GEN_16014; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16016 = 12'h24c == _T_171[11:0] ? image_588 : _GEN_16015; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16017 = 12'h24d == _T_171[11:0] ? image_589 : _GEN_16016; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16018 = 12'h24e == _T_171[11:0] ? image_590 : _GEN_16017; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16019 = 12'h24f == _T_171[11:0] ? image_591 : _GEN_16018; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16020 = 12'h250 == _T_171[11:0] ? image_592 : _GEN_16019; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16021 = 12'h251 == _T_171[11:0] ? image_593 : _GEN_16020; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16022 = 12'h252 == _T_171[11:0] ? image_594 : _GEN_16021; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16023 = 12'h253 == _T_171[11:0] ? image_595 : _GEN_16022; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16024 = 12'h254 == _T_171[11:0] ? image_596 : _GEN_16023; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16025 = 12'h255 == _T_171[11:0] ? image_597 : _GEN_16024; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16026 = 12'h256 == _T_171[11:0] ? image_598 : _GEN_16025; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16027 = 12'h257 == _T_171[11:0] ? image_599 : _GEN_16026; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16028 = 12'h258 == _T_171[11:0] ? image_600 : _GEN_16027; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16029 = 12'h259 == _T_171[11:0] ? image_601 : _GEN_16028; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16030 = 12'h25a == _T_171[11:0] ? image_602 : _GEN_16029; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16031 = 12'h25b == _T_171[11:0] ? image_603 : _GEN_16030; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16032 = 12'h25c == _T_171[11:0] ? image_604 : _GEN_16031; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16033 = 12'h25d == _T_171[11:0] ? image_605 : _GEN_16032; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16034 = 12'h25e == _T_171[11:0] ? image_606 : _GEN_16033; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16035 = 12'h25f == _T_171[11:0] ? image_607 : _GEN_16034; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16036 = 12'h260 == _T_171[11:0] ? 4'h0 : _GEN_16035; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16037 = 12'h261 == _T_171[11:0] ? 4'h0 : _GEN_16036; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16038 = 12'h262 == _T_171[11:0] ? 4'h0 : _GEN_16037; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16039 = 12'h263 == _T_171[11:0] ? 4'h0 : _GEN_16038; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16040 = 12'h264 == _T_171[11:0] ? 4'h0 : _GEN_16039; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16041 = 12'h265 == _T_171[11:0] ? 4'h0 : _GEN_16040; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16042 = 12'h266 == _T_171[11:0] ? image_614 : _GEN_16041; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16043 = 12'h267 == _T_171[11:0] ? image_615 : _GEN_16042; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16044 = 12'h268 == _T_171[11:0] ? image_616 : _GEN_16043; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16045 = 12'h269 == _T_171[11:0] ? image_617 : _GEN_16044; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16046 = 12'h26a == _T_171[11:0] ? image_618 : _GEN_16045; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16047 = 12'h26b == _T_171[11:0] ? image_619 : _GEN_16046; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16048 = 12'h26c == _T_171[11:0] ? image_620 : _GEN_16047; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16049 = 12'h26d == _T_171[11:0] ? image_621 : _GEN_16048; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16050 = 12'h26e == _T_171[11:0] ? image_622 : _GEN_16049; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16051 = 12'h26f == _T_171[11:0] ? image_623 : _GEN_16050; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16052 = 12'h270 == _T_171[11:0] ? image_624 : _GEN_16051; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16053 = 12'h271 == _T_171[11:0] ? image_625 : _GEN_16052; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16054 = 12'h272 == _T_171[11:0] ? image_626 : _GEN_16053; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16055 = 12'h273 == _T_171[11:0] ? image_627 : _GEN_16054; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16056 = 12'h274 == _T_171[11:0] ? image_628 : _GEN_16055; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16057 = 12'h275 == _T_171[11:0] ? 4'h0 : _GEN_16056; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16058 = 12'h276 == _T_171[11:0] ? 4'h0 : _GEN_16057; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16059 = 12'h277 == _T_171[11:0] ? 4'h0 : _GEN_16058; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16060 = 12'h278 == _T_171[11:0] ? 4'h0 : _GEN_16059; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16061 = 12'h279 == _T_171[11:0] ? 4'h0 : _GEN_16060; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16062 = 12'h27a == _T_171[11:0] ? 4'h0 : _GEN_16061; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16063 = 12'h27b == _T_171[11:0] ? 4'h0 : _GEN_16062; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16064 = 12'h27c == _T_171[11:0] ? image_636 : _GEN_16063; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16065 = 12'h27d == _T_171[11:0] ? image_637 : _GEN_16064; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16066 = 12'h27e == _T_171[11:0] ? image_638 : _GEN_16065; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16067 = 12'h27f == _T_171[11:0] ? image_639 : _GEN_16066; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16068 = 12'h280 == _T_171[11:0] ? 4'h0 : _GEN_16067; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16069 = 12'h281 == _T_171[11:0] ? 4'h0 : _GEN_16068; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16070 = 12'h282 == _T_171[11:0] ? image_642 : _GEN_16069; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16071 = 12'h283 == _T_171[11:0] ? image_643 : _GEN_16070; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16072 = 12'h284 == _T_171[11:0] ? image_644 : _GEN_16071; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16073 = 12'h285 == _T_171[11:0] ? image_645 : _GEN_16072; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16074 = 12'h286 == _T_171[11:0] ? image_646 : _GEN_16073; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16075 = 12'h287 == _T_171[11:0] ? image_647 : _GEN_16074; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16076 = 12'h288 == _T_171[11:0] ? image_648 : _GEN_16075; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16077 = 12'h289 == _T_171[11:0] ? image_649 : _GEN_16076; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16078 = 12'h28a == _T_171[11:0] ? image_650 : _GEN_16077; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16079 = 12'h28b == _T_171[11:0] ? image_651 : _GEN_16078; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16080 = 12'h28c == _T_171[11:0] ? image_652 : _GEN_16079; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16081 = 12'h28d == _T_171[11:0] ? image_653 : _GEN_16080; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16082 = 12'h28e == _T_171[11:0] ? image_654 : _GEN_16081; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16083 = 12'h28f == _T_171[11:0] ? image_655 : _GEN_16082; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16084 = 12'h290 == _T_171[11:0] ? image_656 : _GEN_16083; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16085 = 12'h291 == _T_171[11:0] ? image_657 : _GEN_16084; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16086 = 12'h292 == _T_171[11:0] ? image_658 : _GEN_16085; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16087 = 12'h293 == _T_171[11:0] ? image_659 : _GEN_16086; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16088 = 12'h294 == _T_171[11:0] ? image_660 : _GEN_16087; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16089 = 12'h295 == _T_171[11:0] ? image_661 : _GEN_16088; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16090 = 12'h296 == _T_171[11:0] ? image_662 : _GEN_16089; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16091 = 12'h297 == _T_171[11:0] ? image_663 : _GEN_16090; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16092 = 12'h298 == _T_171[11:0] ? image_664 : _GEN_16091; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16093 = 12'h299 == _T_171[11:0] ? image_665 : _GEN_16092; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16094 = 12'h29a == _T_171[11:0] ? image_666 : _GEN_16093; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16095 = 12'h29b == _T_171[11:0] ? image_667 : _GEN_16094; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16096 = 12'h29c == _T_171[11:0] ? image_668 : _GEN_16095; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16097 = 12'h29d == _T_171[11:0] ? image_669 : _GEN_16096; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16098 = 12'h29e == _T_171[11:0] ? image_670 : _GEN_16097; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16099 = 12'h29f == _T_171[11:0] ? 4'h0 : _GEN_16098; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16100 = 12'h2a0 == _T_171[11:0] ? 4'h0 : _GEN_16099; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16101 = 12'h2a1 == _T_171[11:0] ? 4'h0 : _GEN_16100; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16102 = 12'h2a2 == _T_171[11:0] ? 4'h0 : _GEN_16101; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16103 = 12'h2a3 == _T_171[11:0] ? 4'h0 : _GEN_16102; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16104 = 12'h2a4 == _T_171[11:0] ? 4'h0 : _GEN_16103; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16105 = 12'h2a5 == _T_171[11:0] ? 4'h0 : _GEN_16104; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16106 = 12'h2a6 == _T_171[11:0] ? 4'h0 : _GEN_16105; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16107 = 12'h2a7 == _T_171[11:0] ? image_679 : _GEN_16106; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16108 = 12'h2a8 == _T_171[11:0] ? image_680 : _GEN_16107; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16109 = 12'h2a9 == _T_171[11:0] ? image_681 : _GEN_16108; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16110 = 12'h2aa == _T_171[11:0] ? image_682 : _GEN_16109; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16111 = 12'h2ab == _T_171[11:0] ? image_683 : _GEN_16110; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16112 = 12'h2ac == _T_171[11:0] ? image_684 : _GEN_16111; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16113 = 12'h2ad == _T_171[11:0] ? image_685 : _GEN_16112; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16114 = 12'h2ae == _T_171[11:0] ? image_686 : _GEN_16113; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16115 = 12'h2af == _T_171[11:0] ? image_687 : _GEN_16114; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16116 = 12'h2b0 == _T_171[11:0] ? image_688 : _GEN_16115; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16117 = 12'h2b1 == _T_171[11:0] ? image_689 : _GEN_16116; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16118 = 12'h2b2 == _T_171[11:0] ? image_690 : _GEN_16117; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16119 = 12'h2b3 == _T_171[11:0] ? image_691 : _GEN_16118; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16120 = 12'h2b4 == _T_171[11:0] ? image_692 : _GEN_16119; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16121 = 12'h2b5 == _T_171[11:0] ? image_693 : _GEN_16120; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16122 = 12'h2b6 == _T_171[11:0] ? image_694 : _GEN_16121; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16123 = 12'h2b7 == _T_171[11:0] ? image_695 : _GEN_16122; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16124 = 12'h2b8 == _T_171[11:0] ? image_696 : _GEN_16123; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16125 = 12'h2b9 == _T_171[11:0] ? image_697 : _GEN_16124; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16126 = 12'h2ba == _T_171[11:0] ? image_698 : _GEN_16125; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16127 = 12'h2bb == _T_171[11:0] ? 4'h0 : _GEN_16126; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16128 = 12'h2bc == _T_171[11:0] ? 4'h0 : _GEN_16127; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16129 = 12'h2bd == _T_171[11:0] ? image_701 : _GEN_16128; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16130 = 12'h2be == _T_171[11:0] ? image_702 : _GEN_16129; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16131 = 12'h2bf == _T_171[11:0] ? image_703 : _GEN_16130; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16132 = 12'h2c0 == _T_171[11:0] ? 4'h0 : _GEN_16131; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16133 = 12'h2c1 == _T_171[11:0] ? image_705 : _GEN_16132; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16134 = 12'h2c2 == _T_171[11:0] ? image_706 : _GEN_16133; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16135 = 12'h2c3 == _T_171[11:0] ? image_707 : _GEN_16134; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16136 = 12'h2c4 == _T_171[11:0] ? image_708 : _GEN_16135; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16137 = 12'h2c5 == _T_171[11:0] ? image_709 : _GEN_16136; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16138 = 12'h2c6 == _T_171[11:0] ? image_710 : _GEN_16137; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16139 = 12'h2c7 == _T_171[11:0] ? image_711 : _GEN_16138; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16140 = 12'h2c8 == _T_171[11:0] ? image_712 : _GEN_16139; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16141 = 12'h2c9 == _T_171[11:0] ? image_713 : _GEN_16140; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16142 = 12'h2ca == _T_171[11:0] ? image_714 : _GEN_16141; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16143 = 12'h2cb == _T_171[11:0] ? image_715 : _GEN_16142; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16144 = 12'h2cc == _T_171[11:0] ? image_716 : _GEN_16143; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16145 = 12'h2cd == _T_171[11:0] ? image_717 : _GEN_16144; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16146 = 12'h2ce == _T_171[11:0] ? image_718 : _GEN_16145; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16147 = 12'h2cf == _T_171[11:0] ? image_719 : _GEN_16146; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16148 = 12'h2d0 == _T_171[11:0] ? image_720 : _GEN_16147; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16149 = 12'h2d1 == _T_171[11:0] ? image_721 : _GEN_16148; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16150 = 12'h2d2 == _T_171[11:0] ? image_722 : _GEN_16149; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16151 = 12'h2d3 == _T_171[11:0] ? image_723 : _GEN_16150; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16152 = 12'h2d4 == _T_171[11:0] ? image_724 : _GEN_16151; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16153 = 12'h2d5 == _T_171[11:0] ? image_725 : _GEN_16152; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16154 = 12'h2d6 == _T_171[11:0] ? image_726 : _GEN_16153; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16155 = 12'h2d7 == _T_171[11:0] ? image_727 : _GEN_16154; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16156 = 12'h2d8 == _T_171[11:0] ? image_728 : _GEN_16155; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16157 = 12'h2d9 == _T_171[11:0] ? image_729 : _GEN_16156; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16158 = 12'h2da == _T_171[11:0] ? image_730 : _GEN_16157; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16159 = 12'h2db == _T_171[11:0] ? image_731 : _GEN_16158; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16160 = 12'h2dc == _T_171[11:0] ? image_732 : _GEN_16159; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16161 = 12'h2dd == _T_171[11:0] ? image_733 : _GEN_16160; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16162 = 12'h2de == _T_171[11:0] ? image_734 : _GEN_16161; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16163 = 12'h2df == _T_171[11:0] ? 4'h0 : _GEN_16162; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16164 = 12'h2e0 == _T_171[11:0] ? image_736 : _GEN_16163; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16165 = 12'h2e1 == _T_171[11:0] ? image_737 : _GEN_16164; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16166 = 12'h2e2 == _T_171[11:0] ? 4'h0 : _GEN_16165; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16167 = 12'h2e3 == _T_171[11:0] ? image_739 : _GEN_16166; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16168 = 12'h2e4 == _T_171[11:0] ? image_740 : _GEN_16167; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16169 = 12'h2e5 == _T_171[11:0] ? image_741 : _GEN_16168; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16170 = 12'h2e6 == _T_171[11:0] ? 4'h0 : _GEN_16169; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16171 = 12'h2e7 == _T_171[11:0] ? 4'h0 : _GEN_16170; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16172 = 12'h2e8 == _T_171[11:0] ? image_744 : _GEN_16171; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16173 = 12'h2e9 == _T_171[11:0] ? image_745 : _GEN_16172; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16174 = 12'h2ea == _T_171[11:0] ? image_746 : _GEN_16173; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16175 = 12'h2eb == _T_171[11:0] ? image_747 : _GEN_16174; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16176 = 12'h2ec == _T_171[11:0] ? image_748 : _GEN_16175; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16177 = 12'h2ed == _T_171[11:0] ? image_749 : _GEN_16176; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16178 = 12'h2ee == _T_171[11:0] ? image_750 : _GEN_16177; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16179 = 12'h2ef == _T_171[11:0] ? image_751 : _GEN_16178; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16180 = 12'h2f0 == _T_171[11:0] ? image_752 : _GEN_16179; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16181 = 12'h2f1 == _T_171[11:0] ? image_753 : _GEN_16180; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16182 = 12'h2f2 == _T_171[11:0] ? image_754 : _GEN_16181; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16183 = 12'h2f3 == _T_171[11:0] ? image_755 : _GEN_16182; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16184 = 12'h2f4 == _T_171[11:0] ? image_756 : _GEN_16183; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16185 = 12'h2f5 == _T_171[11:0] ? 4'h0 : _GEN_16184; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16186 = 12'h2f6 == _T_171[11:0] ? image_758 : _GEN_16185; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16187 = 12'h2f7 == _T_171[11:0] ? 4'h0 : _GEN_16186; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16188 = 12'h2f8 == _T_171[11:0] ? image_760 : _GEN_16187; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16189 = 12'h2f9 == _T_171[11:0] ? image_761 : _GEN_16188; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16190 = 12'h2fa == _T_171[11:0] ? image_762 : _GEN_16189; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16191 = 12'h2fb == _T_171[11:0] ? image_763 : _GEN_16190; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16192 = 12'h2fc == _T_171[11:0] ? 4'h0 : _GEN_16191; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16193 = 12'h2fd == _T_171[11:0] ? image_765 : _GEN_16192; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16194 = 12'h2fe == _T_171[11:0] ? image_766 : _GEN_16193; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16195 = 12'h2ff == _T_171[11:0] ? image_767 : _GEN_16194; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16196 = 12'h300 == _T_171[11:0] ? image_768 : _GEN_16195; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16197 = 12'h301 == _T_171[11:0] ? image_769 : _GEN_16196; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16198 = 12'h302 == _T_171[11:0] ? image_770 : _GEN_16197; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16199 = 12'h303 == _T_171[11:0] ? image_771 : _GEN_16198; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16200 = 12'h304 == _T_171[11:0] ? image_772 : _GEN_16199; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16201 = 12'h305 == _T_171[11:0] ? image_773 : _GEN_16200; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16202 = 12'h306 == _T_171[11:0] ? image_774 : _GEN_16201; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16203 = 12'h307 == _T_171[11:0] ? image_775 : _GEN_16202; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16204 = 12'h308 == _T_171[11:0] ? image_776 : _GEN_16203; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16205 = 12'h309 == _T_171[11:0] ? image_777 : _GEN_16204; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16206 = 12'h30a == _T_171[11:0] ? image_778 : _GEN_16205; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16207 = 12'h30b == _T_171[11:0] ? image_779 : _GEN_16206; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16208 = 12'h30c == _T_171[11:0] ? image_780 : _GEN_16207; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16209 = 12'h30d == _T_171[11:0] ? image_781 : _GEN_16208; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16210 = 12'h30e == _T_171[11:0] ? image_782 : _GEN_16209; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16211 = 12'h30f == _T_171[11:0] ? image_783 : _GEN_16210; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16212 = 12'h310 == _T_171[11:0] ? image_784 : _GEN_16211; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16213 = 12'h311 == _T_171[11:0] ? image_785 : _GEN_16212; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16214 = 12'h312 == _T_171[11:0] ? image_786 : _GEN_16213; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16215 = 12'h313 == _T_171[11:0] ? image_787 : _GEN_16214; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16216 = 12'h314 == _T_171[11:0] ? image_788 : _GEN_16215; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16217 = 12'h315 == _T_171[11:0] ? image_789 : _GEN_16216; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16218 = 12'h316 == _T_171[11:0] ? image_790 : _GEN_16217; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16219 = 12'h317 == _T_171[11:0] ? image_791 : _GEN_16218; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16220 = 12'h318 == _T_171[11:0] ? image_792 : _GEN_16219; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16221 = 12'h319 == _T_171[11:0] ? image_793 : _GEN_16220; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16222 = 12'h31a == _T_171[11:0] ? image_794 : _GEN_16221; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16223 = 12'h31b == _T_171[11:0] ? image_795 : _GEN_16222; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16224 = 12'h31c == _T_171[11:0] ? image_796 : _GEN_16223; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16225 = 12'h31d == _T_171[11:0] ? image_797 : _GEN_16224; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16226 = 12'h31e == _T_171[11:0] ? 4'h0 : _GEN_16225; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16227 = 12'h31f == _T_171[11:0] ? 4'h0 : _GEN_16226; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16228 = 12'h320 == _T_171[11:0] ? image_800 : _GEN_16227; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16229 = 12'h321 == _T_171[11:0] ? image_801 : _GEN_16228; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16230 = 12'h322 == _T_171[11:0] ? image_802 : _GEN_16229; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16231 = 12'h323 == _T_171[11:0] ? image_803 : _GEN_16230; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16232 = 12'h324 == _T_171[11:0] ? image_804 : _GEN_16231; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16233 = 12'h325 == _T_171[11:0] ? image_805 : _GEN_16232; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16234 = 12'h326 == _T_171[11:0] ? image_806 : _GEN_16233; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16235 = 12'h327 == _T_171[11:0] ? 4'h0 : _GEN_16234; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16236 = 12'h328 == _T_171[11:0] ? image_808 : _GEN_16235; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16237 = 12'h329 == _T_171[11:0] ? image_809 : _GEN_16236; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16238 = 12'h32a == _T_171[11:0] ? image_810 : _GEN_16237; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16239 = 12'h32b == _T_171[11:0] ? image_811 : _GEN_16238; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16240 = 12'h32c == _T_171[11:0] ? image_812 : _GEN_16239; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16241 = 12'h32d == _T_171[11:0] ? image_813 : _GEN_16240; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16242 = 12'h32e == _T_171[11:0] ? image_814 : _GEN_16241; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16243 = 12'h32f == _T_171[11:0] ? image_815 : _GEN_16242; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16244 = 12'h330 == _T_171[11:0] ? image_816 : _GEN_16243; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16245 = 12'h331 == _T_171[11:0] ? image_817 : _GEN_16244; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16246 = 12'h332 == _T_171[11:0] ? image_818 : _GEN_16245; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16247 = 12'h333 == _T_171[11:0] ? image_819 : _GEN_16246; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16248 = 12'h334 == _T_171[11:0] ? image_820 : _GEN_16247; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16249 = 12'h335 == _T_171[11:0] ? 4'h0 : _GEN_16248; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16250 = 12'h336 == _T_171[11:0] ? image_822 : _GEN_16249; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16251 = 12'h337 == _T_171[11:0] ? image_823 : _GEN_16250; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16252 = 12'h338 == _T_171[11:0] ? image_824 : _GEN_16251; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16253 = 12'h339 == _T_171[11:0] ? image_825 : _GEN_16252; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16254 = 12'h33a == _T_171[11:0] ? image_826 : _GEN_16253; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16255 = 12'h33b == _T_171[11:0] ? 4'h0 : _GEN_16254; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16256 = 12'h33c == _T_171[11:0] ? image_828 : _GEN_16255; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16257 = 12'h33d == _T_171[11:0] ? image_829 : _GEN_16256; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16258 = 12'h33e == _T_171[11:0] ? image_830 : _GEN_16257; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16259 = 12'h33f == _T_171[11:0] ? image_831 : _GEN_16258; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16260 = 12'h340 == _T_171[11:0] ? 4'h0 : _GEN_16259; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16261 = 12'h341 == _T_171[11:0] ? image_833 : _GEN_16260; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16262 = 12'h342 == _T_171[11:0] ? image_834 : _GEN_16261; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16263 = 12'h343 == _T_171[11:0] ? image_835 : _GEN_16262; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16264 = 12'h344 == _T_171[11:0] ? image_836 : _GEN_16263; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16265 = 12'h345 == _T_171[11:0] ? image_837 : _GEN_16264; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16266 = 12'h346 == _T_171[11:0] ? image_838 : _GEN_16265; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16267 = 12'h347 == _T_171[11:0] ? image_839 : _GEN_16266; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16268 = 12'h348 == _T_171[11:0] ? image_840 : _GEN_16267; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16269 = 12'h349 == _T_171[11:0] ? image_841 : _GEN_16268; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16270 = 12'h34a == _T_171[11:0] ? image_842 : _GEN_16269; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16271 = 12'h34b == _T_171[11:0] ? image_843 : _GEN_16270; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16272 = 12'h34c == _T_171[11:0] ? image_844 : _GEN_16271; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16273 = 12'h34d == _T_171[11:0] ? image_845 : _GEN_16272; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16274 = 12'h34e == _T_171[11:0] ? image_846 : _GEN_16273; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16275 = 12'h34f == _T_171[11:0] ? image_847 : _GEN_16274; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16276 = 12'h350 == _T_171[11:0] ? image_848 : _GEN_16275; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16277 = 12'h351 == _T_171[11:0] ? image_849 : _GEN_16276; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16278 = 12'h352 == _T_171[11:0] ? image_850 : _GEN_16277; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16279 = 12'h353 == _T_171[11:0] ? image_851 : _GEN_16278; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16280 = 12'h354 == _T_171[11:0] ? image_852 : _GEN_16279; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16281 = 12'h355 == _T_171[11:0] ? image_853 : _GEN_16280; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16282 = 12'h356 == _T_171[11:0] ? image_854 : _GEN_16281; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16283 = 12'h357 == _T_171[11:0] ? image_855 : _GEN_16282; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16284 = 12'h358 == _T_171[11:0] ? image_856 : _GEN_16283; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16285 = 12'h359 == _T_171[11:0] ? image_857 : _GEN_16284; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16286 = 12'h35a == _T_171[11:0] ? image_858 : _GEN_16285; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16287 = 12'h35b == _T_171[11:0] ? image_859 : _GEN_16286; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16288 = 12'h35c == _T_171[11:0] ? image_860 : _GEN_16287; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16289 = 12'h35d == _T_171[11:0] ? image_861 : _GEN_16288; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16290 = 12'h35e == _T_171[11:0] ? image_862 : _GEN_16289; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16291 = 12'h35f == _T_171[11:0] ? 4'h0 : _GEN_16290; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16292 = 12'h360 == _T_171[11:0] ? 4'h0 : _GEN_16291; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16293 = 12'h361 == _T_171[11:0] ? image_865 : _GEN_16292; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16294 = 12'h362 == _T_171[11:0] ? image_866 : _GEN_16293; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16295 = 12'h363 == _T_171[11:0] ? image_867 : _GEN_16294; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16296 = 12'h364 == _T_171[11:0] ? image_868 : _GEN_16295; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16297 = 12'h365 == _T_171[11:0] ? image_869 : _GEN_16296; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16298 = 12'h366 == _T_171[11:0] ? 4'h0 : _GEN_16297; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16299 = 12'h367 == _T_171[11:0] ? 4'h0 : _GEN_16298; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16300 = 12'h368 == _T_171[11:0] ? image_872 : _GEN_16299; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16301 = 12'h369 == _T_171[11:0] ? image_873 : _GEN_16300; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16302 = 12'h36a == _T_171[11:0] ? image_874 : _GEN_16301; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16303 = 12'h36b == _T_171[11:0] ? image_875 : _GEN_16302; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16304 = 12'h36c == _T_171[11:0] ? image_876 : _GEN_16303; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16305 = 12'h36d == _T_171[11:0] ? image_877 : _GEN_16304; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16306 = 12'h36e == _T_171[11:0] ? image_878 : _GEN_16305; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16307 = 12'h36f == _T_171[11:0] ? image_879 : _GEN_16306; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16308 = 12'h370 == _T_171[11:0] ? image_880 : _GEN_16307; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16309 = 12'h371 == _T_171[11:0] ? image_881 : _GEN_16308; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16310 = 12'h372 == _T_171[11:0] ? image_882 : _GEN_16309; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16311 = 12'h373 == _T_171[11:0] ? image_883 : _GEN_16310; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16312 = 12'h374 == _T_171[11:0] ? image_884 : _GEN_16311; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16313 = 12'h375 == _T_171[11:0] ? image_885 : _GEN_16312; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16314 = 12'h376 == _T_171[11:0] ? 4'h0 : _GEN_16313; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16315 = 12'h377 == _T_171[11:0] ? 4'h0 : _GEN_16314; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16316 = 12'h378 == _T_171[11:0] ? 4'h0 : _GEN_16315; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16317 = 12'h379 == _T_171[11:0] ? 4'h0 : _GEN_16316; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16318 = 12'h37a == _T_171[11:0] ? 4'h0 : _GEN_16317; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16319 = 12'h37b == _T_171[11:0] ? image_891 : _GEN_16318; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16320 = 12'h37c == _T_171[11:0] ? image_892 : _GEN_16319; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16321 = 12'h37d == _T_171[11:0] ? image_893 : _GEN_16320; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16322 = 12'h37e == _T_171[11:0] ? image_894 : _GEN_16321; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16323 = 12'h37f == _T_171[11:0] ? image_895 : _GEN_16322; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16324 = 12'h380 == _T_171[11:0] ? 4'h0 : _GEN_16323; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16325 = 12'h381 == _T_171[11:0] ? image_897 : _GEN_16324; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16326 = 12'h382 == _T_171[11:0] ? image_898 : _GEN_16325; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16327 = 12'h383 == _T_171[11:0] ? image_899 : _GEN_16326; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16328 = 12'h384 == _T_171[11:0] ? image_900 : _GEN_16327; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16329 = 12'h385 == _T_171[11:0] ? image_901 : _GEN_16328; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16330 = 12'h386 == _T_171[11:0] ? image_902 : _GEN_16329; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16331 = 12'h387 == _T_171[11:0] ? image_903 : _GEN_16330; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16332 = 12'h388 == _T_171[11:0] ? image_904 : _GEN_16331; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16333 = 12'h389 == _T_171[11:0] ? image_905 : _GEN_16332; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16334 = 12'h38a == _T_171[11:0] ? image_906 : _GEN_16333; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16335 = 12'h38b == _T_171[11:0] ? image_907 : _GEN_16334; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16336 = 12'h38c == _T_171[11:0] ? image_908 : _GEN_16335; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16337 = 12'h38d == _T_171[11:0] ? image_909 : _GEN_16336; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16338 = 12'h38e == _T_171[11:0] ? image_910 : _GEN_16337; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16339 = 12'h38f == _T_171[11:0] ? image_911 : _GEN_16338; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16340 = 12'h390 == _T_171[11:0] ? image_912 : _GEN_16339; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16341 = 12'h391 == _T_171[11:0] ? image_913 : _GEN_16340; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16342 = 12'h392 == _T_171[11:0] ? image_914 : _GEN_16341; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16343 = 12'h393 == _T_171[11:0] ? image_915 : _GEN_16342; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16344 = 12'h394 == _T_171[11:0] ? image_916 : _GEN_16343; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16345 = 12'h395 == _T_171[11:0] ? image_917 : _GEN_16344; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16346 = 12'h396 == _T_171[11:0] ? image_918 : _GEN_16345; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16347 = 12'h397 == _T_171[11:0] ? image_919 : _GEN_16346; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16348 = 12'h398 == _T_171[11:0] ? image_920 : _GEN_16347; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16349 = 12'h399 == _T_171[11:0] ? image_921 : _GEN_16348; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16350 = 12'h39a == _T_171[11:0] ? image_922 : _GEN_16349; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16351 = 12'h39b == _T_171[11:0] ? image_923 : _GEN_16350; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16352 = 12'h39c == _T_171[11:0] ? image_924 : _GEN_16351; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16353 = 12'h39d == _T_171[11:0] ? image_925 : _GEN_16352; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16354 = 12'h39e == _T_171[11:0] ? image_926 : _GEN_16353; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16355 = 12'h39f == _T_171[11:0] ? image_927 : _GEN_16354; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16356 = 12'h3a0 == _T_171[11:0] ? 4'h0 : _GEN_16355; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16357 = 12'h3a1 == _T_171[11:0] ? image_929 : _GEN_16356; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16358 = 12'h3a2 == _T_171[11:0] ? image_930 : _GEN_16357; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16359 = 12'h3a3 == _T_171[11:0] ? 4'h0 : _GEN_16358; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16360 = 12'h3a4 == _T_171[11:0] ? 4'h0 : _GEN_16359; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16361 = 12'h3a5 == _T_171[11:0] ? 4'h0 : _GEN_16360; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16362 = 12'h3a6 == _T_171[11:0] ? 4'h0 : _GEN_16361; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16363 = 12'h3a7 == _T_171[11:0] ? image_935 : _GEN_16362; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16364 = 12'h3a8 == _T_171[11:0] ? image_936 : _GEN_16363; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16365 = 12'h3a9 == _T_171[11:0] ? image_937 : _GEN_16364; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16366 = 12'h3aa == _T_171[11:0] ? image_938 : _GEN_16365; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16367 = 12'h3ab == _T_171[11:0] ? image_939 : _GEN_16366; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16368 = 12'h3ac == _T_171[11:0] ? image_940 : _GEN_16367; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16369 = 12'h3ad == _T_171[11:0] ? image_941 : _GEN_16368; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16370 = 12'h3ae == _T_171[11:0] ? image_942 : _GEN_16369; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16371 = 12'h3af == _T_171[11:0] ? image_943 : _GEN_16370; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16372 = 12'h3b0 == _T_171[11:0] ? image_944 : _GEN_16371; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16373 = 12'h3b1 == _T_171[11:0] ? image_945 : _GEN_16372; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16374 = 12'h3b2 == _T_171[11:0] ? image_946 : _GEN_16373; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16375 = 12'h3b3 == _T_171[11:0] ? image_947 : _GEN_16374; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16376 = 12'h3b4 == _T_171[11:0] ? image_948 : _GEN_16375; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16377 = 12'h3b5 == _T_171[11:0] ? image_949 : _GEN_16376; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16378 = 12'h3b6 == _T_171[11:0] ? image_950 : _GEN_16377; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16379 = 12'h3b7 == _T_171[11:0] ? image_951 : _GEN_16378; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16380 = 12'h3b8 == _T_171[11:0] ? image_952 : _GEN_16379; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16381 = 12'h3b9 == _T_171[11:0] ? image_953 : _GEN_16380; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16382 = 12'h3ba == _T_171[11:0] ? image_954 : _GEN_16381; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16383 = 12'h3bb == _T_171[11:0] ? image_955 : _GEN_16382; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16384 = 12'h3bc == _T_171[11:0] ? image_956 : _GEN_16383; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16385 = 12'h3bd == _T_171[11:0] ? image_957 : _GEN_16384; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16386 = 12'h3be == _T_171[11:0] ? image_958 : _GEN_16385; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16387 = 12'h3bf == _T_171[11:0] ? image_959 : _GEN_16386; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16388 = 12'h3c0 == _T_171[11:0] ? 4'h0 : _GEN_16387; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16389 = 12'h3c1 == _T_171[11:0] ? image_961 : _GEN_16388; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16390 = 12'h3c2 == _T_171[11:0] ? image_962 : _GEN_16389; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16391 = 12'h3c3 == _T_171[11:0] ? image_963 : _GEN_16390; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16392 = 12'h3c4 == _T_171[11:0] ? image_964 : _GEN_16391; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16393 = 12'h3c5 == _T_171[11:0] ? image_965 : _GEN_16392; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16394 = 12'h3c6 == _T_171[11:0] ? image_966 : _GEN_16393; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16395 = 12'h3c7 == _T_171[11:0] ? image_967 : _GEN_16394; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16396 = 12'h3c8 == _T_171[11:0] ? image_968 : _GEN_16395; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16397 = 12'h3c9 == _T_171[11:0] ? image_969 : _GEN_16396; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16398 = 12'h3ca == _T_171[11:0] ? image_970 : _GEN_16397; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16399 = 12'h3cb == _T_171[11:0] ? image_971 : _GEN_16398; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16400 = 12'h3cc == _T_171[11:0] ? image_972 : _GEN_16399; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16401 = 12'h3cd == _T_171[11:0] ? image_973 : _GEN_16400; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16402 = 12'h3ce == _T_171[11:0] ? image_974 : _GEN_16401; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16403 = 12'h3cf == _T_171[11:0] ? image_975 : _GEN_16402; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16404 = 12'h3d0 == _T_171[11:0] ? image_976 : _GEN_16403; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16405 = 12'h3d1 == _T_171[11:0] ? image_977 : _GEN_16404; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16406 = 12'h3d2 == _T_171[11:0] ? image_978 : _GEN_16405; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16407 = 12'h3d3 == _T_171[11:0] ? image_979 : _GEN_16406; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16408 = 12'h3d4 == _T_171[11:0] ? image_980 : _GEN_16407; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16409 = 12'h3d5 == _T_171[11:0] ? image_981 : _GEN_16408; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16410 = 12'h3d6 == _T_171[11:0] ? image_982 : _GEN_16409; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16411 = 12'h3d7 == _T_171[11:0] ? image_983 : _GEN_16410; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16412 = 12'h3d8 == _T_171[11:0] ? image_984 : _GEN_16411; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16413 = 12'h3d9 == _T_171[11:0] ? image_985 : _GEN_16412; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16414 = 12'h3da == _T_171[11:0] ? image_986 : _GEN_16413; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16415 = 12'h3db == _T_171[11:0] ? image_987 : _GEN_16414; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16416 = 12'h3dc == _T_171[11:0] ? image_988 : _GEN_16415; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16417 = 12'h3dd == _T_171[11:0] ? image_989 : _GEN_16416; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16418 = 12'h3de == _T_171[11:0] ? image_990 : _GEN_16417; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16419 = 12'h3df == _T_171[11:0] ? image_991 : _GEN_16418; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16420 = 12'h3e0 == _T_171[11:0] ? image_992 : _GEN_16419; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16421 = 12'h3e1 == _T_171[11:0] ? 4'h0 : _GEN_16420; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16422 = 12'h3e2 == _T_171[11:0] ? 4'h0 : _GEN_16421; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16423 = 12'h3e3 == _T_171[11:0] ? 4'h0 : _GEN_16422; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16424 = 12'h3e4 == _T_171[11:0] ? 4'h0 : _GEN_16423; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16425 = 12'h3e5 == _T_171[11:0] ? image_997 : _GEN_16424; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16426 = 12'h3e6 == _T_171[11:0] ? image_998 : _GEN_16425; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16427 = 12'h3e7 == _T_171[11:0] ? image_999 : _GEN_16426; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16428 = 12'h3e8 == _T_171[11:0] ? image_1000 : _GEN_16427; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16429 = 12'h3e9 == _T_171[11:0] ? image_1001 : _GEN_16428; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16430 = 12'h3ea == _T_171[11:0] ? image_1002 : _GEN_16429; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16431 = 12'h3eb == _T_171[11:0] ? image_1003 : _GEN_16430; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16432 = 12'h3ec == _T_171[11:0] ? image_1004 : _GEN_16431; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16433 = 12'h3ed == _T_171[11:0] ? image_1005 : _GEN_16432; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16434 = 12'h3ee == _T_171[11:0] ? image_1006 : _GEN_16433; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16435 = 12'h3ef == _T_171[11:0] ? image_1007 : _GEN_16434; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16436 = 12'h3f0 == _T_171[11:0] ? image_1008 : _GEN_16435; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16437 = 12'h3f1 == _T_171[11:0] ? image_1009 : _GEN_16436; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16438 = 12'h3f2 == _T_171[11:0] ? image_1010 : _GEN_16437; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16439 = 12'h3f3 == _T_171[11:0] ? image_1011 : _GEN_16438; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16440 = 12'h3f4 == _T_171[11:0] ? image_1012 : _GEN_16439; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16441 = 12'h3f5 == _T_171[11:0] ? image_1013 : _GEN_16440; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16442 = 12'h3f6 == _T_171[11:0] ? image_1014 : _GEN_16441; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16443 = 12'h3f7 == _T_171[11:0] ? image_1015 : _GEN_16442; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16444 = 12'h3f8 == _T_171[11:0] ? image_1016 : _GEN_16443; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16445 = 12'h3f9 == _T_171[11:0] ? image_1017 : _GEN_16444; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16446 = 12'h3fa == _T_171[11:0] ? image_1018 : _GEN_16445; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16447 = 12'h3fb == _T_171[11:0] ? image_1019 : _GEN_16446; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16448 = 12'h3fc == _T_171[11:0] ? image_1020 : _GEN_16447; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16449 = 12'h3fd == _T_171[11:0] ? 4'h0 : _GEN_16448; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16450 = 12'h3fe == _T_171[11:0] ? 4'h0 : _GEN_16449; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16451 = 12'h3ff == _T_171[11:0] ? 4'h0 : _GEN_16450; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16452 = 12'h400 == _T_171[11:0] ? image_1024 : _GEN_16451; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16453 = 12'h401 == _T_171[11:0] ? image_1025 : _GEN_16452; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16454 = 12'h402 == _T_171[11:0] ? image_1026 : _GEN_16453; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16455 = 12'h403 == _T_171[11:0] ? image_1027 : _GEN_16454; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16456 = 12'h404 == _T_171[11:0] ? image_1028 : _GEN_16455; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16457 = 12'h405 == _T_171[11:0] ? image_1029 : _GEN_16456; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16458 = 12'h406 == _T_171[11:0] ? image_1030 : _GEN_16457; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16459 = 12'h407 == _T_171[11:0] ? image_1031 : _GEN_16458; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16460 = 12'h408 == _T_171[11:0] ? image_1032 : _GEN_16459; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16461 = 12'h409 == _T_171[11:0] ? image_1033 : _GEN_16460; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16462 = 12'h40a == _T_171[11:0] ? image_1034 : _GEN_16461; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16463 = 12'h40b == _T_171[11:0] ? image_1035 : _GEN_16462; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16464 = 12'h40c == _T_171[11:0] ? image_1036 : _GEN_16463; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16465 = 12'h40d == _T_171[11:0] ? image_1037 : _GEN_16464; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16466 = 12'h40e == _T_171[11:0] ? image_1038 : _GEN_16465; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16467 = 12'h40f == _T_171[11:0] ? image_1039 : _GEN_16466; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16468 = 12'h410 == _T_171[11:0] ? image_1040 : _GEN_16467; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16469 = 12'h411 == _T_171[11:0] ? image_1041 : _GEN_16468; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16470 = 12'h412 == _T_171[11:0] ? image_1042 : _GEN_16469; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16471 = 12'h413 == _T_171[11:0] ? image_1043 : _GEN_16470; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16472 = 12'h414 == _T_171[11:0] ? image_1044 : _GEN_16471; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16473 = 12'h415 == _T_171[11:0] ? image_1045 : _GEN_16472; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16474 = 12'h416 == _T_171[11:0] ? image_1046 : _GEN_16473; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16475 = 12'h417 == _T_171[11:0] ? image_1047 : _GEN_16474; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16476 = 12'h418 == _T_171[11:0] ? image_1048 : _GEN_16475; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16477 = 12'h419 == _T_171[11:0] ? image_1049 : _GEN_16476; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16478 = 12'h41a == _T_171[11:0] ? image_1050 : _GEN_16477; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16479 = 12'h41b == _T_171[11:0] ? image_1051 : _GEN_16478; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16480 = 12'h41c == _T_171[11:0] ? image_1052 : _GEN_16479; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16481 = 12'h41d == _T_171[11:0] ? image_1053 : _GEN_16480; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16482 = 12'h41e == _T_171[11:0] ? image_1054 : _GEN_16481; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16483 = 12'h41f == _T_171[11:0] ? image_1055 : _GEN_16482; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16484 = 12'h420 == _T_171[11:0] ? image_1056 : _GEN_16483; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16485 = 12'h421 == _T_171[11:0] ? image_1057 : _GEN_16484; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16486 = 12'h422 == _T_171[11:0] ? image_1058 : _GEN_16485; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16487 = 12'h423 == _T_171[11:0] ? image_1059 : _GEN_16486; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16488 = 12'h424 == _T_171[11:0] ? image_1060 : _GEN_16487; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16489 = 12'h425 == _T_171[11:0] ? image_1061 : _GEN_16488; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16490 = 12'h426 == _T_171[11:0] ? image_1062 : _GEN_16489; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16491 = 12'h427 == _T_171[11:0] ? image_1063 : _GEN_16490; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16492 = 12'h428 == _T_171[11:0] ? image_1064 : _GEN_16491; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16493 = 12'h429 == _T_171[11:0] ? image_1065 : _GEN_16492; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16494 = 12'h42a == _T_171[11:0] ? image_1066 : _GEN_16493; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16495 = 12'h42b == _T_171[11:0] ? image_1067 : _GEN_16494; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16496 = 12'h42c == _T_171[11:0] ? image_1068 : _GEN_16495; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16497 = 12'h42d == _T_171[11:0] ? image_1069 : _GEN_16496; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16498 = 12'h42e == _T_171[11:0] ? image_1070 : _GEN_16497; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16499 = 12'h42f == _T_171[11:0] ? image_1071 : _GEN_16498; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16500 = 12'h430 == _T_171[11:0] ? image_1072 : _GEN_16499; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16501 = 12'h431 == _T_171[11:0] ? image_1073 : _GEN_16500; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16502 = 12'h432 == _T_171[11:0] ? image_1074 : _GEN_16501; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16503 = 12'h433 == _T_171[11:0] ? image_1075 : _GEN_16502; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16504 = 12'h434 == _T_171[11:0] ? image_1076 : _GEN_16503; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16505 = 12'h435 == _T_171[11:0] ? image_1077 : _GEN_16504; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16506 = 12'h436 == _T_171[11:0] ? image_1078 : _GEN_16505; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16507 = 12'h437 == _T_171[11:0] ? image_1079 : _GEN_16506; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16508 = 12'h438 == _T_171[11:0] ? image_1080 : _GEN_16507; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16509 = 12'h439 == _T_171[11:0] ? image_1081 : _GEN_16508; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16510 = 12'h43a == _T_171[11:0] ? image_1082 : _GEN_16509; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16511 = 12'h43b == _T_171[11:0] ? image_1083 : _GEN_16510; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16512 = 12'h43c == _T_171[11:0] ? image_1084 : _GEN_16511; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16513 = 12'h43d == _T_171[11:0] ? image_1085 : _GEN_16512; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16514 = 12'h43e == _T_171[11:0] ? 4'h0 : _GEN_16513; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16515 = 12'h43f == _T_171[11:0] ? 4'h0 : _GEN_16514; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16516 = 12'h440 == _T_171[11:0] ? image_1088 : _GEN_16515; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16517 = 12'h441 == _T_171[11:0] ? image_1089 : _GEN_16516; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16518 = 12'h442 == _T_171[11:0] ? image_1090 : _GEN_16517; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16519 = 12'h443 == _T_171[11:0] ? image_1091 : _GEN_16518; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16520 = 12'h444 == _T_171[11:0] ? image_1092 : _GEN_16519; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16521 = 12'h445 == _T_171[11:0] ? image_1093 : _GEN_16520; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16522 = 12'h446 == _T_171[11:0] ? image_1094 : _GEN_16521; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16523 = 12'h447 == _T_171[11:0] ? image_1095 : _GEN_16522; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16524 = 12'h448 == _T_171[11:0] ? image_1096 : _GEN_16523; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16525 = 12'h449 == _T_171[11:0] ? image_1097 : _GEN_16524; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16526 = 12'h44a == _T_171[11:0] ? image_1098 : _GEN_16525; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16527 = 12'h44b == _T_171[11:0] ? image_1099 : _GEN_16526; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16528 = 12'h44c == _T_171[11:0] ? image_1100 : _GEN_16527; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16529 = 12'h44d == _T_171[11:0] ? image_1101 : _GEN_16528; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16530 = 12'h44e == _T_171[11:0] ? image_1102 : _GEN_16529; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16531 = 12'h44f == _T_171[11:0] ? image_1103 : _GEN_16530; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16532 = 12'h450 == _T_171[11:0] ? image_1104 : _GEN_16531; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16533 = 12'h451 == _T_171[11:0] ? image_1105 : _GEN_16532; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16534 = 12'h452 == _T_171[11:0] ? image_1106 : _GEN_16533; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16535 = 12'h453 == _T_171[11:0] ? image_1107 : _GEN_16534; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16536 = 12'h454 == _T_171[11:0] ? image_1108 : _GEN_16535; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16537 = 12'h455 == _T_171[11:0] ? image_1109 : _GEN_16536; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16538 = 12'h456 == _T_171[11:0] ? image_1110 : _GEN_16537; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16539 = 12'h457 == _T_171[11:0] ? image_1111 : _GEN_16538; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16540 = 12'h458 == _T_171[11:0] ? image_1112 : _GEN_16539; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16541 = 12'h459 == _T_171[11:0] ? image_1113 : _GEN_16540; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16542 = 12'h45a == _T_171[11:0] ? image_1114 : _GEN_16541; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16543 = 12'h45b == _T_171[11:0] ? image_1115 : _GEN_16542; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16544 = 12'h45c == _T_171[11:0] ? image_1116 : _GEN_16543; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16545 = 12'h45d == _T_171[11:0] ? image_1117 : _GEN_16544; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16546 = 12'h45e == _T_171[11:0] ? image_1118 : _GEN_16545; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16547 = 12'h45f == _T_171[11:0] ? image_1119 : _GEN_16546; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16548 = 12'h460 == _T_171[11:0] ? image_1120 : _GEN_16547; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16549 = 12'h461 == _T_171[11:0] ? image_1121 : _GEN_16548; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16550 = 12'h462 == _T_171[11:0] ? image_1122 : _GEN_16549; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16551 = 12'h463 == _T_171[11:0] ? image_1123 : _GEN_16550; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16552 = 12'h464 == _T_171[11:0] ? image_1124 : _GEN_16551; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16553 = 12'h465 == _T_171[11:0] ? image_1125 : _GEN_16552; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16554 = 12'h466 == _T_171[11:0] ? image_1126 : _GEN_16553; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16555 = 12'h467 == _T_171[11:0] ? image_1127 : _GEN_16554; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16556 = 12'h468 == _T_171[11:0] ? image_1128 : _GEN_16555; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16557 = 12'h469 == _T_171[11:0] ? image_1129 : _GEN_16556; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16558 = 12'h46a == _T_171[11:0] ? image_1130 : _GEN_16557; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16559 = 12'h46b == _T_171[11:0] ? image_1131 : _GEN_16558; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16560 = 12'h46c == _T_171[11:0] ? image_1132 : _GEN_16559; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16561 = 12'h46d == _T_171[11:0] ? image_1133 : _GEN_16560; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16562 = 12'h46e == _T_171[11:0] ? image_1134 : _GEN_16561; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16563 = 12'h46f == _T_171[11:0] ? image_1135 : _GEN_16562; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16564 = 12'h470 == _T_171[11:0] ? image_1136 : _GEN_16563; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16565 = 12'h471 == _T_171[11:0] ? image_1137 : _GEN_16564; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16566 = 12'h472 == _T_171[11:0] ? image_1138 : _GEN_16565; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16567 = 12'h473 == _T_171[11:0] ? image_1139 : _GEN_16566; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16568 = 12'h474 == _T_171[11:0] ? image_1140 : _GEN_16567; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16569 = 12'h475 == _T_171[11:0] ? image_1141 : _GEN_16568; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16570 = 12'h476 == _T_171[11:0] ? image_1142 : _GEN_16569; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16571 = 12'h477 == _T_171[11:0] ? image_1143 : _GEN_16570; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16572 = 12'h478 == _T_171[11:0] ? image_1144 : _GEN_16571; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16573 = 12'h479 == _T_171[11:0] ? image_1145 : _GEN_16572; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16574 = 12'h47a == _T_171[11:0] ? image_1146 : _GEN_16573; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16575 = 12'h47b == _T_171[11:0] ? image_1147 : _GEN_16574; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16576 = 12'h47c == _T_171[11:0] ? image_1148 : _GEN_16575; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16577 = 12'h47d == _T_171[11:0] ? 4'h0 : _GEN_16576; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16578 = 12'h47e == _T_171[11:0] ? 4'h0 : _GEN_16577; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16579 = 12'h47f == _T_171[11:0] ? 4'h0 : _GEN_16578; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16580 = 12'h480 == _T_171[11:0] ? image_1152 : _GEN_16579; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16581 = 12'h481 == _T_171[11:0] ? image_1153 : _GEN_16580; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16582 = 12'h482 == _T_171[11:0] ? image_1154 : _GEN_16581; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16583 = 12'h483 == _T_171[11:0] ? image_1155 : _GEN_16582; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16584 = 12'h484 == _T_171[11:0] ? image_1156 : _GEN_16583; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16585 = 12'h485 == _T_171[11:0] ? image_1157 : _GEN_16584; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16586 = 12'h486 == _T_171[11:0] ? image_1158 : _GEN_16585; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16587 = 12'h487 == _T_171[11:0] ? image_1159 : _GEN_16586; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16588 = 12'h488 == _T_171[11:0] ? image_1160 : _GEN_16587; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16589 = 12'h489 == _T_171[11:0] ? image_1161 : _GEN_16588; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16590 = 12'h48a == _T_171[11:0] ? image_1162 : _GEN_16589; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16591 = 12'h48b == _T_171[11:0] ? image_1163 : _GEN_16590; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16592 = 12'h48c == _T_171[11:0] ? image_1164 : _GEN_16591; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16593 = 12'h48d == _T_171[11:0] ? image_1165 : _GEN_16592; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16594 = 12'h48e == _T_171[11:0] ? image_1166 : _GEN_16593; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16595 = 12'h48f == _T_171[11:0] ? image_1167 : _GEN_16594; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16596 = 12'h490 == _T_171[11:0] ? image_1168 : _GEN_16595; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16597 = 12'h491 == _T_171[11:0] ? image_1169 : _GEN_16596; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16598 = 12'h492 == _T_171[11:0] ? image_1170 : _GEN_16597; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16599 = 12'h493 == _T_171[11:0] ? image_1171 : _GEN_16598; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16600 = 12'h494 == _T_171[11:0] ? image_1172 : _GEN_16599; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16601 = 12'h495 == _T_171[11:0] ? image_1173 : _GEN_16600; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16602 = 12'h496 == _T_171[11:0] ? image_1174 : _GEN_16601; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16603 = 12'h497 == _T_171[11:0] ? image_1175 : _GEN_16602; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16604 = 12'h498 == _T_171[11:0] ? image_1176 : _GEN_16603; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16605 = 12'h499 == _T_171[11:0] ? image_1177 : _GEN_16604; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16606 = 12'h49a == _T_171[11:0] ? image_1178 : _GEN_16605; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16607 = 12'h49b == _T_171[11:0] ? image_1179 : _GEN_16606; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16608 = 12'h49c == _T_171[11:0] ? image_1180 : _GEN_16607; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16609 = 12'h49d == _T_171[11:0] ? image_1181 : _GEN_16608; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16610 = 12'h49e == _T_171[11:0] ? image_1182 : _GEN_16609; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16611 = 12'h49f == _T_171[11:0] ? image_1183 : _GEN_16610; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16612 = 12'h4a0 == _T_171[11:0] ? image_1184 : _GEN_16611; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16613 = 12'h4a1 == _T_171[11:0] ? image_1185 : _GEN_16612; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16614 = 12'h4a2 == _T_171[11:0] ? image_1186 : _GEN_16613; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16615 = 12'h4a3 == _T_171[11:0] ? image_1187 : _GEN_16614; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16616 = 12'h4a4 == _T_171[11:0] ? image_1188 : _GEN_16615; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16617 = 12'h4a5 == _T_171[11:0] ? image_1189 : _GEN_16616; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16618 = 12'h4a6 == _T_171[11:0] ? image_1190 : _GEN_16617; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16619 = 12'h4a7 == _T_171[11:0] ? image_1191 : _GEN_16618; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16620 = 12'h4a8 == _T_171[11:0] ? image_1192 : _GEN_16619; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16621 = 12'h4a9 == _T_171[11:0] ? image_1193 : _GEN_16620; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16622 = 12'h4aa == _T_171[11:0] ? image_1194 : _GEN_16621; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16623 = 12'h4ab == _T_171[11:0] ? image_1195 : _GEN_16622; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16624 = 12'h4ac == _T_171[11:0] ? image_1196 : _GEN_16623; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16625 = 12'h4ad == _T_171[11:0] ? image_1197 : _GEN_16624; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16626 = 12'h4ae == _T_171[11:0] ? image_1198 : _GEN_16625; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16627 = 12'h4af == _T_171[11:0] ? image_1199 : _GEN_16626; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16628 = 12'h4b0 == _T_171[11:0] ? image_1200 : _GEN_16627; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16629 = 12'h4b1 == _T_171[11:0] ? image_1201 : _GEN_16628; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16630 = 12'h4b2 == _T_171[11:0] ? image_1202 : _GEN_16629; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16631 = 12'h4b3 == _T_171[11:0] ? image_1203 : _GEN_16630; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16632 = 12'h4b4 == _T_171[11:0] ? image_1204 : _GEN_16631; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16633 = 12'h4b5 == _T_171[11:0] ? image_1205 : _GEN_16632; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16634 = 12'h4b6 == _T_171[11:0] ? image_1206 : _GEN_16633; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16635 = 12'h4b7 == _T_171[11:0] ? image_1207 : _GEN_16634; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16636 = 12'h4b8 == _T_171[11:0] ? image_1208 : _GEN_16635; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16637 = 12'h4b9 == _T_171[11:0] ? 4'h0 : _GEN_16636; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16638 = 12'h4ba == _T_171[11:0] ? 4'h0 : _GEN_16637; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16639 = 12'h4bb == _T_171[11:0] ? 4'h0 : _GEN_16638; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16640 = 12'h4bc == _T_171[11:0] ? 4'h0 : _GEN_16639; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16641 = 12'h4bd == _T_171[11:0] ? 4'h0 : _GEN_16640; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16642 = 12'h4be == _T_171[11:0] ? 4'h0 : _GEN_16641; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16643 = 12'h4bf == _T_171[11:0] ? 4'h0 : _GEN_16642; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16644 = 12'h4c0 == _T_171[11:0] ? image_1216 : _GEN_16643; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16645 = 12'h4c1 == _T_171[11:0] ? image_1217 : _GEN_16644; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16646 = 12'h4c2 == _T_171[11:0] ? image_1218 : _GEN_16645; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16647 = 12'h4c3 == _T_171[11:0] ? image_1219 : _GEN_16646; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16648 = 12'h4c4 == _T_171[11:0] ? image_1220 : _GEN_16647; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16649 = 12'h4c5 == _T_171[11:0] ? image_1221 : _GEN_16648; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16650 = 12'h4c6 == _T_171[11:0] ? image_1222 : _GEN_16649; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16651 = 12'h4c7 == _T_171[11:0] ? image_1223 : _GEN_16650; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16652 = 12'h4c8 == _T_171[11:0] ? image_1224 : _GEN_16651; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16653 = 12'h4c9 == _T_171[11:0] ? image_1225 : _GEN_16652; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16654 = 12'h4ca == _T_171[11:0] ? image_1226 : _GEN_16653; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16655 = 12'h4cb == _T_171[11:0] ? image_1227 : _GEN_16654; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16656 = 12'h4cc == _T_171[11:0] ? image_1228 : _GEN_16655; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16657 = 12'h4cd == _T_171[11:0] ? image_1229 : _GEN_16656; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16658 = 12'h4ce == _T_171[11:0] ? image_1230 : _GEN_16657; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16659 = 12'h4cf == _T_171[11:0] ? image_1231 : _GEN_16658; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16660 = 12'h4d0 == _T_171[11:0] ? image_1232 : _GEN_16659; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16661 = 12'h4d1 == _T_171[11:0] ? image_1233 : _GEN_16660; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16662 = 12'h4d2 == _T_171[11:0] ? image_1234 : _GEN_16661; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16663 = 12'h4d3 == _T_171[11:0] ? image_1235 : _GEN_16662; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16664 = 12'h4d4 == _T_171[11:0] ? image_1236 : _GEN_16663; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16665 = 12'h4d5 == _T_171[11:0] ? image_1237 : _GEN_16664; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16666 = 12'h4d6 == _T_171[11:0] ? image_1238 : _GEN_16665; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16667 = 12'h4d7 == _T_171[11:0] ? image_1239 : _GEN_16666; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16668 = 12'h4d8 == _T_171[11:0] ? image_1240 : _GEN_16667; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16669 = 12'h4d9 == _T_171[11:0] ? image_1241 : _GEN_16668; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16670 = 12'h4da == _T_171[11:0] ? image_1242 : _GEN_16669; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16671 = 12'h4db == _T_171[11:0] ? image_1243 : _GEN_16670; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16672 = 12'h4dc == _T_171[11:0] ? image_1244 : _GEN_16671; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16673 = 12'h4dd == _T_171[11:0] ? image_1245 : _GEN_16672; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16674 = 12'h4de == _T_171[11:0] ? image_1246 : _GEN_16673; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16675 = 12'h4df == _T_171[11:0] ? image_1247 : _GEN_16674; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16676 = 12'h4e0 == _T_171[11:0] ? image_1248 : _GEN_16675; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16677 = 12'h4e1 == _T_171[11:0] ? image_1249 : _GEN_16676; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16678 = 12'h4e2 == _T_171[11:0] ? image_1250 : _GEN_16677; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16679 = 12'h4e3 == _T_171[11:0] ? image_1251 : _GEN_16678; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16680 = 12'h4e4 == _T_171[11:0] ? image_1252 : _GEN_16679; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16681 = 12'h4e5 == _T_171[11:0] ? image_1253 : _GEN_16680; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16682 = 12'h4e6 == _T_171[11:0] ? image_1254 : _GEN_16681; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16683 = 12'h4e7 == _T_171[11:0] ? image_1255 : _GEN_16682; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16684 = 12'h4e8 == _T_171[11:0] ? image_1256 : _GEN_16683; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16685 = 12'h4e9 == _T_171[11:0] ? image_1257 : _GEN_16684; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16686 = 12'h4ea == _T_171[11:0] ? image_1258 : _GEN_16685; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16687 = 12'h4eb == _T_171[11:0] ? image_1259 : _GEN_16686; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16688 = 12'h4ec == _T_171[11:0] ? image_1260 : _GEN_16687; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16689 = 12'h4ed == _T_171[11:0] ? image_1261 : _GEN_16688; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16690 = 12'h4ee == _T_171[11:0] ? image_1262 : _GEN_16689; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16691 = 12'h4ef == _T_171[11:0] ? image_1263 : _GEN_16690; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16692 = 12'h4f0 == _T_171[11:0] ? image_1264 : _GEN_16691; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16693 = 12'h4f1 == _T_171[11:0] ? image_1265 : _GEN_16692; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16694 = 12'h4f2 == _T_171[11:0] ? image_1266 : _GEN_16693; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16695 = 12'h4f3 == _T_171[11:0] ? image_1267 : _GEN_16694; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16696 = 12'h4f4 == _T_171[11:0] ? image_1268 : _GEN_16695; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16697 = 12'h4f5 == _T_171[11:0] ? image_1269 : _GEN_16696; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16698 = 12'h4f6 == _T_171[11:0] ? image_1270 : _GEN_16697; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16699 = 12'h4f7 == _T_171[11:0] ? image_1271 : _GEN_16698; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16700 = 12'h4f8 == _T_171[11:0] ? image_1272 : _GEN_16699; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16701 = 12'h4f9 == _T_171[11:0] ? image_1273 : _GEN_16700; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16702 = 12'h4fa == _T_171[11:0] ? image_1274 : _GEN_16701; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16703 = 12'h4fb == _T_171[11:0] ? image_1275 : _GEN_16702; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16704 = 12'h4fc == _T_171[11:0] ? 4'h0 : _GEN_16703; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16705 = 12'h4fd == _T_171[11:0] ? 4'h0 : _GEN_16704; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16706 = 12'h4fe == _T_171[11:0] ? 4'h0 : _GEN_16705; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16707 = 12'h4ff == _T_171[11:0] ? 4'h0 : _GEN_16706; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16708 = 12'h500 == _T_171[11:0] ? image_1280 : _GEN_16707; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16709 = 12'h501 == _T_171[11:0] ? image_1281 : _GEN_16708; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16710 = 12'h502 == _T_171[11:0] ? image_1282 : _GEN_16709; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16711 = 12'h503 == _T_171[11:0] ? image_1283 : _GEN_16710; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16712 = 12'h504 == _T_171[11:0] ? image_1284 : _GEN_16711; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16713 = 12'h505 == _T_171[11:0] ? image_1285 : _GEN_16712; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16714 = 12'h506 == _T_171[11:0] ? image_1286 : _GEN_16713; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16715 = 12'h507 == _T_171[11:0] ? image_1287 : _GEN_16714; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16716 = 12'h508 == _T_171[11:0] ? image_1288 : _GEN_16715; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16717 = 12'h509 == _T_171[11:0] ? image_1289 : _GEN_16716; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16718 = 12'h50a == _T_171[11:0] ? image_1290 : _GEN_16717; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16719 = 12'h50b == _T_171[11:0] ? image_1291 : _GEN_16718; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16720 = 12'h50c == _T_171[11:0] ? image_1292 : _GEN_16719; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16721 = 12'h50d == _T_171[11:0] ? image_1293 : _GEN_16720; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16722 = 12'h50e == _T_171[11:0] ? image_1294 : _GEN_16721; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16723 = 12'h50f == _T_171[11:0] ? image_1295 : _GEN_16722; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16724 = 12'h510 == _T_171[11:0] ? image_1296 : _GEN_16723; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16725 = 12'h511 == _T_171[11:0] ? image_1297 : _GEN_16724; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16726 = 12'h512 == _T_171[11:0] ? image_1298 : _GEN_16725; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16727 = 12'h513 == _T_171[11:0] ? image_1299 : _GEN_16726; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16728 = 12'h514 == _T_171[11:0] ? image_1300 : _GEN_16727; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16729 = 12'h515 == _T_171[11:0] ? image_1301 : _GEN_16728; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16730 = 12'h516 == _T_171[11:0] ? image_1302 : _GEN_16729; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16731 = 12'h517 == _T_171[11:0] ? image_1303 : _GEN_16730; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16732 = 12'h518 == _T_171[11:0] ? image_1304 : _GEN_16731; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16733 = 12'h519 == _T_171[11:0] ? image_1305 : _GEN_16732; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16734 = 12'h51a == _T_171[11:0] ? image_1306 : _GEN_16733; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16735 = 12'h51b == _T_171[11:0] ? image_1307 : _GEN_16734; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16736 = 12'h51c == _T_171[11:0] ? image_1308 : _GEN_16735; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16737 = 12'h51d == _T_171[11:0] ? image_1309 : _GEN_16736; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16738 = 12'h51e == _T_171[11:0] ? image_1310 : _GEN_16737; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16739 = 12'h51f == _T_171[11:0] ? image_1311 : _GEN_16738; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16740 = 12'h520 == _T_171[11:0] ? image_1312 : _GEN_16739; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16741 = 12'h521 == _T_171[11:0] ? image_1313 : _GEN_16740; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16742 = 12'h522 == _T_171[11:0] ? image_1314 : _GEN_16741; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16743 = 12'h523 == _T_171[11:0] ? image_1315 : _GEN_16742; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16744 = 12'h524 == _T_171[11:0] ? image_1316 : _GEN_16743; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16745 = 12'h525 == _T_171[11:0] ? image_1317 : _GEN_16744; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16746 = 12'h526 == _T_171[11:0] ? image_1318 : _GEN_16745; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16747 = 12'h527 == _T_171[11:0] ? image_1319 : _GEN_16746; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16748 = 12'h528 == _T_171[11:0] ? image_1320 : _GEN_16747; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16749 = 12'h529 == _T_171[11:0] ? image_1321 : _GEN_16748; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16750 = 12'h52a == _T_171[11:0] ? image_1322 : _GEN_16749; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16751 = 12'h52b == _T_171[11:0] ? image_1323 : _GEN_16750; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16752 = 12'h52c == _T_171[11:0] ? image_1324 : _GEN_16751; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16753 = 12'h52d == _T_171[11:0] ? image_1325 : _GEN_16752; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16754 = 12'h52e == _T_171[11:0] ? image_1326 : _GEN_16753; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16755 = 12'h52f == _T_171[11:0] ? image_1327 : _GEN_16754; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16756 = 12'h530 == _T_171[11:0] ? image_1328 : _GEN_16755; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16757 = 12'h531 == _T_171[11:0] ? image_1329 : _GEN_16756; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16758 = 12'h532 == _T_171[11:0] ? image_1330 : _GEN_16757; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16759 = 12'h533 == _T_171[11:0] ? image_1331 : _GEN_16758; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16760 = 12'h534 == _T_171[11:0] ? image_1332 : _GEN_16759; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16761 = 12'h535 == _T_171[11:0] ? image_1333 : _GEN_16760; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16762 = 12'h536 == _T_171[11:0] ? image_1334 : _GEN_16761; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16763 = 12'h537 == _T_171[11:0] ? image_1335 : _GEN_16762; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16764 = 12'h538 == _T_171[11:0] ? image_1336 : _GEN_16763; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16765 = 12'h539 == _T_171[11:0] ? image_1337 : _GEN_16764; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16766 = 12'h53a == _T_171[11:0] ? image_1338 : _GEN_16765; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16767 = 12'h53b == _T_171[11:0] ? image_1339 : _GEN_16766; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16768 = 12'h53c == _T_171[11:0] ? image_1340 : _GEN_16767; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16769 = 12'h53d == _T_171[11:0] ? image_1341 : _GEN_16768; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16770 = 12'h53e == _T_171[11:0] ? 4'h0 : _GEN_16769; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16771 = 12'h53f == _T_171[11:0] ? 4'h0 : _GEN_16770; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16772 = 12'h540 == _T_171[11:0] ? image_1344 : _GEN_16771; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16773 = 12'h541 == _T_171[11:0] ? image_1345 : _GEN_16772; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16774 = 12'h542 == _T_171[11:0] ? image_1346 : _GEN_16773; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16775 = 12'h543 == _T_171[11:0] ? image_1347 : _GEN_16774; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16776 = 12'h544 == _T_171[11:0] ? image_1348 : _GEN_16775; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16777 = 12'h545 == _T_171[11:0] ? image_1349 : _GEN_16776; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16778 = 12'h546 == _T_171[11:0] ? image_1350 : _GEN_16777; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16779 = 12'h547 == _T_171[11:0] ? image_1351 : _GEN_16778; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16780 = 12'h548 == _T_171[11:0] ? image_1352 : _GEN_16779; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16781 = 12'h549 == _T_171[11:0] ? image_1353 : _GEN_16780; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16782 = 12'h54a == _T_171[11:0] ? image_1354 : _GEN_16781; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16783 = 12'h54b == _T_171[11:0] ? image_1355 : _GEN_16782; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16784 = 12'h54c == _T_171[11:0] ? image_1356 : _GEN_16783; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16785 = 12'h54d == _T_171[11:0] ? image_1357 : _GEN_16784; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16786 = 12'h54e == _T_171[11:0] ? image_1358 : _GEN_16785; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16787 = 12'h54f == _T_171[11:0] ? image_1359 : _GEN_16786; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16788 = 12'h550 == _T_171[11:0] ? image_1360 : _GEN_16787; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16789 = 12'h551 == _T_171[11:0] ? image_1361 : _GEN_16788; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16790 = 12'h552 == _T_171[11:0] ? image_1362 : _GEN_16789; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16791 = 12'h553 == _T_171[11:0] ? image_1363 : _GEN_16790; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16792 = 12'h554 == _T_171[11:0] ? image_1364 : _GEN_16791; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16793 = 12'h555 == _T_171[11:0] ? image_1365 : _GEN_16792; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16794 = 12'h556 == _T_171[11:0] ? image_1366 : _GEN_16793; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16795 = 12'h557 == _T_171[11:0] ? image_1367 : _GEN_16794; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16796 = 12'h558 == _T_171[11:0] ? image_1368 : _GEN_16795; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16797 = 12'h559 == _T_171[11:0] ? image_1369 : _GEN_16796; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16798 = 12'h55a == _T_171[11:0] ? image_1370 : _GEN_16797; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16799 = 12'h55b == _T_171[11:0] ? image_1371 : _GEN_16798; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16800 = 12'h55c == _T_171[11:0] ? image_1372 : _GEN_16799; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16801 = 12'h55d == _T_171[11:0] ? image_1373 : _GEN_16800; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16802 = 12'h55e == _T_171[11:0] ? image_1374 : _GEN_16801; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16803 = 12'h55f == _T_171[11:0] ? image_1375 : _GEN_16802; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16804 = 12'h560 == _T_171[11:0] ? image_1376 : _GEN_16803; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16805 = 12'h561 == _T_171[11:0] ? image_1377 : _GEN_16804; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16806 = 12'h562 == _T_171[11:0] ? image_1378 : _GEN_16805; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16807 = 12'h563 == _T_171[11:0] ? image_1379 : _GEN_16806; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16808 = 12'h564 == _T_171[11:0] ? image_1380 : _GEN_16807; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16809 = 12'h565 == _T_171[11:0] ? image_1381 : _GEN_16808; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16810 = 12'h566 == _T_171[11:0] ? image_1382 : _GEN_16809; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16811 = 12'h567 == _T_171[11:0] ? image_1383 : _GEN_16810; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16812 = 12'h568 == _T_171[11:0] ? image_1384 : _GEN_16811; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16813 = 12'h569 == _T_171[11:0] ? image_1385 : _GEN_16812; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16814 = 12'h56a == _T_171[11:0] ? image_1386 : _GEN_16813; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16815 = 12'h56b == _T_171[11:0] ? image_1387 : _GEN_16814; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16816 = 12'h56c == _T_171[11:0] ? image_1388 : _GEN_16815; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16817 = 12'h56d == _T_171[11:0] ? image_1389 : _GEN_16816; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16818 = 12'h56e == _T_171[11:0] ? image_1390 : _GEN_16817; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16819 = 12'h56f == _T_171[11:0] ? image_1391 : _GEN_16818; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16820 = 12'h570 == _T_171[11:0] ? image_1392 : _GEN_16819; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16821 = 12'h571 == _T_171[11:0] ? image_1393 : _GEN_16820; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16822 = 12'h572 == _T_171[11:0] ? image_1394 : _GEN_16821; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16823 = 12'h573 == _T_171[11:0] ? image_1395 : _GEN_16822; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16824 = 12'h574 == _T_171[11:0] ? image_1396 : _GEN_16823; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16825 = 12'h575 == _T_171[11:0] ? image_1397 : _GEN_16824; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16826 = 12'h576 == _T_171[11:0] ? image_1398 : _GEN_16825; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16827 = 12'h577 == _T_171[11:0] ? image_1399 : _GEN_16826; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16828 = 12'h578 == _T_171[11:0] ? image_1400 : _GEN_16827; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16829 = 12'h579 == _T_171[11:0] ? image_1401 : _GEN_16828; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16830 = 12'h57a == _T_171[11:0] ? image_1402 : _GEN_16829; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16831 = 12'h57b == _T_171[11:0] ? image_1403 : _GEN_16830; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16832 = 12'h57c == _T_171[11:0] ? image_1404 : _GEN_16831; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16833 = 12'h57d == _T_171[11:0] ? image_1405 : _GEN_16832; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16834 = 12'h57e == _T_171[11:0] ? 4'h0 : _GEN_16833; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16835 = 12'h57f == _T_171[11:0] ? 4'h0 : _GEN_16834; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16836 = 12'h580 == _T_171[11:0] ? image_1408 : _GEN_16835; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16837 = 12'h581 == _T_171[11:0] ? image_1409 : _GEN_16836; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16838 = 12'h582 == _T_171[11:0] ? image_1410 : _GEN_16837; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16839 = 12'h583 == _T_171[11:0] ? image_1411 : _GEN_16838; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16840 = 12'h584 == _T_171[11:0] ? image_1412 : _GEN_16839; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16841 = 12'h585 == _T_171[11:0] ? image_1413 : _GEN_16840; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16842 = 12'h586 == _T_171[11:0] ? image_1414 : _GEN_16841; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16843 = 12'h587 == _T_171[11:0] ? image_1415 : _GEN_16842; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16844 = 12'h588 == _T_171[11:0] ? image_1416 : _GEN_16843; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16845 = 12'h589 == _T_171[11:0] ? image_1417 : _GEN_16844; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16846 = 12'h58a == _T_171[11:0] ? image_1418 : _GEN_16845; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16847 = 12'h58b == _T_171[11:0] ? image_1419 : _GEN_16846; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16848 = 12'h58c == _T_171[11:0] ? image_1420 : _GEN_16847; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16849 = 12'h58d == _T_171[11:0] ? image_1421 : _GEN_16848; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16850 = 12'h58e == _T_171[11:0] ? image_1422 : _GEN_16849; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16851 = 12'h58f == _T_171[11:0] ? image_1423 : _GEN_16850; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16852 = 12'h590 == _T_171[11:0] ? image_1424 : _GEN_16851; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16853 = 12'h591 == _T_171[11:0] ? image_1425 : _GEN_16852; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16854 = 12'h592 == _T_171[11:0] ? image_1426 : _GEN_16853; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16855 = 12'h593 == _T_171[11:0] ? image_1427 : _GEN_16854; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16856 = 12'h594 == _T_171[11:0] ? image_1428 : _GEN_16855; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16857 = 12'h595 == _T_171[11:0] ? image_1429 : _GEN_16856; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16858 = 12'h596 == _T_171[11:0] ? image_1430 : _GEN_16857; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16859 = 12'h597 == _T_171[11:0] ? image_1431 : _GEN_16858; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16860 = 12'h598 == _T_171[11:0] ? image_1432 : _GEN_16859; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16861 = 12'h599 == _T_171[11:0] ? image_1433 : _GEN_16860; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16862 = 12'h59a == _T_171[11:0] ? image_1434 : _GEN_16861; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16863 = 12'h59b == _T_171[11:0] ? image_1435 : _GEN_16862; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16864 = 12'h59c == _T_171[11:0] ? image_1436 : _GEN_16863; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16865 = 12'h59d == _T_171[11:0] ? image_1437 : _GEN_16864; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16866 = 12'h59e == _T_171[11:0] ? image_1438 : _GEN_16865; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16867 = 12'h59f == _T_171[11:0] ? image_1439 : _GEN_16866; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16868 = 12'h5a0 == _T_171[11:0] ? image_1440 : _GEN_16867; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16869 = 12'h5a1 == _T_171[11:0] ? image_1441 : _GEN_16868; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16870 = 12'h5a2 == _T_171[11:0] ? image_1442 : _GEN_16869; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16871 = 12'h5a3 == _T_171[11:0] ? image_1443 : _GEN_16870; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16872 = 12'h5a4 == _T_171[11:0] ? image_1444 : _GEN_16871; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16873 = 12'h5a5 == _T_171[11:0] ? image_1445 : _GEN_16872; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16874 = 12'h5a6 == _T_171[11:0] ? image_1446 : _GEN_16873; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16875 = 12'h5a7 == _T_171[11:0] ? image_1447 : _GEN_16874; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16876 = 12'h5a8 == _T_171[11:0] ? image_1448 : _GEN_16875; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16877 = 12'h5a9 == _T_171[11:0] ? image_1449 : _GEN_16876; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16878 = 12'h5aa == _T_171[11:0] ? image_1450 : _GEN_16877; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16879 = 12'h5ab == _T_171[11:0] ? image_1451 : _GEN_16878; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16880 = 12'h5ac == _T_171[11:0] ? image_1452 : _GEN_16879; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16881 = 12'h5ad == _T_171[11:0] ? image_1453 : _GEN_16880; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16882 = 12'h5ae == _T_171[11:0] ? image_1454 : _GEN_16881; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16883 = 12'h5af == _T_171[11:0] ? image_1455 : _GEN_16882; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16884 = 12'h5b0 == _T_171[11:0] ? image_1456 : _GEN_16883; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16885 = 12'h5b1 == _T_171[11:0] ? image_1457 : _GEN_16884; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16886 = 12'h5b2 == _T_171[11:0] ? image_1458 : _GEN_16885; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16887 = 12'h5b3 == _T_171[11:0] ? image_1459 : _GEN_16886; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16888 = 12'h5b4 == _T_171[11:0] ? image_1460 : _GEN_16887; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16889 = 12'h5b5 == _T_171[11:0] ? image_1461 : _GEN_16888; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16890 = 12'h5b6 == _T_171[11:0] ? image_1462 : _GEN_16889; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16891 = 12'h5b7 == _T_171[11:0] ? image_1463 : _GEN_16890; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16892 = 12'h5b8 == _T_171[11:0] ? image_1464 : _GEN_16891; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16893 = 12'h5b9 == _T_171[11:0] ? image_1465 : _GEN_16892; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16894 = 12'h5ba == _T_171[11:0] ? image_1466 : _GEN_16893; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16895 = 12'h5bb == _T_171[11:0] ? image_1467 : _GEN_16894; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16896 = 12'h5bc == _T_171[11:0] ? image_1468 : _GEN_16895; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16897 = 12'h5bd == _T_171[11:0] ? image_1469 : _GEN_16896; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16898 = 12'h5be == _T_171[11:0] ? 4'h0 : _GEN_16897; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16899 = 12'h5bf == _T_171[11:0] ? 4'h0 : _GEN_16898; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16900 = 12'h5c0 == _T_171[11:0] ? image_1472 : _GEN_16899; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16901 = 12'h5c1 == _T_171[11:0] ? image_1473 : _GEN_16900; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16902 = 12'h5c2 == _T_171[11:0] ? image_1474 : _GEN_16901; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16903 = 12'h5c3 == _T_171[11:0] ? image_1475 : _GEN_16902; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16904 = 12'h5c4 == _T_171[11:0] ? image_1476 : _GEN_16903; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16905 = 12'h5c5 == _T_171[11:0] ? image_1477 : _GEN_16904; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16906 = 12'h5c6 == _T_171[11:0] ? image_1478 : _GEN_16905; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16907 = 12'h5c7 == _T_171[11:0] ? image_1479 : _GEN_16906; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16908 = 12'h5c8 == _T_171[11:0] ? image_1480 : _GEN_16907; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16909 = 12'h5c9 == _T_171[11:0] ? image_1481 : _GEN_16908; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16910 = 12'h5ca == _T_171[11:0] ? image_1482 : _GEN_16909; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16911 = 12'h5cb == _T_171[11:0] ? image_1483 : _GEN_16910; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16912 = 12'h5cc == _T_171[11:0] ? image_1484 : _GEN_16911; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16913 = 12'h5cd == _T_171[11:0] ? image_1485 : _GEN_16912; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16914 = 12'h5ce == _T_171[11:0] ? image_1486 : _GEN_16913; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16915 = 12'h5cf == _T_171[11:0] ? image_1487 : _GEN_16914; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16916 = 12'h5d0 == _T_171[11:0] ? image_1488 : _GEN_16915; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16917 = 12'h5d1 == _T_171[11:0] ? image_1489 : _GEN_16916; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16918 = 12'h5d2 == _T_171[11:0] ? image_1490 : _GEN_16917; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16919 = 12'h5d3 == _T_171[11:0] ? image_1491 : _GEN_16918; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16920 = 12'h5d4 == _T_171[11:0] ? image_1492 : _GEN_16919; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16921 = 12'h5d5 == _T_171[11:0] ? image_1493 : _GEN_16920; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16922 = 12'h5d6 == _T_171[11:0] ? image_1494 : _GEN_16921; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16923 = 12'h5d7 == _T_171[11:0] ? image_1495 : _GEN_16922; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16924 = 12'h5d8 == _T_171[11:0] ? image_1496 : _GEN_16923; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16925 = 12'h5d9 == _T_171[11:0] ? image_1497 : _GEN_16924; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16926 = 12'h5da == _T_171[11:0] ? image_1498 : _GEN_16925; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16927 = 12'h5db == _T_171[11:0] ? image_1499 : _GEN_16926; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16928 = 12'h5dc == _T_171[11:0] ? image_1500 : _GEN_16927; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16929 = 12'h5dd == _T_171[11:0] ? image_1501 : _GEN_16928; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16930 = 12'h5de == _T_171[11:0] ? image_1502 : _GEN_16929; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16931 = 12'h5df == _T_171[11:0] ? image_1503 : _GEN_16930; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16932 = 12'h5e0 == _T_171[11:0] ? image_1504 : _GEN_16931; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16933 = 12'h5e1 == _T_171[11:0] ? image_1505 : _GEN_16932; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16934 = 12'h5e2 == _T_171[11:0] ? image_1506 : _GEN_16933; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16935 = 12'h5e3 == _T_171[11:0] ? image_1507 : _GEN_16934; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16936 = 12'h5e4 == _T_171[11:0] ? image_1508 : _GEN_16935; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16937 = 12'h5e5 == _T_171[11:0] ? image_1509 : _GEN_16936; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16938 = 12'h5e6 == _T_171[11:0] ? image_1510 : _GEN_16937; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16939 = 12'h5e7 == _T_171[11:0] ? image_1511 : _GEN_16938; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16940 = 12'h5e8 == _T_171[11:0] ? image_1512 : _GEN_16939; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16941 = 12'h5e9 == _T_171[11:0] ? image_1513 : _GEN_16940; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16942 = 12'h5ea == _T_171[11:0] ? image_1514 : _GEN_16941; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16943 = 12'h5eb == _T_171[11:0] ? image_1515 : _GEN_16942; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16944 = 12'h5ec == _T_171[11:0] ? image_1516 : _GEN_16943; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16945 = 12'h5ed == _T_171[11:0] ? image_1517 : _GEN_16944; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16946 = 12'h5ee == _T_171[11:0] ? image_1518 : _GEN_16945; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16947 = 12'h5ef == _T_171[11:0] ? image_1519 : _GEN_16946; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16948 = 12'h5f0 == _T_171[11:0] ? image_1520 : _GEN_16947; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16949 = 12'h5f1 == _T_171[11:0] ? image_1521 : _GEN_16948; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16950 = 12'h5f2 == _T_171[11:0] ? image_1522 : _GEN_16949; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16951 = 12'h5f3 == _T_171[11:0] ? image_1523 : _GEN_16950; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16952 = 12'h5f4 == _T_171[11:0] ? image_1524 : _GEN_16951; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16953 = 12'h5f5 == _T_171[11:0] ? image_1525 : _GEN_16952; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16954 = 12'h5f6 == _T_171[11:0] ? image_1526 : _GEN_16953; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16955 = 12'h5f7 == _T_171[11:0] ? image_1527 : _GEN_16954; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16956 = 12'h5f8 == _T_171[11:0] ? image_1528 : _GEN_16955; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16957 = 12'h5f9 == _T_171[11:0] ? image_1529 : _GEN_16956; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16958 = 12'h5fa == _T_171[11:0] ? image_1530 : _GEN_16957; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16959 = 12'h5fb == _T_171[11:0] ? image_1531 : _GEN_16958; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16960 = 12'h5fc == _T_171[11:0] ? image_1532 : _GEN_16959; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16961 = 12'h5fd == _T_171[11:0] ? image_1533 : _GEN_16960; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16962 = 12'h5fe == _T_171[11:0] ? 4'h0 : _GEN_16961; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16963 = 12'h5ff == _T_171[11:0] ? 4'h0 : _GEN_16962; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16964 = 12'h600 == _T_171[11:0] ? image_1536 : _GEN_16963; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16965 = 12'h601 == _T_171[11:0] ? image_1537 : _GEN_16964; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16966 = 12'h602 == _T_171[11:0] ? image_1538 : _GEN_16965; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16967 = 12'h603 == _T_171[11:0] ? image_1539 : _GEN_16966; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16968 = 12'h604 == _T_171[11:0] ? image_1540 : _GEN_16967; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16969 = 12'h605 == _T_171[11:0] ? image_1541 : _GEN_16968; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16970 = 12'h606 == _T_171[11:0] ? image_1542 : _GEN_16969; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16971 = 12'h607 == _T_171[11:0] ? image_1543 : _GEN_16970; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16972 = 12'h608 == _T_171[11:0] ? image_1544 : _GEN_16971; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16973 = 12'h609 == _T_171[11:0] ? image_1545 : _GEN_16972; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16974 = 12'h60a == _T_171[11:0] ? image_1546 : _GEN_16973; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16975 = 12'h60b == _T_171[11:0] ? image_1547 : _GEN_16974; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16976 = 12'h60c == _T_171[11:0] ? image_1548 : _GEN_16975; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16977 = 12'h60d == _T_171[11:0] ? image_1549 : _GEN_16976; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16978 = 12'h60e == _T_171[11:0] ? image_1550 : _GEN_16977; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16979 = 12'h60f == _T_171[11:0] ? image_1551 : _GEN_16978; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16980 = 12'h610 == _T_171[11:0] ? image_1552 : _GEN_16979; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16981 = 12'h611 == _T_171[11:0] ? image_1553 : _GEN_16980; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16982 = 12'h612 == _T_171[11:0] ? image_1554 : _GEN_16981; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16983 = 12'h613 == _T_171[11:0] ? image_1555 : _GEN_16982; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16984 = 12'h614 == _T_171[11:0] ? image_1556 : _GEN_16983; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16985 = 12'h615 == _T_171[11:0] ? image_1557 : _GEN_16984; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16986 = 12'h616 == _T_171[11:0] ? image_1558 : _GEN_16985; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16987 = 12'h617 == _T_171[11:0] ? image_1559 : _GEN_16986; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16988 = 12'h618 == _T_171[11:0] ? image_1560 : _GEN_16987; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16989 = 12'h619 == _T_171[11:0] ? image_1561 : _GEN_16988; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16990 = 12'h61a == _T_171[11:0] ? image_1562 : _GEN_16989; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16991 = 12'h61b == _T_171[11:0] ? image_1563 : _GEN_16990; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16992 = 12'h61c == _T_171[11:0] ? image_1564 : _GEN_16991; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16993 = 12'h61d == _T_171[11:0] ? image_1565 : _GEN_16992; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16994 = 12'h61e == _T_171[11:0] ? image_1566 : _GEN_16993; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16995 = 12'h61f == _T_171[11:0] ? image_1567 : _GEN_16994; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16996 = 12'h620 == _T_171[11:0] ? image_1568 : _GEN_16995; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16997 = 12'h621 == _T_171[11:0] ? image_1569 : _GEN_16996; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16998 = 12'h622 == _T_171[11:0] ? image_1570 : _GEN_16997; // @[Filter.scala 138:46]
  wire [3:0] _GEN_16999 = 12'h623 == _T_171[11:0] ? image_1571 : _GEN_16998; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17000 = 12'h624 == _T_171[11:0] ? image_1572 : _GEN_16999; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17001 = 12'h625 == _T_171[11:0] ? image_1573 : _GEN_17000; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17002 = 12'h626 == _T_171[11:0] ? image_1574 : _GEN_17001; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17003 = 12'h627 == _T_171[11:0] ? image_1575 : _GEN_17002; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17004 = 12'h628 == _T_171[11:0] ? image_1576 : _GEN_17003; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17005 = 12'h629 == _T_171[11:0] ? image_1577 : _GEN_17004; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17006 = 12'h62a == _T_171[11:0] ? image_1578 : _GEN_17005; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17007 = 12'h62b == _T_171[11:0] ? image_1579 : _GEN_17006; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17008 = 12'h62c == _T_171[11:0] ? image_1580 : _GEN_17007; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17009 = 12'h62d == _T_171[11:0] ? image_1581 : _GEN_17008; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17010 = 12'h62e == _T_171[11:0] ? image_1582 : _GEN_17009; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17011 = 12'h62f == _T_171[11:0] ? image_1583 : _GEN_17010; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17012 = 12'h630 == _T_171[11:0] ? image_1584 : _GEN_17011; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17013 = 12'h631 == _T_171[11:0] ? image_1585 : _GEN_17012; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17014 = 12'h632 == _T_171[11:0] ? image_1586 : _GEN_17013; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17015 = 12'h633 == _T_171[11:0] ? image_1587 : _GEN_17014; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17016 = 12'h634 == _T_171[11:0] ? image_1588 : _GEN_17015; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17017 = 12'h635 == _T_171[11:0] ? image_1589 : _GEN_17016; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17018 = 12'h636 == _T_171[11:0] ? image_1590 : _GEN_17017; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17019 = 12'h637 == _T_171[11:0] ? image_1591 : _GEN_17018; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17020 = 12'h638 == _T_171[11:0] ? image_1592 : _GEN_17019; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17021 = 12'h639 == _T_171[11:0] ? image_1593 : _GEN_17020; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17022 = 12'h63a == _T_171[11:0] ? image_1594 : _GEN_17021; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17023 = 12'h63b == _T_171[11:0] ? image_1595 : _GEN_17022; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17024 = 12'h63c == _T_171[11:0] ? image_1596 : _GEN_17023; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17025 = 12'h63d == _T_171[11:0] ? image_1597 : _GEN_17024; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17026 = 12'h63e == _T_171[11:0] ? 4'h0 : _GEN_17025; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17027 = 12'h63f == _T_171[11:0] ? 4'h0 : _GEN_17026; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17028 = 12'h640 == _T_171[11:0] ? image_1600 : _GEN_17027; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17029 = 12'h641 == _T_171[11:0] ? image_1601 : _GEN_17028; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17030 = 12'h642 == _T_171[11:0] ? image_1602 : _GEN_17029; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17031 = 12'h643 == _T_171[11:0] ? image_1603 : _GEN_17030; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17032 = 12'h644 == _T_171[11:0] ? image_1604 : _GEN_17031; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17033 = 12'h645 == _T_171[11:0] ? image_1605 : _GEN_17032; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17034 = 12'h646 == _T_171[11:0] ? image_1606 : _GEN_17033; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17035 = 12'h647 == _T_171[11:0] ? image_1607 : _GEN_17034; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17036 = 12'h648 == _T_171[11:0] ? image_1608 : _GEN_17035; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17037 = 12'h649 == _T_171[11:0] ? image_1609 : _GEN_17036; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17038 = 12'h64a == _T_171[11:0] ? image_1610 : _GEN_17037; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17039 = 12'h64b == _T_171[11:0] ? image_1611 : _GEN_17038; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17040 = 12'h64c == _T_171[11:0] ? image_1612 : _GEN_17039; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17041 = 12'h64d == _T_171[11:0] ? image_1613 : _GEN_17040; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17042 = 12'h64e == _T_171[11:0] ? image_1614 : _GEN_17041; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17043 = 12'h64f == _T_171[11:0] ? image_1615 : _GEN_17042; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17044 = 12'h650 == _T_171[11:0] ? image_1616 : _GEN_17043; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17045 = 12'h651 == _T_171[11:0] ? image_1617 : _GEN_17044; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17046 = 12'h652 == _T_171[11:0] ? image_1618 : _GEN_17045; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17047 = 12'h653 == _T_171[11:0] ? image_1619 : _GEN_17046; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17048 = 12'h654 == _T_171[11:0] ? image_1620 : _GEN_17047; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17049 = 12'h655 == _T_171[11:0] ? image_1621 : _GEN_17048; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17050 = 12'h656 == _T_171[11:0] ? image_1622 : _GEN_17049; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17051 = 12'h657 == _T_171[11:0] ? image_1623 : _GEN_17050; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17052 = 12'h658 == _T_171[11:0] ? image_1624 : _GEN_17051; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17053 = 12'h659 == _T_171[11:0] ? image_1625 : _GEN_17052; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17054 = 12'h65a == _T_171[11:0] ? image_1626 : _GEN_17053; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17055 = 12'h65b == _T_171[11:0] ? image_1627 : _GEN_17054; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17056 = 12'h65c == _T_171[11:0] ? image_1628 : _GEN_17055; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17057 = 12'h65d == _T_171[11:0] ? image_1629 : _GEN_17056; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17058 = 12'h65e == _T_171[11:0] ? image_1630 : _GEN_17057; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17059 = 12'h65f == _T_171[11:0] ? image_1631 : _GEN_17058; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17060 = 12'h660 == _T_171[11:0] ? image_1632 : _GEN_17059; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17061 = 12'h661 == _T_171[11:0] ? image_1633 : _GEN_17060; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17062 = 12'h662 == _T_171[11:0] ? image_1634 : _GEN_17061; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17063 = 12'h663 == _T_171[11:0] ? image_1635 : _GEN_17062; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17064 = 12'h664 == _T_171[11:0] ? image_1636 : _GEN_17063; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17065 = 12'h665 == _T_171[11:0] ? image_1637 : _GEN_17064; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17066 = 12'h666 == _T_171[11:0] ? image_1638 : _GEN_17065; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17067 = 12'h667 == _T_171[11:0] ? image_1639 : _GEN_17066; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17068 = 12'h668 == _T_171[11:0] ? image_1640 : _GEN_17067; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17069 = 12'h669 == _T_171[11:0] ? image_1641 : _GEN_17068; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17070 = 12'h66a == _T_171[11:0] ? image_1642 : _GEN_17069; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17071 = 12'h66b == _T_171[11:0] ? image_1643 : _GEN_17070; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17072 = 12'h66c == _T_171[11:0] ? image_1644 : _GEN_17071; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17073 = 12'h66d == _T_171[11:0] ? image_1645 : _GEN_17072; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17074 = 12'h66e == _T_171[11:0] ? image_1646 : _GEN_17073; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17075 = 12'h66f == _T_171[11:0] ? image_1647 : _GEN_17074; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17076 = 12'h670 == _T_171[11:0] ? image_1648 : _GEN_17075; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17077 = 12'h671 == _T_171[11:0] ? image_1649 : _GEN_17076; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17078 = 12'h672 == _T_171[11:0] ? image_1650 : _GEN_17077; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17079 = 12'h673 == _T_171[11:0] ? image_1651 : _GEN_17078; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17080 = 12'h674 == _T_171[11:0] ? image_1652 : _GEN_17079; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17081 = 12'h675 == _T_171[11:0] ? image_1653 : _GEN_17080; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17082 = 12'h676 == _T_171[11:0] ? image_1654 : _GEN_17081; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17083 = 12'h677 == _T_171[11:0] ? image_1655 : _GEN_17082; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17084 = 12'h678 == _T_171[11:0] ? image_1656 : _GEN_17083; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17085 = 12'h679 == _T_171[11:0] ? image_1657 : _GEN_17084; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17086 = 12'h67a == _T_171[11:0] ? image_1658 : _GEN_17085; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17087 = 12'h67b == _T_171[11:0] ? image_1659 : _GEN_17086; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17088 = 12'h67c == _T_171[11:0] ? image_1660 : _GEN_17087; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17089 = 12'h67d == _T_171[11:0] ? 4'h0 : _GEN_17088; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17090 = 12'h67e == _T_171[11:0] ? 4'h0 : _GEN_17089; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17091 = 12'h67f == _T_171[11:0] ? 4'h0 : _GEN_17090; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17092 = 12'h680 == _T_171[11:0] ? image_1664 : _GEN_17091; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17093 = 12'h681 == _T_171[11:0] ? image_1665 : _GEN_17092; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17094 = 12'h682 == _T_171[11:0] ? image_1666 : _GEN_17093; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17095 = 12'h683 == _T_171[11:0] ? image_1667 : _GEN_17094; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17096 = 12'h684 == _T_171[11:0] ? image_1668 : _GEN_17095; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17097 = 12'h685 == _T_171[11:0] ? image_1669 : _GEN_17096; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17098 = 12'h686 == _T_171[11:0] ? image_1670 : _GEN_17097; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17099 = 12'h687 == _T_171[11:0] ? image_1671 : _GEN_17098; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17100 = 12'h688 == _T_171[11:0] ? image_1672 : _GEN_17099; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17101 = 12'h689 == _T_171[11:0] ? image_1673 : _GEN_17100; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17102 = 12'h68a == _T_171[11:0] ? image_1674 : _GEN_17101; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17103 = 12'h68b == _T_171[11:0] ? image_1675 : _GEN_17102; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17104 = 12'h68c == _T_171[11:0] ? image_1676 : _GEN_17103; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17105 = 12'h68d == _T_171[11:0] ? image_1677 : _GEN_17104; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17106 = 12'h68e == _T_171[11:0] ? image_1678 : _GEN_17105; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17107 = 12'h68f == _T_171[11:0] ? image_1679 : _GEN_17106; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17108 = 12'h690 == _T_171[11:0] ? image_1680 : _GEN_17107; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17109 = 12'h691 == _T_171[11:0] ? image_1681 : _GEN_17108; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17110 = 12'h692 == _T_171[11:0] ? image_1682 : _GEN_17109; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17111 = 12'h693 == _T_171[11:0] ? image_1683 : _GEN_17110; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17112 = 12'h694 == _T_171[11:0] ? image_1684 : _GEN_17111; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17113 = 12'h695 == _T_171[11:0] ? image_1685 : _GEN_17112; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17114 = 12'h696 == _T_171[11:0] ? image_1686 : _GEN_17113; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17115 = 12'h697 == _T_171[11:0] ? image_1687 : _GEN_17114; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17116 = 12'h698 == _T_171[11:0] ? image_1688 : _GEN_17115; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17117 = 12'h699 == _T_171[11:0] ? image_1689 : _GEN_17116; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17118 = 12'h69a == _T_171[11:0] ? image_1690 : _GEN_17117; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17119 = 12'h69b == _T_171[11:0] ? image_1691 : _GEN_17118; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17120 = 12'h69c == _T_171[11:0] ? image_1692 : _GEN_17119; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17121 = 12'h69d == _T_171[11:0] ? image_1693 : _GEN_17120; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17122 = 12'h69e == _T_171[11:0] ? image_1694 : _GEN_17121; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17123 = 12'h69f == _T_171[11:0] ? image_1695 : _GEN_17122; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17124 = 12'h6a0 == _T_171[11:0] ? image_1696 : _GEN_17123; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17125 = 12'h6a1 == _T_171[11:0] ? image_1697 : _GEN_17124; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17126 = 12'h6a2 == _T_171[11:0] ? image_1698 : _GEN_17125; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17127 = 12'h6a3 == _T_171[11:0] ? image_1699 : _GEN_17126; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17128 = 12'h6a4 == _T_171[11:0] ? image_1700 : _GEN_17127; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17129 = 12'h6a5 == _T_171[11:0] ? image_1701 : _GEN_17128; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17130 = 12'h6a6 == _T_171[11:0] ? image_1702 : _GEN_17129; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17131 = 12'h6a7 == _T_171[11:0] ? image_1703 : _GEN_17130; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17132 = 12'h6a8 == _T_171[11:0] ? image_1704 : _GEN_17131; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17133 = 12'h6a9 == _T_171[11:0] ? image_1705 : _GEN_17132; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17134 = 12'h6aa == _T_171[11:0] ? image_1706 : _GEN_17133; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17135 = 12'h6ab == _T_171[11:0] ? image_1707 : _GEN_17134; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17136 = 12'h6ac == _T_171[11:0] ? image_1708 : _GEN_17135; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17137 = 12'h6ad == _T_171[11:0] ? image_1709 : _GEN_17136; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17138 = 12'h6ae == _T_171[11:0] ? image_1710 : _GEN_17137; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17139 = 12'h6af == _T_171[11:0] ? image_1711 : _GEN_17138; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17140 = 12'h6b0 == _T_171[11:0] ? image_1712 : _GEN_17139; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17141 = 12'h6b1 == _T_171[11:0] ? image_1713 : _GEN_17140; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17142 = 12'h6b2 == _T_171[11:0] ? image_1714 : _GEN_17141; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17143 = 12'h6b3 == _T_171[11:0] ? image_1715 : _GEN_17142; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17144 = 12'h6b4 == _T_171[11:0] ? image_1716 : _GEN_17143; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17145 = 12'h6b5 == _T_171[11:0] ? image_1717 : _GEN_17144; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17146 = 12'h6b6 == _T_171[11:0] ? image_1718 : _GEN_17145; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17147 = 12'h6b7 == _T_171[11:0] ? image_1719 : _GEN_17146; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17148 = 12'h6b8 == _T_171[11:0] ? image_1720 : _GEN_17147; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17149 = 12'h6b9 == _T_171[11:0] ? image_1721 : _GEN_17148; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17150 = 12'h6ba == _T_171[11:0] ? image_1722 : _GEN_17149; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17151 = 12'h6bb == _T_171[11:0] ? image_1723 : _GEN_17150; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17152 = 12'h6bc == _T_171[11:0] ? 4'h0 : _GEN_17151; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17153 = 12'h6bd == _T_171[11:0] ? 4'h0 : _GEN_17152; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17154 = 12'h6be == _T_171[11:0] ? 4'h0 : _GEN_17153; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17155 = 12'h6bf == _T_171[11:0] ? 4'h0 : _GEN_17154; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17156 = 12'h6c0 == _T_171[11:0] ? image_1728 : _GEN_17155; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17157 = 12'h6c1 == _T_171[11:0] ? image_1729 : _GEN_17156; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17158 = 12'h6c2 == _T_171[11:0] ? image_1730 : _GEN_17157; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17159 = 12'h6c3 == _T_171[11:0] ? image_1731 : _GEN_17158; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17160 = 12'h6c4 == _T_171[11:0] ? image_1732 : _GEN_17159; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17161 = 12'h6c5 == _T_171[11:0] ? image_1733 : _GEN_17160; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17162 = 12'h6c6 == _T_171[11:0] ? image_1734 : _GEN_17161; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17163 = 12'h6c7 == _T_171[11:0] ? image_1735 : _GEN_17162; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17164 = 12'h6c8 == _T_171[11:0] ? image_1736 : _GEN_17163; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17165 = 12'h6c9 == _T_171[11:0] ? image_1737 : _GEN_17164; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17166 = 12'h6ca == _T_171[11:0] ? image_1738 : _GEN_17165; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17167 = 12'h6cb == _T_171[11:0] ? image_1739 : _GEN_17166; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17168 = 12'h6cc == _T_171[11:0] ? image_1740 : _GEN_17167; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17169 = 12'h6cd == _T_171[11:0] ? image_1741 : _GEN_17168; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17170 = 12'h6ce == _T_171[11:0] ? image_1742 : _GEN_17169; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17171 = 12'h6cf == _T_171[11:0] ? image_1743 : _GEN_17170; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17172 = 12'h6d0 == _T_171[11:0] ? image_1744 : _GEN_17171; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17173 = 12'h6d1 == _T_171[11:0] ? image_1745 : _GEN_17172; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17174 = 12'h6d2 == _T_171[11:0] ? image_1746 : _GEN_17173; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17175 = 12'h6d3 == _T_171[11:0] ? image_1747 : _GEN_17174; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17176 = 12'h6d4 == _T_171[11:0] ? image_1748 : _GEN_17175; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17177 = 12'h6d5 == _T_171[11:0] ? image_1749 : _GEN_17176; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17178 = 12'h6d6 == _T_171[11:0] ? image_1750 : _GEN_17177; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17179 = 12'h6d7 == _T_171[11:0] ? image_1751 : _GEN_17178; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17180 = 12'h6d8 == _T_171[11:0] ? image_1752 : _GEN_17179; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17181 = 12'h6d9 == _T_171[11:0] ? image_1753 : _GEN_17180; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17182 = 12'h6da == _T_171[11:0] ? image_1754 : _GEN_17181; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17183 = 12'h6db == _T_171[11:0] ? image_1755 : _GEN_17182; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17184 = 12'h6dc == _T_171[11:0] ? image_1756 : _GEN_17183; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17185 = 12'h6dd == _T_171[11:0] ? image_1757 : _GEN_17184; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17186 = 12'h6de == _T_171[11:0] ? image_1758 : _GEN_17185; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17187 = 12'h6df == _T_171[11:0] ? image_1759 : _GEN_17186; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17188 = 12'h6e0 == _T_171[11:0] ? image_1760 : _GEN_17187; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17189 = 12'h6e1 == _T_171[11:0] ? image_1761 : _GEN_17188; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17190 = 12'h6e2 == _T_171[11:0] ? image_1762 : _GEN_17189; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17191 = 12'h6e3 == _T_171[11:0] ? image_1763 : _GEN_17190; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17192 = 12'h6e4 == _T_171[11:0] ? image_1764 : _GEN_17191; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17193 = 12'h6e5 == _T_171[11:0] ? image_1765 : _GEN_17192; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17194 = 12'h6e6 == _T_171[11:0] ? image_1766 : _GEN_17193; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17195 = 12'h6e7 == _T_171[11:0] ? image_1767 : _GEN_17194; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17196 = 12'h6e8 == _T_171[11:0] ? image_1768 : _GEN_17195; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17197 = 12'h6e9 == _T_171[11:0] ? image_1769 : _GEN_17196; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17198 = 12'h6ea == _T_171[11:0] ? image_1770 : _GEN_17197; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17199 = 12'h6eb == _T_171[11:0] ? image_1771 : _GEN_17198; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17200 = 12'h6ec == _T_171[11:0] ? image_1772 : _GEN_17199; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17201 = 12'h6ed == _T_171[11:0] ? image_1773 : _GEN_17200; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17202 = 12'h6ee == _T_171[11:0] ? image_1774 : _GEN_17201; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17203 = 12'h6ef == _T_171[11:0] ? image_1775 : _GEN_17202; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17204 = 12'h6f0 == _T_171[11:0] ? image_1776 : _GEN_17203; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17205 = 12'h6f1 == _T_171[11:0] ? image_1777 : _GEN_17204; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17206 = 12'h6f2 == _T_171[11:0] ? image_1778 : _GEN_17205; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17207 = 12'h6f3 == _T_171[11:0] ? image_1779 : _GEN_17206; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17208 = 12'h6f4 == _T_171[11:0] ? image_1780 : _GEN_17207; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17209 = 12'h6f5 == _T_171[11:0] ? image_1781 : _GEN_17208; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17210 = 12'h6f6 == _T_171[11:0] ? image_1782 : _GEN_17209; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17211 = 12'h6f7 == _T_171[11:0] ? image_1783 : _GEN_17210; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17212 = 12'h6f8 == _T_171[11:0] ? image_1784 : _GEN_17211; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17213 = 12'h6f9 == _T_171[11:0] ? image_1785 : _GEN_17212; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17214 = 12'h6fa == _T_171[11:0] ? image_1786 : _GEN_17213; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17215 = 12'h6fb == _T_171[11:0] ? 4'h0 : _GEN_17214; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17216 = 12'h6fc == _T_171[11:0] ? 4'h0 : _GEN_17215; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17217 = 12'h6fd == _T_171[11:0] ? 4'h0 : _GEN_17216; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17218 = 12'h6fe == _T_171[11:0] ? 4'h0 : _GEN_17217; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17219 = 12'h6ff == _T_171[11:0] ? 4'h0 : _GEN_17218; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17220 = 12'h700 == _T_171[11:0] ? 4'h0 : _GEN_17219; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17221 = 12'h701 == _T_171[11:0] ? image_1793 : _GEN_17220; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17222 = 12'h702 == _T_171[11:0] ? image_1794 : _GEN_17221; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17223 = 12'h703 == _T_171[11:0] ? image_1795 : _GEN_17222; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17224 = 12'h704 == _T_171[11:0] ? image_1796 : _GEN_17223; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17225 = 12'h705 == _T_171[11:0] ? image_1797 : _GEN_17224; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17226 = 12'h706 == _T_171[11:0] ? image_1798 : _GEN_17225; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17227 = 12'h707 == _T_171[11:0] ? image_1799 : _GEN_17226; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17228 = 12'h708 == _T_171[11:0] ? image_1800 : _GEN_17227; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17229 = 12'h709 == _T_171[11:0] ? image_1801 : _GEN_17228; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17230 = 12'h70a == _T_171[11:0] ? image_1802 : _GEN_17229; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17231 = 12'h70b == _T_171[11:0] ? image_1803 : _GEN_17230; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17232 = 12'h70c == _T_171[11:0] ? image_1804 : _GEN_17231; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17233 = 12'h70d == _T_171[11:0] ? image_1805 : _GEN_17232; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17234 = 12'h70e == _T_171[11:0] ? image_1806 : _GEN_17233; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17235 = 12'h70f == _T_171[11:0] ? image_1807 : _GEN_17234; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17236 = 12'h710 == _T_171[11:0] ? image_1808 : _GEN_17235; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17237 = 12'h711 == _T_171[11:0] ? image_1809 : _GEN_17236; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17238 = 12'h712 == _T_171[11:0] ? image_1810 : _GEN_17237; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17239 = 12'h713 == _T_171[11:0] ? image_1811 : _GEN_17238; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17240 = 12'h714 == _T_171[11:0] ? image_1812 : _GEN_17239; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17241 = 12'h715 == _T_171[11:0] ? image_1813 : _GEN_17240; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17242 = 12'h716 == _T_171[11:0] ? image_1814 : _GEN_17241; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17243 = 12'h717 == _T_171[11:0] ? image_1815 : _GEN_17242; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17244 = 12'h718 == _T_171[11:0] ? image_1816 : _GEN_17243; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17245 = 12'h719 == _T_171[11:0] ? image_1817 : _GEN_17244; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17246 = 12'h71a == _T_171[11:0] ? image_1818 : _GEN_17245; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17247 = 12'h71b == _T_171[11:0] ? image_1819 : _GEN_17246; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17248 = 12'h71c == _T_171[11:0] ? image_1820 : _GEN_17247; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17249 = 12'h71d == _T_171[11:0] ? image_1821 : _GEN_17248; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17250 = 12'h71e == _T_171[11:0] ? image_1822 : _GEN_17249; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17251 = 12'h71f == _T_171[11:0] ? image_1823 : _GEN_17250; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17252 = 12'h720 == _T_171[11:0] ? image_1824 : _GEN_17251; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17253 = 12'h721 == _T_171[11:0] ? image_1825 : _GEN_17252; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17254 = 12'h722 == _T_171[11:0] ? image_1826 : _GEN_17253; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17255 = 12'h723 == _T_171[11:0] ? image_1827 : _GEN_17254; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17256 = 12'h724 == _T_171[11:0] ? image_1828 : _GEN_17255; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17257 = 12'h725 == _T_171[11:0] ? image_1829 : _GEN_17256; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17258 = 12'h726 == _T_171[11:0] ? image_1830 : _GEN_17257; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17259 = 12'h727 == _T_171[11:0] ? image_1831 : _GEN_17258; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17260 = 12'h728 == _T_171[11:0] ? image_1832 : _GEN_17259; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17261 = 12'h729 == _T_171[11:0] ? image_1833 : _GEN_17260; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17262 = 12'h72a == _T_171[11:0] ? image_1834 : _GEN_17261; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17263 = 12'h72b == _T_171[11:0] ? image_1835 : _GEN_17262; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17264 = 12'h72c == _T_171[11:0] ? image_1836 : _GEN_17263; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17265 = 12'h72d == _T_171[11:0] ? image_1837 : _GEN_17264; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17266 = 12'h72e == _T_171[11:0] ? image_1838 : _GEN_17265; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17267 = 12'h72f == _T_171[11:0] ? image_1839 : _GEN_17266; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17268 = 12'h730 == _T_171[11:0] ? image_1840 : _GEN_17267; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17269 = 12'h731 == _T_171[11:0] ? image_1841 : _GEN_17268; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17270 = 12'h732 == _T_171[11:0] ? image_1842 : _GEN_17269; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17271 = 12'h733 == _T_171[11:0] ? image_1843 : _GEN_17270; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17272 = 12'h734 == _T_171[11:0] ? image_1844 : _GEN_17271; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17273 = 12'h735 == _T_171[11:0] ? image_1845 : _GEN_17272; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17274 = 12'h736 == _T_171[11:0] ? image_1846 : _GEN_17273; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17275 = 12'h737 == _T_171[11:0] ? image_1847 : _GEN_17274; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17276 = 12'h738 == _T_171[11:0] ? image_1848 : _GEN_17275; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17277 = 12'h739 == _T_171[11:0] ? image_1849 : _GEN_17276; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17278 = 12'h73a == _T_171[11:0] ? 4'h0 : _GEN_17277; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17279 = 12'h73b == _T_171[11:0] ? 4'h0 : _GEN_17278; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17280 = 12'h73c == _T_171[11:0] ? 4'h0 : _GEN_17279; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17281 = 12'h73d == _T_171[11:0] ? 4'h0 : _GEN_17280; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17282 = 12'h73e == _T_171[11:0] ? 4'h0 : _GEN_17281; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17283 = 12'h73f == _T_171[11:0] ? 4'h0 : _GEN_17282; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17284 = 12'h740 == _T_171[11:0] ? 4'h0 : _GEN_17283; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17285 = 12'h741 == _T_171[11:0] ? image_1857 : _GEN_17284; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17286 = 12'h742 == _T_171[11:0] ? image_1858 : _GEN_17285; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17287 = 12'h743 == _T_171[11:0] ? image_1859 : _GEN_17286; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17288 = 12'h744 == _T_171[11:0] ? image_1860 : _GEN_17287; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17289 = 12'h745 == _T_171[11:0] ? image_1861 : _GEN_17288; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17290 = 12'h746 == _T_171[11:0] ? image_1862 : _GEN_17289; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17291 = 12'h747 == _T_171[11:0] ? image_1863 : _GEN_17290; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17292 = 12'h748 == _T_171[11:0] ? image_1864 : _GEN_17291; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17293 = 12'h749 == _T_171[11:0] ? image_1865 : _GEN_17292; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17294 = 12'h74a == _T_171[11:0] ? image_1866 : _GEN_17293; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17295 = 12'h74b == _T_171[11:0] ? image_1867 : _GEN_17294; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17296 = 12'h74c == _T_171[11:0] ? image_1868 : _GEN_17295; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17297 = 12'h74d == _T_171[11:0] ? image_1869 : _GEN_17296; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17298 = 12'h74e == _T_171[11:0] ? image_1870 : _GEN_17297; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17299 = 12'h74f == _T_171[11:0] ? image_1871 : _GEN_17298; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17300 = 12'h750 == _T_171[11:0] ? image_1872 : _GEN_17299; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17301 = 12'h751 == _T_171[11:0] ? image_1873 : _GEN_17300; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17302 = 12'h752 == _T_171[11:0] ? image_1874 : _GEN_17301; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17303 = 12'h753 == _T_171[11:0] ? image_1875 : _GEN_17302; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17304 = 12'h754 == _T_171[11:0] ? image_1876 : _GEN_17303; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17305 = 12'h755 == _T_171[11:0] ? image_1877 : _GEN_17304; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17306 = 12'h756 == _T_171[11:0] ? image_1878 : _GEN_17305; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17307 = 12'h757 == _T_171[11:0] ? image_1879 : _GEN_17306; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17308 = 12'h758 == _T_171[11:0] ? image_1880 : _GEN_17307; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17309 = 12'h759 == _T_171[11:0] ? image_1881 : _GEN_17308; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17310 = 12'h75a == _T_171[11:0] ? image_1882 : _GEN_17309; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17311 = 12'h75b == _T_171[11:0] ? image_1883 : _GEN_17310; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17312 = 12'h75c == _T_171[11:0] ? image_1884 : _GEN_17311; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17313 = 12'h75d == _T_171[11:0] ? image_1885 : _GEN_17312; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17314 = 12'h75e == _T_171[11:0] ? image_1886 : _GEN_17313; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17315 = 12'h75f == _T_171[11:0] ? image_1887 : _GEN_17314; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17316 = 12'h760 == _T_171[11:0] ? image_1888 : _GEN_17315; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17317 = 12'h761 == _T_171[11:0] ? image_1889 : _GEN_17316; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17318 = 12'h762 == _T_171[11:0] ? image_1890 : _GEN_17317; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17319 = 12'h763 == _T_171[11:0] ? image_1891 : _GEN_17318; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17320 = 12'h764 == _T_171[11:0] ? image_1892 : _GEN_17319; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17321 = 12'h765 == _T_171[11:0] ? image_1893 : _GEN_17320; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17322 = 12'h766 == _T_171[11:0] ? image_1894 : _GEN_17321; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17323 = 12'h767 == _T_171[11:0] ? image_1895 : _GEN_17322; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17324 = 12'h768 == _T_171[11:0] ? image_1896 : _GEN_17323; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17325 = 12'h769 == _T_171[11:0] ? image_1897 : _GEN_17324; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17326 = 12'h76a == _T_171[11:0] ? image_1898 : _GEN_17325; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17327 = 12'h76b == _T_171[11:0] ? image_1899 : _GEN_17326; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17328 = 12'h76c == _T_171[11:0] ? image_1900 : _GEN_17327; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17329 = 12'h76d == _T_171[11:0] ? image_1901 : _GEN_17328; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17330 = 12'h76e == _T_171[11:0] ? image_1902 : _GEN_17329; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17331 = 12'h76f == _T_171[11:0] ? image_1903 : _GEN_17330; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17332 = 12'h770 == _T_171[11:0] ? image_1904 : _GEN_17331; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17333 = 12'h771 == _T_171[11:0] ? image_1905 : _GEN_17332; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17334 = 12'h772 == _T_171[11:0] ? image_1906 : _GEN_17333; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17335 = 12'h773 == _T_171[11:0] ? image_1907 : _GEN_17334; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17336 = 12'h774 == _T_171[11:0] ? image_1908 : _GEN_17335; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17337 = 12'h775 == _T_171[11:0] ? image_1909 : _GEN_17336; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17338 = 12'h776 == _T_171[11:0] ? image_1910 : _GEN_17337; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17339 = 12'h777 == _T_171[11:0] ? image_1911 : _GEN_17338; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17340 = 12'h778 == _T_171[11:0] ? image_1912 : _GEN_17339; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17341 = 12'h779 == _T_171[11:0] ? image_1913 : _GEN_17340; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17342 = 12'h77a == _T_171[11:0] ? 4'h0 : _GEN_17341; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17343 = 12'h77b == _T_171[11:0] ? 4'h0 : _GEN_17342; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17344 = 12'h77c == _T_171[11:0] ? 4'h0 : _GEN_17343; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17345 = 12'h77d == _T_171[11:0] ? 4'h0 : _GEN_17344; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17346 = 12'h77e == _T_171[11:0] ? 4'h0 : _GEN_17345; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17347 = 12'h77f == _T_171[11:0] ? 4'h0 : _GEN_17346; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17348 = 12'h780 == _T_171[11:0] ? 4'h0 : _GEN_17347; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17349 = 12'h781 == _T_171[11:0] ? image_1921 : _GEN_17348; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17350 = 12'h782 == _T_171[11:0] ? image_1922 : _GEN_17349; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17351 = 12'h783 == _T_171[11:0] ? image_1923 : _GEN_17350; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17352 = 12'h784 == _T_171[11:0] ? image_1924 : _GEN_17351; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17353 = 12'h785 == _T_171[11:0] ? image_1925 : _GEN_17352; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17354 = 12'h786 == _T_171[11:0] ? image_1926 : _GEN_17353; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17355 = 12'h787 == _T_171[11:0] ? image_1927 : _GEN_17354; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17356 = 12'h788 == _T_171[11:0] ? image_1928 : _GEN_17355; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17357 = 12'h789 == _T_171[11:0] ? image_1929 : _GEN_17356; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17358 = 12'h78a == _T_171[11:0] ? image_1930 : _GEN_17357; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17359 = 12'h78b == _T_171[11:0] ? image_1931 : _GEN_17358; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17360 = 12'h78c == _T_171[11:0] ? image_1932 : _GEN_17359; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17361 = 12'h78d == _T_171[11:0] ? image_1933 : _GEN_17360; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17362 = 12'h78e == _T_171[11:0] ? image_1934 : _GEN_17361; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17363 = 12'h78f == _T_171[11:0] ? image_1935 : _GEN_17362; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17364 = 12'h790 == _T_171[11:0] ? image_1936 : _GEN_17363; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17365 = 12'h791 == _T_171[11:0] ? image_1937 : _GEN_17364; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17366 = 12'h792 == _T_171[11:0] ? image_1938 : _GEN_17365; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17367 = 12'h793 == _T_171[11:0] ? image_1939 : _GEN_17366; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17368 = 12'h794 == _T_171[11:0] ? image_1940 : _GEN_17367; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17369 = 12'h795 == _T_171[11:0] ? image_1941 : _GEN_17368; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17370 = 12'h796 == _T_171[11:0] ? image_1942 : _GEN_17369; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17371 = 12'h797 == _T_171[11:0] ? image_1943 : _GEN_17370; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17372 = 12'h798 == _T_171[11:0] ? image_1944 : _GEN_17371; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17373 = 12'h799 == _T_171[11:0] ? image_1945 : _GEN_17372; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17374 = 12'h79a == _T_171[11:0] ? image_1946 : _GEN_17373; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17375 = 12'h79b == _T_171[11:0] ? image_1947 : _GEN_17374; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17376 = 12'h79c == _T_171[11:0] ? image_1948 : _GEN_17375; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17377 = 12'h79d == _T_171[11:0] ? image_1949 : _GEN_17376; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17378 = 12'h79e == _T_171[11:0] ? image_1950 : _GEN_17377; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17379 = 12'h79f == _T_171[11:0] ? image_1951 : _GEN_17378; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17380 = 12'h7a0 == _T_171[11:0] ? image_1952 : _GEN_17379; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17381 = 12'h7a1 == _T_171[11:0] ? image_1953 : _GEN_17380; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17382 = 12'h7a2 == _T_171[11:0] ? image_1954 : _GEN_17381; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17383 = 12'h7a3 == _T_171[11:0] ? image_1955 : _GEN_17382; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17384 = 12'h7a4 == _T_171[11:0] ? image_1956 : _GEN_17383; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17385 = 12'h7a5 == _T_171[11:0] ? image_1957 : _GEN_17384; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17386 = 12'h7a6 == _T_171[11:0] ? image_1958 : _GEN_17385; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17387 = 12'h7a7 == _T_171[11:0] ? image_1959 : _GEN_17386; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17388 = 12'h7a8 == _T_171[11:0] ? image_1960 : _GEN_17387; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17389 = 12'h7a9 == _T_171[11:0] ? image_1961 : _GEN_17388; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17390 = 12'h7aa == _T_171[11:0] ? image_1962 : _GEN_17389; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17391 = 12'h7ab == _T_171[11:0] ? image_1963 : _GEN_17390; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17392 = 12'h7ac == _T_171[11:0] ? image_1964 : _GEN_17391; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17393 = 12'h7ad == _T_171[11:0] ? image_1965 : _GEN_17392; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17394 = 12'h7ae == _T_171[11:0] ? image_1966 : _GEN_17393; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17395 = 12'h7af == _T_171[11:0] ? image_1967 : _GEN_17394; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17396 = 12'h7b0 == _T_171[11:0] ? image_1968 : _GEN_17395; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17397 = 12'h7b1 == _T_171[11:0] ? image_1969 : _GEN_17396; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17398 = 12'h7b2 == _T_171[11:0] ? image_1970 : _GEN_17397; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17399 = 12'h7b3 == _T_171[11:0] ? image_1971 : _GEN_17398; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17400 = 12'h7b4 == _T_171[11:0] ? image_1972 : _GEN_17399; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17401 = 12'h7b5 == _T_171[11:0] ? image_1973 : _GEN_17400; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17402 = 12'h7b6 == _T_171[11:0] ? image_1974 : _GEN_17401; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17403 = 12'h7b7 == _T_171[11:0] ? image_1975 : _GEN_17402; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17404 = 12'h7b8 == _T_171[11:0] ? image_1976 : _GEN_17403; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17405 = 12'h7b9 == _T_171[11:0] ? image_1977 : _GEN_17404; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17406 = 12'h7ba == _T_171[11:0] ? 4'h0 : _GEN_17405; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17407 = 12'h7bb == _T_171[11:0] ? 4'h0 : _GEN_17406; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17408 = 12'h7bc == _T_171[11:0] ? 4'h0 : _GEN_17407; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17409 = 12'h7bd == _T_171[11:0] ? 4'h0 : _GEN_17408; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17410 = 12'h7be == _T_171[11:0] ? 4'h0 : _GEN_17409; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17411 = 12'h7bf == _T_171[11:0] ? 4'h0 : _GEN_17410; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17412 = 12'h7c0 == _T_171[11:0] ? 4'h0 : _GEN_17411; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17413 = 12'h7c1 == _T_171[11:0] ? image_1985 : _GEN_17412; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17414 = 12'h7c2 == _T_171[11:0] ? image_1986 : _GEN_17413; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17415 = 12'h7c3 == _T_171[11:0] ? image_1987 : _GEN_17414; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17416 = 12'h7c4 == _T_171[11:0] ? image_1988 : _GEN_17415; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17417 = 12'h7c5 == _T_171[11:0] ? image_1989 : _GEN_17416; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17418 = 12'h7c6 == _T_171[11:0] ? image_1990 : _GEN_17417; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17419 = 12'h7c7 == _T_171[11:0] ? image_1991 : _GEN_17418; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17420 = 12'h7c8 == _T_171[11:0] ? image_1992 : _GEN_17419; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17421 = 12'h7c9 == _T_171[11:0] ? image_1993 : _GEN_17420; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17422 = 12'h7ca == _T_171[11:0] ? image_1994 : _GEN_17421; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17423 = 12'h7cb == _T_171[11:0] ? image_1995 : _GEN_17422; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17424 = 12'h7cc == _T_171[11:0] ? image_1996 : _GEN_17423; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17425 = 12'h7cd == _T_171[11:0] ? image_1997 : _GEN_17424; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17426 = 12'h7ce == _T_171[11:0] ? image_1998 : _GEN_17425; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17427 = 12'h7cf == _T_171[11:0] ? image_1999 : _GEN_17426; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17428 = 12'h7d0 == _T_171[11:0] ? image_2000 : _GEN_17427; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17429 = 12'h7d1 == _T_171[11:0] ? image_2001 : _GEN_17428; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17430 = 12'h7d2 == _T_171[11:0] ? image_2002 : _GEN_17429; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17431 = 12'h7d3 == _T_171[11:0] ? image_2003 : _GEN_17430; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17432 = 12'h7d4 == _T_171[11:0] ? image_2004 : _GEN_17431; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17433 = 12'h7d5 == _T_171[11:0] ? image_2005 : _GEN_17432; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17434 = 12'h7d6 == _T_171[11:0] ? image_2006 : _GEN_17433; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17435 = 12'h7d7 == _T_171[11:0] ? image_2007 : _GEN_17434; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17436 = 12'h7d8 == _T_171[11:0] ? image_2008 : _GEN_17435; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17437 = 12'h7d9 == _T_171[11:0] ? image_2009 : _GEN_17436; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17438 = 12'h7da == _T_171[11:0] ? image_2010 : _GEN_17437; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17439 = 12'h7db == _T_171[11:0] ? image_2011 : _GEN_17438; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17440 = 12'h7dc == _T_171[11:0] ? image_2012 : _GEN_17439; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17441 = 12'h7dd == _T_171[11:0] ? image_2013 : _GEN_17440; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17442 = 12'h7de == _T_171[11:0] ? image_2014 : _GEN_17441; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17443 = 12'h7df == _T_171[11:0] ? image_2015 : _GEN_17442; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17444 = 12'h7e0 == _T_171[11:0] ? image_2016 : _GEN_17443; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17445 = 12'h7e1 == _T_171[11:0] ? image_2017 : _GEN_17444; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17446 = 12'h7e2 == _T_171[11:0] ? image_2018 : _GEN_17445; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17447 = 12'h7e3 == _T_171[11:0] ? image_2019 : _GEN_17446; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17448 = 12'h7e4 == _T_171[11:0] ? image_2020 : _GEN_17447; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17449 = 12'h7e5 == _T_171[11:0] ? image_2021 : _GEN_17448; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17450 = 12'h7e6 == _T_171[11:0] ? image_2022 : _GEN_17449; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17451 = 12'h7e7 == _T_171[11:0] ? image_2023 : _GEN_17450; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17452 = 12'h7e8 == _T_171[11:0] ? image_2024 : _GEN_17451; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17453 = 12'h7e9 == _T_171[11:0] ? image_2025 : _GEN_17452; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17454 = 12'h7ea == _T_171[11:0] ? image_2026 : _GEN_17453; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17455 = 12'h7eb == _T_171[11:0] ? image_2027 : _GEN_17454; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17456 = 12'h7ec == _T_171[11:0] ? image_2028 : _GEN_17455; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17457 = 12'h7ed == _T_171[11:0] ? image_2029 : _GEN_17456; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17458 = 12'h7ee == _T_171[11:0] ? image_2030 : _GEN_17457; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17459 = 12'h7ef == _T_171[11:0] ? image_2031 : _GEN_17458; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17460 = 12'h7f0 == _T_171[11:0] ? image_2032 : _GEN_17459; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17461 = 12'h7f1 == _T_171[11:0] ? image_2033 : _GEN_17460; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17462 = 12'h7f2 == _T_171[11:0] ? image_2034 : _GEN_17461; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17463 = 12'h7f3 == _T_171[11:0] ? image_2035 : _GEN_17462; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17464 = 12'h7f4 == _T_171[11:0] ? image_2036 : _GEN_17463; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17465 = 12'h7f5 == _T_171[11:0] ? image_2037 : _GEN_17464; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17466 = 12'h7f6 == _T_171[11:0] ? image_2038 : _GEN_17465; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17467 = 12'h7f7 == _T_171[11:0] ? image_2039 : _GEN_17466; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17468 = 12'h7f8 == _T_171[11:0] ? image_2040 : _GEN_17467; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17469 = 12'h7f9 == _T_171[11:0] ? image_2041 : _GEN_17468; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17470 = 12'h7fa == _T_171[11:0] ? 4'h0 : _GEN_17469; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17471 = 12'h7fb == _T_171[11:0] ? 4'h0 : _GEN_17470; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17472 = 12'h7fc == _T_171[11:0] ? 4'h0 : _GEN_17471; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17473 = 12'h7fd == _T_171[11:0] ? 4'h0 : _GEN_17472; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17474 = 12'h7fe == _T_171[11:0] ? 4'h0 : _GEN_17473; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17475 = 12'h7ff == _T_171[11:0] ? 4'h0 : _GEN_17474; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17476 = 12'h800 == _T_171[11:0] ? 4'h0 : _GEN_17475; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17477 = 12'h801 == _T_171[11:0] ? image_2049 : _GEN_17476; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17478 = 12'h802 == _T_171[11:0] ? image_2050 : _GEN_17477; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17479 = 12'h803 == _T_171[11:0] ? image_2051 : _GEN_17478; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17480 = 12'h804 == _T_171[11:0] ? image_2052 : _GEN_17479; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17481 = 12'h805 == _T_171[11:0] ? image_2053 : _GEN_17480; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17482 = 12'h806 == _T_171[11:0] ? image_2054 : _GEN_17481; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17483 = 12'h807 == _T_171[11:0] ? image_2055 : _GEN_17482; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17484 = 12'h808 == _T_171[11:0] ? image_2056 : _GEN_17483; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17485 = 12'h809 == _T_171[11:0] ? image_2057 : _GEN_17484; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17486 = 12'h80a == _T_171[11:0] ? image_2058 : _GEN_17485; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17487 = 12'h80b == _T_171[11:0] ? image_2059 : _GEN_17486; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17488 = 12'h80c == _T_171[11:0] ? image_2060 : _GEN_17487; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17489 = 12'h80d == _T_171[11:0] ? image_2061 : _GEN_17488; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17490 = 12'h80e == _T_171[11:0] ? image_2062 : _GEN_17489; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17491 = 12'h80f == _T_171[11:0] ? image_2063 : _GEN_17490; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17492 = 12'h810 == _T_171[11:0] ? image_2064 : _GEN_17491; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17493 = 12'h811 == _T_171[11:0] ? image_2065 : _GEN_17492; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17494 = 12'h812 == _T_171[11:0] ? image_2066 : _GEN_17493; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17495 = 12'h813 == _T_171[11:0] ? image_2067 : _GEN_17494; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17496 = 12'h814 == _T_171[11:0] ? image_2068 : _GEN_17495; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17497 = 12'h815 == _T_171[11:0] ? image_2069 : _GEN_17496; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17498 = 12'h816 == _T_171[11:0] ? image_2070 : _GEN_17497; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17499 = 12'h817 == _T_171[11:0] ? image_2071 : _GEN_17498; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17500 = 12'h818 == _T_171[11:0] ? image_2072 : _GEN_17499; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17501 = 12'h819 == _T_171[11:0] ? image_2073 : _GEN_17500; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17502 = 12'h81a == _T_171[11:0] ? image_2074 : _GEN_17501; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17503 = 12'h81b == _T_171[11:0] ? image_2075 : _GEN_17502; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17504 = 12'h81c == _T_171[11:0] ? image_2076 : _GEN_17503; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17505 = 12'h81d == _T_171[11:0] ? image_2077 : _GEN_17504; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17506 = 12'h81e == _T_171[11:0] ? image_2078 : _GEN_17505; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17507 = 12'h81f == _T_171[11:0] ? image_2079 : _GEN_17506; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17508 = 12'h820 == _T_171[11:0] ? image_2080 : _GEN_17507; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17509 = 12'h821 == _T_171[11:0] ? image_2081 : _GEN_17508; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17510 = 12'h822 == _T_171[11:0] ? image_2082 : _GEN_17509; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17511 = 12'h823 == _T_171[11:0] ? image_2083 : _GEN_17510; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17512 = 12'h824 == _T_171[11:0] ? image_2084 : _GEN_17511; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17513 = 12'h825 == _T_171[11:0] ? image_2085 : _GEN_17512; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17514 = 12'h826 == _T_171[11:0] ? image_2086 : _GEN_17513; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17515 = 12'h827 == _T_171[11:0] ? image_2087 : _GEN_17514; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17516 = 12'h828 == _T_171[11:0] ? image_2088 : _GEN_17515; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17517 = 12'h829 == _T_171[11:0] ? image_2089 : _GEN_17516; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17518 = 12'h82a == _T_171[11:0] ? image_2090 : _GEN_17517; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17519 = 12'h82b == _T_171[11:0] ? image_2091 : _GEN_17518; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17520 = 12'h82c == _T_171[11:0] ? image_2092 : _GEN_17519; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17521 = 12'h82d == _T_171[11:0] ? image_2093 : _GEN_17520; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17522 = 12'h82e == _T_171[11:0] ? image_2094 : _GEN_17521; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17523 = 12'h82f == _T_171[11:0] ? image_2095 : _GEN_17522; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17524 = 12'h830 == _T_171[11:0] ? image_2096 : _GEN_17523; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17525 = 12'h831 == _T_171[11:0] ? image_2097 : _GEN_17524; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17526 = 12'h832 == _T_171[11:0] ? image_2098 : _GEN_17525; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17527 = 12'h833 == _T_171[11:0] ? image_2099 : _GEN_17526; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17528 = 12'h834 == _T_171[11:0] ? image_2100 : _GEN_17527; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17529 = 12'h835 == _T_171[11:0] ? image_2101 : _GEN_17528; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17530 = 12'h836 == _T_171[11:0] ? image_2102 : _GEN_17529; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17531 = 12'h837 == _T_171[11:0] ? image_2103 : _GEN_17530; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17532 = 12'h838 == _T_171[11:0] ? image_2104 : _GEN_17531; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17533 = 12'h839 == _T_171[11:0] ? image_2105 : _GEN_17532; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17534 = 12'h83a == _T_171[11:0] ? image_2106 : _GEN_17533; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17535 = 12'h83b == _T_171[11:0] ? 4'h0 : _GEN_17534; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17536 = 12'h83c == _T_171[11:0] ? 4'h0 : _GEN_17535; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17537 = 12'h83d == _T_171[11:0] ? 4'h0 : _GEN_17536; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17538 = 12'h83e == _T_171[11:0] ? 4'h0 : _GEN_17537; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17539 = 12'h83f == _T_171[11:0] ? 4'h0 : _GEN_17538; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17540 = 12'h840 == _T_171[11:0] ? 4'h0 : _GEN_17539; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17541 = 12'h841 == _T_171[11:0] ? 4'h0 : _GEN_17540; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17542 = 12'h842 == _T_171[11:0] ? image_2114 : _GEN_17541; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17543 = 12'h843 == _T_171[11:0] ? image_2115 : _GEN_17542; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17544 = 12'h844 == _T_171[11:0] ? image_2116 : _GEN_17543; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17545 = 12'h845 == _T_171[11:0] ? image_2117 : _GEN_17544; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17546 = 12'h846 == _T_171[11:0] ? image_2118 : _GEN_17545; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17547 = 12'h847 == _T_171[11:0] ? image_2119 : _GEN_17546; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17548 = 12'h848 == _T_171[11:0] ? image_2120 : _GEN_17547; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17549 = 12'h849 == _T_171[11:0] ? image_2121 : _GEN_17548; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17550 = 12'h84a == _T_171[11:0] ? image_2122 : _GEN_17549; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17551 = 12'h84b == _T_171[11:0] ? image_2123 : _GEN_17550; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17552 = 12'h84c == _T_171[11:0] ? image_2124 : _GEN_17551; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17553 = 12'h84d == _T_171[11:0] ? image_2125 : _GEN_17552; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17554 = 12'h84e == _T_171[11:0] ? image_2126 : _GEN_17553; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17555 = 12'h84f == _T_171[11:0] ? image_2127 : _GEN_17554; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17556 = 12'h850 == _T_171[11:0] ? image_2128 : _GEN_17555; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17557 = 12'h851 == _T_171[11:0] ? image_2129 : _GEN_17556; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17558 = 12'h852 == _T_171[11:0] ? image_2130 : _GEN_17557; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17559 = 12'h853 == _T_171[11:0] ? image_2131 : _GEN_17558; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17560 = 12'h854 == _T_171[11:0] ? image_2132 : _GEN_17559; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17561 = 12'h855 == _T_171[11:0] ? image_2133 : _GEN_17560; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17562 = 12'h856 == _T_171[11:0] ? image_2134 : _GEN_17561; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17563 = 12'h857 == _T_171[11:0] ? image_2135 : _GEN_17562; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17564 = 12'h858 == _T_171[11:0] ? image_2136 : _GEN_17563; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17565 = 12'h859 == _T_171[11:0] ? image_2137 : _GEN_17564; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17566 = 12'h85a == _T_171[11:0] ? image_2138 : _GEN_17565; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17567 = 12'h85b == _T_171[11:0] ? image_2139 : _GEN_17566; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17568 = 12'h85c == _T_171[11:0] ? image_2140 : _GEN_17567; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17569 = 12'h85d == _T_171[11:0] ? image_2141 : _GEN_17568; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17570 = 12'h85e == _T_171[11:0] ? image_2142 : _GEN_17569; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17571 = 12'h85f == _T_171[11:0] ? image_2143 : _GEN_17570; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17572 = 12'h860 == _T_171[11:0] ? image_2144 : _GEN_17571; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17573 = 12'h861 == _T_171[11:0] ? image_2145 : _GEN_17572; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17574 = 12'h862 == _T_171[11:0] ? image_2146 : _GEN_17573; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17575 = 12'h863 == _T_171[11:0] ? image_2147 : _GEN_17574; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17576 = 12'h864 == _T_171[11:0] ? image_2148 : _GEN_17575; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17577 = 12'h865 == _T_171[11:0] ? image_2149 : _GEN_17576; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17578 = 12'h866 == _T_171[11:0] ? image_2150 : _GEN_17577; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17579 = 12'h867 == _T_171[11:0] ? image_2151 : _GEN_17578; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17580 = 12'h868 == _T_171[11:0] ? image_2152 : _GEN_17579; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17581 = 12'h869 == _T_171[11:0] ? image_2153 : _GEN_17580; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17582 = 12'h86a == _T_171[11:0] ? image_2154 : _GEN_17581; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17583 = 12'h86b == _T_171[11:0] ? image_2155 : _GEN_17582; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17584 = 12'h86c == _T_171[11:0] ? image_2156 : _GEN_17583; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17585 = 12'h86d == _T_171[11:0] ? image_2157 : _GEN_17584; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17586 = 12'h86e == _T_171[11:0] ? image_2158 : _GEN_17585; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17587 = 12'h86f == _T_171[11:0] ? image_2159 : _GEN_17586; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17588 = 12'h870 == _T_171[11:0] ? image_2160 : _GEN_17587; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17589 = 12'h871 == _T_171[11:0] ? image_2161 : _GEN_17588; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17590 = 12'h872 == _T_171[11:0] ? image_2162 : _GEN_17589; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17591 = 12'h873 == _T_171[11:0] ? image_2163 : _GEN_17590; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17592 = 12'h874 == _T_171[11:0] ? image_2164 : _GEN_17591; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17593 = 12'h875 == _T_171[11:0] ? image_2165 : _GEN_17592; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17594 = 12'h876 == _T_171[11:0] ? image_2166 : _GEN_17593; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17595 = 12'h877 == _T_171[11:0] ? image_2167 : _GEN_17594; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17596 = 12'h878 == _T_171[11:0] ? image_2168 : _GEN_17595; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17597 = 12'h879 == _T_171[11:0] ? image_2169 : _GEN_17596; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17598 = 12'h87a == _T_171[11:0] ? image_2170 : _GEN_17597; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17599 = 12'h87b == _T_171[11:0] ? 4'h0 : _GEN_17598; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17600 = 12'h87c == _T_171[11:0] ? 4'h0 : _GEN_17599; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17601 = 12'h87d == _T_171[11:0] ? 4'h0 : _GEN_17600; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17602 = 12'h87e == _T_171[11:0] ? 4'h0 : _GEN_17601; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17603 = 12'h87f == _T_171[11:0] ? 4'h0 : _GEN_17602; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17604 = 12'h880 == _T_171[11:0] ? 4'h0 : _GEN_17603; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17605 = 12'h881 == _T_171[11:0] ? image_2177 : _GEN_17604; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17606 = 12'h882 == _T_171[11:0] ? image_2178 : _GEN_17605; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17607 = 12'h883 == _T_171[11:0] ? image_2179 : _GEN_17606; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17608 = 12'h884 == _T_171[11:0] ? image_2180 : _GEN_17607; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17609 = 12'h885 == _T_171[11:0] ? image_2181 : _GEN_17608; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17610 = 12'h886 == _T_171[11:0] ? image_2182 : _GEN_17609; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17611 = 12'h887 == _T_171[11:0] ? image_2183 : _GEN_17610; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17612 = 12'h888 == _T_171[11:0] ? image_2184 : _GEN_17611; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17613 = 12'h889 == _T_171[11:0] ? image_2185 : _GEN_17612; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17614 = 12'h88a == _T_171[11:0] ? image_2186 : _GEN_17613; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17615 = 12'h88b == _T_171[11:0] ? image_2187 : _GEN_17614; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17616 = 12'h88c == _T_171[11:0] ? image_2188 : _GEN_17615; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17617 = 12'h88d == _T_171[11:0] ? image_2189 : _GEN_17616; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17618 = 12'h88e == _T_171[11:0] ? image_2190 : _GEN_17617; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17619 = 12'h88f == _T_171[11:0] ? image_2191 : _GEN_17618; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17620 = 12'h890 == _T_171[11:0] ? image_2192 : _GEN_17619; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17621 = 12'h891 == _T_171[11:0] ? image_2193 : _GEN_17620; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17622 = 12'h892 == _T_171[11:0] ? image_2194 : _GEN_17621; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17623 = 12'h893 == _T_171[11:0] ? image_2195 : _GEN_17622; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17624 = 12'h894 == _T_171[11:0] ? image_2196 : _GEN_17623; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17625 = 12'h895 == _T_171[11:0] ? image_2197 : _GEN_17624; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17626 = 12'h896 == _T_171[11:0] ? image_2198 : _GEN_17625; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17627 = 12'h897 == _T_171[11:0] ? image_2199 : _GEN_17626; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17628 = 12'h898 == _T_171[11:0] ? image_2200 : _GEN_17627; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17629 = 12'h899 == _T_171[11:0] ? image_2201 : _GEN_17628; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17630 = 12'h89a == _T_171[11:0] ? image_2202 : _GEN_17629; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17631 = 12'h89b == _T_171[11:0] ? image_2203 : _GEN_17630; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17632 = 12'h89c == _T_171[11:0] ? image_2204 : _GEN_17631; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17633 = 12'h89d == _T_171[11:0] ? image_2205 : _GEN_17632; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17634 = 12'h89e == _T_171[11:0] ? image_2206 : _GEN_17633; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17635 = 12'h89f == _T_171[11:0] ? image_2207 : _GEN_17634; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17636 = 12'h8a0 == _T_171[11:0] ? image_2208 : _GEN_17635; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17637 = 12'h8a1 == _T_171[11:0] ? image_2209 : _GEN_17636; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17638 = 12'h8a2 == _T_171[11:0] ? image_2210 : _GEN_17637; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17639 = 12'h8a3 == _T_171[11:0] ? image_2211 : _GEN_17638; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17640 = 12'h8a4 == _T_171[11:0] ? image_2212 : _GEN_17639; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17641 = 12'h8a5 == _T_171[11:0] ? image_2213 : _GEN_17640; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17642 = 12'h8a6 == _T_171[11:0] ? image_2214 : _GEN_17641; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17643 = 12'h8a7 == _T_171[11:0] ? image_2215 : _GEN_17642; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17644 = 12'h8a8 == _T_171[11:0] ? image_2216 : _GEN_17643; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17645 = 12'h8a9 == _T_171[11:0] ? image_2217 : _GEN_17644; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17646 = 12'h8aa == _T_171[11:0] ? image_2218 : _GEN_17645; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17647 = 12'h8ab == _T_171[11:0] ? image_2219 : _GEN_17646; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17648 = 12'h8ac == _T_171[11:0] ? image_2220 : _GEN_17647; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17649 = 12'h8ad == _T_171[11:0] ? image_2221 : _GEN_17648; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17650 = 12'h8ae == _T_171[11:0] ? image_2222 : _GEN_17649; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17651 = 12'h8af == _T_171[11:0] ? image_2223 : _GEN_17650; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17652 = 12'h8b0 == _T_171[11:0] ? image_2224 : _GEN_17651; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17653 = 12'h8b1 == _T_171[11:0] ? image_2225 : _GEN_17652; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17654 = 12'h8b2 == _T_171[11:0] ? image_2226 : _GEN_17653; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17655 = 12'h8b3 == _T_171[11:0] ? image_2227 : _GEN_17654; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17656 = 12'h8b4 == _T_171[11:0] ? image_2228 : _GEN_17655; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17657 = 12'h8b5 == _T_171[11:0] ? image_2229 : _GEN_17656; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17658 = 12'h8b6 == _T_171[11:0] ? image_2230 : _GEN_17657; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17659 = 12'h8b7 == _T_171[11:0] ? image_2231 : _GEN_17658; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17660 = 12'h8b8 == _T_171[11:0] ? image_2232 : _GEN_17659; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17661 = 12'h8b9 == _T_171[11:0] ? image_2233 : _GEN_17660; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17662 = 12'h8ba == _T_171[11:0] ? image_2234 : _GEN_17661; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17663 = 12'h8bb == _T_171[11:0] ? 4'h0 : _GEN_17662; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17664 = 12'h8bc == _T_171[11:0] ? 4'h0 : _GEN_17663; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17665 = 12'h8bd == _T_171[11:0] ? 4'h0 : _GEN_17664; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17666 = 12'h8be == _T_171[11:0] ? 4'h0 : _GEN_17665; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17667 = 12'h8bf == _T_171[11:0] ? 4'h0 : _GEN_17666; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17668 = 12'h8c0 == _T_171[11:0] ? 4'h0 : _GEN_17667; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17669 = 12'h8c1 == _T_171[11:0] ? 4'h0 : _GEN_17668; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17670 = 12'h8c2 == _T_171[11:0] ? 4'h0 : _GEN_17669; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17671 = 12'h8c3 == _T_171[11:0] ? image_2243 : _GEN_17670; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17672 = 12'h8c4 == _T_171[11:0] ? image_2244 : _GEN_17671; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17673 = 12'h8c5 == _T_171[11:0] ? image_2245 : _GEN_17672; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17674 = 12'h8c6 == _T_171[11:0] ? image_2246 : _GEN_17673; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17675 = 12'h8c7 == _T_171[11:0] ? image_2247 : _GEN_17674; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17676 = 12'h8c8 == _T_171[11:0] ? image_2248 : _GEN_17675; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17677 = 12'h8c9 == _T_171[11:0] ? image_2249 : _GEN_17676; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17678 = 12'h8ca == _T_171[11:0] ? image_2250 : _GEN_17677; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17679 = 12'h8cb == _T_171[11:0] ? image_2251 : _GEN_17678; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17680 = 12'h8cc == _T_171[11:0] ? image_2252 : _GEN_17679; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17681 = 12'h8cd == _T_171[11:0] ? image_2253 : _GEN_17680; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17682 = 12'h8ce == _T_171[11:0] ? image_2254 : _GEN_17681; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17683 = 12'h8cf == _T_171[11:0] ? image_2255 : _GEN_17682; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17684 = 12'h8d0 == _T_171[11:0] ? image_2256 : _GEN_17683; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17685 = 12'h8d1 == _T_171[11:0] ? image_2257 : _GEN_17684; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17686 = 12'h8d2 == _T_171[11:0] ? image_2258 : _GEN_17685; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17687 = 12'h8d3 == _T_171[11:0] ? image_2259 : _GEN_17686; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17688 = 12'h8d4 == _T_171[11:0] ? image_2260 : _GEN_17687; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17689 = 12'h8d5 == _T_171[11:0] ? image_2261 : _GEN_17688; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17690 = 12'h8d6 == _T_171[11:0] ? image_2262 : _GEN_17689; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17691 = 12'h8d7 == _T_171[11:0] ? image_2263 : _GEN_17690; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17692 = 12'h8d8 == _T_171[11:0] ? image_2264 : _GEN_17691; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17693 = 12'h8d9 == _T_171[11:0] ? image_2265 : _GEN_17692; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17694 = 12'h8da == _T_171[11:0] ? image_2266 : _GEN_17693; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17695 = 12'h8db == _T_171[11:0] ? image_2267 : _GEN_17694; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17696 = 12'h8dc == _T_171[11:0] ? image_2268 : _GEN_17695; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17697 = 12'h8dd == _T_171[11:0] ? image_2269 : _GEN_17696; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17698 = 12'h8de == _T_171[11:0] ? image_2270 : _GEN_17697; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17699 = 12'h8df == _T_171[11:0] ? image_2271 : _GEN_17698; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17700 = 12'h8e0 == _T_171[11:0] ? image_2272 : _GEN_17699; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17701 = 12'h8e1 == _T_171[11:0] ? image_2273 : _GEN_17700; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17702 = 12'h8e2 == _T_171[11:0] ? image_2274 : _GEN_17701; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17703 = 12'h8e3 == _T_171[11:0] ? image_2275 : _GEN_17702; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17704 = 12'h8e4 == _T_171[11:0] ? image_2276 : _GEN_17703; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17705 = 12'h8e5 == _T_171[11:0] ? image_2277 : _GEN_17704; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17706 = 12'h8e6 == _T_171[11:0] ? image_2278 : _GEN_17705; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17707 = 12'h8e7 == _T_171[11:0] ? image_2279 : _GEN_17706; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17708 = 12'h8e8 == _T_171[11:0] ? image_2280 : _GEN_17707; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17709 = 12'h8e9 == _T_171[11:0] ? image_2281 : _GEN_17708; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17710 = 12'h8ea == _T_171[11:0] ? image_2282 : _GEN_17709; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17711 = 12'h8eb == _T_171[11:0] ? image_2283 : _GEN_17710; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17712 = 12'h8ec == _T_171[11:0] ? image_2284 : _GEN_17711; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17713 = 12'h8ed == _T_171[11:0] ? image_2285 : _GEN_17712; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17714 = 12'h8ee == _T_171[11:0] ? image_2286 : _GEN_17713; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17715 = 12'h8ef == _T_171[11:0] ? image_2287 : _GEN_17714; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17716 = 12'h8f0 == _T_171[11:0] ? image_2288 : _GEN_17715; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17717 = 12'h8f1 == _T_171[11:0] ? image_2289 : _GEN_17716; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17718 = 12'h8f2 == _T_171[11:0] ? image_2290 : _GEN_17717; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17719 = 12'h8f3 == _T_171[11:0] ? image_2291 : _GEN_17718; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17720 = 12'h8f4 == _T_171[11:0] ? image_2292 : _GEN_17719; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17721 = 12'h8f5 == _T_171[11:0] ? image_2293 : _GEN_17720; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17722 = 12'h8f6 == _T_171[11:0] ? image_2294 : _GEN_17721; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17723 = 12'h8f7 == _T_171[11:0] ? image_2295 : _GEN_17722; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17724 = 12'h8f8 == _T_171[11:0] ? image_2296 : _GEN_17723; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17725 = 12'h8f9 == _T_171[11:0] ? image_2297 : _GEN_17724; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17726 = 12'h8fa == _T_171[11:0] ? image_2298 : _GEN_17725; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17727 = 12'h8fb == _T_171[11:0] ? 4'h0 : _GEN_17726; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17728 = 12'h8fc == _T_171[11:0] ? 4'h0 : _GEN_17727; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17729 = 12'h8fd == _T_171[11:0] ? 4'h0 : _GEN_17728; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17730 = 12'h8fe == _T_171[11:0] ? 4'h0 : _GEN_17729; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17731 = 12'h8ff == _T_171[11:0] ? 4'h0 : _GEN_17730; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17732 = 12'h900 == _T_171[11:0] ? 4'h0 : _GEN_17731; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17733 = 12'h901 == _T_171[11:0] ? 4'h0 : _GEN_17732; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17734 = 12'h902 == _T_171[11:0] ? 4'h0 : _GEN_17733; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17735 = 12'h903 == _T_171[11:0] ? image_2307 : _GEN_17734; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17736 = 12'h904 == _T_171[11:0] ? image_2308 : _GEN_17735; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17737 = 12'h905 == _T_171[11:0] ? image_2309 : _GEN_17736; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17738 = 12'h906 == _T_171[11:0] ? image_2310 : _GEN_17737; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17739 = 12'h907 == _T_171[11:0] ? image_2311 : _GEN_17738; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17740 = 12'h908 == _T_171[11:0] ? image_2312 : _GEN_17739; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17741 = 12'h909 == _T_171[11:0] ? image_2313 : _GEN_17740; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17742 = 12'h90a == _T_171[11:0] ? image_2314 : _GEN_17741; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17743 = 12'h90b == _T_171[11:0] ? image_2315 : _GEN_17742; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17744 = 12'h90c == _T_171[11:0] ? image_2316 : _GEN_17743; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17745 = 12'h90d == _T_171[11:0] ? image_2317 : _GEN_17744; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17746 = 12'h90e == _T_171[11:0] ? image_2318 : _GEN_17745; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17747 = 12'h90f == _T_171[11:0] ? image_2319 : _GEN_17746; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17748 = 12'h910 == _T_171[11:0] ? image_2320 : _GEN_17747; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17749 = 12'h911 == _T_171[11:0] ? image_2321 : _GEN_17748; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17750 = 12'h912 == _T_171[11:0] ? image_2322 : _GEN_17749; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17751 = 12'h913 == _T_171[11:0] ? image_2323 : _GEN_17750; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17752 = 12'h914 == _T_171[11:0] ? image_2324 : _GEN_17751; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17753 = 12'h915 == _T_171[11:0] ? image_2325 : _GEN_17752; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17754 = 12'h916 == _T_171[11:0] ? image_2326 : _GEN_17753; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17755 = 12'h917 == _T_171[11:0] ? image_2327 : _GEN_17754; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17756 = 12'h918 == _T_171[11:0] ? image_2328 : _GEN_17755; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17757 = 12'h919 == _T_171[11:0] ? image_2329 : _GEN_17756; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17758 = 12'h91a == _T_171[11:0] ? image_2330 : _GEN_17757; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17759 = 12'h91b == _T_171[11:0] ? image_2331 : _GEN_17758; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17760 = 12'h91c == _T_171[11:0] ? image_2332 : _GEN_17759; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17761 = 12'h91d == _T_171[11:0] ? image_2333 : _GEN_17760; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17762 = 12'h91e == _T_171[11:0] ? image_2334 : _GEN_17761; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17763 = 12'h91f == _T_171[11:0] ? image_2335 : _GEN_17762; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17764 = 12'h920 == _T_171[11:0] ? image_2336 : _GEN_17763; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17765 = 12'h921 == _T_171[11:0] ? image_2337 : _GEN_17764; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17766 = 12'h922 == _T_171[11:0] ? image_2338 : _GEN_17765; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17767 = 12'h923 == _T_171[11:0] ? image_2339 : _GEN_17766; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17768 = 12'h924 == _T_171[11:0] ? image_2340 : _GEN_17767; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17769 = 12'h925 == _T_171[11:0] ? image_2341 : _GEN_17768; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17770 = 12'h926 == _T_171[11:0] ? image_2342 : _GEN_17769; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17771 = 12'h927 == _T_171[11:0] ? image_2343 : _GEN_17770; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17772 = 12'h928 == _T_171[11:0] ? image_2344 : _GEN_17771; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17773 = 12'h929 == _T_171[11:0] ? image_2345 : _GEN_17772; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17774 = 12'h92a == _T_171[11:0] ? image_2346 : _GEN_17773; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17775 = 12'h92b == _T_171[11:0] ? image_2347 : _GEN_17774; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17776 = 12'h92c == _T_171[11:0] ? image_2348 : _GEN_17775; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17777 = 12'h92d == _T_171[11:0] ? image_2349 : _GEN_17776; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17778 = 12'h92e == _T_171[11:0] ? image_2350 : _GEN_17777; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17779 = 12'h92f == _T_171[11:0] ? image_2351 : _GEN_17778; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17780 = 12'h930 == _T_171[11:0] ? image_2352 : _GEN_17779; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17781 = 12'h931 == _T_171[11:0] ? image_2353 : _GEN_17780; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17782 = 12'h932 == _T_171[11:0] ? image_2354 : _GEN_17781; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17783 = 12'h933 == _T_171[11:0] ? image_2355 : _GEN_17782; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17784 = 12'h934 == _T_171[11:0] ? image_2356 : _GEN_17783; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17785 = 12'h935 == _T_171[11:0] ? image_2357 : _GEN_17784; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17786 = 12'h936 == _T_171[11:0] ? image_2358 : _GEN_17785; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17787 = 12'h937 == _T_171[11:0] ? image_2359 : _GEN_17786; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17788 = 12'h938 == _T_171[11:0] ? image_2360 : _GEN_17787; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17789 = 12'h939 == _T_171[11:0] ? image_2361 : _GEN_17788; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17790 = 12'h93a == _T_171[11:0] ? image_2362 : _GEN_17789; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17791 = 12'h93b == _T_171[11:0] ? 4'h0 : _GEN_17790; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17792 = 12'h93c == _T_171[11:0] ? 4'h0 : _GEN_17791; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17793 = 12'h93d == _T_171[11:0] ? 4'h0 : _GEN_17792; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17794 = 12'h93e == _T_171[11:0] ? 4'h0 : _GEN_17793; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17795 = 12'h93f == _T_171[11:0] ? 4'h0 : _GEN_17794; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17796 = 12'h940 == _T_171[11:0] ? 4'h0 : _GEN_17795; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17797 = 12'h941 == _T_171[11:0] ? 4'h0 : _GEN_17796; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17798 = 12'h942 == _T_171[11:0] ? 4'h0 : _GEN_17797; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17799 = 12'h943 == _T_171[11:0] ? 4'h0 : _GEN_17798; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17800 = 12'h944 == _T_171[11:0] ? image_2372 : _GEN_17799; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17801 = 12'h945 == _T_171[11:0] ? image_2373 : _GEN_17800; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17802 = 12'h946 == _T_171[11:0] ? image_2374 : _GEN_17801; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17803 = 12'h947 == _T_171[11:0] ? image_2375 : _GEN_17802; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17804 = 12'h948 == _T_171[11:0] ? image_2376 : _GEN_17803; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17805 = 12'h949 == _T_171[11:0] ? image_2377 : _GEN_17804; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17806 = 12'h94a == _T_171[11:0] ? image_2378 : _GEN_17805; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17807 = 12'h94b == _T_171[11:0] ? image_2379 : _GEN_17806; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17808 = 12'h94c == _T_171[11:0] ? image_2380 : _GEN_17807; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17809 = 12'h94d == _T_171[11:0] ? image_2381 : _GEN_17808; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17810 = 12'h94e == _T_171[11:0] ? image_2382 : _GEN_17809; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17811 = 12'h94f == _T_171[11:0] ? image_2383 : _GEN_17810; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17812 = 12'h950 == _T_171[11:0] ? image_2384 : _GEN_17811; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17813 = 12'h951 == _T_171[11:0] ? image_2385 : _GEN_17812; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17814 = 12'h952 == _T_171[11:0] ? image_2386 : _GEN_17813; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17815 = 12'h953 == _T_171[11:0] ? image_2387 : _GEN_17814; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17816 = 12'h954 == _T_171[11:0] ? image_2388 : _GEN_17815; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17817 = 12'h955 == _T_171[11:0] ? image_2389 : _GEN_17816; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17818 = 12'h956 == _T_171[11:0] ? image_2390 : _GEN_17817; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17819 = 12'h957 == _T_171[11:0] ? image_2391 : _GEN_17818; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17820 = 12'h958 == _T_171[11:0] ? image_2392 : _GEN_17819; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17821 = 12'h959 == _T_171[11:0] ? image_2393 : _GEN_17820; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17822 = 12'h95a == _T_171[11:0] ? image_2394 : _GEN_17821; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17823 = 12'h95b == _T_171[11:0] ? image_2395 : _GEN_17822; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17824 = 12'h95c == _T_171[11:0] ? image_2396 : _GEN_17823; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17825 = 12'h95d == _T_171[11:0] ? image_2397 : _GEN_17824; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17826 = 12'h95e == _T_171[11:0] ? image_2398 : _GEN_17825; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17827 = 12'h95f == _T_171[11:0] ? image_2399 : _GEN_17826; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17828 = 12'h960 == _T_171[11:0] ? image_2400 : _GEN_17827; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17829 = 12'h961 == _T_171[11:0] ? image_2401 : _GEN_17828; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17830 = 12'h962 == _T_171[11:0] ? image_2402 : _GEN_17829; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17831 = 12'h963 == _T_171[11:0] ? image_2403 : _GEN_17830; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17832 = 12'h964 == _T_171[11:0] ? image_2404 : _GEN_17831; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17833 = 12'h965 == _T_171[11:0] ? image_2405 : _GEN_17832; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17834 = 12'h966 == _T_171[11:0] ? image_2406 : _GEN_17833; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17835 = 12'h967 == _T_171[11:0] ? image_2407 : _GEN_17834; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17836 = 12'h968 == _T_171[11:0] ? image_2408 : _GEN_17835; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17837 = 12'h969 == _T_171[11:0] ? image_2409 : _GEN_17836; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17838 = 12'h96a == _T_171[11:0] ? image_2410 : _GEN_17837; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17839 = 12'h96b == _T_171[11:0] ? image_2411 : _GEN_17838; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17840 = 12'h96c == _T_171[11:0] ? image_2412 : _GEN_17839; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17841 = 12'h96d == _T_171[11:0] ? image_2413 : _GEN_17840; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17842 = 12'h96e == _T_171[11:0] ? image_2414 : _GEN_17841; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17843 = 12'h96f == _T_171[11:0] ? image_2415 : _GEN_17842; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17844 = 12'h970 == _T_171[11:0] ? image_2416 : _GEN_17843; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17845 = 12'h971 == _T_171[11:0] ? image_2417 : _GEN_17844; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17846 = 12'h972 == _T_171[11:0] ? image_2418 : _GEN_17845; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17847 = 12'h973 == _T_171[11:0] ? image_2419 : _GEN_17846; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17848 = 12'h974 == _T_171[11:0] ? image_2420 : _GEN_17847; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17849 = 12'h975 == _T_171[11:0] ? image_2421 : _GEN_17848; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17850 = 12'h976 == _T_171[11:0] ? image_2422 : _GEN_17849; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17851 = 12'h977 == _T_171[11:0] ? image_2423 : _GEN_17850; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17852 = 12'h978 == _T_171[11:0] ? image_2424 : _GEN_17851; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17853 = 12'h979 == _T_171[11:0] ? image_2425 : _GEN_17852; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17854 = 12'h97a == _T_171[11:0] ? image_2426 : _GEN_17853; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17855 = 12'h97b == _T_171[11:0] ? 4'h0 : _GEN_17854; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17856 = 12'h97c == _T_171[11:0] ? 4'h0 : _GEN_17855; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17857 = 12'h97d == _T_171[11:0] ? 4'h0 : _GEN_17856; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17858 = 12'h97e == _T_171[11:0] ? 4'h0 : _GEN_17857; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17859 = 12'h97f == _T_171[11:0] ? 4'h0 : _GEN_17858; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17860 = 12'h980 == _T_171[11:0] ? 4'h0 : _GEN_17859; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17861 = 12'h981 == _T_171[11:0] ? 4'h0 : _GEN_17860; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17862 = 12'h982 == _T_171[11:0] ? 4'h0 : _GEN_17861; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17863 = 12'h983 == _T_171[11:0] ? 4'h0 : _GEN_17862; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17864 = 12'h984 == _T_171[11:0] ? 4'h0 : _GEN_17863; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17865 = 12'h985 == _T_171[11:0] ? image_2437 : _GEN_17864; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17866 = 12'h986 == _T_171[11:0] ? image_2438 : _GEN_17865; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17867 = 12'h987 == _T_171[11:0] ? image_2439 : _GEN_17866; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17868 = 12'h988 == _T_171[11:0] ? image_2440 : _GEN_17867; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17869 = 12'h989 == _T_171[11:0] ? image_2441 : _GEN_17868; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17870 = 12'h98a == _T_171[11:0] ? image_2442 : _GEN_17869; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17871 = 12'h98b == _T_171[11:0] ? image_2443 : _GEN_17870; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17872 = 12'h98c == _T_171[11:0] ? image_2444 : _GEN_17871; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17873 = 12'h98d == _T_171[11:0] ? image_2445 : _GEN_17872; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17874 = 12'h98e == _T_171[11:0] ? image_2446 : _GEN_17873; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17875 = 12'h98f == _T_171[11:0] ? image_2447 : _GEN_17874; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17876 = 12'h990 == _T_171[11:0] ? image_2448 : _GEN_17875; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17877 = 12'h991 == _T_171[11:0] ? image_2449 : _GEN_17876; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17878 = 12'h992 == _T_171[11:0] ? image_2450 : _GEN_17877; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17879 = 12'h993 == _T_171[11:0] ? image_2451 : _GEN_17878; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17880 = 12'h994 == _T_171[11:0] ? image_2452 : _GEN_17879; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17881 = 12'h995 == _T_171[11:0] ? image_2453 : _GEN_17880; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17882 = 12'h996 == _T_171[11:0] ? image_2454 : _GEN_17881; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17883 = 12'h997 == _T_171[11:0] ? image_2455 : _GEN_17882; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17884 = 12'h998 == _T_171[11:0] ? image_2456 : _GEN_17883; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17885 = 12'h999 == _T_171[11:0] ? image_2457 : _GEN_17884; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17886 = 12'h99a == _T_171[11:0] ? image_2458 : _GEN_17885; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17887 = 12'h99b == _T_171[11:0] ? image_2459 : _GEN_17886; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17888 = 12'h99c == _T_171[11:0] ? image_2460 : _GEN_17887; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17889 = 12'h99d == _T_171[11:0] ? image_2461 : _GEN_17888; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17890 = 12'h99e == _T_171[11:0] ? image_2462 : _GEN_17889; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17891 = 12'h99f == _T_171[11:0] ? image_2463 : _GEN_17890; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17892 = 12'h9a0 == _T_171[11:0] ? image_2464 : _GEN_17891; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17893 = 12'h9a1 == _T_171[11:0] ? image_2465 : _GEN_17892; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17894 = 12'h9a2 == _T_171[11:0] ? image_2466 : _GEN_17893; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17895 = 12'h9a3 == _T_171[11:0] ? image_2467 : _GEN_17894; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17896 = 12'h9a4 == _T_171[11:0] ? image_2468 : _GEN_17895; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17897 = 12'h9a5 == _T_171[11:0] ? image_2469 : _GEN_17896; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17898 = 12'h9a6 == _T_171[11:0] ? image_2470 : _GEN_17897; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17899 = 12'h9a7 == _T_171[11:0] ? image_2471 : _GEN_17898; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17900 = 12'h9a8 == _T_171[11:0] ? image_2472 : _GEN_17899; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17901 = 12'h9a9 == _T_171[11:0] ? image_2473 : _GEN_17900; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17902 = 12'h9aa == _T_171[11:0] ? image_2474 : _GEN_17901; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17903 = 12'h9ab == _T_171[11:0] ? image_2475 : _GEN_17902; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17904 = 12'h9ac == _T_171[11:0] ? image_2476 : _GEN_17903; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17905 = 12'h9ad == _T_171[11:0] ? image_2477 : _GEN_17904; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17906 = 12'h9ae == _T_171[11:0] ? image_2478 : _GEN_17905; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17907 = 12'h9af == _T_171[11:0] ? image_2479 : _GEN_17906; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17908 = 12'h9b0 == _T_171[11:0] ? image_2480 : _GEN_17907; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17909 = 12'h9b1 == _T_171[11:0] ? image_2481 : _GEN_17908; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17910 = 12'h9b2 == _T_171[11:0] ? image_2482 : _GEN_17909; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17911 = 12'h9b3 == _T_171[11:0] ? image_2483 : _GEN_17910; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17912 = 12'h9b4 == _T_171[11:0] ? image_2484 : _GEN_17911; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17913 = 12'h9b5 == _T_171[11:0] ? image_2485 : _GEN_17912; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17914 = 12'h9b6 == _T_171[11:0] ? image_2486 : _GEN_17913; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17915 = 12'h9b7 == _T_171[11:0] ? image_2487 : _GEN_17914; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17916 = 12'h9b8 == _T_171[11:0] ? image_2488 : _GEN_17915; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17917 = 12'h9b9 == _T_171[11:0] ? image_2489 : _GEN_17916; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17918 = 12'h9ba == _T_171[11:0] ? image_2490 : _GEN_17917; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17919 = 12'h9bb == _T_171[11:0] ? 4'h0 : _GEN_17918; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17920 = 12'h9bc == _T_171[11:0] ? 4'h0 : _GEN_17919; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17921 = 12'h9bd == _T_171[11:0] ? 4'h0 : _GEN_17920; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17922 = 12'h9be == _T_171[11:0] ? 4'h0 : _GEN_17921; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17923 = 12'h9bf == _T_171[11:0] ? 4'h0 : _GEN_17922; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17924 = 12'h9c0 == _T_171[11:0] ? 4'h0 : _GEN_17923; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17925 = 12'h9c1 == _T_171[11:0] ? 4'h0 : _GEN_17924; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17926 = 12'h9c2 == _T_171[11:0] ? 4'h0 : _GEN_17925; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17927 = 12'h9c3 == _T_171[11:0] ? 4'h0 : _GEN_17926; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17928 = 12'h9c4 == _T_171[11:0] ? 4'h0 : _GEN_17927; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17929 = 12'h9c5 == _T_171[11:0] ? 4'h0 : _GEN_17928; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17930 = 12'h9c6 == _T_171[11:0] ? image_2502 : _GEN_17929; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17931 = 12'h9c7 == _T_171[11:0] ? image_2503 : _GEN_17930; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17932 = 12'h9c8 == _T_171[11:0] ? image_2504 : _GEN_17931; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17933 = 12'h9c9 == _T_171[11:0] ? image_2505 : _GEN_17932; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17934 = 12'h9ca == _T_171[11:0] ? image_2506 : _GEN_17933; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17935 = 12'h9cb == _T_171[11:0] ? image_2507 : _GEN_17934; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17936 = 12'h9cc == _T_171[11:0] ? image_2508 : _GEN_17935; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17937 = 12'h9cd == _T_171[11:0] ? image_2509 : _GEN_17936; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17938 = 12'h9ce == _T_171[11:0] ? image_2510 : _GEN_17937; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17939 = 12'h9cf == _T_171[11:0] ? image_2511 : _GEN_17938; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17940 = 12'h9d0 == _T_171[11:0] ? image_2512 : _GEN_17939; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17941 = 12'h9d1 == _T_171[11:0] ? image_2513 : _GEN_17940; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17942 = 12'h9d2 == _T_171[11:0] ? image_2514 : _GEN_17941; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17943 = 12'h9d3 == _T_171[11:0] ? image_2515 : _GEN_17942; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17944 = 12'h9d4 == _T_171[11:0] ? image_2516 : _GEN_17943; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17945 = 12'h9d5 == _T_171[11:0] ? image_2517 : _GEN_17944; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17946 = 12'h9d6 == _T_171[11:0] ? image_2518 : _GEN_17945; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17947 = 12'h9d7 == _T_171[11:0] ? image_2519 : _GEN_17946; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17948 = 12'h9d8 == _T_171[11:0] ? image_2520 : _GEN_17947; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17949 = 12'h9d9 == _T_171[11:0] ? image_2521 : _GEN_17948; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17950 = 12'h9da == _T_171[11:0] ? image_2522 : _GEN_17949; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17951 = 12'h9db == _T_171[11:0] ? image_2523 : _GEN_17950; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17952 = 12'h9dc == _T_171[11:0] ? image_2524 : _GEN_17951; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17953 = 12'h9dd == _T_171[11:0] ? image_2525 : _GEN_17952; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17954 = 12'h9de == _T_171[11:0] ? image_2526 : _GEN_17953; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17955 = 12'h9df == _T_171[11:0] ? image_2527 : _GEN_17954; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17956 = 12'h9e0 == _T_171[11:0] ? image_2528 : _GEN_17955; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17957 = 12'h9e1 == _T_171[11:0] ? image_2529 : _GEN_17956; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17958 = 12'h9e2 == _T_171[11:0] ? image_2530 : _GEN_17957; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17959 = 12'h9e3 == _T_171[11:0] ? image_2531 : _GEN_17958; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17960 = 12'h9e4 == _T_171[11:0] ? image_2532 : _GEN_17959; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17961 = 12'h9e5 == _T_171[11:0] ? image_2533 : _GEN_17960; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17962 = 12'h9e6 == _T_171[11:0] ? image_2534 : _GEN_17961; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17963 = 12'h9e7 == _T_171[11:0] ? image_2535 : _GEN_17962; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17964 = 12'h9e8 == _T_171[11:0] ? image_2536 : _GEN_17963; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17965 = 12'h9e9 == _T_171[11:0] ? image_2537 : _GEN_17964; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17966 = 12'h9ea == _T_171[11:0] ? image_2538 : _GEN_17965; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17967 = 12'h9eb == _T_171[11:0] ? image_2539 : _GEN_17966; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17968 = 12'h9ec == _T_171[11:0] ? image_2540 : _GEN_17967; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17969 = 12'h9ed == _T_171[11:0] ? image_2541 : _GEN_17968; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17970 = 12'h9ee == _T_171[11:0] ? image_2542 : _GEN_17969; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17971 = 12'h9ef == _T_171[11:0] ? image_2543 : _GEN_17970; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17972 = 12'h9f0 == _T_171[11:0] ? image_2544 : _GEN_17971; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17973 = 12'h9f1 == _T_171[11:0] ? image_2545 : _GEN_17972; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17974 = 12'h9f2 == _T_171[11:0] ? image_2546 : _GEN_17973; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17975 = 12'h9f3 == _T_171[11:0] ? image_2547 : _GEN_17974; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17976 = 12'h9f4 == _T_171[11:0] ? image_2548 : _GEN_17975; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17977 = 12'h9f5 == _T_171[11:0] ? image_2549 : _GEN_17976; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17978 = 12'h9f6 == _T_171[11:0] ? image_2550 : _GEN_17977; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17979 = 12'h9f7 == _T_171[11:0] ? image_2551 : _GEN_17978; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17980 = 12'h9f8 == _T_171[11:0] ? image_2552 : _GEN_17979; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17981 = 12'h9f9 == _T_171[11:0] ? image_2553 : _GEN_17980; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17982 = 12'h9fa == _T_171[11:0] ? image_2554 : _GEN_17981; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17983 = 12'h9fb == _T_171[11:0] ? 4'h0 : _GEN_17982; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17984 = 12'h9fc == _T_171[11:0] ? 4'h0 : _GEN_17983; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17985 = 12'h9fd == _T_171[11:0] ? 4'h0 : _GEN_17984; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17986 = 12'h9fe == _T_171[11:0] ? 4'h0 : _GEN_17985; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17987 = 12'h9ff == _T_171[11:0] ? 4'h0 : _GEN_17986; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17988 = 12'ha00 == _T_171[11:0] ? 4'h0 : _GEN_17987; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17989 = 12'ha01 == _T_171[11:0] ? 4'h0 : _GEN_17988; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17990 = 12'ha02 == _T_171[11:0] ? 4'h0 : _GEN_17989; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17991 = 12'ha03 == _T_171[11:0] ? 4'h0 : _GEN_17990; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17992 = 12'ha04 == _T_171[11:0] ? 4'h0 : _GEN_17991; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17993 = 12'ha05 == _T_171[11:0] ? 4'h0 : _GEN_17992; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17994 = 12'ha06 == _T_171[11:0] ? 4'h0 : _GEN_17993; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17995 = 12'ha07 == _T_171[11:0] ? image_2567 : _GEN_17994; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17996 = 12'ha08 == _T_171[11:0] ? image_2568 : _GEN_17995; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17997 = 12'ha09 == _T_171[11:0] ? image_2569 : _GEN_17996; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17998 = 12'ha0a == _T_171[11:0] ? image_2570 : _GEN_17997; // @[Filter.scala 138:46]
  wire [3:0] _GEN_17999 = 12'ha0b == _T_171[11:0] ? image_2571 : _GEN_17998; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18000 = 12'ha0c == _T_171[11:0] ? image_2572 : _GEN_17999; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18001 = 12'ha0d == _T_171[11:0] ? image_2573 : _GEN_18000; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18002 = 12'ha0e == _T_171[11:0] ? image_2574 : _GEN_18001; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18003 = 12'ha0f == _T_171[11:0] ? image_2575 : _GEN_18002; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18004 = 12'ha10 == _T_171[11:0] ? image_2576 : _GEN_18003; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18005 = 12'ha11 == _T_171[11:0] ? image_2577 : _GEN_18004; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18006 = 12'ha12 == _T_171[11:0] ? image_2578 : _GEN_18005; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18007 = 12'ha13 == _T_171[11:0] ? image_2579 : _GEN_18006; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18008 = 12'ha14 == _T_171[11:0] ? image_2580 : _GEN_18007; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18009 = 12'ha15 == _T_171[11:0] ? image_2581 : _GEN_18008; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18010 = 12'ha16 == _T_171[11:0] ? image_2582 : _GEN_18009; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18011 = 12'ha17 == _T_171[11:0] ? image_2583 : _GEN_18010; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18012 = 12'ha18 == _T_171[11:0] ? image_2584 : _GEN_18011; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18013 = 12'ha19 == _T_171[11:0] ? image_2585 : _GEN_18012; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18014 = 12'ha1a == _T_171[11:0] ? image_2586 : _GEN_18013; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18015 = 12'ha1b == _T_171[11:0] ? image_2587 : _GEN_18014; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18016 = 12'ha1c == _T_171[11:0] ? image_2588 : _GEN_18015; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18017 = 12'ha1d == _T_171[11:0] ? image_2589 : _GEN_18016; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18018 = 12'ha1e == _T_171[11:0] ? image_2590 : _GEN_18017; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18019 = 12'ha1f == _T_171[11:0] ? image_2591 : _GEN_18018; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18020 = 12'ha20 == _T_171[11:0] ? image_2592 : _GEN_18019; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18021 = 12'ha21 == _T_171[11:0] ? image_2593 : _GEN_18020; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18022 = 12'ha22 == _T_171[11:0] ? image_2594 : _GEN_18021; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18023 = 12'ha23 == _T_171[11:0] ? image_2595 : _GEN_18022; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18024 = 12'ha24 == _T_171[11:0] ? image_2596 : _GEN_18023; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18025 = 12'ha25 == _T_171[11:0] ? image_2597 : _GEN_18024; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18026 = 12'ha26 == _T_171[11:0] ? image_2598 : _GEN_18025; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18027 = 12'ha27 == _T_171[11:0] ? image_2599 : _GEN_18026; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18028 = 12'ha28 == _T_171[11:0] ? image_2600 : _GEN_18027; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18029 = 12'ha29 == _T_171[11:0] ? image_2601 : _GEN_18028; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18030 = 12'ha2a == _T_171[11:0] ? image_2602 : _GEN_18029; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18031 = 12'ha2b == _T_171[11:0] ? image_2603 : _GEN_18030; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18032 = 12'ha2c == _T_171[11:0] ? image_2604 : _GEN_18031; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18033 = 12'ha2d == _T_171[11:0] ? image_2605 : _GEN_18032; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18034 = 12'ha2e == _T_171[11:0] ? image_2606 : _GEN_18033; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18035 = 12'ha2f == _T_171[11:0] ? image_2607 : _GEN_18034; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18036 = 12'ha30 == _T_171[11:0] ? image_2608 : _GEN_18035; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18037 = 12'ha31 == _T_171[11:0] ? image_2609 : _GEN_18036; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18038 = 12'ha32 == _T_171[11:0] ? image_2610 : _GEN_18037; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18039 = 12'ha33 == _T_171[11:0] ? image_2611 : _GEN_18038; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18040 = 12'ha34 == _T_171[11:0] ? image_2612 : _GEN_18039; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18041 = 12'ha35 == _T_171[11:0] ? image_2613 : _GEN_18040; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18042 = 12'ha36 == _T_171[11:0] ? image_2614 : _GEN_18041; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18043 = 12'ha37 == _T_171[11:0] ? image_2615 : _GEN_18042; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18044 = 12'ha38 == _T_171[11:0] ? image_2616 : _GEN_18043; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18045 = 12'ha39 == _T_171[11:0] ? image_2617 : _GEN_18044; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18046 = 12'ha3a == _T_171[11:0] ? image_2618 : _GEN_18045; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18047 = 12'ha3b == _T_171[11:0] ? 4'h0 : _GEN_18046; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18048 = 12'ha3c == _T_171[11:0] ? 4'h0 : _GEN_18047; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18049 = 12'ha3d == _T_171[11:0] ? 4'h0 : _GEN_18048; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18050 = 12'ha3e == _T_171[11:0] ? 4'h0 : _GEN_18049; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18051 = 12'ha3f == _T_171[11:0] ? 4'h0 : _GEN_18050; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18052 = 12'ha40 == _T_171[11:0] ? 4'h0 : _GEN_18051; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18053 = 12'ha41 == _T_171[11:0] ? 4'h0 : _GEN_18052; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18054 = 12'ha42 == _T_171[11:0] ? 4'h0 : _GEN_18053; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18055 = 12'ha43 == _T_171[11:0] ? 4'h0 : _GEN_18054; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18056 = 12'ha44 == _T_171[11:0] ? 4'h0 : _GEN_18055; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18057 = 12'ha45 == _T_171[11:0] ? 4'h0 : _GEN_18056; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18058 = 12'ha46 == _T_171[11:0] ? 4'h0 : _GEN_18057; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18059 = 12'ha47 == _T_171[11:0] ? 4'h0 : _GEN_18058; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18060 = 12'ha48 == _T_171[11:0] ? image_2632 : _GEN_18059; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18061 = 12'ha49 == _T_171[11:0] ? image_2633 : _GEN_18060; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18062 = 12'ha4a == _T_171[11:0] ? image_2634 : _GEN_18061; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18063 = 12'ha4b == _T_171[11:0] ? image_2635 : _GEN_18062; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18064 = 12'ha4c == _T_171[11:0] ? image_2636 : _GEN_18063; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18065 = 12'ha4d == _T_171[11:0] ? image_2637 : _GEN_18064; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18066 = 12'ha4e == _T_171[11:0] ? image_2638 : _GEN_18065; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18067 = 12'ha4f == _T_171[11:0] ? image_2639 : _GEN_18066; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18068 = 12'ha50 == _T_171[11:0] ? image_2640 : _GEN_18067; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18069 = 12'ha51 == _T_171[11:0] ? image_2641 : _GEN_18068; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18070 = 12'ha52 == _T_171[11:0] ? image_2642 : _GEN_18069; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18071 = 12'ha53 == _T_171[11:0] ? image_2643 : _GEN_18070; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18072 = 12'ha54 == _T_171[11:0] ? image_2644 : _GEN_18071; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18073 = 12'ha55 == _T_171[11:0] ? image_2645 : _GEN_18072; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18074 = 12'ha56 == _T_171[11:0] ? image_2646 : _GEN_18073; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18075 = 12'ha57 == _T_171[11:0] ? image_2647 : _GEN_18074; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18076 = 12'ha58 == _T_171[11:0] ? image_2648 : _GEN_18075; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18077 = 12'ha59 == _T_171[11:0] ? image_2649 : _GEN_18076; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18078 = 12'ha5a == _T_171[11:0] ? image_2650 : _GEN_18077; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18079 = 12'ha5b == _T_171[11:0] ? image_2651 : _GEN_18078; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18080 = 12'ha5c == _T_171[11:0] ? image_2652 : _GEN_18079; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18081 = 12'ha5d == _T_171[11:0] ? image_2653 : _GEN_18080; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18082 = 12'ha5e == _T_171[11:0] ? image_2654 : _GEN_18081; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18083 = 12'ha5f == _T_171[11:0] ? image_2655 : _GEN_18082; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18084 = 12'ha60 == _T_171[11:0] ? image_2656 : _GEN_18083; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18085 = 12'ha61 == _T_171[11:0] ? image_2657 : _GEN_18084; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18086 = 12'ha62 == _T_171[11:0] ? image_2658 : _GEN_18085; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18087 = 12'ha63 == _T_171[11:0] ? image_2659 : _GEN_18086; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18088 = 12'ha64 == _T_171[11:0] ? image_2660 : _GEN_18087; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18089 = 12'ha65 == _T_171[11:0] ? image_2661 : _GEN_18088; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18090 = 12'ha66 == _T_171[11:0] ? image_2662 : _GEN_18089; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18091 = 12'ha67 == _T_171[11:0] ? image_2663 : _GEN_18090; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18092 = 12'ha68 == _T_171[11:0] ? image_2664 : _GEN_18091; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18093 = 12'ha69 == _T_171[11:0] ? image_2665 : _GEN_18092; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18094 = 12'ha6a == _T_171[11:0] ? image_2666 : _GEN_18093; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18095 = 12'ha6b == _T_171[11:0] ? image_2667 : _GEN_18094; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18096 = 12'ha6c == _T_171[11:0] ? image_2668 : _GEN_18095; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18097 = 12'ha6d == _T_171[11:0] ? image_2669 : _GEN_18096; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18098 = 12'ha6e == _T_171[11:0] ? image_2670 : _GEN_18097; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18099 = 12'ha6f == _T_171[11:0] ? image_2671 : _GEN_18098; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18100 = 12'ha70 == _T_171[11:0] ? image_2672 : _GEN_18099; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18101 = 12'ha71 == _T_171[11:0] ? image_2673 : _GEN_18100; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18102 = 12'ha72 == _T_171[11:0] ? image_2674 : _GEN_18101; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18103 = 12'ha73 == _T_171[11:0] ? image_2675 : _GEN_18102; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18104 = 12'ha74 == _T_171[11:0] ? image_2676 : _GEN_18103; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18105 = 12'ha75 == _T_171[11:0] ? image_2677 : _GEN_18104; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18106 = 12'ha76 == _T_171[11:0] ? image_2678 : _GEN_18105; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18107 = 12'ha77 == _T_171[11:0] ? image_2679 : _GEN_18106; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18108 = 12'ha78 == _T_171[11:0] ? image_2680 : _GEN_18107; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18109 = 12'ha79 == _T_171[11:0] ? image_2681 : _GEN_18108; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18110 = 12'ha7a == _T_171[11:0] ? image_2682 : _GEN_18109; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18111 = 12'ha7b == _T_171[11:0] ? 4'h0 : _GEN_18110; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18112 = 12'ha7c == _T_171[11:0] ? 4'h0 : _GEN_18111; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18113 = 12'ha7d == _T_171[11:0] ? 4'h0 : _GEN_18112; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18114 = 12'ha7e == _T_171[11:0] ? 4'h0 : _GEN_18113; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18115 = 12'ha7f == _T_171[11:0] ? 4'h0 : _GEN_18114; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18116 = 12'ha80 == _T_171[11:0] ? 4'h0 : _GEN_18115; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18117 = 12'ha81 == _T_171[11:0] ? 4'h0 : _GEN_18116; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18118 = 12'ha82 == _T_171[11:0] ? 4'h0 : _GEN_18117; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18119 = 12'ha83 == _T_171[11:0] ? 4'h0 : _GEN_18118; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18120 = 12'ha84 == _T_171[11:0] ? 4'h0 : _GEN_18119; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18121 = 12'ha85 == _T_171[11:0] ? 4'h0 : _GEN_18120; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18122 = 12'ha86 == _T_171[11:0] ? 4'h0 : _GEN_18121; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18123 = 12'ha87 == _T_171[11:0] ? 4'h0 : _GEN_18122; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18124 = 12'ha88 == _T_171[11:0] ? 4'h0 : _GEN_18123; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18125 = 12'ha89 == _T_171[11:0] ? image_2697 : _GEN_18124; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18126 = 12'ha8a == _T_171[11:0] ? image_2698 : _GEN_18125; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18127 = 12'ha8b == _T_171[11:0] ? image_2699 : _GEN_18126; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18128 = 12'ha8c == _T_171[11:0] ? image_2700 : _GEN_18127; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18129 = 12'ha8d == _T_171[11:0] ? image_2701 : _GEN_18128; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18130 = 12'ha8e == _T_171[11:0] ? image_2702 : _GEN_18129; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18131 = 12'ha8f == _T_171[11:0] ? image_2703 : _GEN_18130; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18132 = 12'ha90 == _T_171[11:0] ? image_2704 : _GEN_18131; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18133 = 12'ha91 == _T_171[11:0] ? image_2705 : _GEN_18132; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18134 = 12'ha92 == _T_171[11:0] ? image_2706 : _GEN_18133; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18135 = 12'ha93 == _T_171[11:0] ? image_2707 : _GEN_18134; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18136 = 12'ha94 == _T_171[11:0] ? image_2708 : _GEN_18135; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18137 = 12'ha95 == _T_171[11:0] ? image_2709 : _GEN_18136; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18138 = 12'ha96 == _T_171[11:0] ? image_2710 : _GEN_18137; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18139 = 12'ha97 == _T_171[11:0] ? image_2711 : _GEN_18138; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18140 = 12'ha98 == _T_171[11:0] ? image_2712 : _GEN_18139; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18141 = 12'ha99 == _T_171[11:0] ? image_2713 : _GEN_18140; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18142 = 12'ha9a == _T_171[11:0] ? image_2714 : _GEN_18141; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18143 = 12'ha9b == _T_171[11:0] ? image_2715 : _GEN_18142; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18144 = 12'ha9c == _T_171[11:0] ? image_2716 : _GEN_18143; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18145 = 12'ha9d == _T_171[11:0] ? image_2717 : _GEN_18144; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18146 = 12'ha9e == _T_171[11:0] ? image_2718 : _GEN_18145; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18147 = 12'ha9f == _T_171[11:0] ? image_2719 : _GEN_18146; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18148 = 12'haa0 == _T_171[11:0] ? image_2720 : _GEN_18147; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18149 = 12'haa1 == _T_171[11:0] ? image_2721 : _GEN_18148; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18150 = 12'haa2 == _T_171[11:0] ? image_2722 : _GEN_18149; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18151 = 12'haa3 == _T_171[11:0] ? image_2723 : _GEN_18150; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18152 = 12'haa4 == _T_171[11:0] ? image_2724 : _GEN_18151; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18153 = 12'haa5 == _T_171[11:0] ? image_2725 : _GEN_18152; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18154 = 12'haa6 == _T_171[11:0] ? image_2726 : _GEN_18153; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18155 = 12'haa7 == _T_171[11:0] ? image_2727 : _GEN_18154; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18156 = 12'haa8 == _T_171[11:0] ? image_2728 : _GEN_18155; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18157 = 12'haa9 == _T_171[11:0] ? image_2729 : _GEN_18156; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18158 = 12'haaa == _T_171[11:0] ? image_2730 : _GEN_18157; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18159 = 12'haab == _T_171[11:0] ? image_2731 : _GEN_18158; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18160 = 12'haac == _T_171[11:0] ? image_2732 : _GEN_18159; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18161 = 12'haad == _T_171[11:0] ? image_2733 : _GEN_18160; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18162 = 12'haae == _T_171[11:0] ? image_2734 : _GEN_18161; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18163 = 12'haaf == _T_171[11:0] ? image_2735 : _GEN_18162; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18164 = 12'hab0 == _T_171[11:0] ? image_2736 : _GEN_18163; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18165 = 12'hab1 == _T_171[11:0] ? image_2737 : _GEN_18164; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18166 = 12'hab2 == _T_171[11:0] ? image_2738 : _GEN_18165; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18167 = 12'hab3 == _T_171[11:0] ? image_2739 : _GEN_18166; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18168 = 12'hab4 == _T_171[11:0] ? image_2740 : _GEN_18167; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18169 = 12'hab5 == _T_171[11:0] ? image_2741 : _GEN_18168; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18170 = 12'hab6 == _T_171[11:0] ? image_2742 : _GEN_18169; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18171 = 12'hab7 == _T_171[11:0] ? image_2743 : _GEN_18170; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18172 = 12'hab8 == _T_171[11:0] ? image_2744 : _GEN_18171; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18173 = 12'hab9 == _T_171[11:0] ? image_2745 : _GEN_18172; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18174 = 12'haba == _T_171[11:0] ? 4'h0 : _GEN_18173; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18175 = 12'habb == _T_171[11:0] ? 4'h0 : _GEN_18174; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18176 = 12'habc == _T_171[11:0] ? 4'h0 : _GEN_18175; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18177 = 12'habd == _T_171[11:0] ? 4'h0 : _GEN_18176; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18178 = 12'habe == _T_171[11:0] ? 4'h0 : _GEN_18177; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18179 = 12'habf == _T_171[11:0] ? 4'h0 : _GEN_18178; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18180 = 12'hac0 == _T_171[11:0] ? 4'h0 : _GEN_18179; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18181 = 12'hac1 == _T_171[11:0] ? 4'h0 : _GEN_18180; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18182 = 12'hac2 == _T_171[11:0] ? 4'h0 : _GEN_18181; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18183 = 12'hac3 == _T_171[11:0] ? 4'h0 : _GEN_18182; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18184 = 12'hac4 == _T_171[11:0] ? 4'h0 : _GEN_18183; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18185 = 12'hac5 == _T_171[11:0] ? 4'h0 : _GEN_18184; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18186 = 12'hac6 == _T_171[11:0] ? 4'h0 : _GEN_18185; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18187 = 12'hac7 == _T_171[11:0] ? 4'h0 : _GEN_18186; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18188 = 12'hac8 == _T_171[11:0] ? 4'h0 : _GEN_18187; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18189 = 12'hac9 == _T_171[11:0] ? 4'h0 : _GEN_18188; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18190 = 12'haca == _T_171[11:0] ? 4'h0 : _GEN_18189; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18191 = 12'hacb == _T_171[11:0] ? image_2763 : _GEN_18190; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18192 = 12'hacc == _T_171[11:0] ? image_2764 : _GEN_18191; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18193 = 12'hacd == _T_171[11:0] ? image_2765 : _GEN_18192; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18194 = 12'hace == _T_171[11:0] ? image_2766 : _GEN_18193; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18195 = 12'hacf == _T_171[11:0] ? image_2767 : _GEN_18194; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18196 = 12'had0 == _T_171[11:0] ? image_2768 : _GEN_18195; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18197 = 12'had1 == _T_171[11:0] ? image_2769 : _GEN_18196; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18198 = 12'had2 == _T_171[11:0] ? image_2770 : _GEN_18197; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18199 = 12'had3 == _T_171[11:0] ? image_2771 : _GEN_18198; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18200 = 12'had4 == _T_171[11:0] ? image_2772 : _GEN_18199; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18201 = 12'had5 == _T_171[11:0] ? image_2773 : _GEN_18200; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18202 = 12'had6 == _T_171[11:0] ? image_2774 : _GEN_18201; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18203 = 12'had7 == _T_171[11:0] ? image_2775 : _GEN_18202; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18204 = 12'had8 == _T_171[11:0] ? image_2776 : _GEN_18203; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18205 = 12'had9 == _T_171[11:0] ? image_2777 : _GEN_18204; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18206 = 12'hada == _T_171[11:0] ? image_2778 : _GEN_18205; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18207 = 12'hadb == _T_171[11:0] ? image_2779 : _GEN_18206; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18208 = 12'hadc == _T_171[11:0] ? image_2780 : _GEN_18207; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18209 = 12'hadd == _T_171[11:0] ? image_2781 : _GEN_18208; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18210 = 12'hade == _T_171[11:0] ? image_2782 : _GEN_18209; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18211 = 12'hadf == _T_171[11:0] ? image_2783 : _GEN_18210; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18212 = 12'hae0 == _T_171[11:0] ? image_2784 : _GEN_18211; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18213 = 12'hae1 == _T_171[11:0] ? image_2785 : _GEN_18212; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18214 = 12'hae2 == _T_171[11:0] ? image_2786 : _GEN_18213; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18215 = 12'hae3 == _T_171[11:0] ? image_2787 : _GEN_18214; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18216 = 12'hae4 == _T_171[11:0] ? image_2788 : _GEN_18215; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18217 = 12'hae5 == _T_171[11:0] ? image_2789 : _GEN_18216; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18218 = 12'hae6 == _T_171[11:0] ? image_2790 : _GEN_18217; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18219 = 12'hae7 == _T_171[11:0] ? image_2791 : _GEN_18218; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18220 = 12'hae8 == _T_171[11:0] ? image_2792 : _GEN_18219; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18221 = 12'hae9 == _T_171[11:0] ? image_2793 : _GEN_18220; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18222 = 12'haea == _T_171[11:0] ? image_2794 : _GEN_18221; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18223 = 12'haeb == _T_171[11:0] ? image_2795 : _GEN_18222; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18224 = 12'haec == _T_171[11:0] ? image_2796 : _GEN_18223; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18225 = 12'haed == _T_171[11:0] ? image_2797 : _GEN_18224; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18226 = 12'haee == _T_171[11:0] ? image_2798 : _GEN_18225; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18227 = 12'haef == _T_171[11:0] ? image_2799 : _GEN_18226; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18228 = 12'haf0 == _T_171[11:0] ? image_2800 : _GEN_18227; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18229 = 12'haf1 == _T_171[11:0] ? image_2801 : _GEN_18228; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18230 = 12'haf2 == _T_171[11:0] ? image_2802 : _GEN_18229; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18231 = 12'haf3 == _T_171[11:0] ? image_2803 : _GEN_18230; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18232 = 12'haf4 == _T_171[11:0] ? image_2804 : _GEN_18231; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18233 = 12'haf5 == _T_171[11:0] ? image_2805 : _GEN_18232; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18234 = 12'haf6 == _T_171[11:0] ? image_2806 : _GEN_18233; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18235 = 12'haf7 == _T_171[11:0] ? image_2807 : _GEN_18234; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18236 = 12'haf8 == _T_171[11:0] ? image_2808 : _GEN_18235; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18237 = 12'haf9 == _T_171[11:0] ? 4'h0 : _GEN_18236; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18238 = 12'hafa == _T_171[11:0] ? 4'h0 : _GEN_18237; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18239 = 12'hafb == _T_171[11:0] ? 4'h0 : _GEN_18238; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18240 = 12'hafc == _T_171[11:0] ? 4'h0 : _GEN_18239; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18241 = 12'hafd == _T_171[11:0] ? 4'h0 : _GEN_18240; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18242 = 12'hafe == _T_171[11:0] ? 4'h0 : _GEN_18241; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18243 = 12'haff == _T_171[11:0] ? 4'h0 : _GEN_18242; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18244 = 12'hb00 == _T_171[11:0] ? 4'h0 : _GEN_18243; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18245 = 12'hb01 == _T_171[11:0] ? 4'h0 : _GEN_18244; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18246 = 12'hb02 == _T_171[11:0] ? 4'h0 : _GEN_18245; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18247 = 12'hb03 == _T_171[11:0] ? 4'h0 : _GEN_18246; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18248 = 12'hb04 == _T_171[11:0] ? 4'h0 : _GEN_18247; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18249 = 12'hb05 == _T_171[11:0] ? 4'h0 : _GEN_18248; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18250 = 12'hb06 == _T_171[11:0] ? 4'h0 : _GEN_18249; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18251 = 12'hb07 == _T_171[11:0] ? 4'h0 : _GEN_18250; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18252 = 12'hb08 == _T_171[11:0] ? 4'h0 : _GEN_18251; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18253 = 12'hb09 == _T_171[11:0] ? 4'h0 : _GEN_18252; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18254 = 12'hb0a == _T_171[11:0] ? 4'h0 : _GEN_18253; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18255 = 12'hb0b == _T_171[11:0] ? 4'h0 : _GEN_18254; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18256 = 12'hb0c == _T_171[11:0] ? image_2828 : _GEN_18255; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18257 = 12'hb0d == _T_171[11:0] ? image_2829 : _GEN_18256; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18258 = 12'hb0e == _T_171[11:0] ? image_2830 : _GEN_18257; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18259 = 12'hb0f == _T_171[11:0] ? image_2831 : _GEN_18258; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18260 = 12'hb10 == _T_171[11:0] ? image_2832 : _GEN_18259; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18261 = 12'hb11 == _T_171[11:0] ? image_2833 : _GEN_18260; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18262 = 12'hb12 == _T_171[11:0] ? image_2834 : _GEN_18261; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18263 = 12'hb13 == _T_171[11:0] ? image_2835 : _GEN_18262; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18264 = 12'hb14 == _T_171[11:0] ? image_2836 : _GEN_18263; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18265 = 12'hb15 == _T_171[11:0] ? image_2837 : _GEN_18264; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18266 = 12'hb16 == _T_171[11:0] ? image_2838 : _GEN_18265; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18267 = 12'hb17 == _T_171[11:0] ? image_2839 : _GEN_18266; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18268 = 12'hb18 == _T_171[11:0] ? image_2840 : _GEN_18267; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18269 = 12'hb19 == _T_171[11:0] ? image_2841 : _GEN_18268; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18270 = 12'hb1a == _T_171[11:0] ? image_2842 : _GEN_18269; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18271 = 12'hb1b == _T_171[11:0] ? image_2843 : _GEN_18270; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18272 = 12'hb1c == _T_171[11:0] ? image_2844 : _GEN_18271; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18273 = 12'hb1d == _T_171[11:0] ? image_2845 : _GEN_18272; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18274 = 12'hb1e == _T_171[11:0] ? image_2846 : _GEN_18273; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18275 = 12'hb1f == _T_171[11:0] ? image_2847 : _GEN_18274; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18276 = 12'hb20 == _T_171[11:0] ? image_2848 : _GEN_18275; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18277 = 12'hb21 == _T_171[11:0] ? image_2849 : _GEN_18276; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18278 = 12'hb22 == _T_171[11:0] ? image_2850 : _GEN_18277; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18279 = 12'hb23 == _T_171[11:0] ? image_2851 : _GEN_18278; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18280 = 12'hb24 == _T_171[11:0] ? image_2852 : _GEN_18279; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18281 = 12'hb25 == _T_171[11:0] ? image_2853 : _GEN_18280; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18282 = 12'hb26 == _T_171[11:0] ? image_2854 : _GEN_18281; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18283 = 12'hb27 == _T_171[11:0] ? image_2855 : _GEN_18282; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18284 = 12'hb28 == _T_171[11:0] ? image_2856 : _GEN_18283; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18285 = 12'hb29 == _T_171[11:0] ? image_2857 : _GEN_18284; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18286 = 12'hb2a == _T_171[11:0] ? image_2858 : _GEN_18285; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18287 = 12'hb2b == _T_171[11:0] ? image_2859 : _GEN_18286; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18288 = 12'hb2c == _T_171[11:0] ? image_2860 : _GEN_18287; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18289 = 12'hb2d == _T_171[11:0] ? image_2861 : _GEN_18288; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18290 = 12'hb2e == _T_171[11:0] ? image_2862 : _GEN_18289; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18291 = 12'hb2f == _T_171[11:0] ? image_2863 : _GEN_18290; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18292 = 12'hb30 == _T_171[11:0] ? image_2864 : _GEN_18291; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18293 = 12'hb31 == _T_171[11:0] ? image_2865 : _GEN_18292; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18294 = 12'hb32 == _T_171[11:0] ? image_2866 : _GEN_18293; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18295 = 12'hb33 == _T_171[11:0] ? image_2867 : _GEN_18294; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18296 = 12'hb34 == _T_171[11:0] ? image_2868 : _GEN_18295; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18297 = 12'hb35 == _T_171[11:0] ? image_2869 : _GEN_18296; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18298 = 12'hb36 == _T_171[11:0] ? image_2870 : _GEN_18297; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18299 = 12'hb37 == _T_171[11:0] ? image_2871 : _GEN_18298; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18300 = 12'hb38 == _T_171[11:0] ? 4'h0 : _GEN_18299; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18301 = 12'hb39 == _T_171[11:0] ? 4'h0 : _GEN_18300; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18302 = 12'hb3a == _T_171[11:0] ? 4'h0 : _GEN_18301; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18303 = 12'hb3b == _T_171[11:0] ? 4'h0 : _GEN_18302; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18304 = 12'hb3c == _T_171[11:0] ? 4'h0 : _GEN_18303; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18305 = 12'hb3d == _T_171[11:0] ? 4'h0 : _GEN_18304; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18306 = 12'hb3e == _T_171[11:0] ? 4'h0 : _GEN_18305; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18307 = 12'hb3f == _T_171[11:0] ? 4'h0 : _GEN_18306; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18308 = 12'hb40 == _T_171[11:0] ? 4'h0 : _GEN_18307; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18309 = 12'hb41 == _T_171[11:0] ? 4'h0 : _GEN_18308; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18310 = 12'hb42 == _T_171[11:0] ? 4'h0 : _GEN_18309; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18311 = 12'hb43 == _T_171[11:0] ? 4'h0 : _GEN_18310; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18312 = 12'hb44 == _T_171[11:0] ? 4'h0 : _GEN_18311; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18313 = 12'hb45 == _T_171[11:0] ? 4'h0 : _GEN_18312; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18314 = 12'hb46 == _T_171[11:0] ? 4'h0 : _GEN_18313; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18315 = 12'hb47 == _T_171[11:0] ? 4'h0 : _GEN_18314; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18316 = 12'hb48 == _T_171[11:0] ? 4'h0 : _GEN_18315; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18317 = 12'hb49 == _T_171[11:0] ? 4'h0 : _GEN_18316; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18318 = 12'hb4a == _T_171[11:0] ? 4'h0 : _GEN_18317; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18319 = 12'hb4b == _T_171[11:0] ? 4'h0 : _GEN_18318; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18320 = 12'hb4c == _T_171[11:0] ? 4'h0 : _GEN_18319; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18321 = 12'hb4d == _T_171[11:0] ? 4'h0 : _GEN_18320; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18322 = 12'hb4e == _T_171[11:0] ? 4'h0 : _GEN_18321; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18323 = 12'hb4f == _T_171[11:0] ? image_2895 : _GEN_18322; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18324 = 12'hb50 == _T_171[11:0] ? image_2896 : _GEN_18323; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18325 = 12'hb51 == _T_171[11:0] ? image_2897 : _GEN_18324; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18326 = 12'hb52 == _T_171[11:0] ? image_2898 : _GEN_18325; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18327 = 12'hb53 == _T_171[11:0] ? image_2899 : _GEN_18326; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18328 = 12'hb54 == _T_171[11:0] ? image_2900 : _GEN_18327; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18329 = 12'hb55 == _T_171[11:0] ? image_2901 : _GEN_18328; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18330 = 12'hb56 == _T_171[11:0] ? image_2902 : _GEN_18329; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18331 = 12'hb57 == _T_171[11:0] ? image_2903 : _GEN_18330; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18332 = 12'hb58 == _T_171[11:0] ? image_2904 : _GEN_18331; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18333 = 12'hb59 == _T_171[11:0] ? image_2905 : _GEN_18332; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18334 = 12'hb5a == _T_171[11:0] ? image_2906 : _GEN_18333; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18335 = 12'hb5b == _T_171[11:0] ? image_2907 : _GEN_18334; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18336 = 12'hb5c == _T_171[11:0] ? image_2908 : _GEN_18335; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18337 = 12'hb5d == _T_171[11:0] ? image_2909 : _GEN_18336; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18338 = 12'hb5e == _T_171[11:0] ? image_2910 : _GEN_18337; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18339 = 12'hb5f == _T_171[11:0] ? image_2911 : _GEN_18338; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18340 = 12'hb60 == _T_171[11:0] ? image_2912 : _GEN_18339; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18341 = 12'hb61 == _T_171[11:0] ? image_2913 : _GEN_18340; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18342 = 12'hb62 == _T_171[11:0] ? image_2914 : _GEN_18341; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18343 = 12'hb63 == _T_171[11:0] ? image_2915 : _GEN_18342; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18344 = 12'hb64 == _T_171[11:0] ? image_2916 : _GEN_18343; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18345 = 12'hb65 == _T_171[11:0] ? image_2917 : _GEN_18344; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18346 = 12'hb66 == _T_171[11:0] ? image_2918 : _GEN_18345; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18347 = 12'hb67 == _T_171[11:0] ? image_2919 : _GEN_18346; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18348 = 12'hb68 == _T_171[11:0] ? image_2920 : _GEN_18347; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18349 = 12'hb69 == _T_171[11:0] ? image_2921 : _GEN_18348; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18350 = 12'hb6a == _T_171[11:0] ? image_2922 : _GEN_18349; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18351 = 12'hb6b == _T_171[11:0] ? image_2923 : _GEN_18350; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18352 = 12'hb6c == _T_171[11:0] ? image_2924 : _GEN_18351; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18353 = 12'hb6d == _T_171[11:0] ? image_2925 : _GEN_18352; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18354 = 12'hb6e == _T_171[11:0] ? image_2926 : _GEN_18353; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18355 = 12'hb6f == _T_171[11:0] ? image_2927 : _GEN_18354; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18356 = 12'hb70 == _T_171[11:0] ? image_2928 : _GEN_18355; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18357 = 12'hb71 == _T_171[11:0] ? image_2929 : _GEN_18356; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18358 = 12'hb72 == _T_171[11:0] ? image_2930 : _GEN_18357; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18359 = 12'hb73 == _T_171[11:0] ? image_2931 : _GEN_18358; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18360 = 12'hb74 == _T_171[11:0] ? image_2932 : _GEN_18359; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18361 = 12'hb75 == _T_171[11:0] ? image_2933 : _GEN_18360; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18362 = 12'hb76 == _T_171[11:0] ? image_2934 : _GEN_18361; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18363 = 12'hb77 == _T_171[11:0] ? 4'h0 : _GEN_18362; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18364 = 12'hb78 == _T_171[11:0] ? 4'h0 : _GEN_18363; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18365 = 12'hb79 == _T_171[11:0] ? 4'h0 : _GEN_18364; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18366 = 12'hb7a == _T_171[11:0] ? 4'h0 : _GEN_18365; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18367 = 12'hb7b == _T_171[11:0] ? 4'h0 : _GEN_18366; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18368 = 12'hb7c == _T_171[11:0] ? 4'h0 : _GEN_18367; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18369 = 12'hb7d == _T_171[11:0] ? 4'h0 : _GEN_18368; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18370 = 12'hb7e == _T_171[11:0] ? 4'h0 : _GEN_18369; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18371 = 12'hb7f == _T_171[11:0] ? 4'h0 : _GEN_18370; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18372 = 12'hb80 == _T_171[11:0] ? 4'h0 : _GEN_18371; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18373 = 12'hb81 == _T_171[11:0] ? 4'h0 : _GEN_18372; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18374 = 12'hb82 == _T_171[11:0] ? 4'h0 : _GEN_18373; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18375 = 12'hb83 == _T_171[11:0] ? 4'h0 : _GEN_18374; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18376 = 12'hb84 == _T_171[11:0] ? 4'h0 : _GEN_18375; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18377 = 12'hb85 == _T_171[11:0] ? 4'h0 : _GEN_18376; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18378 = 12'hb86 == _T_171[11:0] ? 4'h0 : _GEN_18377; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18379 = 12'hb87 == _T_171[11:0] ? 4'h0 : _GEN_18378; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18380 = 12'hb88 == _T_171[11:0] ? 4'h0 : _GEN_18379; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18381 = 12'hb89 == _T_171[11:0] ? 4'h0 : _GEN_18380; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18382 = 12'hb8a == _T_171[11:0] ? 4'h0 : _GEN_18381; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18383 = 12'hb8b == _T_171[11:0] ? 4'h0 : _GEN_18382; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18384 = 12'hb8c == _T_171[11:0] ? 4'h0 : _GEN_18383; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18385 = 12'hb8d == _T_171[11:0] ? 4'h0 : _GEN_18384; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18386 = 12'hb8e == _T_171[11:0] ? 4'h0 : _GEN_18385; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18387 = 12'hb8f == _T_171[11:0] ? 4'h0 : _GEN_18386; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18388 = 12'hb90 == _T_171[11:0] ? 4'h0 : _GEN_18387; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18389 = 12'hb91 == _T_171[11:0] ? 4'h0 : _GEN_18388; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18390 = 12'hb92 == _T_171[11:0] ? 4'h0 : _GEN_18389; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18391 = 12'hb93 == _T_171[11:0] ? 4'h0 : _GEN_18390; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18392 = 12'hb94 == _T_171[11:0] ? 4'h0 : _GEN_18391; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18393 = 12'hb95 == _T_171[11:0] ? image_2965 : _GEN_18392; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18394 = 12'hb96 == _T_171[11:0] ? image_2966 : _GEN_18393; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18395 = 12'hb97 == _T_171[11:0] ? image_2967 : _GEN_18394; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18396 = 12'hb98 == _T_171[11:0] ? image_2968 : _GEN_18395; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18397 = 12'hb99 == _T_171[11:0] ? image_2969 : _GEN_18396; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18398 = 12'hb9a == _T_171[11:0] ? image_2970 : _GEN_18397; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18399 = 12'hb9b == _T_171[11:0] ? image_2971 : _GEN_18398; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18400 = 12'hb9c == _T_171[11:0] ? image_2972 : _GEN_18399; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18401 = 12'hb9d == _T_171[11:0] ? image_2973 : _GEN_18400; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18402 = 12'hb9e == _T_171[11:0] ? image_2974 : _GEN_18401; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18403 = 12'hb9f == _T_171[11:0] ? image_2975 : _GEN_18402; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18404 = 12'hba0 == _T_171[11:0] ? image_2976 : _GEN_18403; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18405 = 12'hba1 == _T_171[11:0] ? image_2977 : _GEN_18404; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18406 = 12'hba2 == _T_171[11:0] ? image_2978 : _GEN_18405; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18407 = 12'hba3 == _T_171[11:0] ? image_2979 : _GEN_18406; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18408 = 12'hba4 == _T_171[11:0] ? image_2980 : _GEN_18407; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18409 = 12'hba5 == _T_171[11:0] ? image_2981 : _GEN_18408; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18410 = 12'hba6 == _T_171[11:0] ? image_2982 : _GEN_18409; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18411 = 12'hba7 == _T_171[11:0] ? image_2983 : _GEN_18410; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18412 = 12'hba8 == _T_171[11:0] ? image_2984 : _GEN_18411; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18413 = 12'hba9 == _T_171[11:0] ? image_2985 : _GEN_18412; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18414 = 12'hbaa == _T_171[11:0] ? image_2986 : _GEN_18413; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18415 = 12'hbab == _T_171[11:0] ? image_2987 : _GEN_18414; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18416 = 12'hbac == _T_171[11:0] ? image_2988 : _GEN_18415; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18417 = 12'hbad == _T_171[11:0] ? image_2989 : _GEN_18416; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18418 = 12'hbae == _T_171[11:0] ? image_2990 : _GEN_18417; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18419 = 12'hbaf == _T_171[11:0] ? image_2991 : _GEN_18418; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18420 = 12'hbb0 == _T_171[11:0] ? image_2992 : _GEN_18419; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18421 = 12'hbb1 == _T_171[11:0] ? image_2993 : _GEN_18420; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18422 = 12'hbb2 == _T_171[11:0] ? image_2994 : _GEN_18421; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18423 = 12'hbb3 == _T_171[11:0] ? image_2995 : _GEN_18422; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18424 = 12'hbb4 == _T_171[11:0] ? image_2996 : _GEN_18423; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18425 = 12'hbb5 == _T_171[11:0] ? 4'h0 : _GEN_18424; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18426 = 12'hbb6 == _T_171[11:0] ? 4'h0 : _GEN_18425; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18427 = 12'hbb7 == _T_171[11:0] ? 4'h0 : _GEN_18426; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18428 = 12'hbb8 == _T_171[11:0] ? 4'h0 : _GEN_18427; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18429 = 12'hbb9 == _T_171[11:0] ? 4'h0 : _GEN_18428; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18430 = 12'hbba == _T_171[11:0] ? 4'h0 : _GEN_18429; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18431 = 12'hbbb == _T_171[11:0] ? 4'h0 : _GEN_18430; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18432 = 12'hbbc == _T_171[11:0] ? 4'h0 : _GEN_18431; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18433 = 12'hbbd == _T_171[11:0] ? 4'h0 : _GEN_18432; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18434 = 12'hbbe == _T_171[11:0] ? 4'h0 : _GEN_18433; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18435 = 12'hbbf == _T_171[11:0] ? 4'h0 : _GEN_18434; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18436 = 12'hbc0 == _T_171[11:0] ? 4'h0 : _GEN_18435; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18437 = 12'hbc1 == _T_171[11:0] ? 4'h0 : _GEN_18436; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18438 = 12'hbc2 == _T_171[11:0] ? 4'h0 : _GEN_18437; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18439 = 12'hbc3 == _T_171[11:0] ? 4'h0 : _GEN_18438; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18440 = 12'hbc4 == _T_171[11:0] ? 4'h0 : _GEN_18439; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18441 = 12'hbc5 == _T_171[11:0] ? 4'h0 : _GEN_18440; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18442 = 12'hbc6 == _T_171[11:0] ? 4'h0 : _GEN_18441; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18443 = 12'hbc7 == _T_171[11:0] ? 4'h0 : _GEN_18442; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18444 = 12'hbc8 == _T_171[11:0] ? 4'h0 : _GEN_18443; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18445 = 12'hbc9 == _T_171[11:0] ? 4'h0 : _GEN_18444; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18446 = 12'hbca == _T_171[11:0] ? 4'h0 : _GEN_18445; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18447 = 12'hbcb == _T_171[11:0] ? 4'h0 : _GEN_18446; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18448 = 12'hbcc == _T_171[11:0] ? 4'h0 : _GEN_18447; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18449 = 12'hbcd == _T_171[11:0] ? 4'h0 : _GEN_18448; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18450 = 12'hbce == _T_171[11:0] ? 4'h0 : _GEN_18449; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18451 = 12'hbcf == _T_171[11:0] ? 4'h0 : _GEN_18450; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18452 = 12'hbd0 == _T_171[11:0] ? 4'h0 : _GEN_18451; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18453 = 12'hbd1 == _T_171[11:0] ? 4'h0 : _GEN_18452; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18454 = 12'hbd2 == _T_171[11:0] ? 4'h0 : _GEN_18453; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18455 = 12'hbd3 == _T_171[11:0] ? 4'h0 : _GEN_18454; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18456 = 12'hbd4 == _T_171[11:0] ? 4'h0 : _GEN_18455; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18457 = 12'hbd5 == _T_171[11:0] ? 4'h0 : _GEN_18456; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18458 = 12'hbd6 == _T_171[11:0] ? 4'h0 : _GEN_18457; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18459 = 12'hbd7 == _T_171[11:0] ? 4'h0 : _GEN_18458; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18460 = 12'hbd8 == _T_171[11:0] ? 4'h0 : _GEN_18459; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18461 = 12'hbd9 == _T_171[11:0] ? 4'h0 : _GEN_18460; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18462 = 12'hbda == _T_171[11:0] ? 4'h0 : _GEN_18461; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18463 = 12'hbdb == _T_171[11:0] ? image_3035 : _GEN_18462; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18464 = 12'hbdc == _T_171[11:0] ? image_3036 : _GEN_18463; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18465 = 12'hbdd == _T_171[11:0] ? image_3037 : _GEN_18464; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18466 = 12'hbde == _T_171[11:0] ? image_3038 : _GEN_18465; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18467 = 12'hbdf == _T_171[11:0] ? image_3039 : _GEN_18466; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18468 = 12'hbe0 == _T_171[11:0] ? image_3040 : _GEN_18467; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18469 = 12'hbe1 == _T_171[11:0] ? image_3041 : _GEN_18468; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18470 = 12'hbe2 == _T_171[11:0] ? image_3042 : _GEN_18469; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18471 = 12'hbe3 == _T_171[11:0] ? image_3043 : _GEN_18470; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18472 = 12'hbe4 == _T_171[11:0] ? image_3044 : _GEN_18471; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18473 = 12'hbe5 == _T_171[11:0] ? image_3045 : _GEN_18472; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18474 = 12'hbe6 == _T_171[11:0] ? image_3046 : _GEN_18473; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18475 = 12'hbe7 == _T_171[11:0] ? image_3047 : _GEN_18474; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18476 = 12'hbe8 == _T_171[11:0] ? image_3048 : _GEN_18475; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18477 = 12'hbe9 == _T_171[11:0] ? image_3049 : _GEN_18476; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18478 = 12'hbea == _T_171[11:0] ? image_3050 : _GEN_18477; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18479 = 12'hbeb == _T_171[11:0] ? image_3051 : _GEN_18478; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18480 = 12'hbec == _T_171[11:0] ? image_3052 : _GEN_18479; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18481 = 12'hbed == _T_171[11:0] ? image_3053 : _GEN_18480; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18482 = 12'hbee == _T_171[11:0] ? image_3054 : _GEN_18481; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18483 = 12'hbef == _T_171[11:0] ? image_3055 : _GEN_18482; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18484 = 12'hbf0 == _T_171[11:0] ? image_3056 : _GEN_18483; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18485 = 12'hbf1 == _T_171[11:0] ? 4'h0 : _GEN_18484; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18486 = 12'hbf2 == _T_171[11:0] ? 4'h0 : _GEN_18485; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18487 = 12'hbf3 == _T_171[11:0] ? 4'h0 : _GEN_18486; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18488 = 12'hbf4 == _T_171[11:0] ? 4'h0 : _GEN_18487; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18489 = 12'hbf5 == _T_171[11:0] ? 4'h0 : _GEN_18488; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18490 = 12'hbf6 == _T_171[11:0] ? 4'h0 : _GEN_18489; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18491 = 12'hbf7 == _T_171[11:0] ? 4'h0 : _GEN_18490; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18492 = 12'hbf8 == _T_171[11:0] ? 4'h0 : _GEN_18491; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18493 = 12'hbf9 == _T_171[11:0] ? 4'h0 : _GEN_18492; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18494 = 12'hbfa == _T_171[11:0] ? 4'h0 : _GEN_18493; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18495 = 12'hbfb == _T_171[11:0] ? 4'h0 : _GEN_18494; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18496 = 12'hbfc == _T_171[11:0] ? 4'h0 : _GEN_18495; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18497 = 12'hbfd == _T_171[11:0] ? 4'h0 : _GEN_18496; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18498 = 12'hbfe == _T_171[11:0] ? 4'h0 : _GEN_18497; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18499 = 12'hbff == _T_171[11:0] ? 4'h0 : _GEN_18498; // @[Filter.scala 138:46]
  wire [31:0] _T_174 = pixelIndex + 32'h6; // @[Filter.scala 133:29]
  wire [31:0] _T_175 = _T_174 / 32'h40; // @[Filter.scala 133:36]
  wire [31:0] _T_177 = _T_175 + _GEN_24805; // @[Filter.scala 133:51]
  wire [31:0] _T_179 = _T_177 - 32'h1; // @[Filter.scala 133:67]
  wire [31:0] _GEN_6 = _T_174 % 32'h40; // @[Filter.scala 134:36]
  wire [6:0] _T_182 = _GEN_6[6:0]; // @[Filter.scala 134:36]
  wire [6:0] _T_184 = _T_182 + _GEN_24806; // @[Filter.scala 134:51]
  wire [6:0] _T_186 = _T_184 - 7'h1; // @[Filter.scala 134:67]
  wire  _T_188 = _T_179 >= 32'h40; // @[Filter.scala 135:27]
  wire  _T_192 = _T_186 >= 7'h30; // @[Filter.scala 135:59]
  wire  _T_193 = _T_188 | _T_192; // @[Filter.scala 135:54]
  wire [13:0] _T_194 = _T_186 * 7'h40; // @[Filter.scala 138:57]
  wire [31:0] _GEN_24825 = {{18'd0}, _T_194}; // @[Filter.scala 138:72]
  wire [31:0] _T_196 = _GEN_24825 + _T_179; // @[Filter.scala 138:72]
  wire [3:0] _GEN_18513 = 12'hc == _T_196[11:0] ? image_12 : 4'h0; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18514 = 12'hd == _T_196[11:0] ? 4'h0 : _GEN_18513; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18515 = 12'he == _T_196[11:0] ? image_14 : _GEN_18514; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18516 = 12'hf == _T_196[11:0] ? image_15 : _GEN_18515; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18517 = 12'h10 == _T_196[11:0] ? image_16 : _GEN_18516; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18518 = 12'h11 == _T_196[11:0] ? image_17 : _GEN_18517; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18519 = 12'h12 == _T_196[11:0] ? image_18 : _GEN_18518; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18520 = 12'h13 == _T_196[11:0] ? image_19 : _GEN_18519; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18521 = 12'h14 == _T_196[11:0] ? image_20 : _GEN_18520; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18522 = 12'h15 == _T_196[11:0] ? image_21 : _GEN_18521; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18523 = 12'h16 == _T_196[11:0] ? image_22 : _GEN_18522; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18524 = 12'h17 == _T_196[11:0] ? image_23 : _GEN_18523; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18525 = 12'h18 == _T_196[11:0] ? 4'h0 : _GEN_18524; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18526 = 12'h19 == _T_196[11:0] ? 4'h0 : _GEN_18525; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18527 = 12'h1a == _T_196[11:0] ? 4'h0 : _GEN_18526; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18528 = 12'h1b == _T_196[11:0] ? 4'h0 : _GEN_18527; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18529 = 12'h1c == _T_196[11:0] ? 4'h0 : _GEN_18528; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18530 = 12'h1d == _T_196[11:0] ? 4'h0 : _GEN_18529; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18531 = 12'h1e == _T_196[11:0] ? 4'h0 : _GEN_18530; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18532 = 12'h1f == _T_196[11:0] ? 4'h0 : _GEN_18531; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18533 = 12'h20 == _T_196[11:0] ? 4'h0 : _GEN_18532; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18534 = 12'h21 == _T_196[11:0] ? 4'h0 : _GEN_18533; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18535 = 12'h22 == _T_196[11:0] ? 4'h0 : _GEN_18534; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18536 = 12'h23 == _T_196[11:0] ? image_35 : _GEN_18535; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18537 = 12'h24 == _T_196[11:0] ? image_36 : _GEN_18536; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18538 = 12'h25 == _T_196[11:0] ? image_37 : _GEN_18537; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18539 = 12'h26 == _T_196[11:0] ? image_38 : _GEN_18538; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18540 = 12'h27 == _T_196[11:0] ? image_39 : _GEN_18539; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18541 = 12'h28 == _T_196[11:0] ? image_40 : _GEN_18540; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18542 = 12'h29 == _T_196[11:0] ? image_41 : _GEN_18541; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18543 = 12'h2a == _T_196[11:0] ? image_42 : _GEN_18542; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18544 = 12'h2b == _T_196[11:0] ? 4'h0 : _GEN_18543; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18545 = 12'h2c == _T_196[11:0] ? 4'h0 : _GEN_18544; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18546 = 12'h2d == _T_196[11:0] ? 4'h0 : _GEN_18545; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18547 = 12'h2e == _T_196[11:0] ? 4'h0 : _GEN_18546; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18548 = 12'h2f == _T_196[11:0] ? 4'h0 : _GEN_18547; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18549 = 12'h30 == _T_196[11:0] ? 4'h0 : _GEN_18548; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18550 = 12'h31 == _T_196[11:0] ? 4'h0 : _GEN_18549; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18551 = 12'h32 == _T_196[11:0] ? 4'h0 : _GEN_18550; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18552 = 12'h33 == _T_196[11:0] ? 4'h0 : _GEN_18551; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18553 = 12'h34 == _T_196[11:0] ? 4'h0 : _GEN_18552; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18554 = 12'h35 == _T_196[11:0] ? 4'h0 : _GEN_18553; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18555 = 12'h36 == _T_196[11:0] ? 4'h0 : _GEN_18554; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18556 = 12'h37 == _T_196[11:0] ? 4'h0 : _GEN_18555; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18557 = 12'h38 == _T_196[11:0] ? 4'h0 : _GEN_18556; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18558 = 12'h39 == _T_196[11:0] ? 4'h0 : _GEN_18557; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18559 = 12'h3a == _T_196[11:0] ? 4'h0 : _GEN_18558; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18560 = 12'h3b == _T_196[11:0] ? 4'h0 : _GEN_18559; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18561 = 12'h3c == _T_196[11:0] ? 4'h0 : _GEN_18560; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18562 = 12'h3d == _T_196[11:0] ? 4'h0 : _GEN_18561; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18563 = 12'h3e == _T_196[11:0] ? 4'h0 : _GEN_18562; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18564 = 12'h3f == _T_196[11:0] ? 4'h0 : _GEN_18563; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18565 = 12'h40 == _T_196[11:0] ? 4'h0 : _GEN_18564; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18566 = 12'h41 == _T_196[11:0] ? 4'h0 : _GEN_18565; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18567 = 12'h42 == _T_196[11:0] ? 4'h0 : _GEN_18566; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18568 = 12'h43 == _T_196[11:0] ? 4'h0 : _GEN_18567; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18569 = 12'h44 == _T_196[11:0] ? 4'h0 : _GEN_18568; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18570 = 12'h45 == _T_196[11:0] ? 4'h0 : _GEN_18569; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18571 = 12'h46 == _T_196[11:0] ? 4'h0 : _GEN_18570; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18572 = 12'h47 == _T_196[11:0] ? 4'h0 : _GEN_18571; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18573 = 12'h48 == _T_196[11:0] ? 4'h0 : _GEN_18572; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18574 = 12'h49 == _T_196[11:0] ? 4'h0 : _GEN_18573; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18575 = 12'h4a == _T_196[11:0] ? 4'h0 : _GEN_18574; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18576 = 12'h4b == _T_196[11:0] ? image_75 : _GEN_18575; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18577 = 12'h4c == _T_196[11:0] ? image_76 : _GEN_18576; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18578 = 12'h4d == _T_196[11:0] ? image_77 : _GEN_18577; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18579 = 12'h4e == _T_196[11:0] ? image_78 : _GEN_18578; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18580 = 12'h4f == _T_196[11:0] ? image_79 : _GEN_18579; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18581 = 12'h50 == _T_196[11:0] ? image_80 : _GEN_18580; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18582 = 12'h51 == _T_196[11:0] ? image_81 : _GEN_18581; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18583 = 12'h52 == _T_196[11:0] ? image_82 : _GEN_18582; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18584 = 12'h53 == _T_196[11:0] ? image_83 : _GEN_18583; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18585 = 12'h54 == _T_196[11:0] ? image_84 : _GEN_18584; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18586 = 12'h55 == _T_196[11:0] ? image_85 : _GEN_18585; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18587 = 12'h56 == _T_196[11:0] ? image_86 : _GEN_18586; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18588 = 12'h57 == _T_196[11:0] ? image_87 : _GEN_18587; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18589 = 12'h58 == _T_196[11:0] ? image_88 : _GEN_18588; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18590 = 12'h59 == _T_196[11:0] ? image_89 : _GEN_18589; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18591 = 12'h5a == _T_196[11:0] ? image_90 : _GEN_18590; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18592 = 12'h5b == _T_196[11:0] ? 4'h0 : _GEN_18591; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18593 = 12'h5c == _T_196[11:0] ? 4'h0 : _GEN_18592; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18594 = 12'h5d == _T_196[11:0] ? image_93 : _GEN_18593; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18595 = 12'h5e == _T_196[11:0] ? 4'h0 : _GEN_18594; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18596 = 12'h5f == _T_196[11:0] ? image_95 : _GEN_18595; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18597 = 12'h60 == _T_196[11:0] ? image_96 : _GEN_18596; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18598 = 12'h61 == _T_196[11:0] ? image_97 : _GEN_18597; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18599 = 12'h62 == _T_196[11:0] ? image_98 : _GEN_18598; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18600 = 12'h63 == _T_196[11:0] ? image_99 : _GEN_18599; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18601 = 12'h64 == _T_196[11:0] ? image_100 : _GEN_18600; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18602 = 12'h65 == _T_196[11:0] ? image_101 : _GEN_18601; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18603 = 12'h66 == _T_196[11:0] ? image_102 : _GEN_18602; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18604 = 12'h67 == _T_196[11:0] ? image_103 : _GEN_18603; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18605 = 12'h68 == _T_196[11:0] ? image_104 : _GEN_18604; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18606 = 12'h69 == _T_196[11:0] ? image_105 : _GEN_18605; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18607 = 12'h6a == _T_196[11:0] ? image_106 : _GEN_18606; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18608 = 12'h6b == _T_196[11:0] ? image_107 : _GEN_18607; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18609 = 12'h6c == _T_196[11:0] ? image_108 : _GEN_18608; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18610 = 12'h6d == _T_196[11:0] ? 4'h0 : _GEN_18609; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18611 = 12'h6e == _T_196[11:0] ? 4'h0 : _GEN_18610; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18612 = 12'h6f == _T_196[11:0] ? 4'h0 : _GEN_18611; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18613 = 12'h70 == _T_196[11:0] ? 4'h0 : _GEN_18612; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18614 = 12'h71 == _T_196[11:0] ? 4'h0 : _GEN_18613; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18615 = 12'h72 == _T_196[11:0] ? 4'h0 : _GEN_18614; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18616 = 12'h73 == _T_196[11:0] ? 4'h0 : _GEN_18615; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18617 = 12'h74 == _T_196[11:0] ? 4'h0 : _GEN_18616; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18618 = 12'h75 == _T_196[11:0] ? 4'h0 : _GEN_18617; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18619 = 12'h76 == _T_196[11:0] ? 4'h0 : _GEN_18618; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18620 = 12'h77 == _T_196[11:0] ? 4'h0 : _GEN_18619; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18621 = 12'h78 == _T_196[11:0] ? 4'h0 : _GEN_18620; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18622 = 12'h79 == _T_196[11:0] ? 4'h0 : _GEN_18621; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18623 = 12'h7a == _T_196[11:0] ? 4'h0 : _GEN_18622; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18624 = 12'h7b == _T_196[11:0] ? 4'h0 : _GEN_18623; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18625 = 12'h7c == _T_196[11:0] ? 4'h0 : _GEN_18624; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18626 = 12'h7d == _T_196[11:0] ? 4'h0 : _GEN_18625; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18627 = 12'h7e == _T_196[11:0] ? 4'h0 : _GEN_18626; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18628 = 12'h7f == _T_196[11:0] ? 4'h0 : _GEN_18627; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18629 = 12'h80 == _T_196[11:0] ? 4'h0 : _GEN_18628; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18630 = 12'h81 == _T_196[11:0] ? 4'h0 : _GEN_18629; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18631 = 12'h82 == _T_196[11:0] ? 4'h0 : _GEN_18630; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18632 = 12'h83 == _T_196[11:0] ? 4'h0 : _GEN_18631; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18633 = 12'h84 == _T_196[11:0] ? 4'h0 : _GEN_18632; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18634 = 12'h85 == _T_196[11:0] ? 4'h0 : _GEN_18633; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18635 = 12'h86 == _T_196[11:0] ? 4'h0 : _GEN_18634; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18636 = 12'h87 == _T_196[11:0] ? 4'h0 : _GEN_18635; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18637 = 12'h88 == _T_196[11:0] ? image_136 : _GEN_18636; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18638 = 12'h89 == _T_196[11:0] ? image_137 : _GEN_18637; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18639 = 12'h8a == _T_196[11:0] ? image_138 : _GEN_18638; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18640 = 12'h8b == _T_196[11:0] ? image_139 : _GEN_18639; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18641 = 12'h8c == _T_196[11:0] ? image_140 : _GEN_18640; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18642 = 12'h8d == _T_196[11:0] ? image_141 : _GEN_18641; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18643 = 12'h8e == _T_196[11:0] ? image_142 : _GEN_18642; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18644 = 12'h8f == _T_196[11:0] ? image_143 : _GEN_18643; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18645 = 12'h90 == _T_196[11:0] ? image_144 : _GEN_18644; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18646 = 12'h91 == _T_196[11:0] ? image_145 : _GEN_18645; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18647 = 12'h92 == _T_196[11:0] ? image_146 : _GEN_18646; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18648 = 12'h93 == _T_196[11:0] ? image_147 : _GEN_18647; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18649 = 12'h94 == _T_196[11:0] ? image_148 : _GEN_18648; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18650 = 12'h95 == _T_196[11:0] ? image_149 : _GEN_18649; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18651 = 12'h96 == _T_196[11:0] ? image_150 : _GEN_18650; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18652 = 12'h97 == _T_196[11:0] ? image_151 : _GEN_18651; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18653 = 12'h98 == _T_196[11:0] ? image_152 : _GEN_18652; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18654 = 12'h99 == _T_196[11:0] ? image_153 : _GEN_18653; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18655 = 12'h9a == _T_196[11:0] ? image_154 : _GEN_18654; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18656 = 12'h9b == _T_196[11:0] ? image_155 : _GEN_18655; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18657 = 12'h9c == _T_196[11:0] ? 4'h0 : _GEN_18656; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18658 = 12'h9d == _T_196[11:0] ? image_157 : _GEN_18657; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18659 = 12'h9e == _T_196[11:0] ? image_158 : _GEN_18658; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18660 = 12'h9f == _T_196[11:0] ? image_159 : _GEN_18659; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18661 = 12'ha0 == _T_196[11:0] ? image_160 : _GEN_18660; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18662 = 12'ha1 == _T_196[11:0] ? image_161 : _GEN_18661; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18663 = 12'ha2 == _T_196[11:0] ? image_162 : _GEN_18662; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18664 = 12'ha3 == _T_196[11:0] ? image_163 : _GEN_18663; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18665 = 12'ha4 == _T_196[11:0] ? image_164 : _GEN_18664; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18666 = 12'ha5 == _T_196[11:0] ? image_165 : _GEN_18665; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18667 = 12'ha6 == _T_196[11:0] ? image_166 : _GEN_18666; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18668 = 12'ha7 == _T_196[11:0] ? image_167 : _GEN_18667; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18669 = 12'ha8 == _T_196[11:0] ? image_168 : _GEN_18668; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18670 = 12'ha9 == _T_196[11:0] ? image_169 : _GEN_18669; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18671 = 12'haa == _T_196[11:0] ? image_170 : _GEN_18670; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18672 = 12'hab == _T_196[11:0] ? image_171 : _GEN_18671; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18673 = 12'hac == _T_196[11:0] ? image_172 : _GEN_18672; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18674 = 12'had == _T_196[11:0] ? image_173 : _GEN_18673; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18675 = 12'hae == _T_196[11:0] ? image_174 : _GEN_18674; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18676 = 12'haf == _T_196[11:0] ? image_175 : _GEN_18675; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18677 = 12'hb0 == _T_196[11:0] ? image_176 : _GEN_18676; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18678 = 12'hb1 == _T_196[11:0] ? image_177 : _GEN_18677; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18679 = 12'hb2 == _T_196[11:0] ? image_178 : _GEN_18678; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18680 = 12'hb3 == _T_196[11:0] ? image_179 : _GEN_18679; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18681 = 12'hb4 == _T_196[11:0] ? 4'h0 : _GEN_18680; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18682 = 12'hb5 == _T_196[11:0] ? 4'h0 : _GEN_18681; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18683 = 12'hb6 == _T_196[11:0] ? 4'h0 : _GEN_18682; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18684 = 12'hb7 == _T_196[11:0] ? 4'h0 : _GEN_18683; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18685 = 12'hb8 == _T_196[11:0] ? 4'h0 : _GEN_18684; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18686 = 12'hb9 == _T_196[11:0] ? 4'h0 : _GEN_18685; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18687 = 12'hba == _T_196[11:0] ? 4'h0 : _GEN_18686; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18688 = 12'hbb == _T_196[11:0] ? 4'h0 : _GEN_18687; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18689 = 12'hbc == _T_196[11:0] ? 4'h0 : _GEN_18688; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18690 = 12'hbd == _T_196[11:0] ? 4'h0 : _GEN_18689; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18691 = 12'hbe == _T_196[11:0] ? 4'h0 : _GEN_18690; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18692 = 12'hbf == _T_196[11:0] ? 4'h0 : _GEN_18691; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18693 = 12'hc0 == _T_196[11:0] ? 4'h0 : _GEN_18692; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18694 = 12'hc1 == _T_196[11:0] ? 4'h0 : _GEN_18693; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18695 = 12'hc2 == _T_196[11:0] ? 4'h0 : _GEN_18694; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18696 = 12'hc3 == _T_196[11:0] ? 4'h0 : _GEN_18695; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18697 = 12'hc4 == _T_196[11:0] ? 4'h0 : _GEN_18696; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18698 = 12'hc5 == _T_196[11:0] ? 4'h0 : _GEN_18697; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18699 = 12'hc6 == _T_196[11:0] ? 4'h0 : _GEN_18698; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18700 = 12'hc7 == _T_196[11:0] ? image_199 : _GEN_18699; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18701 = 12'hc8 == _T_196[11:0] ? image_200 : _GEN_18700; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18702 = 12'hc9 == _T_196[11:0] ? image_201 : _GEN_18701; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18703 = 12'hca == _T_196[11:0] ? image_202 : _GEN_18702; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18704 = 12'hcb == _T_196[11:0] ? image_203 : _GEN_18703; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18705 = 12'hcc == _T_196[11:0] ? image_204 : _GEN_18704; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18706 = 12'hcd == _T_196[11:0] ? image_205 : _GEN_18705; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18707 = 12'hce == _T_196[11:0] ? image_206 : _GEN_18706; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18708 = 12'hcf == _T_196[11:0] ? image_207 : _GEN_18707; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18709 = 12'hd0 == _T_196[11:0] ? image_208 : _GEN_18708; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18710 = 12'hd1 == _T_196[11:0] ? image_209 : _GEN_18709; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18711 = 12'hd2 == _T_196[11:0] ? image_210 : _GEN_18710; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18712 = 12'hd3 == _T_196[11:0] ? image_211 : _GEN_18711; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18713 = 12'hd4 == _T_196[11:0] ? image_212 : _GEN_18712; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18714 = 12'hd5 == _T_196[11:0] ? image_213 : _GEN_18713; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18715 = 12'hd6 == _T_196[11:0] ? image_214 : _GEN_18714; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18716 = 12'hd7 == _T_196[11:0] ? image_215 : _GEN_18715; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18717 = 12'hd8 == _T_196[11:0] ? image_216 : _GEN_18716; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18718 = 12'hd9 == _T_196[11:0] ? image_217 : _GEN_18717; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18719 = 12'hda == _T_196[11:0] ? image_218 : _GEN_18718; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18720 = 12'hdb == _T_196[11:0] ? image_219 : _GEN_18719; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18721 = 12'hdc == _T_196[11:0] ? image_220 : _GEN_18720; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18722 = 12'hdd == _T_196[11:0] ? image_221 : _GEN_18721; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18723 = 12'hde == _T_196[11:0] ? image_222 : _GEN_18722; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18724 = 12'hdf == _T_196[11:0] ? image_223 : _GEN_18723; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18725 = 12'he0 == _T_196[11:0] ? image_224 : _GEN_18724; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18726 = 12'he1 == _T_196[11:0] ? image_225 : _GEN_18725; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18727 = 12'he2 == _T_196[11:0] ? image_226 : _GEN_18726; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18728 = 12'he3 == _T_196[11:0] ? image_227 : _GEN_18727; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18729 = 12'he4 == _T_196[11:0] ? image_228 : _GEN_18728; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18730 = 12'he5 == _T_196[11:0] ? image_229 : _GEN_18729; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18731 = 12'he6 == _T_196[11:0] ? image_230 : _GEN_18730; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18732 = 12'he7 == _T_196[11:0] ? image_231 : _GEN_18731; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18733 = 12'he8 == _T_196[11:0] ? image_232 : _GEN_18732; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18734 = 12'he9 == _T_196[11:0] ? image_233 : _GEN_18733; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18735 = 12'hea == _T_196[11:0] ? image_234 : _GEN_18734; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18736 = 12'heb == _T_196[11:0] ? image_235 : _GEN_18735; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18737 = 12'hec == _T_196[11:0] ? image_236 : _GEN_18736; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18738 = 12'hed == _T_196[11:0] ? image_237 : _GEN_18737; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18739 = 12'hee == _T_196[11:0] ? image_238 : _GEN_18738; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18740 = 12'hef == _T_196[11:0] ? image_239 : _GEN_18739; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18741 = 12'hf0 == _T_196[11:0] ? image_240 : _GEN_18740; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18742 = 12'hf1 == _T_196[11:0] ? image_241 : _GEN_18741; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18743 = 12'hf2 == _T_196[11:0] ? image_242 : _GEN_18742; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18744 = 12'hf3 == _T_196[11:0] ? image_243 : _GEN_18743; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18745 = 12'hf4 == _T_196[11:0] ? image_244 : _GEN_18744; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18746 = 12'hf5 == _T_196[11:0] ? image_245 : _GEN_18745; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18747 = 12'hf6 == _T_196[11:0] ? image_246 : _GEN_18746; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18748 = 12'hf7 == _T_196[11:0] ? 4'h0 : _GEN_18747; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18749 = 12'hf8 == _T_196[11:0] ? 4'h0 : _GEN_18748; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18750 = 12'hf9 == _T_196[11:0] ? 4'h0 : _GEN_18749; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18751 = 12'hfa == _T_196[11:0] ? 4'h0 : _GEN_18750; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18752 = 12'hfb == _T_196[11:0] ? 4'h0 : _GEN_18751; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18753 = 12'hfc == _T_196[11:0] ? 4'h0 : _GEN_18752; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18754 = 12'hfd == _T_196[11:0] ? 4'h0 : _GEN_18753; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18755 = 12'hfe == _T_196[11:0] ? 4'h0 : _GEN_18754; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18756 = 12'hff == _T_196[11:0] ? 4'h0 : _GEN_18755; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18757 = 12'h100 == _T_196[11:0] ? 4'h0 : _GEN_18756; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18758 = 12'h101 == _T_196[11:0] ? 4'h0 : _GEN_18757; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18759 = 12'h102 == _T_196[11:0] ? 4'h0 : _GEN_18758; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18760 = 12'h103 == _T_196[11:0] ? 4'h0 : _GEN_18759; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18761 = 12'h104 == _T_196[11:0] ? 4'h0 : _GEN_18760; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18762 = 12'h105 == _T_196[11:0] ? 4'h0 : _GEN_18761; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18763 = 12'h106 == _T_196[11:0] ? image_262 : _GEN_18762; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18764 = 12'h107 == _T_196[11:0] ? image_263 : _GEN_18763; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18765 = 12'h108 == _T_196[11:0] ? image_264 : _GEN_18764; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18766 = 12'h109 == _T_196[11:0] ? image_265 : _GEN_18765; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18767 = 12'h10a == _T_196[11:0] ? image_266 : _GEN_18766; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18768 = 12'h10b == _T_196[11:0] ? image_267 : _GEN_18767; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18769 = 12'h10c == _T_196[11:0] ? image_268 : _GEN_18768; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18770 = 12'h10d == _T_196[11:0] ? image_269 : _GEN_18769; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18771 = 12'h10e == _T_196[11:0] ? image_270 : _GEN_18770; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18772 = 12'h10f == _T_196[11:0] ? image_271 : _GEN_18771; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18773 = 12'h110 == _T_196[11:0] ? image_272 : _GEN_18772; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18774 = 12'h111 == _T_196[11:0] ? image_273 : _GEN_18773; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18775 = 12'h112 == _T_196[11:0] ? image_274 : _GEN_18774; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18776 = 12'h113 == _T_196[11:0] ? image_275 : _GEN_18775; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18777 = 12'h114 == _T_196[11:0] ? image_276 : _GEN_18776; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18778 = 12'h115 == _T_196[11:0] ? image_277 : _GEN_18777; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18779 = 12'h116 == _T_196[11:0] ? image_278 : _GEN_18778; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18780 = 12'h117 == _T_196[11:0] ? image_279 : _GEN_18779; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18781 = 12'h118 == _T_196[11:0] ? image_280 : _GEN_18780; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18782 = 12'h119 == _T_196[11:0] ? image_281 : _GEN_18781; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18783 = 12'h11a == _T_196[11:0] ? image_282 : _GEN_18782; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18784 = 12'h11b == _T_196[11:0] ? image_283 : _GEN_18783; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18785 = 12'h11c == _T_196[11:0] ? image_284 : _GEN_18784; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18786 = 12'h11d == _T_196[11:0] ? image_285 : _GEN_18785; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18787 = 12'h11e == _T_196[11:0] ? image_286 : _GEN_18786; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18788 = 12'h11f == _T_196[11:0] ? image_287 : _GEN_18787; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18789 = 12'h120 == _T_196[11:0] ? image_288 : _GEN_18788; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18790 = 12'h121 == _T_196[11:0] ? image_289 : _GEN_18789; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18791 = 12'h122 == _T_196[11:0] ? image_290 : _GEN_18790; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18792 = 12'h123 == _T_196[11:0] ? image_291 : _GEN_18791; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18793 = 12'h124 == _T_196[11:0] ? image_292 : _GEN_18792; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18794 = 12'h125 == _T_196[11:0] ? image_293 : _GEN_18793; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18795 = 12'h126 == _T_196[11:0] ? image_294 : _GEN_18794; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18796 = 12'h127 == _T_196[11:0] ? image_295 : _GEN_18795; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18797 = 12'h128 == _T_196[11:0] ? image_296 : _GEN_18796; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18798 = 12'h129 == _T_196[11:0] ? image_297 : _GEN_18797; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18799 = 12'h12a == _T_196[11:0] ? image_298 : _GEN_18798; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18800 = 12'h12b == _T_196[11:0] ? image_299 : _GEN_18799; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18801 = 12'h12c == _T_196[11:0] ? image_300 : _GEN_18800; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18802 = 12'h12d == _T_196[11:0] ? image_301 : _GEN_18801; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18803 = 12'h12e == _T_196[11:0] ? image_302 : _GEN_18802; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18804 = 12'h12f == _T_196[11:0] ? image_303 : _GEN_18803; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18805 = 12'h130 == _T_196[11:0] ? image_304 : _GEN_18804; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18806 = 12'h131 == _T_196[11:0] ? image_305 : _GEN_18805; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18807 = 12'h132 == _T_196[11:0] ? image_306 : _GEN_18806; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18808 = 12'h133 == _T_196[11:0] ? image_307 : _GEN_18807; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18809 = 12'h134 == _T_196[11:0] ? image_308 : _GEN_18808; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18810 = 12'h135 == _T_196[11:0] ? image_309 : _GEN_18809; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18811 = 12'h136 == _T_196[11:0] ? image_310 : _GEN_18810; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18812 = 12'h137 == _T_196[11:0] ? image_311 : _GEN_18811; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18813 = 12'h138 == _T_196[11:0] ? image_312 : _GEN_18812; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18814 = 12'h139 == _T_196[11:0] ? image_313 : _GEN_18813; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18815 = 12'h13a == _T_196[11:0] ? image_314 : _GEN_18814; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18816 = 12'h13b == _T_196[11:0] ? image_315 : _GEN_18815; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18817 = 12'h13c == _T_196[11:0] ? 4'h0 : _GEN_18816; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18818 = 12'h13d == _T_196[11:0] ? 4'h0 : _GEN_18817; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18819 = 12'h13e == _T_196[11:0] ? 4'h0 : _GEN_18818; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18820 = 12'h13f == _T_196[11:0] ? 4'h0 : _GEN_18819; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18821 = 12'h140 == _T_196[11:0] ? 4'h0 : _GEN_18820; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18822 = 12'h141 == _T_196[11:0] ? 4'h0 : _GEN_18821; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18823 = 12'h142 == _T_196[11:0] ? 4'h0 : _GEN_18822; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18824 = 12'h143 == _T_196[11:0] ? 4'h0 : _GEN_18823; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18825 = 12'h144 == _T_196[11:0] ? 4'h0 : _GEN_18824; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18826 = 12'h145 == _T_196[11:0] ? image_325 : _GEN_18825; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18827 = 12'h146 == _T_196[11:0] ? image_326 : _GEN_18826; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18828 = 12'h147 == _T_196[11:0] ? image_327 : _GEN_18827; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18829 = 12'h148 == _T_196[11:0] ? image_328 : _GEN_18828; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18830 = 12'h149 == _T_196[11:0] ? image_329 : _GEN_18829; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18831 = 12'h14a == _T_196[11:0] ? image_330 : _GEN_18830; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18832 = 12'h14b == _T_196[11:0] ? image_331 : _GEN_18831; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18833 = 12'h14c == _T_196[11:0] ? image_332 : _GEN_18832; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18834 = 12'h14d == _T_196[11:0] ? image_333 : _GEN_18833; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18835 = 12'h14e == _T_196[11:0] ? image_334 : _GEN_18834; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18836 = 12'h14f == _T_196[11:0] ? image_335 : _GEN_18835; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18837 = 12'h150 == _T_196[11:0] ? image_336 : _GEN_18836; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18838 = 12'h151 == _T_196[11:0] ? image_337 : _GEN_18837; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18839 = 12'h152 == _T_196[11:0] ? image_338 : _GEN_18838; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18840 = 12'h153 == _T_196[11:0] ? image_339 : _GEN_18839; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18841 = 12'h154 == _T_196[11:0] ? image_340 : _GEN_18840; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18842 = 12'h155 == _T_196[11:0] ? image_341 : _GEN_18841; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18843 = 12'h156 == _T_196[11:0] ? image_342 : _GEN_18842; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18844 = 12'h157 == _T_196[11:0] ? image_343 : _GEN_18843; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18845 = 12'h158 == _T_196[11:0] ? image_344 : _GEN_18844; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18846 = 12'h159 == _T_196[11:0] ? image_345 : _GEN_18845; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18847 = 12'h15a == _T_196[11:0] ? image_346 : _GEN_18846; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18848 = 12'h15b == _T_196[11:0] ? image_347 : _GEN_18847; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18849 = 12'h15c == _T_196[11:0] ? image_348 : _GEN_18848; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18850 = 12'h15d == _T_196[11:0] ? image_349 : _GEN_18849; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18851 = 12'h15e == _T_196[11:0] ? image_350 : _GEN_18850; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18852 = 12'h15f == _T_196[11:0] ? image_351 : _GEN_18851; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18853 = 12'h160 == _T_196[11:0] ? image_352 : _GEN_18852; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18854 = 12'h161 == _T_196[11:0] ? image_353 : _GEN_18853; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18855 = 12'h162 == _T_196[11:0] ? image_354 : _GEN_18854; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18856 = 12'h163 == _T_196[11:0] ? image_355 : _GEN_18855; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18857 = 12'h164 == _T_196[11:0] ? image_356 : _GEN_18856; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18858 = 12'h165 == _T_196[11:0] ? image_357 : _GEN_18857; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18859 = 12'h166 == _T_196[11:0] ? image_358 : _GEN_18858; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18860 = 12'h167 == _T_196[11:0] ? image_359 : _GEN_18859; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18861 = 12'h168 == _T_196[11:0] ? image_360 : _GEN_18860; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18862 = 12'h169 == _T_196[11:0] ? image_361 : _GEN_18861; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18863 = 12'h16a == _T_196[11:0] ? image_362 : _GEN_18862; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18864 = 12'h16b == _T_196[11:0] ? image_363 : _GEN_18863; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18865 = 12'h16c == _T_196[11:0] ? image_364 : _GEN_18864; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18866 = 12'h16d == _T_196[11:0] ? image_365 : _GEN_18865; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18867 = 12'h16e == _T_196[11:0] ? image_366 : _GEN_18866; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18868 = 12'h16f == _T_196[11:0] ? image_367 : _GEN_18867; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18869 = 12'h170 == _T_196[11:0] ? image_368 : _GEN_18868; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18870 = 12'h171 == _T_196[11:0] ? image_369 : _GEN_18869; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18871 = 12'h172 == _T_196[11:0] ? image_370 : _GEN_18870; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18872 = 12'h173 == _T_196[11:0] ? image_371 : _GEN_18871; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18873 = 12'h174 == _T_196[11:0] ? image_372 : _GEN_18872; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18874 = 12'h175 == _T_196[11:0] ? image_373 : _GEN_18873; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18875 = 12'h176 == _T_196[11:0] ? image_374 : _GEN_18874; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18876 = 12'h177 == _T_196[11:0] ? image_375 : _GEN_18875; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18877 = 12'h178 == _T_196[11:0] ? image_376 : _GEN_18876; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18878 = 12'h179 == _T_196[11:0] ? image_377 : _GEN_18877; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18879 = 12'h17a == _T_196[11:0] ? image_378 : _GEN_18878; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18880 = 12'h17b == _T_196[11:0] ? image_379 : _GEN_18879; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18881 = 12'h17c == _T_196[11:0] ? 4'h0 : _GEN_18880; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18882 = 12'h17d == _T_196[11:0] ? 4'h0 : _GEN_18881; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18883 = 12'h17e == _T_196[11:0] ? 4'h0 : _GEN_18882; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18884 = 12'h17f == _T_196[11:0] ? 4'h0 : _GEN_18883; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18885 = 12'h180 == _T_196[11:0] ? 4'h0 : _GEN_18884; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18886 = 12'h181 == _T_196[11:0] ? 4'h0 : _GEN_18885; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18887 = 12'h182 == _T_196[11:0] ? 4'h0 : _GEN_18886; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18888 = 12'h183 == _T_196[11:0] ? 4'h0 : _GEN_18887; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18889 = 12'h184 == _T_196[11:0] ? image_388 : _GEN_18888; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18890 = 12'h185 == _T_196[11:0] ? image_389 : _GEN_18889; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18891 = 12'h186 == _T_196[11:0] ? image_390 : _GEN_18890; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18892 = 12'h187 == _T_196[11:0] ? image_391 : _GEN_18891; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18893 = 12'h188 == _T_196[11:0] ? image_392 : _GEN_18892; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18894 = 12'h189 == _T_196[11:0] ? image_393 : _GEN_18893; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18895 = 12'h18a == _T_196[11:0] ? image_394 : _GEN_18894; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18896 = 12'h18b == _T_196[11:0] ? image_395 : _GEN_18895; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18897 = 12'h18c == _T_196[11:0] ? image_396 : _GEN_18896; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18898 = 12'h18d == _T_196[11:0] ? image_397 : _GEN_18897; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18899 = 12'h18e == _T_196[11:0] ? image_398 : _GEN_18898; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18900 = 12'h18f == _T_196[11:0] ? image_399 : _GEN_18899; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18901 = 12'h190 == _T_196[11:0] ? image_400 : _GEN_18900; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18902 = 12'h191 == _T_196[11:0] ? image_401 : _GEN_18901; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18903 = 12'h192 == _T_196[11:0] ? image_402 : _GEN_18902; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18904 = 12'h193 == _T_196[11:0] ? image_403 : _GEN_18903; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18905 = 12'h194 == _T_196[11:0] ? image_404 : _GEN_18904; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18906 = 12'h195 == _T_196[11:0] ? image_405 : _GEN_18905; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18907 = 12'h196 == _T_196[11:0] ? image_406 : _GEN_18906; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18908 = 12'h197 == _T_196[11:0] ? image_407 : _GEN_18907; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18909 = 12'h198 == _T_196[11:0] ? image_408 : _GEN_18908; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18910 = 12'h199 == _T_196[11:0] ? image_409 : _GEN_18909; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18911 = 12'h19a == _T_196[11:0] ? image_410 : _GEN_18910; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18912 = 12'h19b == _T_196[11:0] ? image_411 : _GEN_18911; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18913 = 12'h19c == _T_196[11:0] ? image_412 : _GEN_18912; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18914 = 12'h19d == _T_196[11:0] ? image_413 : _GEN_18913; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18915 = 12'h19e == _T_196[11:0] ? image_414 : _GEN_18914; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18916 = 12'h19f == _T_196[11:0] ? image_415 : _GEN_18915; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18917 = 12'h1a0 == _T_196[11:0] ? image_416 : _GEN_18916; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18918 = 12'h1a1 == _T_196[11:0] ? image_417 : _GEN_18917; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18919 = 12'h1a2 == _T_196[11:0] ? image_418 : _GEN_18918; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18920 = 12'h1a3 == _T_196[11:0] ? image_419 : _GEN_18919; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18921 = 12'h1a4 == _T_196[11:0] ? image_420 : _GEN_18920; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18922 = 12'h1a5 == _T_196[11:0] ? image_421 : _GEN_18921; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18923 = 12'h1a6 == _T_196[11:0] ? image_422 : _GEN_18922; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18924 = 12'h1a7 == _T_196[11:0] ? image_423 : _GEN_18923; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18925 = 12'h1a8 == _T_196[11:0] ? image_424 : _GEN_18924; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18926 = 12'h1a9 == _T_196[11:0] ? image_425 : _GEN_18925; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18927 = 12'h1aa == _T_196[11:0] ? image_426 : _GEN_18926; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18928 = 12'h1ab == _T_196[11:0] ? image_427 : _GEN_18927; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18929 = 12'h1ac == _T_196[11:0] ? image_428 : _GEN_18928; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18930 = 12'h1ad == _T_196[11:0] ? image_429 : _GEN_18929; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18931 = 12'h1ae == _T_196[11:0] ? image_430 : _GEN_18930; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18932 = 12'h1af == _T_196[11:0] ? image_431 : _GEN_18931; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18933 = 12'h1b0 == _T_196[11:0] ? image_432 : _GEN_18932; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18934 = 12'h1b1 == _T_196[11:0] ? image_433 : _GEN_18933; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18935 = 12'h1b2 == _T_196[11:0] ? image_434 : _GEN_18934; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18936 = 12'h1b3 == _T_196[11:0] ? image_435 : _GEN_18935; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18937 = 12'h1b4 == _T_196[11:0] ? image_436 : _GEN_18936; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18938 = 12'h1b5 == _T_196[11:0] ? image_437 : _GEN_18937; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18939 = 12'h1b6 == _T_196[11:0] ? image_438 : _GEN_18938; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18940 = 12'h1b7 == _T_196[11:0] ? image_439 : _GEN_18939; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18941 = 12'h1b8 == _T_196[11:0] ? image_440 : _GEN_18940; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18942 = 12'h1b9 == _T_196[11:0] ? image_441 : _GEN_18941; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18943 = 12'h1ba == _T_196[11:0] ? image_442 : _GEN_18942; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18944 = 12'h1bb == _T_196[11:0] ? image_443 : _GEN_18943; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18945 = 12'h1bc == _T_196[11:0] ? image_444 : _GEN_18944; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18946 = 12'h1bd == _T_196[11:0] ? 4'h0 : _GEN_18945; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18947 = 12'h1be == _T_196[11:0] ? 4'h0 : _GEN_18946; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18948 = 12'h1bf == _T_196[11:0] ? 4'h0 : _GEN_18947; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18949 = 12'h1c0 == _T_196[11:0] ? 4'h0 : _GEN_18948; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18950 = 12'h1c1 == _T_196[11:0] ? 4'h0 : _GEN_18949; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18951 = 12'h1c2 == _T_196[11:0] ? 4'h0 : _GEN_18950; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18952 = 12'h1c3 == _T_196[11:0] ? image_451 : _GEN_18951; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18953 = 12'h1c4 == _T_196[11:0] ? image_452 : _GEN_18952; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18954 = 12'h1c5 == _T_196[11:0] ? image_453 : _GEN_18953; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18955 = 12'h1c6 == _T_196[11:0] ? image_454 : _GEN_18954; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18956 = 12'h1c7 == _T_196[11:0] ? image_455 : _GEN_18955; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18957 = 12'h1c8 == _T_196[11:0] ? image_456 : _GEN_18956; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18958 = 12'h1c9 == _T_196[11:0] ? image_457 : _GEN_18957; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18959 = 12'h1ca == _T_196[11:0] ? image_458 : _GEN_18958; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18960 = 12'h1cb == _T_196[11:0] ? image_459 : _GEN_18959; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18961 = 12'h1cc == _T_196[11:0] ? image_460 : _GEN_18960; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18962 = 12'h1cd == _T_196[11:0] ? image_461 : _GEN_18961; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18963 = 12'h1ce == _T_196[11:0] ? image_462 : _GEN_18962; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18964 = 12'h1cf == _T_196[11:0] ? image_463 : _GEN_18963; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18965 = 12'h1d0 == _T_196[11:0] ? image_464 : _GEN_18964; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18966 = 12'h1d1 == _T_196[11:0] ? image_465 : _GEN_18965; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18967 = 12'h1d2 == _T_196[11:0] ? image_466 : _GEN_18966; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18968 = 12'h1d3 == _T_196[11:0] ? image_467 : _GEN_18967; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18969 = 12'h1d4 == _T_196[11:0] ? image_468 : _GEN_18968; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18970 = 12'h1d5 == _T_196[11:0] ? image_469 : _GEN_18969; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18971 = 12'h1d6 == _T_196[11:0] ? image_470 : _GEN_18970; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18972 = 12'h1d7 == _T_196[11:0] ? image_471 : _GEN_18971; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18973 = 12'h1d8 == _T_196[11:0] ? image_472 : _GEN_18972; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18974 = 12'h1d9 == _T_196[11:0] ? image_473 : _GEN_18973; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18975 = 12'h1da == _T_196[11:0] ? image_474 : _GEN_18974; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18976 = 12'h1db == _T_196[11:0] ? image_475 : _GEN_18975; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18977 = 12'h1dc == _T_196[11:0] ? image_476 : _GEN_18976; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18978 = 12'h1dd == _T_196[11:0] ? image_477 : _GEN_18977; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18979 = 12'h1de == _T_196[11:0] ? image_478 : _GEN_18978; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18980 = 12'h1df == _T_196[11:0] ? image_479 : _GEN_18979; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18981 = 12'h1e0 == _T_196[11:0] ? image_480 : _GEN_18980; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18982 = 12'h1e1 == _T_196[11:0] ? image_481 : _GEN_18981; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18983 = 12'h1e2 == _T_196[11:0] ? image_482 : _GEN_18982; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18984 = 12'h1e3 == _T_196[11:0] ? image_483 : _GEN_18983; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18985 = 12'h1e4 == _T_196[11:0] ? image_484 : _GEN_18984; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18986 = 12'h1e5 == _T_196[11:0] ? image_485 : _GEN_18985; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18987 = 12'h1e6 == _T_196[11:0] ? image_486 : _GEN_18986; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18988 = 12'h1e7 == _T_196[11:0] ? image_487 : _GEN_18987; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18989 = 12'h1e8 == _T_196[11:0] ? image_488 : _GEN_18988; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18990 = 12'h1e9 == _T_196[11:0] ? image_489 : _GEN_18989; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18991 = 12'h1ea == _T_196[11:0] ? image_490 : _GEN_18990; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18992 = 12'h1eb == _T_196[11:0] ? image_491 : _GEN_18991; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18993 = 12'h1ec == _T_196[11:0] ? image_492 : _GEN_18992; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18994 = 12'h1ed == _T_196[11:0] ? image_493 : _GEN_18993; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18995 = 12'h1ee == _T_196[11:0] ? image_494 : _GEN_18994; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18996 = 12'h1ef == _T_196[11:0] ? image_495 : _GEN_18995; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18997 = 12'h1f0 == _T_196[11:0] ? image_496 : _GEN_18996; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18998 = 12'h1f1 == _T_196[11:0] ? image_497 : _GEN_18997; // @[Filter.scala 138:46]
  wire [3:0] _GEN_18999 = 12'h1f2 == _T_196[11:0] ? image_498 : _GEN_18998; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19000 = 12'h1f3 == _T_196[11:0] ? image_499 : _GEN_18999; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19001 = 12'h1f4 == _T_196[11:0] ? image_500 : _GEN_19000; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19002 = 12'h1f5 == _T_196[11:0] ? image_501 : _GEN_19001; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19003 = 12'h1f6 == _T_196[11:0] ? image_502 : _GEN_19002; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19004 = 12'h1f7 == _T_196[11:0] ? image_503 : _GEN_19003; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19005 = 12'h1f8 == _T_196[11:0] ? image_504 : _GEN_19004; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19006 = 12'h1f9 == _T_196[11:0] ? image_505 : _GEN_19005; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19007 = 12'h1fa == _T_196[11:0] ? image_506 : _GEN_19006; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19008 = 12'h1fb == _T_196[11:0] ? image_507 : _GEN_19007; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19009 = 12'h1fc == _T_196[11:0] ? image_508 : _GEN_19008; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19010 = 12'h1fd == _T_196[11:0] ? image_509 : _GEN_19009; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19011 = 12'h1fe == _T_196[11:0] ? 4'h0 : _GEN_19010; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19012 = 12'h1ff == _T_196[11:0] ? 4'h0 : _GEN_19011; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19013 = 12'h200 == _T_196[11:0] ? 4'h0 : _GEN_19012; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19014 = 12'h201 == _T_196[11:0] ? 4'h0 : _GEN_19013; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19015 = 12'h202 == _T_196[11:0] ? 4'h0 : _GEN_19014; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19016 = 12'h203 == _T_196[11:0] ? image_515 : _GEN_19015; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19017 = 12'h204 == _T_196[11:0] ? image_516 : _GEN_19016; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19018 = 12'h205 == _T_196[11:0] ? image_517 : _GEN_19017; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19019 = 12'h206 == _T_196[11:0] ? image_518 : _GEN_19018; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19020 = 12'h207 == _T_196[11:0] ? image_519 : _GEN_19019; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19021 = 12'h208 == _T_196[11:0] ? image_520 : _GEN_19020; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19022 = 12'h209 == _T_196[11:0] ? image_521 : _GEN_19021; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19023 = 12'h20a == _T_196[11:0] ? image_522 : _GEN_19022; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19024 = 12'h20b == _T_196[11:0] ? image_523 : _GEN_19023; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19025 = 12'h20c == _T_196[11:0] ? image_524 : _GEN_19024; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19026 = 12'h20d == _T_196[11:0] ? image_525 : _GEN_19025; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19027 = 12'h20e == _T_196[11:0] ? image_526 : _GEN_19026; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19028 = 12'h20f == _T_196[11:0] ? image_527 : _GEN_19027; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19029 = 12'h210 == _T_196[11:0] ? image_528 : _GEN_19028; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19030 = 12'h211 == _T_196[11:0] ? image_529 : _GEN_19029; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19031 = 12'h212 == _T_196[11:0] ? image_530 : _GEN_19030; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19032 = 12'h213 == _T_196[11:0] ? image_531 : _GEN_19031; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19033 = 12'h214 == _T_196[11:0] ? image_532 : _GEN_19032; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19034 = 12'h215 == _T_196[11:0] ? image_533 : _GEN_19033; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19035 = 12'h216 == _T_196[11:0] ? image_534 : _GEN_19034; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19036 = 12'h217 == _T_196[11:0] ? image_535 : _GEN_19035; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19037 = 12'h218 == _T_196[11:0] ? image_536 : _GEN_19036; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19038 = 12'h219 == _T_196[11:0] ? image_537 : _GEN_19037; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19039 = 12'h21a == _T_196[11:0] ? image_538 : _GEN_19038; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19040 = 12'h21b == _T_196[11:0] ? image_539 : _GEN_19039; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19041 = 12'h21c == _T_196[11:0] ? image_540 : _GEN_19040; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19042 = 12'h21d == _T_196[11:0] ? image_541 : _GEN_19041; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19043 = 12'h21e == _T_196[11:0] ? image_542 : _GEN_19042; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19044 = 12'h21f == _T_196[11:0] ? image_543 : _GEN_19043; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19045 = 12'h220 == _T_196[11:0] ? image_544 : _GEN_19044; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19046 = 12'h221 == _T_196[11:0] ? image_545 : _GEN_19045; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19047 = 12'h222 == _T_196[11:0] ? image_546 : _GEN_19046; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19048 = 12'h223 == _T_196[11:0] ? image_547 : _GEN_19047; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19049 = 12'h224 == _T_196[11:0] ? image_548 : _GEN_19048; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19050 = 12'h225 == _T_196[11:0] ? image_549 : _GEN_19049; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19051 = 12'h226 == _T_196[11:0] ? image_550 : _GEN_19050; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19052 = 12'h227 == _T_196[11:0] ? image_551 : _GEN_19051; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19053 = 12'h228 == _T_196[11:0] ? image_552 : _GEN_19052; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19054 = 12'h229 == _T_196[11:0] ? image_553 : _GEN_19053; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19055 = 12'h22a == _T_196[11:0] ? image_554 : _GEN_19054; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19056 = 12'h22b == _T_196[11:0] ? image_555 : _GEN_19055; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19057 = 12'h22c == _T_196[11:0] ? image_556 : _GEN_19056; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19058 = 12'h22d == _T_196[11:0] ? image_557 : _GEN_19057; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19059 = 12'h22e == _T_196[11:0] ? image_558 : _GEN_19058; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19060 = 12'h22f == _T_196[11:0] ? image_559 : _GEN_19059; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19061 = 12'h230 == _T_196[11:0] ? image_560 : _GEN_19060; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19062 = 12'h231 == _T_196[11:0] ? image_561 : _GEN_19061; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19063 = 12'h232 == _T_196[11:0] ? image_562 : _GEN_19062; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19064 = 12'h233 == _T_196[11:0] ? image_563 : _GEN_19063; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19065 = 12'h234 == _T_196[11:0] ? image_564 : _GEN_19064; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19066 = 12'h235 == _T_196[11:0] ? image_565 : _GEN_19065; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19067 = 12'h236 == _T_196[11:0] ? image_566 : _GEN_19066; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19068 = 12'h237 == _T_196[11:0] ? 4'h0 : _GEN_19067; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19069 = 12'h238 == _T_196[11:0] ? 4'h0 : _GEN_19068; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19070 = 12'h239 == _T_196[11:0] ? 4'h0 : _GEN_19069; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19071 = 12'h23a == _T_196[11:0] ? 4'h0 : _GEN_19070; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19072 = 12'h23b == _T_196[11:0] ? image_571 : _GEN_19071; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19073 = 12'h23c == _T_196[11:0] ? image_572 : _GEN_19072; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19074 = 12'h23d == _T_196[11:0] ? image_573 : _GEN_19073; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19075 = 12'h23e == _T_196[11:0] ? image_574 : _GEN_19074; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19076 = 12'h23f == _T_196[11:0] ? 4'h0 : _GEN_19075; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19077 = 12'h240 == _T_196[11:0] ? 4'h0 : _GEN_19076; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19078 = 12'h241 == _T_196[11:0] ? 4'h0 : _GEN_19077; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19079 = 12'h242 == _T_196[11:0] ? image_578 : _GEN_19078; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19080 = 12'h243 == _T_196[11:0] ? image_579 : _GEN_19079; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19081 = 12'h244 == _T_196[11:0] ? image_580 : _GEN_19080; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19082 = 12'h245 == _T_196[11:0] ? image_581 : _GEN_19081; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19083 = 12'h246 == _T_196[11:0] ? image_582 : _GEN_19082; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19084 = 12'h247 == _T_196[11:0] ? image_583 : _GEN_19083; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19085 = 12'h248 == _T_196[11:0] ? image_584 : _GEN_19084; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19086 = 12'h249 == _T_196[11:0] ? image_585 : _GEN_19085; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19087 = 12'h24a == _T_196[11:0] ? image_586 : _GEN_19086; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19088 = 12'h24b == _T_196[11:0] ? image_587 : _GEN_19087; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19089 = 12'h24c == _T_196[11:0] ? image_588 : _GEN_19088; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19090 = 12'h24d == _T_196[11:0] ? image_589 : _GEN_19089; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19091 = 12'h24e == _T_196[11:0] ? image_590 : _GEN_19090; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19092 = 12'h24f == _T_196[11:0] ? image_591 : _GEN_19091; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19093 = 12'h250 == _T_196[11:0] ? image_592 : _GEN_19092; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19094 = 12'h251 == _T_196[11:0] ? image_593 : _GEN_19093; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19095 = 12'h252 == _T_196[11:0] ? image_594 : _GEN_19094; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19096 = 12'h253 == _T_196[11:0] ? image_595 : _GEN_19095; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19097 = 12'h254 == _T_196[11:0] ? image_596 : _GEN_19096; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19098 = 12'h255 == _T_196[11:0] ? image_597 : _GEN_19097; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19099 = 12'h256 == _T_196[11:0] ? image_598 : _GEN_19098; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19100 = 12'h257 == _T_196[11:0] ? image_599 : _GEN_19099; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19101 = 12'h258 == _T_196[11:0] ? image_600 : _GEN_19100; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19102 = 12'h259 == _T_196[11:0] ? image_601 : _GEN_19101; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19103 = 12'h25a == _T_196[11:0] ? image_602 : _GEN_19102; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19104 = 12'h25b == _T_196[11:0] ? image_603 : _GEN_19103; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19105 = 12'h25c == _T_196[11:0] ? image_604 : _GEN_19104; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19106 = 12'h25d == _T_196[11:0] ? image_605 : _GEN_19105; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19107 = 12'h25e == _T_196[11:0] ? image_606 : _GEN_19106; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19108 = 12'h25f == _T_196[11:0] ? image_607 : _GEN_19107; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19109 = 12'h260 == _T_196[11:0] ? 4'h0 : _GEN_19108; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19110 = 12'h261 == _T_196[11:0] ? 4'h0 : _GEN_19109; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19111 = 12'h262 == _T_196[11:0] ? 4'h0 : _GEN_19110; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19112 = 12'h263 == _T_196[11:0] ? 4'h0 : _GEN_19111; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19113 = 12'h264 == _T_196[11:0] ? 4'h0 : _GEN_19112; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19114 = 12'h265 == _T_196[11:0] ? 4'h0 : _GEN_19113; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19115 = 12'h266 == _T_196[11:0] ? image_614 : _GEN_19114; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19116 = 12'h267 == _T_196[11:0] ? image_615 : _GEN_19115; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19117 = 12'h268 == _T_196[11:0] ? image_616 : _GEN_19116; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19118 = 12'h269 == _T_196[11:0] ? image_617 : _GEN_19117; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19119 = 12'h26a == _T_196[11:0] ? image_618 : _GEN_19118; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19120 = 12'h26b == _T_196[11:0] ? image_619 : _GEN_19119; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19121 = 12'h26c == _T_196[11:0] ? image_620 : _GEN_19120; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19122 = 12'h26d == _T_196[11:0] ? image_621 : _GEN_19121; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19123 = 12'h26e == _T_196[11:0] ? image_622 : _GEN_19122; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19124 = 12'h26f == _T_196[11:0] ? image_623 : _GEN_19123; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19125 = 12'h270 == _T_196[11:0] ? image_624 : _GEN_19124; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19126 = 12'h271 == _T_196[11:0] ? image_625 : _GEN_19125; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19127 = 12'h272 == _T_196[11:0] ? image_626 : _GEN_19126; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19128 = 12'h273 == _T_196[11:0] ? image_627 : _GEN_19127; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19129 = 12'h274 == _T_196[11:0] ? image_628 : _GEN_19128; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19130 = 12'h275 == _T_196[11:0] ? 4'h0 : _GEN_19129; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19131 = 12'h276 == _T_196[11:0] ? 4'h0 : _GEN_19130; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19132 = 12'h277 == _T_196[11:0] ? 4'h0 : _GEN_19131; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19133 = 12'h278 == _T_196[11:0] ? 4'h0 : _GEN_19132; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19134 = 12'h279 == _T_196[11:0] ? 4'h0 : _GEN_19133; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19135 = 12'h27a == _T_196[11:0] ? 4'h0 : _GEN_19134; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19136 = 12'h27b == _T_196[11:0] ? 4'h0 : _GEN_19135; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19137 = 12'h27c == _T_196[11:0] ? image_636 : _GEN_19136; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19138 = 12'h27d == _T_196[11:0] ? image_637 : _GEN_19137; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19139 = 12'h27e == _T_196[11:0] ? image_638 : _GEN_19138; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19140 = 12'h27f == _T_196[11:0] ? image_639 : _GEN_19139; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19141 = 12'h280 == _T_196[11:0] ? 4'h0 : _GEN_19140; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19142 = 12'h281 == _T_196[11:0] ? 4'h0 : _GEN_19141; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19143 = 12'h282 == _T_196[11:0] ? image_642 : _GEN_19142; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19144 = 12'h283 == _T_196[11:0] ? image_643 : _GEN_19143; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19145 = 12'h284 == _T_196[11:0] ? image_644 : _GEN_19144; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19146 = 12'h285 == _T_196[11:0] ? image_645 : _GEN_19145; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19147 = 12'h286 == _T_196[11:0] ? image_646 : _GEN_19146; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19148 = 12'h287 == _T_196[11:0] ? image_647 : _GEN_19147; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19149 = 12'h288 == _T_196[11:0] ? image_648 : _GEN_19148; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19150 = 12'h289 == _T_196[11:0] ? image_649 : _GEN_19149; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19151 = 12'h28a == _T_196[11:0] ? image_650 : _GEN_19150; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19152 = 12'h28b == _T_196[11:0] ? image_651 : _GEN_19151; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19153 = 12'h28c == _T_196[11:0] ? image_652 : _GEN_19152; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19154 = 12'h28d == _T_196[11:0] ? image_653 : _GEN_19153; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19155 = 12'h28e == _T_196[11:0] ? image_654 : _GEN_19154; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19156 = 12'h28f == _T_196[11:0] ? image_655 : _GEN_19155; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19157 = 12'h290 == _T_196[11:0] ? image_656 : _GEN_19156; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19158 = 12'h291 == _T_196[11:0] ? image_657 : _GEN_19157; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19159 = 12'h292 == _T_196[11:0] ? image_658 : _GEN_19158; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19160 = 12'h293 == _T_196[11:0] ? image_659 : _GEN_19159; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19161 = 12'h294 == _T_196[11:0] ? image_660 : _GEN_19160; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19162 = 12'h295 == _T_196[11:0] ? image_661 : _GEN_19161; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19163 = 12'h296 == _T_196[11:0] ? image_662 : _GEN_19162; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19164 = 12'h297 == _T_196[11:0] ? image_663 : _GEN_19163; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19165 = 12'h298 == _T_196[11:0] ? image_664 : _GEN_19164; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19166 = 12'h299 == _T_196[11:0] ? image_665 : _GEN_19165; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19167 = 12'h29a == _T_196[11:0] ? image_666 : _GEN_19166; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19168 = 12'h29b == _T_196[11:0] ? image_667 : _GEN_19167; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19169 = 12'h29c == _T_196[11:0] ? image_668 : _GEN_19168; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19170 = 12'h29d == _T_196[11:0] ? image_669 : _GEN_19169; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19171 = 12'h29e == _T_196[11:0] ? image_670 : _GEN_19170; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19172 = 12'h29f == _T_196[11:0] ? 4'h0 : _GEN_19171; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19173 = 12'h2a0 == _T_196[11:0] ? 4'h0 : _GEN_19172; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19174 = 12'h2a1 == _T_196[11:0] ? 4'h0 : _GEN_19173; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19175 = 12'h2a2 == _T_196[11:0] ? 4'h0 : _GEN_19174; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19176 = 12'h2a3 == _T_196[11:0] ? 4'h0 : _GEN_19175; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19177 = 12'h2a4 == _T_196[11:0] ? 4'h0 : _GEN_19176; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19178 = 12'h2a5 == _T_196[11:0] ? 4'h0 : _GEN_19177; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19179 = 12'h2a6 == _T_196[11:0] ? 4'h0 : _GEN_19178; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19180 = 12'h2a7 == _T_196[11:0] ? image_679 : _GEN_19179; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19181 = 12'h2a8 == _T_196[11:0] ? image_680 : _GEN_19180; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19182 = 12'h2a9 == _T_196[11:0] ? image_681 : _GEN_19181; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19183 = 12'h2aa == _T_196[11:0] ? image_682 : _GEN_19182; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19184 = 12'h2ab == _T_196[11:0] ? image_683 : _GEN_19183; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19185 = 12'h2ac == _T_196[11:0] ? image_684 : _GEN_19184; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19186 = 12'h2ad == _T_196[11:0] ? image_685 : _GEN_19185; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19187 = 12'h2ae == _T_196[11:0] ? image_686 : _GEN_19186; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19188 = 12'h2af == _T_196[11:0] ? image_687 : _GEN_19187; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19189 = 12'h2b0 == _T_196[11:0] ? image_688 : _GEN_19188; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19190 = 12'h2b1 == _T_196[11:0] ? image_689 : _GEN_19189; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19191 = 12'h2b2 == _T_196[11:0] ? image_690 : _GEN_19190; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19192 = 12'h2b3 == _T_196[11:0] ? image_691 : _GEN_19191; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19193 = 12'h2b4 == _T_196[11:0] ? image_692 : _GEN_19192; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19194 = 12'h2b5 == _T_196[11:0] ? image_693 : _GEN_19193; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19195 = 12'h2b6 == _T_196[11:0] ? image_694 : _GEN_19194; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19196 = 12'h2b7 == _T_196[11:0] ? image_695 : _GEN_19195; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19197 = 12'h2b8 == _T_196[11:0] ? image_696 : _GEN_19196; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19198 = 12'h2b9 == _T_196[11:0] ? image_697 : _GEN_19197; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19199 = 12'h2ba == _T_196[11:0] ? image_698 : _GEN_19198; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19200 = 12'h2bb == _T_196[11:0] ? 4'h0 : _GEN_19199; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19201 = 12'h2bc == _T_196[11:0] ? 4'h0 : _GEN_19200; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19202 = 12'h2bd == _T_196[11:0] ? image_701 : _GEN_19201; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19203 = 12'h2be == _T_196[11:0] ? image_702 : _GEN_19202; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19204 = 12'h2bf == _T_196[11:0] ? image_703 : _GEN_19203; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19205 = 12'h2c0 == _T_196[11:0] ? 4'h0 : _GEN_19204; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19206 = 12'h2c1 == _T_196[11:0] ? image_705 : _GEN_19205; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19207 = 12'h2c2 == _T_196[11:0] ? image_706 : _GEN_19206; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19208 = 12'h2c3 == _T_196[11:0] ? image_707 : _GEN_19207; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19209 = 12'h2c4 == _T_196[11:0] ? image_708 : _GEN_19208; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19210 = 12'h2c5 == _T_196[11:0] ? image_709 : _GEN_19209; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19211 = 12'h2c6 == _T_196[11:0] ? image_710 : _GEN_19210; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19212 = 12'h2c7 == _T_196[11:0] ? image_711 : _GEN_19211; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19213 = 12'h2c8 == _T_196[11:0] ? image_712 : _GEN_19212; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19214 = 12'h2c9 == _T_196[11:0] ? image_713 : _GEN_19213; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19215 = 12'h2ca == _T_196[11:0] ? image_714 : _GEN_19214; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19216 = 12'h2cb == _T_196[11:0] ? image_715 : _GEN_19215; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19217 = 12'h2cc == _T_196[11:0] ? image_716 : _GEN_19216; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19218 = 12'h2cd == _T_196[11:0] ? image_717 : _GEN_19217; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19219 = 12'h2ce == _T_196[11:0] ? image_718 : _GEN_19218; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19220 = 12'h2cf == _T_196[11:0] ? image_719 : _GEN_19219; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19221 = 12'h2d0 == _T_196[11:0] ? image_720 : _GEN_19220; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19222 = 12'h2d1 == _T_196[11:0] ? image_721 : _GEN_19221; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19223 = 12'h2d2 == _T_196[11:0] ? image_722 : _GEN_19222; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19224 = 12'h2d3 == _T_196[11:0] ? image_723 : _GEN_19223; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19225 = 12'h2d4 == _T_196[11:0] ? image_724 : _GEN_19224; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19226 = 12'h2d5 == _T_196[11:0] ? image_725 : _GEN_19225; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19227 = 12'h2d6 == _T_196[11:0] ? image_726 : _GEN_19226; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19228 = 12'h2d7 == _T_196[11:0] ? image_727 : _GEN_19227; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19229 = 12'h2d8 == _T_196[11:0] ? image_728 : _GEN_19228; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19230 = 12'h2d9 == _T_196[11:0] ? image_729 : _GEN_19229; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19231 = 12'h2da == _T_196[11:0] ? image_730 : _GEN_19230; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19232 = 12'h2db == _T_196[11:0] ? image_731 : _GEN_19231; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19233 = 12'h2dc == _T_196[11:0] ? image_732 : _GEN_19232; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19234 = 12'h2dd == _T_196[11:0] ? image_733 : _GEN_19233; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19235 = 12'h2de == _T_196[11:0] ? image_734 : _GEN_19234; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19236 = 12'h2df == _T_196[11:0] ? 4'h0 : _GEN_19235; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19237 = 12'h2e0 == _T_196[11:0] ? image_736 : _GEN_19236; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19238 = 12'h2e1 == _T_196[11:0] ? image_737 : _GEN_19237; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19239 = 12'h2e2 == _T_196[11:0] ? 4'h0 : _GEN_19238; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19240 = 12'h2e3 == _T_196[11:0] ? image_739 : _GEN_19239; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19241 = 12'h2e4 == _T_196[11:0] ? image_740 : _GEN_19240; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19242 = 12'h2e5 == _T_196[11:0] ? image_741 : _GEN_19241; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19243 = 12'h2e6 == _T_196[11:0] ? 4'h0 : _GEN_19242; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19244 = 12'h2e7 == _T_196[11:0] ? 4'h0 : _GEN_19243; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19245 = 12'h2e8 == _T_196[11:0] ? image_744 : _GEN_19244; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19246 = 12'h2e9 == _T_196[11:0] ? image_745 : _GEN_19245; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19247 = 12'h2ea == _T_196[11:0] ? image_746 : _GEN_19246; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19248 = 12'h2eb == _T_196[11:0] ? image_747 : _GEN_19247; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19249 = 12'h2ec == _T_196[11:0] ? image_748 : _GEN_19248; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19250 = 12'h2ed == _T_196[11:0] ? image_749 : _GEN_19249; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19251 = 12'h2ee == _T_196[11:0] ? image_750 : _GEN_19250; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19252 = 12'h2ef == _T_196[11:0] ? image_751 : _GEN_19251; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19253 = 12'h2f0 == _T_196[11:0] ? image_752 : _GEN_19252; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19254 = 12'h2f1 == _T_196[11:0] ? image_753 : _GEN_19253; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19255 = 12'h2f2 == _T_196[11:0] ? image_754 : _GEN_19254; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19256 = 12'h2f3 == _T_196[11:0] ? image_755 : _GEN_19255; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19257 = 12'h2f4 == _T_196[11:0] ? image_756 : _GEN_19256; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19258 = 12'h2f5 == _T_196[11:0] ? 4'h0 : _GEN_19257; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19259 = 12'h2f6 == _T_196[11:0] ? image_758 : _GEN_19258; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19260 = 12'h2f7 == _T_196[11:0] ? 4'h0 : _GEN_19259; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19261 = 12'h2f8 == _T_196[11:0] ? image_760 : _GEN_19260; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19262 = 12'h2f9 == _T_196[11:0] ? image_761 : _GEN_19261; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19263 = 12'h2fa == _T_196[11:0] ? image_762 : _GEN_19262; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19264 = 12'h2fb == _T_196[11:0] ? image_763 : _GEN_19263; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19265 = 12'h2fc == _T_196[11:0] ? 4'h0 : _GEN_19264; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19266 = 12'h2fd == _T_196[11:0] ? image_765 : _GEN_19265; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19267 = 12'h2fe == _T_196[11:0] ? image_766 : _GEN_19266; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19268 = 12'h2ff == _T_196[11:0] ? image_767 : _GEN_19267; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19269 = 12'h300 == _T_196[11:0] ? image_768 : _GEN_19268; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19270 = 12'h301 == _T_196[11:0] ? image_769 : _GEN_19269; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19271 = 12'h302 == _T_196[11:0] ? image_770 : _GEN_19270; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19272 = 12'h303 == _T_196[11:0] ? image_771 : _GEN_19271; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19273 = 12'h304 == _T_196[11:0] ? image_772 : _GEN_19272; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19274 = 12'h305 == _T_196[11:0] ? image_773 : _GEN_19273; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19275 = 12'h306 == _T_196[11:0] ? image_774 : _GEN_19274; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19276 = 12'h307 == _T_196[11:0] ? image_775 : _GEN_19275; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19277 = 12'h308 == _T_196[11:0] ? image_776 : _GEN_19276; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19278 = 12'h309 == _T_196[11:0] ? image_777 : _GEN_19277; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19279 = 12'h30a == _T_196[11:0] ? image_778 : _GEN_19278; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19280 = 12'h30b == _T_196[11:0] ? image_779 : _GEN_19279; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19281 = 12'h30c == _T_196[11:0] ? image_780 : _GEN_19280; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19282 = 12'h30d == _T_196[11:0] ? image_781 : _GEN_19281; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19283 = 12'h30e == _T_196[11:0] ? image_782 : _GEN_19282; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19284 = 12'h30f == _T_196[11:0] ? image_783 : _GEN_19283; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19285 = 12'h310 == _T_196[11:0] ? image_784 : _GEN_19284; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19286 = 12'h311 == _T_196[11:0] ? image_785 : _GEN_19285; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19287 = 12'h312 == _T_196[11:0] ? image_786 : _GEN_19286; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19288 = 12'h313 == _T_196[11:0] ? image_787 : _GEN_19287; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19289 = 12'h314 == _T_196[11:0] ? image_788 : _GEN_19288; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19290 = 12'h315 == _T_196[11:0] ? image_789 : _GEN_19289; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19291 = 12'h316 == _T_196[11:0] ? image_790 : _GEN_19290; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19292 = 12'h317 == _T_196[11:0] ? image_791 : _GEN_19291; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19293 = 12'h318 == _T_196[11:0] ? image_792 : _GEN_19292; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19294 = 12'h319 == _T_196[11:0] ? image_793 : _GEN_19293; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19295 = 12'h31a == _T_196[11:0] ? image_794 : _GEN_19294; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19296 = 12'h31b == _T_196[11:0] ? image_795 : _GEN_19295; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19297 = 12'h31c == _T_196[11:0] ? image_796 : _GEN_19296; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19298 = 12'h31d == _T_196[11:0] ? image_797 : _GEN_19297; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19299 = 12'h31e == _T_196[11:0] ? 4'h0 : _GEN_19298; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19300 = 12'h31f == _T_196[11:0] ? 4'h0 : _GEN_19299; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19301 = 12'h320 == _T_196[11:0] ? image_800 : _GEN_19300; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19302 = 12'h321 == _T_196[11:0] ? image_801 : _GEN_19301; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19303 = 12'h322 == _T_196[11:0] ? image_802 : _GEN_19302; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19304 = 12'h323 == _T_196[11:0] ? image_803 : _GEN_19303; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19305 = 12'h324 == _T_196[11:0] ? image_804 : _GEN_19304; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19306 = 12'h325 == _T_196[11:0] ? image_805 : _GEN_19305; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19307 = 12'h326 == _T_196[11:0] ? image_806 : _GEN_19306; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19308 = 12'h327 == _T_196[11:0] ? 4'h0 : _GEN_19307; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19309 = 12'h328 == _T_196[11:0] ? image_808 : _GEN_19308; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19310 = 12'h329 == _T_196[11:0] ? image_809 : _GEN_19309; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19311 = 12'h32a == _T_196[11:0] ? image_810 : _GEN_19310; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19312 = 12'h32b == _T_196[11:0] ? image_811 : _GEN_19311; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19313 = 12'h32c == _T_196[11:0] ? image_812 : _GEN_19312; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19314 = 12'h32d == _T_196[11:0] ? image_813 : _GEN_19313; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19315 = 12'h32e == _T_196[11:0] ? image_814 : _GEN_19314; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19316 = 12'h32f == _T_196[11:0] ? image_815 : _GEN_19315; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19317 = 12'h330 == _T_196[11:0] ? image_816 : _GEN_19316; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19318 = 12'h331 == _T_196[11:0] ? image_817 : _GEN_19317; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19319 = 12'h332 == _T_196[11:0] ? image_818 : _GEN_19318; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19320 = 12'h333 == _T_196[11:0] ? image_819 : _GEN_19319; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19321 = 12'h334 == _T_196[11:0] ? image_820 : _GEN_19320; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19322 = 12'h335 == _T_196[11:0] ? 4'h0 : _GEN_19321; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19323 = 12'h336 == _T_196[11:0] ? image_822 : _GEN_19322; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19324 = 12'h337 == _T_196[11:0] ? image_823 : _GEN_19323; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19325 = 12'h338 == _T_196[11:0] ? image_824 : _GEN_19324; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19326 = 12'h339 == _T_196[11:0] ? image_825 : _GEN_19325; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19327 = 12'h33a == _T_196[11:0] ? image_826 : _GEN_19326; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19328 = 12'h33b == _T_196[11:0] ? 4'h0 : _GEN_19327; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19329 = 12'h33c == _T_196[11:0] ? image_828 : _GEN_19328; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19330 = 12'h33d == _T_196[11:0] ? image_829 : _GEN_19329; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19331 = 12'h33e == _T_196[11:0] ? image_830 : _GEN_19330; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19332 = 12'h33f == _T_196[11:0] ? image_831 : _GEN_19331; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19333 = 12'h340 == _T_196[11:0] ? 4'h0 : _GEN_19332; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19334 = 12'h341 == _T_196[11:0] ? image_833 : _GEN_19333; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19335 = 12'h342 == _T_196[11:0] ? image_834 : _GEN_19334; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19336 = 12'h343 == _T_196[11:0] ? image_835 : _GEN_19335; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19337 = 12'h344 == _T_196[11:0] ? image_836 : _GEN_19336; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19338 = 12'h345 == _T_196[11:0] ? image_837 : _GEN_19337; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19339 = 12'h346 == _T_196[11:0] ? image_838 : _GEN_19338; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19340 = 12'h347 == _T_196[11:0] ? image_839 : _GEN_19339; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19341 = 12'h348 == _T_196[11:0] ? image_840 : _GEN_19340; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19342 = 12'h349 == _T_196[11:0] ? image_841 : _GEN_19341; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19343 = 12'h34a == _T_196[11:0] ? image_842 : _GEN_19342; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19344 = 12'h34b == _T_196[11:0] ? image_843 : _GEN_19343; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19345 = 12'h34c == _T_196[11:0] ? image_844 : _GEN_19344; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19346 = 12'h34d == _T_196[11:0] ? image_845 : _GEN_19345; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19347 = 12'h34e == _T_196[11:0] ? image_846 : _GEN_19346; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19348 = 12'h34f == _T_196[11:0] ? image_847 : _GEN_19347; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19349 = 12'h350 == _T_196[11:0] ? image_848 : _GEN_19348; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19350 = 12'h351 == _T_196[11:0] ? image_849 : _GEN_19349; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19351 = 12'h352 == _T_196[11:0] ? image_850 : _GEN_19350; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19352 = 12'h353 == _T_196[11:0] ? image_851 : _GEN_19351; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19353 = 12'h354 == _T_196[11:0] ? image_852 : _GEN_19352; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19354 = 12'h355 == _T_196[11:0] ? image_853 : _GEN_19353; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19355 = 12'h356 == _T_196[11:0] ? image_854 : _GEN_19354; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19356 = 12'h357 == _T_196[11:0] ? image_855 : _GEN_19355; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19357 = 12'h358 == _T_196[11:0] ? image_856 : _GEN_19356; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19358 = 12'h359 == _T_196[11:0] ? image_857 : _GEN_19357; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19359 = 12'h35a == _T_196[11:0] ? image_858 : _GEN_19358; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19360 = 12'h35b == _T_196[11:0] ? image_859 : _GEN_19359; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19361 = 12'h35c == _T_196[11:0] ? image_860 : _GEN_19360; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19362 = 12'h35d == _T_196[11:0] ? image_861 : _GEN_19361; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19363 = 12'h35e == _T_196[11:0] ? image_862 : _GEN_19362; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19364 = 12'h35f == _T_196[11:0] ? 4'h0 : _GEN_19363; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19365 = 12'h360 == _T_196[11:0] ? 4'h0 : _GEN_19364; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19366 = 12'h361 == _T_196[11:0] ? image_865 : _GEN_19365; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19367 = 12'h362 == _T_196[11:0] ? image_866 : _GEN_19366; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19368 = 12'h363 == _T_196[11:0] ? image_867 : _GEN_19367; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19369 = 12'h364 == _T_196[11:0] ? image_868 : _GEN_19368; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19370 = 12'h365 == _T_196[11:0] ? image_869 : _GEN_19369; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19371 = 12'h366 == _T_196[11:0] ? 4'h0 : _GEN_19370; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19372 = 12'h367 == _T_196[11:0] ? 4'h0 : _GEN_19371; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19373 = 12'h368 == _T_196[11:0] ? image_872 : _GEN_19372; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19374 = 12'h369 == _T_196[11:0] ? image_873 : _GEN_19373; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19375 = 12'h36a == _T_196[11:0] ? image_874 : _GEN_19374; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19376 = 12'h36b == _T_196[11:0] ? image_875 : _GEN_19375; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19377 = 12'h36c == _T_196[11:0] ? image_876 : _GEN_19376; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19378 = 12'h36d == _T_196[11:0] ? image_877 : _GEN_19377; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19379 = 12'h36e == _T_196[11:0] ? image_878 : _GEN_19378; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19380 = 12'h36f == _T_196[11:0] ? image_879 : _GEN_19379; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19381 = 12'h370 == _T_196[11:0] ? image_880 : _GEN_19380; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19382 = 12'h371 == _T_196[11:0] ? image_881 : _GEN_19381; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19383 = 12'h372 == _T_196[11:0] ? image_882 : _GEN_19382; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19384 = 12'h373 == _T_196[11:0] ? image_883 : _GEN_19383; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19385 = 12'h374 == _T_196[11:0] ? image_884 : _GEN_19384; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19386 = 12'h375 == _T_196[11:0] ? image_885 : _GEN_19385; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19387 = 12'h376 == _T_196[11:0] ? 4'h0 : _GEN_19386; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19388 = 12'h377 == _T_196[11:0] ? 4'h0 : _GEN_19387; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19389 = 12'h378 == _T_196[11:0] ? 4'h0 : _GEN_19388; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19390 = 12'h379 == _T_196[11:0] ? 4'h0 : _GEN_19389; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19391 = 12'h37a == _T_196[11:0] ? 4'h0 : _GEN_19390; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19392 = 12'h37b == _T_196[11:0] ? image_891 : _GEN_19391; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19393 = 12'h37c == _T_196[11:0] ? image_892 : _GEN_19392; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19394 = 12'h37d == _T_196[11:0] ? image_893 : _GEN_19393; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19395 = 12'h37e == _T_196[11:0] ? image_894 : _GEN_19394; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19396 = 12'h37f == _T_196[11:0] ? image_895 : _GEN_19395; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19397 = 12'h380 == _T_196[11:0] ? 4'h0 : _GEN_19396; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19398 = 12'h381 == _T_196[11:0] ? image_897 : _GEN_19397; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19399 = 12'h382 == _T_196[11:0] ? image_898 : _GEN_19398; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19400 = 12'h383 == _T_196[11:0] ? image_899 : _GEN_19399; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19401 = 12'h384 == _T_196[11:0] ? image_900 : _GEN_19400; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19402 = 12'h385 == _T_196[11:0] ? image_901 : _GEN_19401; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19403 = 12'h386 == _T_196[11:0] ? image_902 : _GEN_19402; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19404 = 12'h387 == _T_196[11:0] ? image_903 : _GEN_19403; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19405 = 12'h388 == _T_196[11:0] ? image_904 : _GEN_19404; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19406 = 12'h389 == _T_196[11:0] ? image_905 : _GEN_19405; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19407 = 12'h38a == _T_196[11:0] ? image_906 : _GEN_19406; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19408 = 12'h38b == _T_196[11:0] ? image_907 : _GEN_19407; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19409 = 12'h38c == _T_196[11:0] ? image_908 : _GEN_19408; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19410 = 12'h38d == _T_196[11:0] ? image_909 : _GEN_19409; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19411 = 12'h38e == _T_196[11:0] ? image_910 : _GEN_19410; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19412 = 12'h38f == _T_196[11:0] ? image_911 : _GEN_19411; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19413 = 12'h390 == _T_196[11:0] ? image_912 : _GEN_19412; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19414 = 12'h391 == _T_196[11:0] ? image_913 : _GEN_19413; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19415 = 12'h392 == _T_196[11:0] ? image_914 : _GEN_19414; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19416 = 12'h393 == _T_196[11:0] ? image_915 : _GEN_19415; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19417 = 12'h394 == _T_196[11:0] ? image_916 : _GEN_19416; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19418 = 12'h395 == _T_196[11:0] ? image_917 : _GEN_19417; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19419 = 12'h396 == _T_196[11:0] ? image_918 : _GEN_19418; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19420 = 12'h397 == _T_196[11:0] ? image_919 : _GEN_19419; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19421 = 12'h398 == _T_196[11:0] ? image_920 : _GEN_19420; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19422 = 12'h399 == _T_196[11:0] ? image_921 : _GEN_19421; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19423 = 12'h39a == _T_196[11:0] ? image_922 : _GEN_19422; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19424 = 12'h39b == _T_196[11:0] ? image_923 : _GEN_19423; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19425 = 12'h39c == _T_196[11:0] ? image_924 : _GEN_19424; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19426 = 12'h39d == _T_196[11:0] ? image_925 : _GEN_19425; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19427 = 12'h39e == _T_196[11:0] ? image_926 : _GEN_19426; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19428 = 12'h39f == _T_196[11:0] ? image_927 : _GEN_19427; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19429 = 12'h3a0 == _T_196[11:0] ? 4'h0 : _GEN_19428; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19430 = 12'h3a1 == _T_196[11:0] ? image_929 : _GEN_19429; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19431 = 12'h3a2 == _T_196[11:0] ? image_930 : _GEN_19430; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19432 = 12'h3a3 == _T_196[11:0] ? 4'h0 : _GEN_19431; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19433 = 12'h3a4 == _T_196[11:0] ? 4'h0 : _GEN_19432; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19434 = 12'h3a5 == _T_196[11:0] ? 4'h0 : _GEN_19433; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19435 = 12'h3a6 == _T_196[11:0] ? 4'h0 : _GEN_19434; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19436 = 12'h3a7 == _T_196[11:0] ? image_935 : _GEN_19435; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19437 = 12'h3a8 == _T_196[11:0] ? image_936 : _GEN_19436; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19438 = 12'h3a9 == _T_196[11:0] ? image_937 : _GEN_19437; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19439 = 12'h3aa == _T_196[11:0] ? image_938 : _GEN_19438; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19440 = 12'h3ab == _T_196[11:0] ? image_939 : _GEN_19439; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19441 = 12'h3ac == _T_196[11:0] ? image_940 : _GEN_19440; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19442 = 12'h3ad == _T_196[11:0] ? image_941 : _GEN_19441; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19443 = 12'h3ae == _T_196[11:0] ? image_942 : _GEN_19442; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19444 = 12'h3af == _T_196[11:0] ? image_943 : _GEN_19443; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19445 = 12'h3b0 == _T_196[11:0] ? image_944 : _GEN_19444; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19446 = 12'h3b1 == _T_196[11:0] ? image_945 : _GEN_19445; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19447 = 12'h3b2 == _T_196[11:0] ? image_946 : _GEN_19446; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19448 = 12'h3b3 == _T_196[11:0] ? image_947 : _GEN_19447; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19449 = 12'h3b4 == _T_196[11:0] ? image_948 : _GEN_19448; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19450 = 12'h3b5 == _T_196[11:0] ? image_949 : _GEN_19449; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19451 = 12'h3b6 == _T_196[11:0] ? image_950 : _GEN_19450; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19452 = 12'h3b7 == _T_196[11:0] ? image_951 : _GEN_19451; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19453 = 12'h3b8 == _T_196[11:0] ? image_952 : _GEN_19452; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19454 = 12'h3b9 == _T_196[11:0] ? image_953 : _GEN_19453; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19455 = 12'h3ba == _T_196[11:0] ? image_954 : _GEN_19454; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19456 = 12'h3bb == _T_196[11:0] ? image_955 : _GEN_19455; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19457 = 12'h3bc == _T_196[11:0] ? image_956 : _GEN_19456; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19458 = 12'h3bd == _T_196[11:0] ? image_957 : _GEN_19457; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19459 = 12'h3be == _T_196[11:0] ? image_958 : _GEN_19458; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19460 = 12'h3bf == _T_196[11:0] ? image_959 : _GEN_19459; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19461 = 12'h3c0 == _T_196[11:0] ? 4'h0 : _GEN_19460; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19462 = 12'h3c1 == _T_196[11:0] ? image_961 : _GEN_19461; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19463 = 12'h3c2 == _T_196[11:0] ? image_962 : _GEN_19462; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19464 = 12'h3c3 == _T_196[11:0] ? image_963 : _GEN_19463; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19465 = 12'h3c4 == _T_196[11:0] ? image_964 : _GEN_19464; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19466 = 12'h3c5 == _T_196[11:0] ? image_965 : _GEN_19465; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19467 = 12'h3c6 == _T_196[11:0] ? image_966 : _GEN_19466; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19468 = 12'h3c7 == _T_196[11:0] ? image_967 : _GEN_19467; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19469 = 12'h3c8 == _T_196[11:0] ? image_968 : _GEN_19468; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19470 = 12'h3c9 == _T_196[11:0] ? image_969 : _GEN_19469; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19471 = 12'h3ca == _T_196[11:0] ? image_970 : _GEN_19470; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19472 = 12'h3cb == _T_196[11:0] ? image_971 : _GEN_19471; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19473 = 12'h3cc == _T_196[11:0] ? image_972 : _GEN_19472; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19474 = 12'h3cd == _T_196[11:0] ? image_973 : _GEN_19473; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19475 = 12'h3ce == _T_196[11:0] ? image_974 : _GEN_19474; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19476 = 12'h3cf == _T_196[11:0] ? image_975 : _GEN_19475; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19477 = 12'h3d0 == _T_196[11:0] ? image_976 : _GEN_19476; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19478 = 12'h3d1 == _T_196[11:0] ? image_977 : _GEN_19477; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19479 = 12'h3d2 == _T_196[11:0] ? image_978 : _GEN_19478; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19480 = 12'h3d3 == _T_196[11:0] ? image_979 : _GEN_19479; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19481 = 12'h3d4 == _T_196[11:0] ? image_980 : _GEN_19480; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19482 = 12'h3d5 == _T_196[11:0] ? image_981 : _GEN_19481; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19483 = 12'h3d6 == _T_196[11:0] ? image_982 : _GEN_19482; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19484 = 12'h3d7 == _T_196[11:0] ? image_983 : _GEN_19483; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19485 = 12'h3d8 == _T_196[11:0] ? image_984 : _GEN_19484; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19486 = 12'h3d9 == _T_196[11:0] ? image_985 : _GEN_19485; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19487 = 12'h3da == _T_196[11:0] ? image_986 : _GEN_19486; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19488 = 12'h3db == _T_196[11:0] ? image_987 : _GEN_19487; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19489 = 12'h3dc == _T_196[11:0] ? image_988 : _GEN_19488; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19490 = 12'h3dd == _T_196[11:0] ? image_989 : _GEN_19489; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19491 = 12'h3de == _T_196[11:0] ? image_990 : _GEN_19490; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19492 = 12'h3df == _T_196[11:0] ? image_991 : _GEN_19491; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19493 = 12'h3e0 == _T_196[11:0] ? image_992 : _GEN_19492; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19494 = 12'h3e1 == _T_196[11:0] ? 4'h0 : _GEN_19493; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19495 = 12'h3e2 == _T_196[11:0] ? 4'h0 : _GEN_19494; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19496 = 12'h3e3 == _T_196[11:0] ? 4'h0 : _GEN_19495; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19497 = 12'h3e4 == _T_196[11:0] ? 4'h0 : _GEN_19496; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19498 = 12'h3e5 == _T_196[11:0] ? image_997 : _GEN_19497; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19499 = 12'h3e6 == _T_196[11:0] ? image_998 : _GEN_19498; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19500 = 12'h3e7 == _T_196[11:0] ? image_999 : _GEN_19499; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19501 = 12'h3e8 == _T_196[11:0] ? image_1000 : _GEN_19500; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19502 = 12'h3e9 == _T_196[11:0] ? image_1001 : _GEN_19501; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19503 = 12'h3ea == _T_196[11:0] ? image_1002 : _GEN_19502; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19504 = 12'h3eb == _T_196[11:0] ? image_1003 : _GEN_19503; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19505 = 12'h3ec == _T_196[11:0] ? image_1004 : _GEN_19504; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19506 = 12'h3ed == _T_196[11:0] ? image_1005 : _GEN_19505; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19507 = 12'h3ee == _T_196[11:0] ? image_1006 : _GEN_19506; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19508 = 12'h3ef == _T_196[11:0] ? image_1007 : _GEN_19507; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19509 = 12'h3f0 == _T_196[11:0] ? image_1008 : _GEN_19508; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19510 = 12'h3f1 == _T_196[11:0] ? image_1009 : _GEN_19509; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19511 = 12'h3f2 == _T_196[11:0] ? image_1010 : _GEN_19510; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19512 = 12'h3f3 == _T_196[11:0] ? image_1011 : _GEN_19511; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19513 = 12'h3f4 == _T_196[11:0] ? image_1012 : _GEN_19512; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19514 = 12'h3f5 == _T_196[11:0] ? image_1013 : _GEN_19513; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19515 = 12'h3f6 == _T_196[11:0] ? image_1014 : _GEN_19514; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19516 = 12'h3f7 == _T_196[11:0] ? image_1015 : _GEN_19515; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19517 = 12'h3f8 == _T_196[11:0] ? image_1016 : _GEN_19516; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19518 = 12'h3f9 == _T_196[11:0] ? image_1017 : _GEN_19517; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19519 = 12'h3fa == _T_196[11:0] ? image_1018 : _GEN_19518; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19520 = 12'h3fb == _T_196[11:0] ? image_1019 : _GEN_19519; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19521 = 12'h3fc == _T_196[11:0] ? image_1020 : _GEN_19520; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19522 = 12'h3fd == _T_196[11:0] ? 4'h0 : _GEN_19521; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19523 = 12'h3fe == _T_196[11:0] ? 4'h0 : _GEN_19522; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19524 = 12'h3ff == _T_196[11:0] ? 4'h0 : _GEN_19523; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19525 = 12'h400 == _T_196[11:0] ? image_1024 : _GEN_19524; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19526 = 12'h401 == _T_196[11:0] ? image_1025 : _GEN_19525; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19527 = 12'h402 == _T_196[11:0] ? image_1026 : _GEN_19526; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19528 = 12'h403 == _T_196[11:0] ? image_1027 : _GEN_19527; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19529 = 12'h404 == _T_196[11:0] ? image_1028 : _GEN_19528; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19530 = 12'h405 == _T_196[11:0] ? image_1029 : _GEN_19529; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19531 = 12'h406 == _T_196[11:0] ? image_1030 : _GEN_19530; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19532 = 12'h407 == _T_196[11:0] ? image_1031 : _GEN_19531; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19533 = 12'h408 == _T_196[11:0] ? image_1032 : _GEN_19532; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19534 = 12'h409 == _T_196[11:0] ? image_1033 : _GEN_19533; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19535 = 12'h40a == _T_196[11:0] ? image_1034 : _GEN_19534; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19536 = 12'h40b == _T_196[11:0] ? image_1035 : _GEN_19535; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19537 = 12'h40c == _T_196[11:0] ? image_1036 : _GEN_19536; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19538 = 12'h40d == _T_196[11:0] ? image_1037 : _GEN_19537; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19539 = 12'h40e == _T_196[11:0] ? image_1038 : _GEN_19538; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19540 = 12'h40f == _T_196[11:0] ? image_1039 : _GEN_19539; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19541 = 12'h410 == _T_196[11:0] ? image_1040 : _GEN_19540; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19542 = 12'h411 == _T_196[11:0] ? image_1041 : _GEN_19541; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19543 = 12'h412 == _T_196[11:0] ? image_1042 : _GEN_19542; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19544 = 12'h413 == _T_196[11:0] ? image_1043 : _GEN_19543; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19545 = 12'h414 == _T_196[11:0] ? image_1044 : _GEN_19544; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19546 = 12'h415 == _T_196[11:0] ? image_1045 : _GEN_19545; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19547 = 12'h416 == _T_196[11:0] ? image_1046 : _GEN_19546; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19548 = 12'h417 == _T_196[11:0] ? image_1047 : _GEN_19547; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19549 = 12'h418 == _T_196[11:0] ? image_1048 : _GEN_19548; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19550 = 12'h419 == _T_196[11:0] ? image_1049 : _GEN_19549; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19551 = 12'h41a == _T_196[11:0] ? image_1050 : _GEN_19550; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19552 = 12'h41b == _T_196[11:0] ? image_1051 : _GEN_19551; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19553 = 12'h41c == _T_196[11:0] ? image_1052 : _GEN_19552; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19554 = 12'h41d == _T_196[11:0] ? image_1053 : _GEN_19553; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19555 = 12'h41e == _T_196[11:0] ? image_1054 : _GEN_19554; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19556 = 12'h41f == _T_196[11:0] ? image_1055 : _GEN_19555; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19557 = 12'h420 == _T_196[11:0] ? image_1056 : _GEN_19556; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19558 = 12'h421 == _T_196[11:0] ? image_1057 : _GEN_19557; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19559 = 12'h422 == _T_196[11:0] ? image_1058 : _GEN_19558; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19560 = 12'h423 == _T_196[11:0] ? image_1059 : _GEN_19559; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19561 = 12'h424 == _T_196[11:0] ? image_1060 : _GEN_19560; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19562 = 12'h425 == _T_196[11:0] ? image_1061 : _GEN_19561; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19563 = 12'h426 == _T_196[11:0] ? image_1062 : _GEN_19562; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19564 = 12'h427 == _T_196[11:0] ? image_1063 : _GEN_19563; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19565 = 12'h428 == _T_196[11:0] ? image_1064 : _GEN_19564; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19566 = 12'h429 == _T_196[11:0] ? image_1065 : _GEN_19565; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19567 = 12'h42a == _T_196[11:0] ? image_1066 : _GEN_19566; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19568 = 12'h42b == _T_196[11:0] ? image_1067 : _GEN_19567; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19569 = 12'h42c == _T_196[11:0] ? image_1068 : _GEN_19568; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19570 = 12'h42d == _T_196[11:0] ? image_1069 : _GEN_19569; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19571 = 12'h42e == _T_196[11:0] ? image_1070 : _GEN_19570; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19572 = 12'h42f == _T_196[11:0] ? image_1071 : _GEN_19571; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19573 = 12'h430 == _T_196[11:0] ? image_1072 : _GEN_19572; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19574 = 12'h431 == _T_196[11:0] ? image_1073 : _GEN_19573; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19575 = 12'h432 == _T_196[11:0] ? image_1074 : _GEN_19574; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19576 = 12'h433 == _T_196[11:0] ? image_1075 : _GEN_19575; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19577 = 12'h434 == _T_196[11:0] ? image_1076 : _GEN_19576; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19578 = 12'h435 == _T_196[11:0] ? image_1077 : _GEN_19577; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19579 = 12'h436 == _T_196[11:0] ? image_1078 : _GEN_19578; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19580 = 12'h437 == _T_196[11:0] ? image_1079 : _GEN_19579; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19581 = 12'h438 == _T_196[11:0] ? image_1080 : _GEN_19580; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19582 = 12'h439 == _T_196[11:0] ? image_1081 : _GEN_19581; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19583 = 12'h43a == _T_196[11:0] ? image_1082 : _GEN_19582; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19584 = 12'h43b == _T_196[11:0] ? image_1083 : _GEN_19583; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19585 = 12'h43c == _T_196[11:0] ? image_1084 : _GEN_19584; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19586 = 12'h43d == _T_196[11:0] ? image_1085 : _GEN_19585; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19587 = 12'h43e == _T_196[11:0] ? 4'h0 : _GEN_19586; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19588 = 12'h43f == _T_196[11:0] ? 4'h0 : _GEN_19587; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19589 = 12'h440 == _T_196[11:0] ? image_1088 : _GEN_19588; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19590 = 12'h441 == _T_196[11:0] ? image_1089 : _GEN_19589; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19591 = 12'h442 == _T_196[11:0] ? image_1090 : _GEN_19590; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19592 = 12'h443 == _T_196[11:0] ? image_1091 : _GEN_19591; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19593 = 12'h444 == _T_196[11:0] ? image_1092 : _GEN_19592; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19594 = 12'h445 == _T_196[11:0] ? image_1093 : _GEN_19593; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19595 = 12'h446 == _T_196[11:0] ? image_1094 : _GEN_19594; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19596 = 12'h447 == _T_196[11:0] ? image_1095 : _GEN_19595; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19597 = 12'h448 == _T_196[11:0] ? image_1096 : _GEN_19596; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19598 = 12'h449 == _T_196[11:0] ? image_1097 : _GEN_19597; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19599 = 12'h44a == _T_196[11:0] ? image_1098 : _GEN_19598; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19600 = 12'h44b == _T_196[11:0] ? image_1099 : _GEN_19599; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19601 = 12'h44c == _T_196[11:0] ? image_1100 : _GEN_19600; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19602 = 12'h44d == _T_196[11:0] ? image_1101 : _GEN_19601; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19603 = 12'h44e == _T_196[11:0] ? image_1102 : _GEN_19602; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19604 = 12'h44f == _T_196[11:0] ? image_1103 : _GEN_19603; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19605 = 12'h450 == _T_196[11:0] ? image_1104 : _GEN_19604; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19606 = 12'h451 == _T_196[11:0] ? image_1105 : _GEN_19605; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19607 = 12'h452 == _T_196[11:0] ? image_1106 : _GEN_19606; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19608 = 12'h453 == _T_196[11:0] ? image_1107 : _GEN_19607; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19609 = 12'h454 == _T_196[11:0] ? image_1108 : _GEN_19608; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19610 = 12'h455 == _T_196[11:0] ? image_1109 : _GEN_19609; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19611 = 12'h456 == _T_196[11:0] ? image_1110 : _GEN_19610; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19612 = 12'h457 == _T_196[11:0] ? image_1111 : _GEN_19611; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19613 = 12'h458 == _T_196[11:0] ? image_1112 : _GEN_19612; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19614 = 12'h459 == _T_196[11:0] ? image_1113 : _GEN_19613; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19615 = 12'h45a == _T_196[11:0] ? image_1114 : _GEN_19614; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19616 = 12'h45b == _T_196[11:0] ? image_1115 : _GEN_19615; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19617 = 12'h45c == _T_196[11:0] ? image_1116 : _GEN_19616; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19618 = 12'h45d == _T_196[11:0] ? image_1117 : _GEN_19617; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19619 = 12'h45e == _T_196[11:0] ? image_1118 : _GEN_19618; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19620 = 12'h45f == _T_196[11:0] ? image_1119 : _GEN_19619; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19621 = 12'h460 == _T_196[11:0] ? image_1120 : _GEN_19620; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19622 = 12'h461 == _T_196[11:0] ? image_1121 : _GEN_19621; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19623 = 12'h462 == _T_196[11:0] ? image_1122 : _GEN_19622; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19624 = 12'h463 == _T_196[11:0] ? image_1123 : _GEN_19623; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19625 = 12'h464 == _T_196[11:0] ? image_1124 : _GEN_19624; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19626 = 12'h465 == _T_196[11:0] ? image_1125 : _GEN_19625; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19627 = 12'h466 == _T_196[11:0] ? image_1126 : _GEN_19626; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19628 = 12'h467 == _T_196[11:0] ? image_1127 : _GEN_19627; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19629 = 12'h468 == _T_196[11:0] ? image_1128 : _GEN_19628; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19630 = 12'h469 == _T_196[11:0] ? image_1129 : _GEN_19629; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19631 = 12'h46a == _T_196[11:0] ? image_1130 : _GEN_19630; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19632 = 12'h46b == _T_196[11:0] ? image_1131 : _GEN_19631; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19633 = 12'h46c == _T_196[11:0] ? image_1132 : _GEN_19632; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19634 = 12'h46d == _T_196[11:0] ? image_1133 : _GEN_19633; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19635 = 12'h46e == _T_196[11:0] ? image_1134 : _GEN_19634; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19636 = 12'h46f == _T_196[11:0] ? image_1135 : _GEN_19635; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19637 = 12'h470 == _T_196[11:0] ? image_1136 : _GEN_19636; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19638 = 12'h471 == _T_196[11:0] ? image_1137 : _GEN_19637; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19639 = 12'h472 == _T_196[11:0] ? image_1138 : _GEN_19638; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19640 = 12'h473 == _T_196[11:0] ? image_1139 : _GEN_19639; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19641 = 12'h474 == _T_196[11:0] ? image_1140 : _GEN_19640; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19642 = 12'h475 == _T_196[11:0] ? image_1141 : _GEN_19641; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19643 = 12'h476 == _T_196[11:0] ? image_1142 : _GEN_19642; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19644 = 12'h477 == _T_196[11:0] ? image_1143 : _GEN_19643; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19645 = 12'h478 == _T_196[11:0] ? image_1144 : _GEN_19644; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19646 = 12'h479 == _T_196[11:0] ? image_1145 : _GEN_19645; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19647 = 12'h47a == _T_196[11:0] ? image_1146 : _GEN_19646; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19648 = 12'h47b == _T_196[11:0] ? image_1147 : _GEN_19647; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19649 = 12'h47c == _T_196[11:0] ? image_1148 : _GEN_19648; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19650 = 12'h47d == _T_196[11:0] ? 4'h0 : _GEN_19649; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19651 = 12'h47e == _T_196[11:0] ? 4'h0 : _GEN_19650; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19652 = 12'h47f == _T_196[11:0] ? 4'h0 : _GEN_19651; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19653 = 12'h480 == _T_196[11:0] ? image_1152 : _GEN_19652; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19654 = 12'h481 == _T_196[11:0] ? image_1153 : _GEN_19653; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19655 = 12'h482 == _T_196[11:0] ? image_1154 : _GEN_19654; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19656 = 12'h483 == _T_196[11:0] ? image_1155 : _GEN_19655; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19657 = 12'h484 == _T_196[11:0] ? image_1156 : _GEN_19656; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19658 = 12'h485 == _T_196[11:0] ? image_1157 : _GEN_19657; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19659 = 12'h486 == _T_196[11:0] ? image_1158 : _GEN_19658; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19660 = 12'h487 == _T_196[11:0] ? image_1159 : _GEN_19659; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19661 = 12'h488 == _T_196[11:0] ? image_1160 : _GEN_19660; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19662 = 12'h489 == _T_196[11:0] ? image_1161 : _GEN_19661; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19663 = 12'h48a == _T_196[11:0] ? image_1162 : _GEN_19662; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19664 = 12'h48b == _T_196[11:0] ? image_1163 : _GEN_19663; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19665 = 12'h48c == _T_196[11:0] ? image_1164 : _GEN_19664; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19666 = 12'h48d == _T_196[11:0] ? image_1165 : _GEN_19665; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19667 = 12'h48e == _T_196[11:0] ? image_1166 : _GEN_19666; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19668 = 12'h48f == _T_196[11:0] ? image_1167 : _GEN_19667; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19669 = 12'h490 == _T_196[11:0] ? image_1168 : _GEN_19668; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19670 = 12'h491 == _T_196[11:0] ? image_1169 : _GEN_19669; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19671 = 12'h492 == _T_196[11:0] ? image_1170 : _GEN_19670; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19672 = 12'h493 == _T_196[11:0] ? image_1171 : _GEN_19671; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19673 = 12'h494 == _T_196[11:0] ? image_1172 : _GEN_19672; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19674 = 12'h495 == _T_196[11:0] ? image_1173 : _GEN_19673; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19675 = 12'h496 == _T_196[11:0] ? image_1174 : _GEN_19674; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19676 = 12'h497 == _T_196[11:0] ? image_1175 : _GEN_19675; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19677 = 12'h498 == _T_196[11:0] ? image_1176 : _GEN_19676; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19678 = 12'h499 == _T_196[11:0] ? image_1177 : _GEN_19677; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19679 = 12'h49a == _T_196[11:0] ? image_1178 : _GEN_19678; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19680 = 12'h49b == _T_196[11:0] ? image_1179 : _GEN_19679; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19681 = 12'h49c == _T_196[11:0] ? image_1180 : _GEN_19680; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19682 = 12'h49d == _T_196[11:0] ? image_1181 : _GEN_19681; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19683 = 12'h49e == _T_196[11:0] ? image_1182 : _GEN_19682; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19684 = 12'h49f == _T_196[11:0] ? image_1183 : _GEN_19683; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19685 = 12'h4a0 == _T_196[11:0] ? image_1184 : _GEN_19684; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19686 = 12'h4a1 == _T_196[11:0] ? image_1185 : _GEN_19685; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19687 = 12'h4a2 == _T_196[11:0] ? image_1186 : _GEN_19686; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19688 = 12'h4a3 == _T_196[11:0] ? image_1187 : _GEN_19687; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19689 = 12'h4a4 == _T_196[11:0] ? image_1188 : _GEN_19688; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19690 = 12'h4a5 == _T_196[11:0] ? image_1189 : _GEN_19689; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19691 = 12'h4a6 == _T_196[11:0] ? image_1190 : _GEN_19690; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19692 = 12'h4a7 == _T_196[11:0] ? image_1191 : _GEN_19691; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19693 = 12'h4a8 == _T_196[11:0] ? image_1192 : _GEN_19692; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19694 = 12'h4a9 == _T_196[11:0] ? image_1193 : _GEN_19693; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19695 = 12'h4aa == _T_196[11:0] ? image_1194 : _GEN_19694; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19696 = 12'h4ab == _T_196[11:0] ? image_1195 : _GEN_19695; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19697 = 12'h4ac == _T_196[11:0] ? image_1196 : _GEN_19696; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19698 = 12'h4ad == _T_196[11:0] ? image_1197 : _GEN_19697; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19699 = 12'h4ae == _T_196[11:0] ? image_1198 : _GEN_19698; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19700 = 12'h4af == _T_196[11:0] ? image_1199 : _GEN_19699; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19701 = 12'h4b0 == _T_196[11:0] ? image_1200 : _GEN_19700; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19702 = 12'h4b1 == _T_196[11:0] ? image_1201 : _GEN_19701; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19703 = 12'h4b2 == _T_196[11:0] ? image_1202 : _GEN_19702; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19704 = 12'h4b3 == _T_196[11:0] ? image_1203 : _GEN_19703; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19705 = 12'h4b4 == _T_196[11:0] ? image_1204 : _GEN_19704; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19706 = 12'h4b5 == _T_196[11:0] ? image_1205 : _GEN_19705; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19707 = 12'h4b6 == _T_196[11:0] ? image_1206 : _GEN_19706; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19708 = 12'h4b7 == _T_196[11:0] ? image_1207 : _GEN_19707; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19709 = 12'h4b8 == _T_196[11:0] ? image_1208 : _GEN_19708; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19710 = 12'h4b9 == _T_196[11:0] ? 4'h0 : _GEN_19709; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19711 = 12'h4ba == _T_196[11:0] ? 4'h0 : _GEN_19710; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19712 = 12'h4bb == _T_196[11:0] ? 4'h0 : _GEN_19711; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19713 = 12'h4bc == _T_196[11:0] ? 4'h0 : _GEN_19712; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19714 = 12'h4bd == _T_196[11:0] ? 4'h0 : _GEN_19713; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19715 = 12'h4be == _T_196[11:0] ? 4'h0 : _GEN_19714; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19716 = 12'h4bf == _T_196[11:0] ? 4'h0 : _GEN_19715; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19717 = 12'h4c0 == _T_196[11:0] ? image_1216 : _GEN_19716; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19718 = 12'h4c1 == _T_196[11:0] ? image_1217 : _GEN_19717; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19719 = 12'h4c2 == _T_196[11:0] ? image_1218 : _GEN_19718; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19720 = 12'h4c3 == _T_196[11:0] ? image_1219 : _GEN_19719; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19721 = 12'h4c4 == _T_196[11:0] ? image_1220 : _GEN_19720; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19722 = 12'h4c5 == _T_196[11:0] ? image_1221 : _GEN_19721; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19723 = 12'h4c6 == _T_196[11:0] ? image_1222 : _GEN_19722; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19724 = 12'h4c7 == _T_196[11:0] ? image_1223 : _GEN_19723; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19725 = 12'h4c8 == _T_196[11:0] ? image_1224 : _GEN_19724; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19726 = 12'h4c9 == _T_196[11:0] ? image_1225 : _GEN_19725; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19727 = 12'h4ca == _T_196[11:0] ? image_1226 : _GEN_19726; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19728 = 12'h4cb == _T_196[11:0] ? image_1227 : _GEN_19727; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19729 = 12'h4cc == _T_196[11:0] ? image_1228 : _GEN_19728; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19730 = 12'h4cd == _T_196[11:0] ? image_1229 : _GEN_19729; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19731 = 12'h4ce == _T_196[11:0] ? image_1230 : _GEN_19730; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19732 = 12'h4cf == _T_196[11:0] ? image_1231 : _GEN_19731; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19733 = 12'h4d0 == _T_196[11:0] ? image_1232 : _GEN_19732; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19734 = 12'h4d1 == _T_196[11:0] ? image_1233 : _GEN_19733; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19735 = 12'h4d2 == _T_196[11:0] ? image_1234 : _GEN_19734; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19736 = 12'h4d3 == _T_196[11:0] ? image_1235 : _GEN_19735; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19737 = 12'h4d4 == _T_196[11:0] ? image_1236 : _GEN_19736; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19738 = 12'h4d5 == _T_196[11:0] ? image_1237 : _GEN_19737; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19739 = 12'h4d6 == _T_196[11:0] ? image_1238 : _GEN_19738; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19740 = 12'h4d7 == _T_196[11:0] ? image_1239 : _GEN_19739; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19741 = 12'h4d8 == _T_196[11:0] ? image_1240 : _GEN_19740; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19742 = 12'h4d9 == _T_196[11:0] ? image_1241 : _GEN_19741; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19743 = 12'h4da == _T_196[11:0] ? image_1242 : _GEN_19742; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19744 = 12'h4db == _T_196[11:0] ? image_1243 : _GEN_19743; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19745 = 12'h4dc == _T_196[11:0] ? image_1244 : _GEN_19744; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19746 = 12'h4dd == _T_196[11:0] ? image_1245 : _GEN_19745; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19747 = 12'h4de == _T_196[11:0] ? image_1246 : _GEN_19746; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19748 = 12'h4df == _T_196[11:0] ? image_1247 : _GEN_19747; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19749 = 12'h4e0 == _T_196[11:0] ? image_1248 : _GEN_19748; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19750 = 12'h4e1 == _T_196[11:0] ? image_1249 : _GEN_19749; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19751 = 12'h4e2 == _T_196[11:0] ? image_1250 : _GEN_19750; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19752 = 12'h4e3 == _T_196[11:0] ? image_1251 : _GEN_19751; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19753 = 12'h4e4 == _T_196[11:0] ? image_1252 : _GEN_19752; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19754 = 12'h4e5 == _T_196[11:0] ? image_1253 : _GEN_19753; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19755 = 12'h4e6 == _T_196[11:0] ? image_1254 : _GEN_19754; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19756 = 12'h4e7 == _T_196[11:0] ? image_1255 : _GEN_19755; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19757 = 12'h4e8 == _T_196[11:0] ? image_1256 : _GEN_19756; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19758 = 12'h4e9 == _T_196[11:0] ? image_1257 : _GEN_19757; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19759 = 12'h4ea == _T_196[11:0] ? image_1258 : _GEN_19758; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19760 = 12'h4eb == _T_196[11:0] ? image_1259 : _GEN_19759; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19761 = 12'h4ec == _T_196[11:0] ? image_1260 : _GEN_19760; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19762 = 12'h4ed == _T_196[11:0] ? image_1261 : _GEN_19761; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19763 = 12'h4ee == _T_196[11:0] ? image_1262 : _GEN_19762; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19764 = 12'h4ef == _T_196[11:0] ? image_1263 : _GEN_19763; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19765 = 12'h4f0 == _T_196[11:0] ? image_1264 : _GEN_19764; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19766 = 12'h4f1 == _T_196[11:0] ? image_1265 : _GEN_19765; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19767 = 12'h4f2 == _T_196[11:0] ? image_1266 : _GEN_19766; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19768 = 12'h4f3 == _T_196[11:0] ? image_1267 : _GEN_19767; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19769 = 12'h4f4 == _T_196[11:0] ? image_1268 : _GEN_19768; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19770 = 12'h4f5 == _T_196[11:0] ? image_1269 : _GEN_19769; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19771 = 12'h4f6 == _T_196[11:0] ? image_1270 : _GEN_19770; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19772 = 12'h4f7 == _T_196[11:0] ? image_1271 : _GEN_19771; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19773 = 12'h4f8 == _T_196[11:0] ? image_1272 : _GEN_19772; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19774 = 12'h4f9 == _T_196[11:0] ? image_1273 : _GEN_19773; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19775 = 12'h4fa == _T_196[11:0] ? image_1274 : _GEN_19774; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19776 = 12'h4fb == _T_196[11:0] ? image_1275 : _GEN_19775; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19777 = 12'h4fc == _T_196[11:0] ? 4'h0 : _GEN_19776; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19778 = 12'h4fd == _T_196[11:0] ? 4'h0 : _GEN_19777; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19779 = 12'h4fe == _T_196[11:0] ? 4'h0 : _GEN_19778; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19780 = 12'h4ff == _T_196[11:0] ? 4'h0 : _GEN_19779; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19781 = 12'h500 == _T_196[11:0] ? image_1280 : _GEN_19780; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19782 = 12'h501 == _T_196[11:0] ? image_1281 : _GEN_19781; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19783 = 12'h502 == _T_196[11:0] ? image_1282 : _GEN_19782; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19784 = 12'h503 == _T_196[11:0] ? image_1283 : _GEN_19783; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19785 = 12'h504 == _T_196[11:0] ? image_1284 : _GEN_19784; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19786 = 12'h505 == _T_196[11:0] ? image_1285 : _GEN_19785; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19787 = 12'h506 == _T_196[11:0] ? image_1286 : _GEN_19786; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19788 = 12'h507 == _T_196[11:0] ? image_1287 : _GEN_19787; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19789 = 12'h508 == _T_196[11:0] ? image_1288 : _GEN_19788; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19790 = 12'h509 == _T_196[11:0] ? image_1289 : _GEN_19789; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19791 = 12'h50a == _T_196[11:0] ? image_1290 : _GEN_19790; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19792 = 12'h50b == _T_196[11:0] ? image_1291 : _GEN_19791; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19793 = 12'h50c == _T_196[11:0] ? image_1292 : _GEN_19792; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19794 = 12'h50d == _T_196[11:0] ? image_1293 : _GEN_19793; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19795 = 12'h50e == _T_196[11:0] ? image_1294 : _GEN_19794; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19796 = 12'h50f == _T_196[11:0] ? image_1295 : _GEN_19795; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19797 = 12'h510 == _T_196[11:0] ? image_1296 : _GEN_19796; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19798 = 12'h511 == _T_196[11:0] ? image_1297 : _GEN_19797; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19799 = 12'h512 == _T_196[11:0] ? image_1298 : _GEN_19798; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19800 = 12'h513 == _T_196[11:0] ? image_1299 : _GEN_19799; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19801 = 12'h514 == _T_196[11:0] ? image_1300 : _GEN_19800; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19802 = 12'h515 == _T_196[11:0] ? image_1301 : _GEN_19801; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19803 = 12'h516 == _T_196[11:0] ? image_1302 : _GEN_19802; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19804 = 12'h517 == _T_196[11:0] ? image_1303 : _GEN_19803; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19805 = 12'h518 == _T_196[11:0] ? image_1304 : _GEN_19804; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19806 = 12'h519 == _T_196[11:0] ? image_1305 : _GEN_19805; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19807 = 12'h51a == _T_196[11:0] ? image_1306 : _GEN_19806; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19808 = 12'h51b == _T_196[11:0] ? image_1307 : _GEN_19807; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19809 = 12'h51c == _T_196[11:0] ? image_1308 : _GEN_19808; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19810 = 12'h51d == _T_196[11:0] ? image_1309 : _GEN_19809; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19811 = 12'h51e == _T_196[11:0] ? image_1310 : _GEN_19810; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19812 = 12'h51f == _T_196[11:0] ? image_1311 : _GEN_19811; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19813 = 12'h520 == _T_196[11:0] ? image_1312 : _GEN_19812; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19814 = 12'h521 == _T_196[11:0] ? image_1313 : _GEN_19813; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19815 = 12'h522 == _T_196[11:0] ? image_1314 : _GEN_19814; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19816 = 12'h523 == _T_196[11:0] ? image_1315 : _GEN_19815; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19817 = 12'h524 == _T_196[11:0] ? image_1316 : _GEN_19816; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19818 = 12'h525 == _T_196[11:0] ? image_1317 : _GEN_19817; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19819 = 12'h526 == _T_196[11:0] ? image_1318 : _GEN_19818; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19820 = 12'h527 == _T_196[11:0] ? image_1319 : _GEN_19819; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19821 = 12'h528 == _T_196[11:0] ? image_1320 : _GEN_19820; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19822 = 12'h529 == _T_196[11:0] ? image_1321 : _GEN_19821; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19823 = 12'h52a == _T_196[11:0] ? image_1322 : _GEN_19822; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19824 = 12'h52b == _T_196[11:0] ? image_1323 : _GEN_19823; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19825 = 12'h52c == _T_196[11:0] ? image_1324 : _GEN_19824; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19826 = 12'h52d == _T_196[11:0] ? image_1325 : _GEN_19825; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19827 = 12'h52e == _T_196[11:0] ? image_1326 : _GEN_19826; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19828 = 12'h52f == _T_196[11:0] ? image_1327 : _GEN_19827; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19829 = 12'h530 == _T_196[11:0] ? image_1328 : _GEN_19828; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19830 = 12'h531 == _T_196[11:0] ? image_1329 : _GEN_19829; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19831 = 12'h532 == _T_196[11:0] ? image_1330 : _GEN_19830; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19832 = 12'h533 == _T_196[11:0] ? image_1331 : _GEN_19831; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19833 = 12'h534 == _T_196[11:0] ? image_1332 : _GEN_19832; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19834 = 12'h535 == _T_196[11:0] ? image_1333 : _GEN_19833; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19835 = 12'h536 == _T_196[11:0] ? image_1334 : _GEN_19834; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19836 = 12'h537 == _T_196[11:0] ? image_1335 : _GEN_19835; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19837 = 12'h538 == _T_196[11:0] ? image_1336 : _GEN_19836; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19838 = 12'h539 == _T_196[11:0] ? image_1337 : _GEN_19837; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19839 = 12'h53a == _T_196[11:0] ? image_1338 : _GEN_19838; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19840 = 12'h53b == _T_196[11:0] ? image_1339 : _GEN_19839; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19841 = 12'h53c == _T_196[11:0] ? image_1340 : _GEN_19840; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19842 = 12'h53d == _T_196[11:0] ? image_1341 : _GEN_19841; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19843 = 12'h53e == _T_196[11:0] ? 4'h0 : _GEN_19842; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19844 = 12'h53f == _T_196[11:0] ? 4'h0 : _GEN_19843; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19845 = 12'h540 == _T_196[11:0] ? image_1344 : _GEN_19844; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19846 = 12'h541 == _T_196[11:0] ? image_1345 : _GEN_19845; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19847 = 12'h542 == _T_196[11:0] ? image_1346 : _GEN_19846; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19848 = 12'h543 == _T_196[11:0] ? image_1347 : _GEN_19847; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19849 = 12'h544 == _T_196[11:0] ? image_1348 : _GEN_19848; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19850 = 12'h545 == _T_196[11:0] ? image_1349 : _GEN_19849; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19851 = 12'h546 == _T_196[11:0] ? image_1350 : _GEN_19850; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19852 = 12'h547 == _T_196[11:0] ? image_1351 : _GEN_19851; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19853 = 12'h548 == _T_196[11:0] ? image_1352 : _GEN_19852; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19854 = 12'h549 == _T_196[11:0] ? image_1353 : _GEN_19853; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19855 = 12'h54a == _T_196[11:0] ? image_1354 : _GEN_19854; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19856 = 12'h54b == _T_196[11:0] ? image_1355 : _GEN_19855; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19857 = 12'h54c == _T_196[11:0] ? image_1356 : _GEN_19856; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19858 = 12'h54d == _T_196[11:0] ? image_1357 : _GEN_19857; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19859 = 12'h54e == _T_196[11:0] ? image_1358 : _GEN_19858; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19860 = 12'h54f == _T_196[11:0] ? image_1359 : _GEN_19859; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19861 = 12'h550 == _T_196[11:0] ? image_1360 : _GEN_19860; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19862 = 12'h551 == _T_196[11:0] ? image_1361 : _GEN_19861; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19863 = 12'h552 == _T_196[11:0] ? image_1362 : _GEN_19862; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19864 = 12'h553 == _T_196[11:0] ? image_1363 : _GEN_19863; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19865 = 12'h554 == _T_196[11:0] ? image_1364 : _GEN_19864; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19866 = 12'h555 == _T_196[11:0] ? image_1365 : _GEN_19865; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19867 = 12'h556 == _T_196[11:0] ? image_1366 : _GEN_19866; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19868 = 12'h557 == _T_196[11:0] ? image_1367 : _GEN_19867; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19869 = 12'h558 == _T_196[11:0] ? image_1368 : _GEN_19868; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19870 = 12'h559 == _T_196[11:0] ? image_1369 : _GEN_19869; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19871 = 12'h55a == _T_196[11:0] ? image_1370 : _GEN_19870; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19872 = 12'h55b == _T_196[11:0] ? image_1371 : _GEN_19871; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19873 = 12'h55c == _T_196[11:0] ? image_1372 : _GEN_19872; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19874 = 12'h55d == _T_196[11:0] ? image_1373 : _GEN_19873; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19875 = 12'h55e == _T_196[11:0] ? image_1374 : _GEN_19874; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19876 = 12'h55f == _T_196[11:0] ? image_1375 : _GEN_19875; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19877 = 12'h560 == _T_196[11:0] ? image_1376 : _GEN_19876; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19878 = 12'h561 == _T_196[11:0] ? image_1377 : _GEN_19877; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19879 = 12'h562 == _T_196[11:0] ? image_1378 : _GEN_19878; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19880 = 12'h563 == _T_196[11:0] ? image_1379 : _GEN_19879; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19881 = 12'h564 == _T_196[11:0] ? image_1380 : _GEN_19880; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19882 = 12'h565 == _T_196[11:0] ? image_1381 : _GEN_19881; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19883 = 12'h566 == _T_196[11:0] ? image_1382 : _GEN_19882; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19884 = 12'h567 == _T_196[11:0] ? image_1383 : _GEN_19883; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19885 = 12'h568 == _T_196[11:0] ? image_1384 : _GEN_19884; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19886 = 12'h569 == _T_196[11:0] ? image_1385 : _GEN_19885; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19887 = 12'h56a == _T_196[11:0] ? image_1386 : _GEN_19886; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19888 = 12'h56b == _T_196[11:0] ? image_1387 : _GEN_19887; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19889 = 12'h56c == _T_196[11:0] ? image_1388 : _GEN_19888; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19890 = 12'h56d == _T_196[11:0] ? image_1389 : _GEN_19889; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19891 = 12'h56e == _T_196[11:0] ? image_1390 : _GEN_19890; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19892 = 12'h56f == _T_196[11:0] ? image_1391 : _GEN_19891; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19893 = 12'h570 == _T_196[11:0] ? image_1392 : _GEN_19892; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19894 = 12'h571 == _T_196[11:0] ? image_1393 : _GEN_19893; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19895 = 12'h572 == _T_196[11:0] ? image_1394 : _GEN_19894; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19896 = 12'h573 == _T_196[11:0] ? image_1395 : _GEN_19895; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19897 = 12'h574 == _T_196[11:0] ? image_1396 : _GEN_19896; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19898 = 12'h575 == _T_196[11:0] ? image_1397 : _GEN_19897; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19899 = 12'h576 == _T_196[11:0] ? image_1398 : _GEN_19898; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19900 = 12'h577 == _T_196[11:0] ? image_1399 : _GEN_19899; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19901 = 12'h578 == _T_196[11:0] ? image_1400 : _GEN_19900; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19902 = 12'h579 == _T_196[11:0] ? image_1401 : _GEN_19901; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19903 = 12'h57a == _T_196[11:0] ? image_1402 : _GEN_19902; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19904 = 12'h57b == _T_196[11:0] ? image_1403 : _GEN_19903; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19905 = 12'h57c == _T_196[11:0] ? image_1404 : _GEN_19904; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19906 = 12'h57d == _T_196[11:0] ? image_1405 : _GEN_19905; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19907 = 12'h57e == _T_196[11:0] ? 4'h0 : _GEN_19906; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19908 = 12'h57f == _T_196[11:0] ? 4'h0 : _GEN_19907; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19909 = 12'h580 == _T_196[11:0] ? image_1408 : _GEN_19908; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19910 = 12'h581 == _T_196[11:0] ? image_1409 : _GEN_19909; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19911 = 12'h582 == _T_196[11:0] ? image_1410 : _GEN_19910; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19912 = 12'h583 == _T_196[11:0] ? image_1411 : _GEN_19911; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19913 = 12'h584 == _T_196[11:0] ? image_1412 : _GEN_19912; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19914 = 12'h585 == _T_196[11:0] ? image_1413 : _GEN_19913; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19915 = 12'h586 == _T_196[11:0] ? image_1414 : _GEN_19914; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19916 = 12'h587 == _T_196[11:0] ? image_1415 : _GEN_19915; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19917 = 12'h588 == _T_196[11:0] ? image_1416 : _GEN_19916; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19918 = 12'h589 == _T_196[11:0] ? image_1417 : _GEN_19917; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19919 = 12'h58a == _T_196[11:0] ? image_1418 : _GEN_19918; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19920 = 12'h58b == _T_196[11:0] ? image_1419 : _GEN_19919; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19921 = 12'h58c == _T_196[11:0] ? image_1420 : _GEN_19920; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19922 = 12'h58d == _T_196[11:0] ? image_1421 : _GEN_19921; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19923 = 12'h58e == _T_196[11:0] ? image_1422 : _GEN_19922; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19924 = 12'h58f == _T_196[11:0] ? image_1423 : _GEN_19923; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19925 = 12'h590 == _T_196[11:0] ? image_1424 : _GEN_19924; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19926 = 12'h591 == _T_196[11:0] ? image_1425 : _GEN_19925; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19927 = 12'h592 == _T_196[11:0] ? image_1426 : _GEN_19926; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19928 = 12'h593 == _T_196[11:0] ? image_1427 : _GEN_19927; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19929 = 12'h594 == _T_196[11:0] ? image_1428 : _GEN_19928; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19930 = 12'h595 == _T_196[11:0] ? image_1429 : _GEN_19929; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19931 = 12'h596 == _T_196[11:0] ? image_1430 : _GEN_19930; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19932 = 12'h597 == _T_196[11:0] ? image_1431 : _GEN_19931; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19933 = 12'h598 == _T_196[11:0] ? image_1432 : _GEN_19932; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19934 = 12'h599 == _T_196[11:0] ? image_1433 : _GEN_19933; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19935 = 12'h59a == _T_196[11:0] ? image_1434 : _GEN_19934; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19936 = 12'h59b == _T_196[11:0] ? image_1435 : _GEN_19935; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19937 = 12'h59c == _T_196[11:0] ? image_1436 : _GEN_19936; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19938 = 12'h59d == _T_196[11:0] ? image_1437 : _GEN_19937; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19939 = 12'h59e == _T_196[11:0] ? image_1438 : _GEN_19938; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19940 = 12'h59f == _T_196[11:0] ? image_1439 : _GEN_19939; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19941 = 12'h5a0 == _T_196[11:0] ? image_1440 : _GEN_19940; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19942 = 12'h5a1 == _T_196[11:0] ? image_1441 : _GEN_19941; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19943 = 12'h5a2 == _T_196[11:0] ? image_1442 : _GEN_19942; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19944 = 12'h5a3 == _T_196[11:0] ? image_1443 : _GEN_19943; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19945 = 12'h5a4 == _T_196[11:0] ? image_1444 : _GEN_19944; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19946 = 12'h5a5 == _T_196[11:0] ? image_1445 : _GEN_19945; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19947 = 12'h5a6 == _T_196[11:0] ? image_1446 : _GEN_19946; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19948 = 12'h5a7 == _T_196[11:0] ? image_1447 : _GEN_19947; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19949 = 12'h5a8 == _T_196[11:0] ? image_1448 : _GEN_19948; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19950 = 12'h5a9 == _T_196[11:0] ? image_1449 : _GEN_19949; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19951 = 12'h5aa == _T_196[11:0] ? image_1450 : _GEN_19950; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19952 = 12'h5ab == _T_196[11:0] ? image_1451 : _GEN_19951; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19953 = 12'h5ac == _T_196[11:0] ? image_1452 : _GEN_19952; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19954 = 12'h5ad == _T_196[11:0] ? image_1453 : _GEN_19953; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19955 = 12'h5ae == _T_196[11:0] ? image_1454 : _GEN_19954; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19956 = 12'h5af == _T_196[11:0] ? image_1455 : _GEN_19955; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19957 = 12'h5b0 == _T_196[11:0] ? image_1456 : _GEN_19956; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19958 = 12'h5b1 == _T_196[11:0] ? image_1457 : _GEN_19957; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19959 = 12'h5b2 == _T_196[11:0] ? image_1458 : _GEN_19958; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19960 = 12'h5b3 == _T_196[11:0] ? image_1459 : _GEN_19959; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19961 = 12'h5b4 == _T_196[11:0] ? image_1460 : _GEN_19960; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19962 = 12'h5b5 == _T_196[11:0] ? image_1461 : _GEN_19961; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19963 = 12'h5b6 == _T_196[11:0] ? image_1462 : _GEN_19962; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19964 = 12'h5b7 == _T_196[11:0] ? image_1463 : _GEN_19963; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19965 = 12'h5b8 == _T_196[11:0] ? image_1464 : _GEN_19964; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19966 = 12'h5b9 == _T_196[11:0] ? image_1465 : _GEN_19965; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19967 = 12'h5ba == _T_196[11:0] ? image_1466 : _GEN_19966; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19968 = 12'h5bb == _T_196[11:0] ? image_1467 : _GEN_19967; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19969 = 12'h5bc == _T_196[11:0] ? image_1468 : _GEN_19968; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19970 = 12'h5bd == _T_196[11:0] ? image_1469 : _GEN_19969; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19971 = 12'h5be == _T_196[11:0] ? 4'h0 : _GEN_19970; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19972 = 12'h5bf == _T_196[11:0] ? 4'h0 : _GEN_19971; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19973 = 12'h5c0 == _T_196[11:0] ? image_1472 : _GEN_19972; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19974 = 12'h5c1 == _T_196[11:0] ? image_1473 : _GEN_19973; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19975 = 12'h5c2 == _T_196[11:0] ? image_1474 : _GEN_19974; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19976 = 12'h5c3 == _T_196[11:0] ? image_1475 : _GEN_19975; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19977 = 12'h5c4 == _T_196[11:0] ? image_1476 : _GEN_19976; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19978 = 12'h5c5 == _T_196[11:0] ? image_1477 : _GEN_19977; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19979 = 12'h5c6 == _T_196[11:0] ? image_1478 : _GEN_19978; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19980 = 12'h5c7 == _T_196[11:0] ? image_1479 : _GEN_19979; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19981 = 12'h5c8 == _T_196[11:0] ? image_1480 : _GEN_19980; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19982 = 12'h5c9 == _T_196[11:0] ? image_1481 : _GEN_19981; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19983 = 12'h5ca == _T_196[11:0] ? image_1482 : _GEN_19982; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19984 = 12'h5cb == _T_196[11:0] ? image_1483 : _GEN_19983; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19985 = 12'h5cc == _T_196[11:0] ? image_1484 : _GEN_19984; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19986 = 12'h5cd == _T_196[11:0] ? image_1485 : _GEN_19985; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19987 = 12'h5ce == _T_196[11:0] ? image_1486 : _GEN_19986; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19988 = 12'h5cf == _T_196[11:0] ? image_1487 : _GEN_19987; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19989 = 12'h5d0 == _T_196[11:0] ? image_1488 : _GEN_19988; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19990 = 12'h5d1 == _T_196[11:0] ? image_1489 : _GEN_19989; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19991 = 12'h5d2 == _T_196[11:0] ? image_1490 : _GEN_19990; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19992 = 12'h5d3 == _T_196[11:0] ? image_1491 : _GEN_19991; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19993 = 12'h5d4 == _T_196[11:0] ? image_1492 : _GEN_19992; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19994 = 12'h5d5 == _T_196[11:0] ? image_1493 : _GEN_19993; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19995 = 12'h5d6 == _T_196[11:0] ? image_1494 : _GEN_19994; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19996 = 12'h5d7 == _T_196[11:0] ? image_1495 : _GEN_19995; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19997 = 12'h5d8 == _T_196[11:0] ? image_1496 : _GEN_19996; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19998 = 12'h5d9 == _T_196[11:0] ? image_1497 : _GEN_19997; // @[Filter.scala 138:46]
  wire [3:0] _GEN_19999 = 12'h5da == _T_196[11:0] ? image_1498 : _GEN_19998; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20000 = 12'h5db == _T_196[11:0] ? image_1499 : _GEN_19999; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20001 = 12'h5dc == _T_196[11:0] ? image_1500 : _GEN_20000; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20002 = 12'h5dd == _T_196[11:0] ? image_1501 : _GEN_20001; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20003 = 12'h5de == _T_196[11:0] ? image_1502 : _GEN_20002; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20004 = 12'h5df == _T_196[11:0] ? image_1503 : _GEN_20003; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20005 = 12'h5e0 == _T_196[11:0] ? image_1504 : _GEN_20004; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20006 = 12'h5e1 == _T_196[11:0] ? image_1505 : _GEN_20005; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20007 = 12'h5e2 == _T_196[11:0] ? image_1506 : _GEN_20006; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20008 = 12'h5e3 == _T_196[11:0] ? image_1507 : _GEN_20007; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20009 = 12'h5e4 == _T_196[11:0] ? image_1508 : _GEN_20008; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20010 = 12'h5e5 == _T_196[11:0] ? image_1509 : _GEN_20009; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20011 = 12'h5e6 == _T_196[11:0] ? image_1510 : _GEN_20010; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20012 = 12'h5e7 == _T_196[11:0] ? image_1511 : _GEN_20011; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20013 = 12'h5e8 == _T_196[11:0] ? image_1512 : _GEN_20012; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20014 = 12'h5e9 == _T_196[11:0] ? image_1513 : _GEN_20013; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20015 = 12'h5ea == _T_196[11:0] ? image_1514 : _GEN_20014; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20016 = 12'h5eb == _T_196[11:0] ? image_1515 : _GEN_20015; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20017 = 12'h5ec == _T_196[11:0] ? image_1516 : _GEN_20016; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20018 = 12'h5ed == _T_196[11:0] ? image_1517 : _GEN_20017; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20019 = 12'h5ee == _T_196[11:0] ? image_1518 : _GEN_20018; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20020 = 12'h5ef == _T_196[11:0] ? image_1519 : _GEN_20019; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20021 = 12'h5f0 == _T_196[11:0] ? image_1520 : _GEN_20020; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20022 = 12'h5f1 == _T_196[11:0] ? image_1521 : _GEN_20021; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20023 = 12'h5f2 == _T_196[11:0] ? image_1522 : _GEN_20022; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20024 = 12'h5f3 == _T_196[11:0] ? image_1523 : _GEN_20023; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20025 = 12'h5f4 == _T_196[11:0] ? image_1524 : _GEN_20024; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20026 = 12'h5f5 == _T_196[11:0] ? image_1525 : _GEN_20025; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20027 = 12'h5f6 == _T_196[11:0] ? image_1526 : _GEN_20026; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20028 = 12'h5f7 == _T_196[11:0] ? image_1527 : _GEN_20027; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20029 = 12'h5f8 == _T_196[11:0] ? image_1528 : _GEN_20028; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20030 = 12'h5f9 == _T_196[11:0] ? image_1529 : _GEN_20029; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20031 = 12'h5fa == _T_196[11:0] ? image_1530 : _GEN_20030; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20032 = 12'h5fb == _T_196[11:0] ? image_1531 : _GEN_20031; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20033 = 12'h5fc == _T_196[11:0] ? image_1532 : _GEN_20032; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20034 = 12'h5fd == _T_196[11:0] ? image_1533 : _GEN_20033; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20035 = 12'h5fe == _T_196[11:0] ? 4'h0 : _GEN_20034; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20036 = 12'h5ff == _T_196[11:0] ? 4'h0 : _GEN_20035; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20037 = 12'h600 == _T_196[11:0] ? image_1536 : _GEN_20036; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20038 = 12'h601 == _T_196[11:0] ? image_1537 : _GEN_20037; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20039 = 12'h602 == _T_196[11:0] ? image_1538 : _GEN_20038; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20040 = 12'h603 == _T_196[11:0] ? image_1539 : _GEN_20039; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20041 = 12'h604 == _T_196[11:0] ? image_1540 : _GEN_20040; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20042 = 12'h605 == _T_196[11:0] ? image_1541 : _GEN_20041; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20043 = 12'h606 == _T_196[11:0] ? image_1542 : _GEN_20042; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20044 = 12'h607 == _T_196[11:0] ? image_1543 : _GEN_20043; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20045 = 12'h608 == _T_196[11:0] ? image_1544 : _GEN_20044; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20046 = 12'h609 == _T_196[11:0] ? image_1545 : _GEN_20045; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20047 = 12'h60a == _T_196[11:0] ? image_1546 : _GEN_20046; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20048 = 12'h60b == _T_196[11:0] ? image_1547 : _GEN_20047; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20049 = 12'h60c == _T_196[11:0] ? image_1548 : _GEN_20048; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20050 = 12'h60d == _T_196[11:0] ? image_1549 : _GEN_20049; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20051 = 12'h60e == _T_196[11:0] ? image_1550 : _GEN_20050; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20052 = 12'h60f == _T_196[11:0] ? image_1551 : _GEN_20051; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20053 = 12'h610 == _T_196[11:0] ? image_1552 : _GEN_20052; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20054 = 12'h611 == _T_196[11:0] ? image_1553 : _GEN_20053; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20055 = 12'h612 == _T_196[11:0] ? image_1554 : _GEN_20054; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20056 = 12'h613 == _T_196[11:0] ? image_1555 : _GEN_20055; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20057 = 12'h614 == _T_196[11:0] ? image_1556 : _GEN_20056; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20058 = 12'h615 == _T_196[11:0] ? image_1557 : _GEN_20057; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20059 = 12'h616 == _T_196[11:0] ? image_1558 : _GEN_20058; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20060 = 12'h617 == _T_196[11:0] ? image_1559 : _GEN_20059; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20061 = 12'h618 == _T_196[11:0] ? image_1560 : _GEN_20060; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20062 = 12'h619 == _T_196[11:0] ? image_1561 : _GEN_20061; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20063 = 12'h61a == _T_196[11:0] ? image_1562 : _GEN_20062; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20064 = 12'h61b == _T_196[11:0] ? image_1563 : _GEN_20063; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20065 = 12'h61c == _T_196[11:0] ? image_1564 : _GEN_20064; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20066 = 12'h61d == _T_196[11:0] ? image_1565 : _GEN_20065; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20067 = 12'h61e == _T_196[11:0] ? image_1566 : _GEN_20066; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20068 = 12'h61f == _T_196[11:0] ? image_1567 : _GEN_20067; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20069 = 12'h620 == _T_196[11:0] ? image_1568 : _GEN_20068; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20070 = 12'h621 == _T_196[11:0] ? image_1569 : _GEN_20069; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20071 = 12'h622 == _T_196[11:0] ? image_1570 : _GEN_20070; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20072 = 12'h623 == _T_196[11:0] ? image_1571 : _GEN_20071; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20073 = 12'h624 == _T_196[11:0] ? image_1572 : _GEN_20072; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20074 = 12'h625 == _T_196[11:0] ? image_1573 : _GEN_20073; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20075 = 12'h626 == _T_196[11:0] ? image_1574 : _GEN_20074; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20076 = 12'h627 == _T_196[11:0] ? image_1575 : _GEN_20075; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20077 = 12'h628 == _T_196[11:0] ? image_1576 : _GEN_20076; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20078 = 12'h629 == _T_196[11:0] ? image_1577 : _GEN_20077; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20079 = 12'h62a == _T_196[11:0] ? image_1578 : _GEN_20078; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20080 = 12'h62b == _T_196[11:0] ? image_1579 : _GEN_20079; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20081 = 12'h62c == _T_196[11:0] ? image_1580 : _GEN_20080; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20082 = 12'h62d == _T_196[11:0] ? image_1581 : _GEN_20081; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20083 = 12'h62e == _T_196[11:0] ? image_1582 : _GEN_20082; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20084 = 12'h62f == _T_196[11:0] ? image_1583 : _GEN_20083; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20085 = 12'h630 == _T_196[11:0] ? image_1584 : _GEN_20084; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20086 = 12'h631 == _T_196[11:0] ? image_1585 : _GEN_20085; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20087 = 12'h632 == _T_196[11:0] ? image_1586 : _GEN_20086; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20088 = 12'h633 == _T_196[11:0] ? image_1587 : _GEN_20087; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20089 = 12'h634 == _T_196[11:0] ? image_1588 : _GEN_20088; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20090 = 12'h635 == _T_196[11:0] ? image_1589 : _GEN_20089; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20091 = 12'h636 == _T_196[11:0] ? image_1590 : _GEN_20090; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20092 = 12'h637 == _T_196[11:0] ? image_1591 : _GEN_20091; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20093 = 12'h638 == _T_196[11:0] ? image_1592 : _GEN_20092; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20094 = 12'h639 == _T_196[11:0] ? image_1593 : _GEN_20093; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20095 = 12'h63a == _T_196[11:0] ? image_1594 : _GEN_20094; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20096 = 12'h63b == _T_196[11:0] ? image_1595 : _GEN_20095; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20097 = 12'h63c == _T_196[11:0] ? image_1596 : _GEN_20096; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20098 = 12'h63d == _T_196[11:0] ? image_1597 : _GEN_20097; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20099 = 12'h63e == _T_196[11:0] ? 4'h0 : _GEN_20098; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20100 = 12'h63f == _T_196[11:0] ? 4'h0 : _GEN_20099; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20101 = 12'h640 == _T_196[11:0] ? image_1600 : _GEN_20100; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20102 = 12'h641 == _T_196[11:0] ? image_1601 : _GEN_20101; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20103 = 12'h642 == _T_196[11:0] ? image_1602 : _GEN_20102; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20104 = 12'h643 == _T_196[11:0] ? image_1603 : _GEN_20103; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20105 = 12'h644 == _T_196[11:0] ? image_1604 : _GEN_20104; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20106 = 12'h645 == _T_196[11:0] ? image_1605 : _GEN_20105; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20107 = 12'h646 == _T_196[11:0] ? image_1606 : _GEN_20106; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20108 = 12'h647 == _T_196[11:0] ? image_1607 : _GEN_20107; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20109 = 12'h648 == _T_196[11:0] ? image_1608 : _GEN_20108; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20110 = 12'h649 == _T_196[11:0] ? image_1609 : _GEN_20109; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20111 = 12'h64a == _T_196[11:0] ? image_1610 : _GEN_20110; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20112 = 12'h64b == _T_196[11:0] ? image_1611 : _GEN_20111; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20113 = 12'h64c == _T_196[11:0] ? image_1612 : _GEN_20112; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20114 = 12'h64d == _T_196[11:0] ? image_1613 : _GEN_20113; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20115 = 12'h64e == _T_196[11:0] ? image_1614 : _GEN_20114; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20116 = 12'h64f == _T_196[11:0] ? image_1615 : _GEN_20115; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20117 = 12'h650 == _T_196[11:0] ? image_1616 : _GEN_20116; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20118 = 12'h651 == _T_196[11:0] ? image_1617 : _GEN_20117; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20119 = 12'h652 == _T_196[11:0] ? image_1618 : _GEN_20118; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20120 = 12'h653 == _T_196[11:0] ? image_1619 : _GEN_20119; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20121 = 12'h654 == _T_196[11:0] ? image_1620 : _GEN_20120; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20122 = 12'h655 == _T_196[11:0] ? image_1621 : _GEN_20121; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20123 = 12'h656 == _T_196[11:0] ? image_1622 : _GEN_20122; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20124 = 12'h657 == _T_196[11:0] ? image_1623 : _GEN_20123; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20125 = 12'h658 == _T_196[11:0] ? image_1624 : _GEN_20124; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20126 = 12'h659 == _T_196[11:0] ? image_1625 : _GEN_20125; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20127 = 12'h65a == _T_196[11:0] ? image_1626 : _GEN_20126; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20128 = 12'h65b == _T_196[11:0] ? image_1627 : _GEN_20127; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20129 = 12'h65c == _T_196[11:0] ? image_1628 : _GEN_20128; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20130 = 12'h65d == _T_196[11:0] ? image_1629 : _GEN_20129; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20131 = 12'h65e == _T_196[11:0] ? image_1630 : _GEN_20130; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20132 = 12'h65f == _T_196[11:0] ? image_1631 : _GEN_20131; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20133 = 12'h660 == _T_196[11:0] ? image_1632 : _GEN_20132; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20134 = 12'h661 == _T_196[11:0] ? image_1633 : _GEN_20133; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20135 = 12'h662 == _T_196[11:0] ? image_1634 : _GEN_20134; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20136 = 12'h663 == _T_196[11:0] ? image_1635 : _GEN_20135; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20137 = 12'h664 == _T_196[11:0] ? image_1636 : _GEN_20136; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20138 = 12'h665 == _T_196[11:0] ? image_1637 : _GEN_20137; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20139 = 12'h666 == _T_196[11:0] ? image_1638 : _GEN_20138; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20140 = 12'h667 == _T_196[11:0] ? image_1639 : _GEN_20139; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20141 = 12'h668 == _T_196[11:0] ? image_1640 : _GEN_20140; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20142 = 12'h669 == _T_196[11:0] ? image_1641 : _GEN_20141; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20143 = 12'h66a == _T_196[11:0] ? image_1642 : _GEN_20142; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20144 = 12'h66b == _T_196[11:0] ? image_1643 : _GEN_20143; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20145 = 12'h66c == _T_196[11:0] ? image_1644 : _GEN_20144; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20146 = 12'h66d == _T_196[11:0] ? image_1645 : _GEN_20145; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20147 = 12'h66e == _T_196[11:0] ? image_1646 : _GEN_20146; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20148 = 12'h66f == _T_196[11:0] ? image_1647 : _GEN_20147; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20149 = 12'h670 == _T_196[11:0] ? image_1648 : _GEN_20148; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20150 = 12'h671 == _T_196[11:0] ? image_1649 : _GEN_20149; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20151 = 12'h672 == _T_196[11:0] ? image_1650 : _GEN_20150; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20152 = 12'h673 == _T_196[11:0] ? image_1651 : _GEN_20151; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20153 = 12'h674 == _T_196[11:0] ? image_1652 : _GEN_20152; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20154 = 12'h675 == _T_196[11:0] ? image_1653 : _GEN_20153; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20155 = 12'h676 == _T_196[11:0] ? image_1654 : _GEN_20154; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20156 = 12'h677 == _T_196[11:0] ? image_1655 : _GEN_20155; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20157 = 12'h678 == _T_196[11:0] ? image_1656 : _GEN_20156; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20158 = 12'h679 == _T_196[11:0] ? image_1657 : _GEN_20157; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20159 = 12'h67a == _T_196[11:0] ? image_1658 : _GEN_20158; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20160 = 12'h67b == _T_196[11:0] ? image_1659 : _GEN_20159; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20161 = 12'h67c == _T_196[11:0] ? image_1660 : _GEN_20160; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20162 = 12'h67d == _T_196[11:0] ? 4'h0 : _GEN_20161; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20163 = 12'h67e == _T_196[11:0] ? 4'h0 : _GEN_20162; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20164 = 12'h67f == _T_196[11:0] ? 4'h0 : _GEN_20163; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20165 = 12'h680 == _T_196[11:0] ? image_1664 : _GEN_20164; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20166 = 12'h681 == _T_196[11:0] ? image_1665 : _GEN_20165; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20167 = 12'h682 == _T_196[11:0] ? image_1666 : _GEN_20166; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20168 = 12'h683 == _T_196[11:0] ? image_1667 : _GEN_20167; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20169 = 12'h684 == _T_196[11:0] ? image_1668 : _GEN_20168; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20170 = 12'h685 == _T_196[11:0] ? image_1669 : _GEN_20169; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20171 = 12'h686 == _T_196[11:0] ? image_1670 : _GEN_20170; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20172 = 12'h687 == _T_196[11:0] ? image_1671 : _GEN_20171; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20173 = 12'h688 == _T_196[11:0] ? image_1672 : _GEN_20172; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20174 = 12'h689 == _T_196[11:0] ? image_1673 : _GEN_20173; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20175 = 12'h68a == _T_196[11:0] ? image_1674 : _GEN_20174; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20176 = 12'h68b == _T_196[11:0] ? image_1675 : _GEN_20175; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20177 = 12'h68c == _T_196[11:0] ? image_1676 : _GEN_20176; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20178 = 12'h68d == _T_196[11:0] ? image_1677 : _GEN_20177; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20179 = 12'h68e == _T_196[11:0] ? image_1678 : _GEN_20178; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20180 = 12'h68f == _T_196[11:0] ? image_1679 : _GEN_20179; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20181 = 12'h690 == _T_196[11:0] ? image_1680 : _GEN_20180; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20182 = 12'h691 == _T_196[11:0] ? image_1681 : _GEN_20181; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20183 = 12'h692 == _T_196[11:0] ? image_1682 : _GEN_20182; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20184 = 12'h693 == _T_196[11:0] ? image_1683 : _GEN_20183; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20185 = 12'h694 == _T_196[11:0] ? image_1684 : _GEN_20184; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20186 = 12'h695 == _T_196[11:0] ? image_1685 : _GEN_20185; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20187 = 12'h696 == _T_196[11:0] ? image_1686 : _GEN_20186; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20188 = 12'h697 == _T_196[11:0] ? image_1687 : _GEN_20187; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20189 = 12'h698 == _T_196[11:0] ? image_1688 : _GEN_20188; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20190 = 12'h699 == _T_196[11:0] ? image_1689 : _GEN_20189; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20191 = 12'h69a == _T_196[11:0] ? image_1690 : _GEN_20190; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20192 = 12'h69b == _T_196[11:0] ? image_1691 : _GEN_20191; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20193 = 12'h69c == _T_196[11:0] ? image_1692 : _GEN_20192; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20194 = 12'h69d == _T_196[11:0] ? image_1693 : _GEN_20193; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20195 = 12'h69e == _T_196[11:0] ? image_1694 : _GEN_20194; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20196 = 12'h69f == _T_196[11:0] ? image_1695 : _GEN_20195; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20197 = 12'h6a0 == _T_196[11:0] ? image_1696 : _GEN_20196; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20198 = 12'h6a1 == _T_196[11:0] ? image_1697 : _GEN_20197; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20199 = 12'h6a2 == _T_196[11:0] ? image_1698 : _GEN_20198; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20200 = 12'h6a3 == _T_196[11:0] ? image_1699 : _GEN_20199; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20201 = 12'h6a4 == _T_196[11:0] ? image_1700 : _GEN_20200; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20202 = 12'h6a5 == _T_196[11:0] ? image_1701 : _GEN_20201; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20203 = 12'h6a6 == _T_196[11:0] ? image_1702 : _GEN_20202; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20204 = 12'h6a7 == _T_196[11:0] ? image_1703 : _GEN_20203; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20205 = 12'h6a8 == _T_196[11:0] ? image_1704 : _GEN_20204; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20206 = 12'h6a9 == _T_196[11:0] ? image_1705 : _GEN_20205; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20207 = 12'h6aa == _T_196[11:0] ? image_1706 : _GEN_20206; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20208 = 12'h6ab == _T_196[11:0] ? image_1707 : _GEN_20207; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20209 = 12'h6ac == _T_196[11:0] ? image_1708 : _GEN_20208; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20210 = 12'h6ad == _T_196[11:0] ? image_1709 : _GEN_20209; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20211 = 12'h6ae == _T_196[11:0] ? image_1710 : _GEN_20210; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20212 = 12'h6af == _T_196[11:0] ? image_1711 : _GEN_20211; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20213 = 12'h6b0 == _T_196[11:0] ? image_1712 : _GEN_20212; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20214 = 12'h6b1 == _T_196[11:0] ? image_1713 : _GEN_20213; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20215 = 12'h6b2 == _T_196[11:0] ? image_1714 : _GEN_20214; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20216 = 12'h6b3 == _T_196[11:0] ? image_1715 : _GEN_20215; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20217 = 12'h6b4 == _T_196[11:0] ? image_1716 : _GEN_20216; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20218 = 12'h6b5 == _T_196[11:0] ? image_1717 : _GEN_20217; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20219 = 12'h6b6 == _T_196[11:0] ? image_1718 : _GEN_20218; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20220 = 12'h6b7 == _T_196[11:0] ? image_1719 : _GEN_20219; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20221 = 12'h6b8 == _T_196[11:0] ? image_1720 : _GEN_20220; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20222 = 12'h6b9 == _T_196[11:0] ? image_1721 : _GEN_20221; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20223 = 12'h6ba == _T_196[11:0] ? image_1722 : _GEN_20222; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20224 = 12'h6bb == _T_196[11:0] ? image_1723 : _GEN_20223; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20225 = 12'h6bc == _T_196[11:0] ? 4'h0 : _GEN_20224; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20226 = 12'h6bd == _T_196[11:0] ? 4'h0 : _GEN_20225; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20227 = 12'h6be == _T_196[11:0] ? 4'h0 : _GEN_20226; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20228 = 12'h6bf == _T_196[11:0] ? 4'h0 : _GEN_20227; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20229 = 12'h6c0 == _T_196[11:0] ? image_1728 : _GEN_20228; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20230 = 12'h6c1 == _T_196[11:0] ? image_1729 : _GEN_20229; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20231 = 12'h6c2 == _T_196[11:0] ? image_1730 : _GEN_20230; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20232 = 12'h6c3 == _T_196[11:0] ? image_1731 : _GEN_20231; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20233 = 12'h6c4 == _T_196[11:0] ? image_1732 : _GEN_20232; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20234 = 12'h6c5 == _T_196[11:0] ? image_1733 : _GEN_20233; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20235 = 12'h6c6 == _T_196[11:0] ? image_1734 : _GEN_20234; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20236 = 12'h6c7 == _T_196[11:0] ? image_1735 : _GEN_20235; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20237 = 12'h6c8 == _T_196[11:0] ? image_1736 : _GEN_20236; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20238 = 12'h6c9 == _T_196[11:0] ? image_1737 : _GEN_20237; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20239 = 12'h6ca == _T_196[11:0] ? image_1738 : _GEN_20238; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20240 = 12'h6cb == _T_196[11:0] ? image_1739 : _GEN_20239; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20241 = 12'h6cc == _T_196[11:0] ? image_1740 : _GEN_20240; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20242 = 12'h6cd == _T_196[11:0] ? image_1741 : _GEN_20241; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20243 = 12'h6ce == _T_196[11:0] ? image_1742 : _GEN_20242; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20244 = 12'h6cf == _T_196[11:0] ? image_1743 : _GEN_20243; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20245 = 12'h6d0 == _T_196[11:0] ? image_1744 : _GEN_20244; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20246 = 12'h6d1 == _T_196[11:0] ? image_1745 : _GEN_20245; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20247 = 12'h6d2 == _T_196[11:0] ? image_1746 : _GEN_20246; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20248 = 12'h6d3 == _T_196[11:0] ? image_1747 : _GEN_20247; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20249 = 12'h6d4 == _T_196[11:0] ? image_1748 : _GEN_20248; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20250 = 12'h6d5 == _T_196[11:0] ? image_1749 : _GEN_20249; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20251 = 12'h6d6 == _T_196[11:0] ? image_1750 : _GEN_20250; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20252 = 12'h6d7 == _T_196[11:0] ? image_1751 : _GEN_20251; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20253 = 12'h6d8 == _T_196[11:0] ? image_1752 : _GEN_20252; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20254 = 12'h6d9 == _T_196[11:0] ? image_1753 : _GEN_20253; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20255 = 12'h6da == _T_196[11:0] ? image_1754 : _GEN_20254; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20256 = 12'h6db == _T_196[11:0] ? image_1755 : _GEN_20255; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20257 = 12'h6dc == _T_196[11:0] ? image_1756 : _GEN_20256; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20258 = 12'h6dd == _T_196[11:0] ? image_1757 : _GEN_20257; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20259 = 12'h6de == _T_196[11:0] ? image_1758 : _GEN_20258; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20260 = 12'h6df == _T_196[11:0] ? image_1759 : _GEN_20259; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20261 = 12'h6e0 == _T_196[11:0] ? image_1760 : _GEN_20260; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20262 = 12'h6e1 == _T_196[11:0] ? image_1761 : _GEN_20261; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20263 = 12'h6e2 == _T_196[11:0] ? image_1762 : _GEN_20262; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20264 = 12'h6e3 == _T_196[11:0] ? image_1763 : _GEN_20263; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20265 = 12'h6e4 == _T_196[11:0] ? image_1764 : _GEN_20264; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20266 = 12'h6e5 == _T_196[11:0] ? image_1765 : _GEN_20265; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20267 = 12'h6e6 == _T_196[11:0] ? image_1766 : _GEN_20266; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20268 = 12'h6e7 == _T_196[11:0] ? image_1767 : _GEN_20267; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20269 = 12'h6e8 == _T_196[11:0] ? image_1768 : _GEN_20268; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20270 = 12'h6e9 == _T_196[11:0] ? image_1769 : _GEN_20269; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20271 = 12'h6ea == _T_196[11:0] ? image_1770 : _GEN_20270; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20272 = 12'h6eb == _T_196[11:0] ? image_1771 : _GEN_20271; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20273 = 12'h6ec == _T_196[11:0] ? image_1772 : _GEN_20272; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20274 = 12'h6ed == _T_196[11:0] ? image_1773 : _GEN_20273; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20275 = 12'h6ee == _T_196[11:0] ? image_1774 : _GEN_20274; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20276 = 12'h6ef == _T_196[11:0] ? image_1775 : _GEN_20275; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20277 = 12'h6f0 == _T_196[11:0] ? image_1776 : _GEN_20276; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20278 = 12'h6f1 == _T_196[11:0] ? image_1777 : _GEN_20277; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20279 = 12'h6f2 == _T_196[11:0] ? image_1778 : _GEN_20278; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20280 = 12'h6f3 == _T_196[11:0] ? image_1779 : _GEN_20279; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20281 = 12'h6f4 == _T_196[11:0] ? image_1780 : _GEN_20280; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20282 = 12'h6f5 == _T_196[11:0] ? image_1781 : _GEN_20281; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20283 = 12'h6f6 == _T_196[11:0] ? image_1782 : _GEN_20282; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20284 = 12'h6f7 == _T_196[11:0] ? image_1783 : _GEN_20283; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20285 = 12'h6f8 == _T_196[11:0] ? image_1784 : _GEN_20284; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20286 = 12'h6f9 == _T_196[11:0] ? image_1785 : _GEN_20285; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20287 = 12'h6fa == _T_196[11:0] ? image_1786 : _GEN_20286; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20288 = 12'h6fb == _T_196[11:0] ? 4'h0 : _GEN_20287; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20289 = 12'h6fc == _T_196[11:0] ? 4'h0 : _GEN_20288; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20290 = 12'h6fd == _T_196[11:0] ? 4'h0 : _GEN_20289; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20291 = 12'h6fe == _T_196[11:0] ? 4'h0 : _GEN_20290; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20292 = 12'h6ff == _T_196[11:0] ? 4'h0 : _GEN_20291; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20293 = 12'h700 == _T_196[11:0] ? 4'h0 : _GEN_20292; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20294 = 12'h701 == _T_196[11:0] ? image_1793 : _GEN_20293; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20295 = 12'h702 == _T_196[11:0] ? image_1794 : _GEN_20294; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20296 = 12'h703 == _T_196[11:0] ? image_1795 : _GEN_20295; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20297 = 12'h704 == _T_196[11:0] ? image_1796 : _GEN_20296; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20298 = 12'h705 == _T_196[11:0] ? image_1797 : _GEN_20297; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20299 = 12'h706 == _T_196[11:0] ? image_1798 : _GEN_20298; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20300 = 12'h707 == _T_196[11:0] ? image_1799 : _GEN_20299; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20301 = 12'h708 == _T_196[11:0] ? image_1800 : _GEN_20300; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20302 = 12'h709 == _T_196[11:0] ? image_1801 : _GEN_20301; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20303 = 12'h70a == _T_196[11:0] ? image_1802 : _GEN_20302; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20304 = 12'h70b == _T_196[11:0] ? image_1803 : _GEN_20303; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20305 = 12'h70c == _T_196[11:0] ? image_1804 : _GEN_20304; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20306 = 12'h70d == _T_196[11:0] ? image_1805 : _GEN_20305; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20307 = 12'h70e == _T_196[11:0] ? image_1806 : _GEN_20306; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20308 = 12'h70f == _T_196[11:0] ? image_1807 : _GEN_20307; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20309 = 12'h710 == _T_196[11:0] ? image_1808 : _GEN_20308; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20310 = 12'h711 == _T_196[11:0] ? image_1809 : _GEN_20309; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20311 = 12'h712 == _T_196[11:0] ? image_1810 : _GEN_20310; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20312 = 12'h713 == _T_196[11:0] ? image_1811 : _GEN_20311; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20313 = 12'h714 == _T_196[11:0] ? image_1812 : _GEN_20312; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20314 = 12'h715 == _T_196[11:0] ? image_1813 : _GEN_20313; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20315 = 12'h716 == _T_196[11:0] ? image_1814 : _GEN_20314; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20316 = 12'h717 == _T_196[11:0] ? image_1815 : _GEN_20315; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20317 = 12'h718 == _T_196[11:0] ? image_1816 : _GEN_20316; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20318 = 12'h719 == _T_196[11:0] ? image_1817 : _GEN_20317; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20319 = 12'h71a == _T_196[11:0] ? image_1818 : _GEN_20318; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20320 = 12'h71b == _T_196[11:0] ? image_1819 : _GEN_20319; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20321 = 12'h71c == _T_196[11:0] ? image_1820 : _GEN_20320; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20322 = 12'h71d == _T_196[11:0] ? image_1821 : _GEN_20321; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20323 = 12'h71e == _T_196[11:0] ? image_1822 : _GEN_20322; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20324 = 12'h71f == _T_196[11:0] ? image_1823 : _GEN_20323; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20325 = 12'h720 == _T_196[11:0] ? image_1824 : _GEN_20324; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20326 = 12'h721 == _T_196[11:0] ? image_1825 : _GEN_20325; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20327 = 12'h722 == _T_196[11:0] ? image_1826 : _GEN_20326; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20328 = 12'h723 == _T_196[11:0] ? image_1827 : _GEN_20327; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20329 = 12'h724 == _T_196[11:0] ? image_1828 : _GEN_20328; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20330 = 12'h725 == _T_196[11:0] ? image_1829 : _GEN_20329; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20331 = 12'h726 == _T_196[11:0] ? image_1830 : _GEN_20330; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20332 = 12'h727 == _T_196[11:0] ? image_1831 : _GEN_20331; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20333 = 12'h728 == _T_196[11:0] ? image_1832 : _GEN_20332; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20334 = 12'h729 == _T_196[11:0] ? image_1833 : _GEN_20333; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20335 = 12'h72a == _T_196[11:0] ? image_1834 : _GEN_20334; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20336 = 12'h72b == _T_196[11:0] ? image_1835 : _GEN_20335; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20337 = 12'h72c == _T_196[11:0] ? image_1836 : _GEN_20336; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20338 = 12'h72d == _T_196[11:0] ? image_1837 : _GEN_20337; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20339 = 12'h72e == _T_196[11:0] ? image_1838 : _GEN_20338; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20340 = 12'h72f == _T_196[11:0] ? image_1839 : _GEN_20339; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20341 = 12'h730 == _T_196[11:0] ? image_1840 : _GEN_20340; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20342 = 12'h731 == _T_196[11:0] ? image_1841 : _GEN_20341; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20343 = 12'h732 == _T_196[11:0] ? image_1842 : _GEN_20342; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20344 = 12'h733 == _T_196[11:0] ? image_1843 : _GEN_20343; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20345 = 12'h734 == _T_196[11:0] ? image_1844 : _GEN_20344; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20346 = 12'h735 == _T_196[11:0] ? image_1845 : _GEN_20345; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20347 = 12'h736 == _T_196[11:0] ? image_1846 : _GEN_20346; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20348 = 12'h737 == _T_196[11:0] ? image_1847 : _GEN_20347; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20349 = 12'h738 == _T_196[11:0] ? image_1848 : _GEN_20348; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20350 = 12'h739 == _T_196[11:0] ? image_1849 : _GEN_20349; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20351 = 12'h73a == _T_196[11:0] ? 4'h0 : _GEN_20350; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20352 = 12'h73b == _T_196[11:0] ? 4'h0 : _GEN_20351; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20353 = 12'h73c == _T_196[11:0] ? 4'h0 : _GEN_20352; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20354 = 12'h73d == _T_196[11:0] ? 4'h0 : _GEN_20353; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20355 = 12'h73e == _T_196[11:0] ? 4'h0 : _GEN_20354; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20356 = 12'h73f == _T_196[11:0] ? 4'h0 : _GEN_20355; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20357 = 12'h740 == _T_196[11:0] ? 4'h0 : _GEN_20356; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20358 = 12'h741 == _T_196[11:0] ? image_1857 : _GEN_20357; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20359 = 12'h742 == _T_196[11:0] ? image_1858 : _GEN_20358; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20360 = 12'h743 == _T_196[11:0] ? image_1859 : _GEN_20359; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20361 = 12'h744 == _T_196[11:0] ? image_1860 : _GEN_20360; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20362 = 12'h745 == _T_196[11:0] ? image_1861 : _GEN_20361; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20363 = 12'h746 == _T_196[11:0] ? image_1862 : _GEN_20362; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20364 = 12'h747 == _T_196[11:0] ? image_1863 : _GEN_20363; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20365 = 12'h748 == _T_196[11:0] ? image_1864 : _GEN_20364; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20366 = 12'h749 == _T_196[11:0] ? image_1865 : _GEN_20365; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20367 = 12'h74a == _T_196[11:0] ? image_1866 : _GEN_20366; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20368 = 12'h74b == _T_196[11:0] ? image_1867 : _GEN_20367; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20369 = 12'h74c == _T_196[11:0] ? image_1868 : _GEN_20368; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20370 = 12'h74d == _T_196[11:0] ? image_1869 : _GEN_20369; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20371 = 12'h74e == _T_196[11:0] ? image_1870 : _GEN_20370; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20372 = 12'h74f == _T_196[11:0] ? image_1871 : _GEN_20371; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20373 = 12'h750 == _T_196[11:0] ? image_1872 : _GEN_20372; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20374 = 12'h751 == _T_196[11:0] ? image_1873 : _GEN_20373; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20375 = 12'h752 == _T_196[11:0] ? image_1874 : _GEN_20374; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20376 = 12'h753 == _T_196[11:0] ? image_1875 : _GEN_20375; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20377 = 12'h754 == _T_196[11:0] ? image_1876 : _GEN_20376; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20378 = 12'h755 == _T_196[11:0] ? image_1877 : _GEN_20377; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20379 = 12'h756 == _T_196[11:0] ? image_1878 : _GEN_20378; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20380 = 12'h757 == _T_196[11:0] ? image_1879 : _GEN_20379; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20381 = 12'h758 == _T_196[11:0] ? image_1880 : _GEN_20380; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20382 = 12'h759 == _T_196[11:0] ? image_1881 : _GEN_20381; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20383 = 12'h75a == _T_196[11:0] ? image_1882 : _GEN_20382; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20384 = 12'h75b == _T_196[11:0] ? image_1883 : _GEN_20383; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20385 = 12'h75c == _T_196[11:0] ? image_1884 : _GEN_20384; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20386 = 12'h75d == _T_196[11:0] ? image_1885 : _GEN_20385; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20387 = 12'h75e == _T_196[11:0] ? image_1886 : _GEN_20386; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20388 = 12'h75f == _T_196[11:0] ? image_1887 : _GEN_20387; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20389 = 12'h760 == _T_196[11:0] ? image_1888 : _GEN_20388; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20390 = 12'h761 == _T_196[11:0] ? image_1889 : _GEN_20389; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20391 = 12'h762 == _T_196[11:0] ? image_1890 : _GEN_20390; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20392 = 12'h763 == _T_196[11:0] ? image_1891 : _GEN_20391; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20393 = 12'h764 == _T_196[11:0] ? image_1892 : _GEN_20392; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20394 = 12'h765 == _T_196[11:0] ? image_1893 : _GEN_20393; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20395 = 12'h766 == _T_196[11:0] ? image_1894 : _GEN_20394; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20396 = 12'h767 == _T_196[11:0] ? image_1895 : _GEN_20395; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20397 = 12'h768 == _T_196[11:0] ? image_1896 : _GEN_20396; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20398 = 12'h769 == _T_196[11:0] ? image_1897 : _GEN_20397; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20399 = 12'h76a == _T_196[11:0] ? image_1898 : _GEN_20398; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20400 = 12'h76b == _T_196[11:0] ? image_1899 : _GEN_20399; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20401 = 12'h76c == _T_196[11:0] ? image_1900 : _GEN_20400; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20402 = 12'h76d == _T_196[11:0] ? image_1901 : _GEN_20401; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20403 = 12'h76e == _T_196[11:0] ? image_1902 : _GEN_20402; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20404 = 12'h76f == _T_196[11:0] ? image_1903 : _GEN_20403; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20405 = 12'h770 == _T_196[11:0] ? image_1904 : _GEN_20404; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20406 = 12'h771 == _T_196[11:0] ? image_1905 : _GEN_20405; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20407 = 12'h772 == _T_196[11:0] ? image_1906 : _GEN_20406; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20408 = 12'h773 == _T_196[11:0] ? image_1907 : _GEN_20407; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20409 = 12'h774 == _T_196[11:0] ? image_1908 : _GEN_20408; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20410 = 12'h775 == _T_196[11:0] ? image_1909 : _GEN_20409; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20411 = 12'h776 == _T_196[11:0] ? image_1910 : _GEN_20410; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20412 = 12'h777 == _T_196[11:0] ? image_1911 : _GEN_20411; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20413 = 12'h778 == _T_196[11:0] ? image_1912 : _GEN_20412; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20414 = 12'h779 == _T_196[11:0] ? image_1913 : _GEN_20413; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20415 = 12'h77a == _T_196[11:0] ? 4'h0 : _GEN_20414; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20416 = 12'h77b == _T_196[11:0] ? 4'h0 : _GEN_20415; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20417 = 12'h77c == _T_196[11:0] ? 4'h0 : _GEN_20416; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20418 = 12'h77d == _T_196[11:0] ? 4'h0 : _GEN_20417; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20419 = 12'h77e == _T_196[11:0] ? 4'h0 : _GEN_20418; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20420 = 12'h77f == _T_196[11:0] ? 4'h0 : _GEN_20419; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20421 = 12'h780 == _T_196[11:0] ? 4'h0 : _GEN_20420; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20422 = 12'h781 == _T_196[11:0] ? image_1921 : _GEN_20421; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20423 = 12'h782 == _T_196[11:0] ? image_1922 : _GEN_20422; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20424 = 12'h783 == _T_196[11:0] ? image_1923 : _GEN_20423; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20425 = 12'h784 == _T_196[11:0] ? image_1924 : _GEN_20424; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20426 = 12'h785 == _T_196[11:0] ? image_1925 : _GEN_20425; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20427 = 12'h786 == _T_196[11:0] ? image_1926 : _GEN_20426; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20428 = 12'h787 == _T_196[11:0] ? image_1927 : _GEN_20427; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20429 = 12'h788 == _T_196[11:0] ? image_1928 : _GEN_20428; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20430 = 12'h789 == _T_196[11:0] ? image_1929 : _GEN_20429; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20431 = 12'h78a == _T_196[11:0] ? image_1930 : _GEN_20430; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20432 = 12'h78b == _T_196[11:0] ? image_1931 : _GEN_20431; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20433 = 12'h78c == _T_196[11:0] ? image_1932 : _GEN_20432; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20434 = 12'h78d == _T_196[11:0] ? image_1933 : _GEN_20433; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20435 = 12'h78e == _T_196[11:0] ? image_1934 : _GEN_20434; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20436 = 12'h78f == _T_196[11:0] ? image_1935 : _GEN_20435; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20437 = 12'h790 == _T_196[11:0] ? image_1936 : _GEN_20436; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20438 = 12'h791 == _T_196[11:0] ? image_1937 : _GEN_20437; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20439 = 12'h792 == _T_196[11:0] ? image_1938 : _GEN_20438; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20440 = 12'h793 == _T_196[11:0] ? image_1939 : _GEN_20439; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20441 = 12'h794 == _T_196[11:0] ? image_1940 : _GEN_20440; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20442 = 12'h795 == _T_196[11:0] ? image_1941 : _GEN_20441; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20443 = 12'h796 == _T_196[11:0] ? image_1942 : _GEN_20442; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20444 = 12'h797 == _T_196[11:0] ? image_1943 : _GEN_20443; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20445 = 12'h798 == _T_196[11:0] ? image_1944 : _GEN_20444; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20446 = 12'h799 == _T_196[11:0] ? image_1945 : _GEN_20445; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20447 = 12'h79a == _T_196[11:0] ? image_1946 : _GEN_20446; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20448 = 12'h79b == _T_196[11:0] ? image_1947 : _GEN_20447; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20449 = 12'h79c == _T_196[11:0] ? image_1948 : _GEN_20448; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20450 = 12'h79d == _T_196[11:0] ? image_1949 : _GEN_20449; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20451 = 12'h79e == _T_196[11:0] ? image_1950 : _GEN_20450; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20452 = 12'h79f == _T_196[11:0] ? image_1951 : _GEN_20451; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20453 = 12'h7a0 == _T_196[11:0] ? image_1952 : _GEN_20452; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20454 = 12'h7a1 == _T_196[11:0] ? image_1953 : _GEN_20453; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20455 = 12'h7a2 == _T_196[11:0] ? image_1954 : _GEN_20454; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20456 = 12'h7a3 == _T_196[11:0] ? image_1955 : _GEN_20455; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20457 = 12'h7a4 == _T_196[11:0] ? image_1956 : _GEN_20456; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20458 = 12'h7a5 == _T_196[11:0] ? image_1957 : _GEN_20457; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20459 = 12'h7a6 == _T_196[11:0] ? image_1958 : _GEN_20458; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20460 = 12'h7a7 == _T_196[11:0] ? image_1959 : _GEN_20459; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20461 = 12'h7a8 == _T_196[11:0] ? image_1960 : _GEN_20460; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20462 = 12'h7a9 == _T_196[11:0] ? image_1961 : _GEN_20461; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20463 = 12'h7aa == _T_196[11:0] ? image_1962 : _GEN_20462; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20464 = 12'h7ab == _T_196[11:0] ? image_1963 : _GEN_20463; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20465 = 12'h7ac == _T_196[11:0] ? image_1964 : _GEN_20464; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20466 = 12'h7ad == _T_196[11:0] ? image_1965 : _GEN_20465; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20467 = 12'h7ae == _T_196[11:0] ? image_1966 : _GEN_20466; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20468 = 12'h7af == _T_196[11:0] ? image_1967 : _GEN_20467; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20469 = 12'h7b0 == _T_196[11:0] ? image_1968 : _GEN_20468; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20470 = 12'h7b1 == _T_196[11:0] ? image_1969 : _GEN_20469; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20471 = 12'h7b2 == _T_196[11:0] ? image_1970 : _GEN_20470; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20472 = 12'h7b3 == _T_196[11:0] ? image_1971 : _GEN_20471; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20473 = 12'h7b4 == _T_196[11:0] ? image_1972 : _GEN_20472; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20474 = 12'h7b5 == _T_196[11:0] ? image_1973 : _GEN_20473; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20475 = 12'h7b6 == _T_196[11:0] ? image_1974 : _GEN_20474; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20476 = 12'h7b7 == _T_196[11:0] ? image_1975 : _GEN_20475; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20477 = 12'h7b8 == _T_196[11:0] ? image_1976 : _GEN_20476; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20478 = 12'h7b9 == _T_196[11:0] ? image_1977 : _GEN_20477; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20479 = 12'h7ba == _T_196[11:0] ? 4'h0 : _GEN_20478; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20480 = 12'h7bb == _T_196[11:0] ? 4'h0 : _GEN_20479; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20481 = 12'h7bc == _T_196[11:0] ? 4'h0 : _GEN_20480; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20482 = 12'h7bd == _T_196[11:0] ? 4'h0 : _GEN_20481; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20483 = 12'h7be == _T_196[11:0] ? 4'h0 : _GEN_20482; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20484 = 12'h7bf == _T_196[11:0] ? 4'h0 : _GEN_20483; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20485 = 12'h7c0 == _T_196[11:0] ? 4'h0 : _GEN_20484; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20486 = 12'h7c1 == _T_196[11:0] ? image_1985 : _GEN_20485; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20487 = 12'h7c2 == _T_196[11:0] ? image_1986 : _GEN_20486; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20488 = 12'h7c3 == _T_196[11:0] ? image_1987 : _GEN_20487; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20489 = 12'h7c4 == _T_196[11:0] ? image_1988 : _GEN_20488; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20490 = 12'h7c5 == _T_196[11:0] ? image_1989 : _GEN_20489; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20491 = 12'h7c6 == _T_196[11:0] ? image_1990 : _GEN_20490; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20492 = 12'h7c7 == _T_196[11:0] ? image_1991 : _GEN_20491; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20493 = 12'h7c8 == _T_196[11:0] ? image_1992 : _GEN_20492; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20494 = 12'h7c9 == _T_196[11:0] ? image_1993 : _GEN_20493; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20495 = 12'h7ca == _T_196[11:0] ? image_1994 : _GEN_20494; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20496 = 12'h7cb == _T_196[11:0] ? image_1995 : _GEN_20495; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20497 = 12'h7cc == _T_196[11:0] ? image_1996 : _GEN_20496; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20498 = 12'h7cd == _T_196[11:0] ? image_1997 : _GEN_20497; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20499 = 12'h7ce == _T_196[11:0] ? image_1998 : _GEN_20498; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20500 = 12'h7cf == _T_196[11:0] ? image_1999 : _GEN_20499; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20501 = 12'h7d0 == _T_196[11:0] ? image_2000 : _GEN_20500; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20502 = 12'h7d1 == _T_196[11:0] ? image_2001 : _GEN_20501; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20503 = 12'h7d2 == _T_196[11:0] ? image_2002 : _GEN_20502; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20504 = 12'h7d3 == _T_196[11:0] ? image_2003 : _GEN_20503; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20505 = 12'h7d4 == _T_196[11:0] ? image_2004 : _GEN_20504; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20506 = 12'h7d5 == _T_196[11:0] ? image_2005 : _GEN_20505; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20507 = 12'h7d6 == _T_196[11:0] ? image_2006 : _GEN_20506; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20508 = 12'h7d7 == _T_196[11:0] ? image_2007 : _GEN_20507; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20509 = 12'h7d8 == _T_196[11:0] ? image_2008 : _GEN_20508; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20510 = 12'h7d9 == _T_196[11:0] ? image_2009 : _GEN_20509; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20511 = 12'h7da == _T_196[11:0] ? image_2010 : _GEN_20510; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20512 = 12'h7db == _T_196[11:0] ? image_2011 : _GEN_20511; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20513 = 12'h7dc == _T_196[11:0] ? image_2012 : _GEN_20512; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20514 = 12'h7dd == _T_196[11:0] ? image_2013 : _GEN_20513; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20515 = 12'h7de == _T_196[11:0] ? image_2014 : _GEN_20514; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20516 = 12'h7df == _T_196[11:0] ? image_2015 : _GEN_20515; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20517 = 12'h7e0 == _T_196[11:0] ? image_2016 : _GEN_20516; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20518 = 12'h7e1 == _T_196[11:0] ? image_2017 : _GEN_20517; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20519 = 12'h7e2 == _T_196[11:0] ? image_2018 : _GEN_20518; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20520 = 12'h7e3 == _T_196[11:0] ? image_2019 : _GEN_20519; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20521 = 12'h7e4 == _T_196[11:0] ? image_2020 : _GEN_20520; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20522 = 12'h7e5 == _T_196[11:0] ? image_2021 : _GEN_20521; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20523 = 12'h7e6 == _T_196[11:0] ? image_2022 : _GEN_20522; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20524 = 12'h7e7 == _T_196[11:0] ? image_2023 : _GEN_20523; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20525 = 12'h7e8 == _T_196[11:0] ? image_2024 : _GEN_20524; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20526 = 12'h7e9 == _T_196[11:0] ? image_2025 : _GEN_20525; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20527 = 12'h7ea == _T_196[11:0] ? image_2026 : _GEN_20526; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20528 = 12'h7eb == _T_196[11:0] ? image_2027 : _GEN_20527; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20529 = 12'h7ec == _T_196[11:0] ? image_2028 : _GEN_20528; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20530 = 12'h7ed == _T_196[11:0] ? image_2029 : _GEN_20529; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20531 = 12'h7ee == _T_196[11:0] ? image_2030 : _GEN_20530; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20532 = 12'h7ef == _T_196[11:0] ? image_2031 : _GEN_20531; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20533 = 12'h7f0 == _T_196[11:0] ? image_2032 : _GEN_20532; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20534 = 12'h7f1 == _T_196[11:0] ? image_2033 : _GEN_20533; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20535 = 12'h7f2 == _T_196[11:0] ? image_2034 : _GEN_20534; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20536 = 12'h7f3 == _T_196[11:0] ? image_2035 : _GEN_20535; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20537 = 12'h7f4 == _T_196[11:0] ? image_2036 : _GEN_20536; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20538 = 12'h7f5 == _T_196[11:0] ? image_2037 : _GEN_20537; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20539 = 12'h7f6 == _T_196[11:0] ? image_2038 : _GEN_20538; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20540 = 12'h7f7 == _T_196[11:0] ? image_2039 : _GEN_20539; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20541 = 12'h7f8 == _T_196[11:0] ? image_2040 : _GEN_20540; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20542 = 12'h7f9 == _T_196[11:0] ? image_2041 : _GEN_20541; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20543 = 12'h7fa == _T_196[11:0] ? 4'h0 : _GEN_20542; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20544 = 12'h7fb == _T_196[11:0] ? 4'h0 : _GEN_20543; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20545 = 12'h7fc == _T_196[11:0] ? 4'h0 : _GEN_20544; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20546 = 12'h7fd == _T_196[11:0] ? 4'h0 : _GEN_20545; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20547 = 12'h7fe == _T_196[11:0] ? 4'h0 : _GEN_20546; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20548 = 12'h7ff == _T_196[11:0] ? 4'h0 : _GEN_20547; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20549 = 12'h800 == _T_196[11:0] ? 4'h0 : _GEN_20548; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20550 = 12'h801 == _T_196[11:0] ? image_2049 : _GEN_20549; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20551 = 12'h802 == _T_196[11:0] ? image_2050 : _GEN_20550; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20552 = 12'h803 == _T_196[11:0] ? image_2051 : _GEN_20551; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20553 = 12'h804 == _T_196[11:0] ? image_2052 : _GEN_20552; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20554 = 12'h805 == _T_196[11:0] ? image_2053 : _GEN_20553; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20555 = 12'h806 == _T_196[11:0] ? image_2054 : _GEN_20554; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20556 = 12'h807 == _T_196[11:0] ? image_2055 : _GEN_20555; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20557 = 12'h808 == _T_196[11:0] ? image_2056 : _GEN_20556; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20558 = 12'h809 == _T_196[11:0] ? image_2057 : _GEN_20557; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20559 = 12'h80a == _T_196[11:0] ? image_2058 : _GEN_20558; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20560 = 12'h80b == _T_196[11:0] ? image_2059 : _GEN_20559; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20561 = 12'h80c == _T_196[11:0] ? image_2060 : _GEN_20560; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20562 = 12'h80d == _T_196[11:0] ? image_2061 : _GEN_20561; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20563 = 12'h80e == _T_196[11:0] ? image_2062 : _GEN_20562; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20564 = 12'h80f == _T_196[11:0] ? image_2063 : _GEN_20563; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20565 = 12'h810 == _T_196[11:0] ? image_2064 : _GEN_20564; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20566 = 12'h811 == _T_196[11:0] ? image_2065 : _GEN_20565; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20567 = 12'h812 == _T_196[11:0] ? image_2066 : _GEN_20566; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20568 = 12'h813 == _T_196[11:0] ? image_2067 : _GEN_20567; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20569 = 12'h814 == _T_196[11:0] ? image_2068 : _GEN_20568; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20570 = 12'h815 == _T_196[11:0] ? image_2069 : _GEN_20569; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20571 = 12'h816 == _T_196[11:0] ? image_2070 : _GEN_20570; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20572 = 12'h817 == _T_196[11:0] ? image_2071 : _GEN_20571; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20573 = 12'h818 == _T_196[11:0] ? image_2072 : _GEN_20572; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20574 = 12'h819 == _T_196[11:0] ? image_2073 : _GEN_20573; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20575 = 12'h81a == _T_196[11:0] ? image_2074 : _GEN_20574; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20576 = 12'h81b == _T_196[11:0] ? image_2075 : _GEN_20575; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20577 = 12'h81c == _T_196[11:0] ? image_2076 : _GEN_20576; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20578 = 12'h81d == _T_196[11:0] ? image_2077 : _GEN_20577; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20579 = 12'h81e == _T_196[11:0] ? image_2078 : _GEN_20578; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20580 = 12'h81f == _T_196[11:0] ? image_2079 : _GEN_20579; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20581 = 12'h820 == _T_196[11:0] ? image_2080 : _GEN_20580; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20582 = 12'h821 == _T_196[11:0] ? image_2081 : _GEN_20581; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20583 = 12'h822 == _T_196[11:0] ? image_2082 : _GEN_20582; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20584 = 12'h823 == _T_196[11:0] ? image_2083 : _GEN_20583; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20585 = 12'h824 == _T_196[11:0] ? image_2084 : _GEN_20584; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20586 = 12'h825 == _T_196[11:0] ? image_2085 : _GEN_20585; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20587 = 12'h826 == _T_196[11:0] ? image_2086 : _GEN_20586; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20588 = 12'h827 == _T_196[11:0] ? image_2087 : _GEN_20587; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20589 = 12'h828 == _T_196[11:0] ? image_2088 : _GEN_20588; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20590 = 12'h829 == _T_196[11:0] ? image_2089 : _GEN_20589; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20591 = 12'h82a == _T_196[11:0] ? image_2090 : _GEN_20590; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20592 = 12'h82b == _T_196[11:0] ? image_2091 : _GEN_20591; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20593 = 12'h82c == _T_196[11:0] ? image_2092 : _GEN_20592; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20594 = 12'h82d == _T_196[11:0] ? image_2093 : _GEN_20593; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20595 = 12'h82e == _T_196[11:0] ? image_2094 : _GEN_20594; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20596 = 12'h82f == _T_196[11:0] ? image_2095 : _GEN_20595; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20597 = 12'h830 == _T_196[11:0] ? image_2096 : _GEN_20596; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20598 = 12'h831 == _T_196[11:0] ? image_2097 : _GEN_20597; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20599 = 12'h832 == _T_196[11:0] ? image_2098 : _GEN_20598; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20600 = 12'h833 == _T_196[11:0] ? image_2099 : _GEN_20599; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20601 = 12'h834 == _T_196[11:0] ? image_2100 : _GEN_20600; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20602 = 12'h835 == _T_196[11:0] ? image_2101 : _GEN_20601; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20603 = 12'h836 == _T_196[11:0] ? image_2102 : _GEN_20602; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20604 = 12'h837 == _T_196[11:0] ? image_2103 : _GEN_20603; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20605 = 12'h838 == _T_196[11:0] ? image_2104 : _GEN_20604; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20606 = 12'h839 == _T_196[11:0] ? image_2105 : _GEN_20605; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20607 = 12'h83a == _T_196[11:0] ? image_2106 : _GEN_20606; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20608 = 12'h83b == _T_196[11:0] ? 4'h0 : _GEN_20607; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20609 = 12'h83c == _T_196[11:0] ? 4'h0 : _GEN_20608; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20610 = 12'h83d == _T_196[11:0] ? 4'h0 : _GEN_20609; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20611 = 12'h83e == _T_196[11:0] ? 4'h0 : _GEN_20610; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20612 = 12'h83f == _T_196[11:0] ? 4'h0 : _GEN_20611; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20613 = 12'h840 == _T_196[11:0] ? 4'h0 : _GEN_20612; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20614 = 12'h841 == _T_196[11:0] ? 4'h0 : _GEN_20613; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20615 = 12'h842 == _T_196[11:0] ? image_2114 : _GEN_20614; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20616 = 12'h843 == _T_196[11:0] ? image_2115 : _GEN_20615; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20617 = 12'h844 == _T_196[11:0] ? image_2116 : _GEN_20616; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20618 = 12'h845 == _T_196[11:0] ? image_2117 : _GEN_20617; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20619 = 12'h846 == _T_196[11:0] ? image_2118 : _GEN_20618; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20620 = 12'h847 == _T_196[11:0] ? image_2119 : _GEN_20619; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20621 = 12'h848 == _T_196[11:0] ? image_2120 : _GEN_20620; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20622 = 12'h849 == _T_196[11:0] ? image_2121 : _GEN_20621; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20623 = 12'h84a == _T_196[11:0] ? image_2122 : _GEN_20622; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20624 = 12'h84b == _T_196[11:0] ? image_2123 : _GEN_20623; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20625 = 12'h84c == _T_196[11:0] ? image_2124 : _GEN_20624; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20626 = 12'h84d == _T_196[11:0] ? image_2125 : _GEN_20625; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20627 = 12'h84e == _T_196[11:0] ? image_2126 : _GEN_20626; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20628 = 12'h84f == _T_196[11:0] ? image_2127 : _GEN_20627; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20629 = 12'h850 == _T_196[11:0] ? image_2128 : _GEN_20628; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20630 = 12'h851 == _T_196[11:0] ? image_2129 : _GEN_20629; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20631 = 12'h852 == _T_196[11:0] ? image_2130 : _GEN_20630; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20632 = 12'h853 == _T_196[11:0] ? image_2131 : _GEN_20631; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20633 = 12'h854 == _T_196[11:0] ? image_2132 : _GEN_20632; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20634 = 12'h855 == _T_196[11:0] ? image_2133 : _GEN_20633; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20635 = 12'h856 == _T_196[11:0] ? image_2134 : _GEN_20634; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20636 = 12'h857 == _T_196[11:0] ? image_2135 : _GEN_20635; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20637 = 12'h858 == _T_196[11:0] ? image_2136 : _GEN_20636; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20638 = 12'h859 == _T_196[11:0] ? image_2137 : _GEN_20637; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20639 = 12'h85a == _T_196[11:0] ? image_2138 : _GEN_20638; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20640 = 12'h85b == _T_196[11:0] ? image_2139 : _GEN_20639; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20641 = 12'h85c == _T_196[11:0] ? image_2140 : _GEN_20640; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20642 = 12'h85d == _T_196[11:0] ? image_2141 : _GEN_20641; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20643 = 12'h85e == _T_196[11:0] ? image_2142 : _GEN_20642; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20644 = 12'h85f == _T_196[11:0] ? image_2143 : _GEN_20643; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20645 = 12'h860 == _T_196[11:0] ? image_2144 : _GEN_20644; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20646 = 12'h861 == _T_196[11:0] ? image_2145 : _GEN_20645; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20647 = 12'h862 == _T_196[11:0] ? image_2146 : _GEN_20646; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20648 = 12'h863 == _T_196[11:0] ? image_2147 : _GEN_20647; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20649 = 12'h864 == _T_196[11:0] ? image_2148 : _GEN_20648; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20650 = 12'h865 == _T_196[11:0] ? image_2149 : _GEN_20649; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20651 = 12'h866 == _T_196[11:0] ? image_2150 : _GEN_20650; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20652 = 12'h867 == _T_196[11:0] ? image_2151 : _GEN_20651; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20653 = 12'h868 == _T_196[11:0] ? image_2152 : _GEN_20652; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20654 = 12'h869 == _T_196[11:0] ? image_2153 : _GEN_20653; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20655 = 12'h86a == _T_196[11:0] ? image_2154 : _GEN_20654; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20656 = 12'h86b == _T_196[11:0] ? image_2155 : _GEN_20655; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20657 = 12'h86c == _T_196[11:0] ? image_2156 : _GEN_20656; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20658 = 12'h86d == _T_196[11:0] ? image_2157 : _GEN_20657; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20659 = 12'h86e == _T_196[11:0] ? image_2158 : _GEN_20658; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20660 = 12'h86f == _T_196[11:0] ? image_2159 : _GEN_20659; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20661 = 12'h870 == _T_196[11:0] ? image_2160 : _GEN_20660; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20662 = 12'h871 == _T_196[11:0] ? image_2161 : _GEN_20661; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20663 = 12'h872 == _T_196[11:0] ? image_2162 : _GEN_20662; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20664 = 12'h873 == _T_196[11:0] ? image_2163 : _GEN_20663; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20665 = 12'h874 == _T_196[11:0] ? image_2164 : _GEN_20664; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20666 = 12'h875 == _T_196[11:0] ? image_2165 : _GEN_20665; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20667 = 12'h876 == _T_196[11:0] ? image_2166 : _GEN_20666; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20668 = 12'h877 == _T_196[11:0] ? image_2167 : _GEN_20667; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20669 = 12'h878 == _T_196[11:0] ? image_2168 : _GEN_20668; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20670 = 12'h879 == _T_196[11:0] ? image_2169 : _GEN_20669; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20671 = 12'h87a == _T_196[11:0] ? image_2170 : _GEN_20670; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20672 = 12'h87b == _T_196[11:0] ? 4'h0 : _GEN_20671; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20673 = 12'h87c == _T_196[11:0] ? 4'h0 : _GEN_20672; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20674 = 12'h87d == _T_196[11:0] ? 4'h0 : _GEN_20673; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20675 = 12'h87e == _T_196[11:0] ? 4'h0 : _GEN_20674; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20676 = 12'h87f == _T_196[11:0] ? 4'h0 : _GEN_20675; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20677 = 12'h880 == _T_196[11:0] ? 4'h0 : _GEN_20676; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20678 = 12'h881 == _T_196[11:0] ? image_2177 : _GEN_20677; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20679 = 12'h882 == _T_196[11:0] ? image_2178 : _GEN_20678; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20680 = 12'h883 == _T_196[11:0] ? image_2179 : _GEN_20679; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20681 = 12'h884 == _T_196[11:0] ? image_2180 : _GEN_20680; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20682 = 12'h885 == _T_196[11:0] ? image_2181 : _GEN_20681; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20683 = 12'h886 == _T_196[11:0] ? image_2182 : _GEN_20682; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20684 = 12'h887 == _T_196[11:0] ? image_2183 : _GEN_20683; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20685 = 12'h888 == _T_196[11:0] ? image_2184 : _GEN_20684; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20686 = 12'h889 == _T_196[11:0] ? image_2185 : _GEN_20685; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20687 = 12'h88a == _T_196[11:0] ? image_2186 : _GEN_20686; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20688 = 12'h88b == _T_196[11:0] ? image_2187 : _GEN_20687; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20689 = 12'h88c == _T_196[11:0] ? image_2188 : _GEN_20688; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20690 = 12'h88d == _T_196[11:0] ? image_2189 : _GEN_20689; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20691 = 12'h88e == _T_196[11:0] ? image_2190 : _GEN_20690; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20692 = 12'h88f == _T_196[11:0] ? image_2191 : _GEN_20691; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20693 = 12'h890 == _T_196[11:0] ? image_2192 : _GEN_20692; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20694 = 12'h891 == _T_196[11:0] ? image_2193 : _GEN_20693; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20695 = 12'h892 == _T_196[11:0] ? image_2194 : _GEN_20694; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20696 = 12'h893 == _T_196[11:0] ? image_2195 : _GEN_20695; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20697 = 12'h894 == _T_196[11:0] ? image_2196 : _GEN_20696; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20698 = 12'h895 == _T_196[11:0] ? image_2197 : _GEN_20697; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20699 = 12'h896 == _T_196[11:0] ? image_2198 : _GEN_20698; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20700 = 12'h897 == _T_196[11:0] ? image_2199 : _GEN_20699; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20701 = 12'h898 == _T_196[11:0] ? image_2200 : _GEN_20700; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20702 = 12'h899 == _T_196[11:0] ? image_2201 : _GEN_20701; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20703 = 12'h89a == _T_196[11:0] ? image_2202 : _GEN_20702; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20704 = 12'h89b == _T_196[11:0] ? image_2203 : _GEN_20703; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20705 = 12'h89c == _T_196[11:0] ? image_2204 : _GEN_20704; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20706 = 12'h89d == _T_196[11:0] ? image_2205 : _GEN_20705; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20707 = 12'h89e == _T_196[11:0] ? image_2206 : _GEN_20706; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20708 = 12'h89f == _T_196[11:0] ? image_2207 : _GEN_20707; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20709 = 12'h8a0 == _T_196[11:0] ? image_2208 : _GEN_20708; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20710 = 12'h8a1 == _T_196[11:0] ? image_2209 : _GEN_20709; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20711 = 12'h8a2 == _T_196[11:0] ? image_2210 : _GEN_20710; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20712 = 12'h8a3 == _T_196[11:0] ? image_2211 : _GEN_20711; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20713 = 12'h8a4 == _T_196[11:0] ? image_2212 : _GEN_20712; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20714 = 12'h8a5 == _T_196[11:0] ? image_2213 : _GEN_20713; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20715 = 12'h8a6 == _T_196[11:0] ? image_2214 : _GEN_20714; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20716 = 12'h8a7 == _T_196[11:0] ? image_2215 : _GEN_20715; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20717 = 12'h8a8 == _T_196[11:0] ? image_2216 : _GEN_20716; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20718 = 12'h8a9 == _T_196[11:0] ? image_2217 : _GEN_20717; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20719 = 12'h8aa == _T_196[11:0] ? image_2218 : _GEN_20718; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20720 = 12'h8ab == _T_196[11:0] ? image_2219 : _GEN_20719; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20721 = 12'h8ac == _T_196[11:0] ? image_2220 : _GEN_20720; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20722 = 12'h8ad == _T_196[11:0] ? image_2221 : _GEN_20721; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20723 = 12'h8ae == _T_196[11:0] ? image_2222 : _GEN_20722; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20724 = 12'h8af == _T_196[11:0] ? image_2223 : _GEN_20723; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20725 = 12'h8b0 == _T_196[11:0] ? image_2224 : _GEN_20724; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20726 = 12'h8b1 == _T_196[11:0] ? image_2225 : _GEN_20725; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20727 = 12'h8b2 == _T_196[11:0] ? image_2226 : _GEN_20726; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20728 = 12'h8b3 == _T_196[11:0] ? image_2227 : _GEN_20727; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20729 = 12'h8b4 == _T_196[11:0] ? image_2228 : _GEN_20728; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20730 = 12'h8b5 == _T_196[11:0] ? image_2229 : _GEN_20729; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20731 = 12'h8b6 == _T_196[11:0] ? image_2230 : _GEN_20730; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20732 = 12'h8b7 == _T_196[11:0] ? image_2231 : _GEN_20731; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20733 = 12'h8b8 == _T_196[11:0] ? image_2232 : _GEN_20732; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20734 = 12'h8b9 == _T_196[11:0] ? image_2233 : _GEN_20733; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20735 = 12'h8ba == _T_196[11:0] ? image_2234 : _GEN_20734; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20736 = 12'h8bb == _T_196[11:0] ? 4'h0 : _GEN_20735; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20737 = 12'h8bc == _T_196[11:0] ? 4'h0 : _GEN_20736; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20738 = 12'h8bd == _T_196[11:0] ? 4'h0 : _GEN_20737; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20739 = 12'h8be == _T_196[11:0] ? 4'h0 : _GEN_20738; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20740 = 12'h8bf == _T_196[11:0] ? 4'h0 : _GEN_20739; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20741 = 12'h8c0 == _T_196[11:0] ? 4'h0 : _GEN_20740; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20742 = 12'h8c1 == _T_196[11:0] ? 4'h0 : _GEN_20741; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20743 = 12'h8c2 == _T_196[11:0] ? 4'h0 : _GEN_20742; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20744 = 12'h8c3 == _T_196[11:0] ? image_2243 : _GEN_20743; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20745 = 12'h8c4 == _T_196[11:0] ? image_2244 : _GEN_20744; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20746 = 12'h8c5 == _T_196[11:0] ? image_2245 : _GEN_20745; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20747 = 12'h8c6 == _T_196[11:0] ? image_2246 : _GEN_20746; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20748 = 12'h8c7 == _T_196[11:0] ? image_2247 : _GEN_20747; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20749 = 12'h8c8 == _T_196[11:0] ? image_2248 : _GEN_20748; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20750 = 12'h8c9 == _T_196[11:0] ? image_2249 : _GEN_20749; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20751 = 12'h8ca == _T_196[11:0] ? image_2250 : _GEN_20750; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20752 = 12'h8cb == _T_196[11:0] ? image_2251 : _GEN_20751; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20753 = 12'h8cc == _T_196[11:0] ? image_2252 : _GEN_20752; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20754 = 12'h8cd == _T_196[11:0] ? image_2253 : _GEN_20753; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20755 = 12'h8ce == _T_196[11:0] ? image_2254 : _GEN_20754; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20756 = 12'h8cf == _T_196[11:0] ? image_2255 : _GEN_20755; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20757 = 12'h8d0 == _T_196[11:0] ? image_2256 : _GEN_20756; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20758 = 12'h8d1 == _T_196[11:0] ? image_2257 : _GEN_20757; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20759 = 12'h8d2 == _T_196[11:0] ? image_2258 : _GEN_20758; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20760 = 12'h8d3 == _T_196[11:0] ? image_2259 : _GEN_20759; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20761 = 12'h8d4 == _T_196[11:0] ? image_2260 : _GEN_20760; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20762 = 12'h8d5 == _T_196[11:0] ? image_2261 : _GEN_20761; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20763 = 12'h8d6 == _T_196[11:0] ? image_2262 : _GEN_20762; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20764 = 12'h8d7 == _T_196[11:0] ? image_2263 : _GEN_20763; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20765 = 12'h8d8 == _T_196[11:0] ? image_2264 : _GEN_20764; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20766 = 12'h8d9 == _T_196[11:0] ? image_2265 : _GEN_20765; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20767 = 12'h8da == _T_196[11:0] ? image_2266 : _GEN_20766; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20768 = 12'h8db == _T_196[11:0] ? image_2267 : _GEN_20767; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20769 = 12'h8dc == _T_196[11:0] ? image_2268 : _GEN_20768; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20770 = 12'h8dd == _T_196[11:0] ? image_2269 : _GEN_20769; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20771 = 12'h8de == _T_196[11:0] ? image_2270 : _GEN_20770; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20772 = 12'h8df == _T_196[11:0] ? image_2271 : _GEN_20771; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20773 = 12'h8e0 == _T_196[11:0] ? image_2272 : _GEN_20772; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20774 = 12'h8e1 == _T_196[11:0] ? image_2273 : _GEN_20773; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20775 = 12'h8e2 == _T_196[11:0] ? image_2274 : _GEN_20774; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20776 = 12'h8e3 == _T_196[11:0] ? image_2275 : _GEN_20775; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20777 = 12'h8e4 == _T_196[11:0] ? image_2276 : _GEN_20776; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20778 = 12'h8e5 == _T_196[11:0] ? image_2277 : _GEN_20777; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20779 = 12'h8e6 == _T_196[11:0] ? image_2278 : _GEN_20778; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20780 = 12'h8e7 == _T_196[11:0] ? image_2279 : _GEN_20779; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20781 = 12'h8e8 == _T_196[11:0] ? image_2280 : _GEN_20780; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20782 = 12'h8e9 == _T_196[11:0] ? image_2281 : _GEN_20781; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20783 = 12'h8ea == _T_196[11:0] ? image_2282 : _GEN_20782; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20784 = 12'h8eb == _T_196[11:0] ? image_2283 : _GEN_20783; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20785 = 12'h8ec == _T_196[11:0] ? image_2284 : _GEN_20784; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20786 = 12'h8ed == _T_196[11:0] ? image_2285 : _GEN_20785; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20787 = 12'h8ee == _T_196[11:0] ? image_2286 : _GEN_20786; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20788 = 12'h8ef == _T_196[11:0] ? image_2287 : _GEN_20787; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20789 = 12'h8f0 == _T_196[11:0] ? image_2288 : _GEN_20788; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20790 = 12'h8f1 == _T_196[11:0] ? image_2289 : _GEN_20789; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20791 = 12'h8f2 == _T_196[11:0] ? image_2290 : _GEN_20790; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20792 = 12'h8f3 == _T_196[11:0] ? image_2291 : _GEN_20791; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20793 = 12'h8f4 == _T_196[11:0] ? image_2292 : _GEN_20792; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20794 = 12'h8f5 == _T_196[11:0] ? image_2293 : _GEN_20793; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20795 = 12'h8f6 == _T_196[11:0] ? image_2294 : _GEN_20794; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20796 = 12'h8f7 == _T_196[11:0] ? image_2295 : _GEN_20795; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20797 = 12'h8f8 == _T_196[11:0] ? image_2296 : _GEN_20796; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20798 = 12'h8f9 == _T_196[11:0] ? image_2297 : _GEN_20797; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20799 = 12'h8fa == _T_196[11:0] ? image_2298 : _GEN_20798; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20800 = 12'h8fb == _T_196[11:0] ? 4'h0 : _GEN_20799; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20801 = 12'h8fc == _T_196[11:0] ? 4'h0 : _GEN_20800; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20802 = 12'h8fd == _T_196[11:0] ? 4'h0 : _GEN_20801; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20803 = 12'h8fe == _T_196[11:0] ? 4'h0 : _GEN_20802; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20804 = 12'h8ff == _T_196[11:0] ? 4'h0 : _GEN_20803; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20805 = 12'h900 == _T_196[11:0] ? 4'h0 : _GEN_20804; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20806 = 12'h901 == _T_196[11:0] ? 4'h0 : _GEN_20805; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20807 = 12'h902 == _T_196[11:0] ? 4'h0 : _GEN_20806; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20808 = 12'h903 == _T_196[11:0] ? image_2307 : _GEN_20807; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20809 = 12'h904 == _T_196[11:0] ? image_2308 : _GEN_20808; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20810 = 12'h905 == _T_196[11:0] ? image_2309 : _GEN_20809; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20811 = 12'h906 == _T_196[11:0] ? image_2310 : _GEN_20810; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20812 = 12'h907 == _T_196[11:0] ? image_2311 : _GEN_20811; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20813 = 12'h908 == _T_196[11:0] ? image_2312 : _GEN_20812; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20814 = 12'h909 == _T_196[11:0] ? image_2313 : _GEN_20813; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20815 = 12'h90a == _T_196[11:0] ? image_2314 : _GEN_20814; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20816 = 12'h90b == _T_196[11:0] ? image_2315 : _GEN_20815; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20817 = 12'h90c == _T_196[11:0] ? image_2316 : _GEN_20816; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20818 = 12'h90d == _T_196[11:0] ? image_2317 : _GEN_20817; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20819 = 12'h90e == _T_196[11:0] ? image_2318 : _GEN_20818; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20820 = 12'h90f == _T_196[11:0] ? image_2319 : _GEN_20819; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20821 = 12'h910 == _T_196[11:0] ? image_2320 : _GEN_20820; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20822 = 12'h911 == _T_196[11:0] ? image_2321 : _GEN_20821; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20823 = 12'h912 == _T_196[11:0] ? image_2322 : _GEN_20822; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20824 = 12'h913 == _T_196[11:0] ? image_2323 : _GEN_20823; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20825 = 12'h914 == _T_196[11:0] ? image_2324 : _GEN_20824; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20826 = 12'h915 == _T_196[11:0] ? image_2325 : _GEN_20825; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20827 = 12'h916 == _T_196[11:0] ? image_2326 : _GEN_20826; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20828 = 12'h917 == _T_196[11:0] ? image_2327 : _GEN_20827; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20829 = 12'h918 == _T_196[11:0] ? image_2328 : _GEN_20828; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20830 = 12'h919 == _T_196[11:0] ? image_2329 : _GEN_20829; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20831 = 12'h91a == _T_196[11:0] ? image_2330 : _GEN_20830; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20832 = 12'h91b == _T_196[11:0] ? image_2331 : _GEN_20831; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20833 = 12'h91c == _T_196[11:0] ? image_2332 : _GEN_20832; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20834 = 12'h91d == _T_196[11:0] ? image_2333 : _GEN_20833; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20835 = 12'h91e == _T_196[11:0] ? image_2334 : _GEN_20834; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20836 = 12'h91f == _T_196[11:0] ? image_2335 : _GEN_20835; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20837 = 12'h920 == _T_196[11:0] ? image_2336 : _GEN_20836; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20838 = 12'h921 == _T_196[11:0] ? image_2337 : _GEN_20837; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20839 = 12'h922 == _T_196[11:0] ? image_2338 : _GEN_20838; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20840 = 12'h923 == _T_196[11:0] ? image_2339 : _GEN_20839; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20841 = 12'h924 == _T_196[11:0] ? image_2340 : _GEN_20840; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20842 = 12'h925 == _T_196[11:0] ? image_2341 : _GEN_20841; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20843 = 12'h926 == _T_196[11:0] ? image_2342 : _GEN_20842; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20844 = 12'h927 == _T_196[11:0] ? image_2343 : _GEN_20843; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20845 = 12'h928 == _T_196[11:0] ? image_2344 : _GEN_20844; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20846 = 12'h929 == _T_196[11:0] ? image_2345 : _GEN_20845; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20847 = 12'h92a == _T_196[11:0] ? image_2346 : _GEN_20846; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20848 = 12'h92b == _T_196[11:0] ? image_2347 : _GEN_20847; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20849 = 12'h92c == _T_196[11:0] ? image_2348 : _GEN_20848; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20850 = 12'h92d == _T_196[11:0] ? image_2349 : _GEN_20849; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20851 = 12'h92e == _T_196[11:0] ? image_2350 : _GEN_20850; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20852 = 12'h92f == _T_196[11:0] ? image_2351 : _GEN_20851; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20853 = 12'h930 == _T_196[11:0] ? image_2352 : _GEN_20852; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20854 = 12'h931 == _T_196[11:0] ? image_2353 : _GEN_20853; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20855 = 12'h932 == _T_196[11:0] ? image_2354 : _GEN_20854; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20856 = 12'h933 == _T_196[11:0] ? image_2355 : _GEN_20855; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20857 = 12'h934 == _T_196[11:0] ? image_2356 : _GEN_20856; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20858 = 12'h935 == _T_196[11:0] ? image_2357 : _GEN_20857; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20859 = 12'h936 == _T_196[11:0] ? image_2358 : _GEN_20858; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20860 = 12'h937 == _T_196[11:0] ? image_2359 : _GEN_20859; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20861 = 12'h938 == _T_196[11:0] ? image_2360 : _GEN_20860; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20862 = 12'h939 == _T_196[11:0] ? image_2361 : _GEN_20861; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20863 = 12'h93a == _T_196[11:0] ? image_2362 : _GEN_20862; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20864 = 12'h93b == _T_196[11:0] ? 4'h0 : _GEN_20863; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20865 = 12'h93c == _T_196[11:0] ? 4'h0 : _GEN_20864; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20866 = 12'h93d == _T_196[11:0] ? 4'h0 : _GEN_20865; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20867 = 12'h93e == _T_196[11:0] ? 4'h0 : _GEN_20866; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20868 = 12'h93f == _T_196[11:0] ? 4'h0 : _GEN_20867; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20869 = 12'h940 == _T_196[11:0] ? 4'h0 : _GEN_20868; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20870 = 12'h941 == _T_196[11:0] ? 4'h0 : _GEN_20869; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20871 = 12'h942 == _T_196[11:0] ? 4'h0 : _GEN_20870; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20872 = 12'h943 == _T_196[11:0] ? 4'h0 : _GEN_20871; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20873 = 12'h944 == _T_196[11:0] ? image_2372 : _GEN_20872; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20874 = 12'h945 == _T_196[11:0] ? image_2373 : _GEN_20873; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20875 = 12'h946 == _T_196[11:0] ? image_2374 : _GEN_20874; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20876 = 12'h947 == _T_196[11:0] ? image_2375 : _GEN_20875; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20877 = 12'h948 == _T_196[11:0] ? image_2376 : _GEN_20876; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20878 = 12'h949 == _T_196[11:0] ? image_2377 : _GEN_20877; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20879 = 12'h94a == _T_196[11:0] ? image_2378 : _GEN_20878; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20880 = 12'h94b == _T_196[11:0] ? image_2379 : _GEN_20879; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20881 = 12'h94c == _T_196[11:0] ? image_2380 : _GEN_20880; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20882 = 12'h94d == _T_196[11:0] ? image_2381 : _GEN_20881; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20883 = 12'h94e == _T_196[11:0] ? image_2382 : _GEN_20882; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20884 = 12'h94f == _T_196[11:0] ? image_2383 : _GEN_20883; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20885 = 12'h950 == _T_196[11:0] ? image_2384 : _GEN_20884; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20886 = 12'h951 == _T_196[11:0] ? image_2385 : _GEN_20885; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20887 = 12'h952 == _T_196[11:0] ? image_2386 : _GEN_20886; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20888 = 12'h953 == _T_196[11:0] ? image_2387 : _GEN_20887; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20889 = 12'h954 == _T_196[11:0] ? image_2388 : _GEN_20888; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20890 = 12'h955 == _T_196[11:0] ? image_2389 : _GEN_20889; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20891 = 12'h956 == _T_196[11:0] ? image_2390 : _GEN_20890; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20892 = 12'h957 == _T_196[11:0] ? image_2391 : _GEN_20891; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20893 = 12'h958 == _T_196[11:0] ? image_2392 : _GEN_20892; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20894 = 12'h959 == _T_196[11:0] ? image_2393 : _GEN_20893; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20895 = 12'h95a == _T_196[11:0] ? image_2394 : _GEN_20894; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20896 = 12'h95b == _T_196[11:0] ? image_2395 : _GEN_20895; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20897 = 12'h95c == _T_196[11:0] ? image_2396 : _GEN_20896; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20898 = 12'h95d == _T_196[11:0] ? image_2397 : _GEN_20897; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20899 = 12'h95e == _T_196[11:0] ? image_2398 : _GEN_20898; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20900 = 12'h95f == _T_196[11:0] ? image_2399 : _GEN_20899; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20901 = 12'h960 == _T_196[11:0] ? image_2400 : _GEN_20900; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20902 = 12'h961 == _T_196[11:0] ? image_2401 : _GEN_20901; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20903 = 12'h962 == _T_196[11:0] ? image_2402 : _GEN_20902; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20904 = 12'h963 == _T_196[11:0] ? image_2403 : _GEN_20903; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20905 = 12'h964 == _T_196[11:0] ? image_2404 : _GEN_20904; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20906 = 12'h965 == _T_196[11:0] ? image_2405 : _GEN_20905; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20907 = 12'h966 == _T_196[11:0] ? image_2406 : _GEN_20906; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20908 = 12'h967 == _T_196[11:0] ? image_2407 : _GEN_20907; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20909 = 12'h968 == _T_196[11:0] ? image_2408 : _GEN_20908; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20910 = 12'h969 == _T_196[11:0] ? image_2409 : _GEN_20909; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20911 = 12'h96a == _T_196[11:0] ? image_2410 : _GEN_20910; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20912 = 12'h96b == _T_196[11:0] ? image_2411 : _GEN_20911; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20913 = 12'h96c == _T_196[11:0] ? image_2412 : _GEN_20912; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20914 = 12'h96d == _T_196[11:0] ? image_2413 : _GEN_20913; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20915 = 12'h96e == _T_196[11:0] ? image_2414 : _GEN_20914; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20916 = 12'h96f == _T_196[11:0] ? image_2415 : _GEN_20915; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20917 = 12'h970 == _T_196[11:0] ? image_2416 : _GEN_20916; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20918 = 12'h971 == _T_196[11:0] ? image_2417 : _GEN_20917; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20919 = 12'h972 == _T_196[11:0] ? image_2418 : _GEN_20918; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20920 = 12'h973 == _T_196[11:0] ? image_2419 : _GEN_20919; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20921 = 12'h974 == _T_196[11:0] ? image_2420 : _GEN_20920; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20922 = 12'h975 == _T_196[11:0] ? image_2421 : _GEN_20921; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20923 = 12'h976 == _T_196[11:0] ? image_2422 : _GEN_20922; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20924 = 12'h977 == _T_196[11:0] ? image_2423 : _GEN_20923; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20925 = 12'h978 == _T_196[11:0] ? image_2424 : _GEN_20924; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20926 = 12'h979 == _T_196[11:0] ? image_2425 : _GEN_20925; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20927 = 12'h97a == _T_196[11:0] ? image_2426 : _GEN_20926; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20928 = 12'h97b == _T_196[11:0] ? 4'h0 : _GEN_20927; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20929 = 12'h97c == _T_196[11:0] ? 4'h0 : _GEN_20928; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20930 = 12'h97d == _T_196[11:0] ? 4'h0 : _GEN_20929; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20931 = 12'h97e == _T_196[11:0] ? 4'h0 : _GEN_20930; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20932 = 12'h97f == _T_196[11:0] ? 4'h0 : _GEN_20931; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20933 = 12'h980 == _T_196[11:0] ? 4'h0 : _GEN_20932; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20934 = 12'h981 == _T_196[11:0] ? 4'h0 : _GEN_20933; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20935 = 12'h982 == _T_196[11:0] ? 4'h0 : _GEN_20934; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20936 = 12'h983 == _T_196[11:0] ? 4'h0 : _GEN_20935; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20937 = 12'h984 == _T_196[11:0] ? 4'h0 : _GEN_20936; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20938 = 12'h985 == _T_196[11:0] ? image_2437 : _GEN_20937; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20939 = 12'h986 == _T_196[11:0] ? image_2438 : _GEN_20938; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20940 = 12'h987 == _T_196[11:0] ? image_2439 : _GEN_20939; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20941 = 12'h988 == _T_196[11:0] ? image_2440 : _GEN_20940; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20942 = 12'h989 == _T_196[11:0] ? image_2441 : _GEN_20941; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20943 = 12'h98a == _T_196[11:0] ? image_2442 : _GEN_20942; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20944 = 12'h98b == _T_196[11:0] ? image_2443 : _GEN_20943; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20945 = 12'h98c == _T_196[11:0] ? image_2444 : _GEN_20944; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20946 = 12'h98d == _T_196[11:0] ? image_2445 : _GEN_20945; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20947 = 12'h98e == _T_196[11:0] ? image_2446 : _GEN_20946; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20948 = 12'h98f == _T_196[11:0] ? image_2447 : _GEN_20947; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20949 = 12'h990 == _T_196[11:0] ? image_2448 : _GEN_20948; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20950 = 12'h991 == _T_196[11:0] ? image_2449 : _GEN_20949; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20951 = 12'h992 == _T_196[11:0] ? image_2450 : _GEN_20950; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20952 = 12'h993 == _T_196[11:0] ? image_2451 : _GEN_20951; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20953 = 12'h994 == _T_196[11:0] ? image_2452 : _GEN_20952; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20954 = 12'h995 == _T_196[11:0] ? image_2453 : _GEN_20953; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20955 = 12'h996 == _T_196[11:0] ? image_2454 : _GEN_20954; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20956 = 12'h997 == _T_196[11:0] ? image_2455 : _GEN_20955; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20957 = 12'h998 == _T_196[11:0] ? image_2456 : _GEN_20956; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20958 = 12'h999 == _T_196[11:0] ? image_2457 : _GEN_20957; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20959 = 12'h99a == _T_196[11:0] ? image_2458 : _GEN_20958; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20960 = 12'h99b == _T_196[11:0] ? image_2459 : _GEN_20959; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20961 = 12'h99c == _T_196[11:0] ? image_2460 : _GEN_20960; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20962 = 12'h99d == _T_196[11:0] ? image_2461 : _GEN_20961; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20963 = 12'h99e == _T_196[11:0] ? image_2462 : _GEN_20962; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20964 = 12'h99f == _T_196[11:0] ? image_2463 : _GEN_20963; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20965 = 12'h9a0 == _T_196[11:0] ? image_2464 : _GEN_20964; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20966 = 12'h9a1 == _T_196[11:0] ? image_2465 : _GEN_20965; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20967 = 12'h9a2 == _T_196[11:0] ? image_2466 : _GEN_20966; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20968 = 12'h9a3 == _T_196[11:0] ? image_2467 : _GEN_20967; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20969 = 12'h9a4 == _T_196[11:0] ? image_2468 : _GEN_20968; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20970 = 12'h9a5 == _T_196[11:0] ? image_2469 : _GEN_20969; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20971 = 12'h9a6 == _T_196[11:0] ? image_2470 : _GEN_20970; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20972 = 12'h9a7 == _T_196[11:0] ? image_2471 : _GEN_20971; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20973 = 12'h9a8 == _T_196[11:0] ? image_2472 : _GEN_20972; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20974 = 12'h9a9 == _T_196[11:0] ? image_2473 : _GEN_20973; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20975 = 12'h9aa == _T_196[11:0] ? image_2474 : _GEN_20974; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20976 = 12'h9ab == _T_196[11:0] ? image_2475 : _GEN_20975; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20977 = 12'h9ac == _T_196[11:0] ? image_2476 : _GEN_20976; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20978 = 12'h9ad == _T_196[11:0] ? image_2477 : _GEN_20977; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20979 = 12'h9ae == _T_196[11:0] ? image_2478 : _GEN_20978; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20980 = 12'h9af == _T_196[11:0] ? image_2479 : _GEN_20979; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20981 = 12'h9b0 == _T_196[11:0] ? image_2480 : _GEN_20980; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20982 = 12'h9b1 == _T_196[11:0] ? image_2481 : _GEN_20981; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20983 = 12'h9b2 == _T_196[11:0] ? image_2482 : _GEN_20982; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20984 = 12'h9b3 == _T_196[11:0] ? image_2483 : _GEN_20983; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20985 = 12'h9b4 == _T_196[11:0] ? image_2484 : _GEN_20984; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20986 = 12'h9b5 == _T_196[11:0] ? image_2485 : _GEN_20985; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20987 = 12'h9b6 == _T_196[11:0] ? image_2486 : _GEN_20986; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20988 = 12'h9b7 == _T_196[11:0] ? image_2487 : _GEN_20987; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20989 = 12'h9b8 == _T_196[11:0] ? image_2488 : _GEN_20988; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20990 = 12'h9b9 == _T_196[11:0] ? image_2489 : _GEN_20989; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20991 = 12'h9ba == _T_196[11:0] ? image_2490 : _GEN_20990; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20992 = 12'h9bb == _T_196[11:0] ? 4'h0 : _GEN_20991; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20993 = 12'h9bc == _T_196[11:0] ? 4'h0 : _GEN_20992; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20994 = 12'h9bd == _T_196[11:0] ? 4'h0 : _GEN_20993; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20995 = 12'h9be == _T_196[11:0] ? 4'h0 : _GEN_20994; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20996 = 12'h9bf == _T_196[11:0] ? 4'h0 : _GEN_20995; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20997 = 12'h9c0 == _T_196[11:0] ? 4'h0 : _GEN_20996; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20998 = 12'h9c1 == _T_196[11:0] ? 4'h0 : _GEN_20997; // @[Filter.scala 138:46]
  wire [3:0] _GEN_20999 = 12'h9c2 == _T_196[11:0] ? 4'h0 : _GEN_20998; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21000 = 12'h9c3 == _T_196[11:0] ? 4'h0 : _GEN_20999; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21001 = 12'h9c4 == _T_196[11:0] ? 4'h0 : _GEN_21000; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21002 = 12'h9c5 == _T_196[11:0] ? 4'h0 : _GEN_21001; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21003 = 12'h9c6 == _T_196[11:0] ? image_2502 : _GEN_21002; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21004 = 12'h9c7 == _T_196[11:0] ? image_2503 : _GEN_21003; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21005 = 12'h9c8 == _T_196[11:0] ? image_2504 : _GEN_21004; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21006 = 12'h9c9 == _T_196[11:0] ? image_2505 : _GEN_21005; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21007 = 12'h9ca == _T_196[11:0] ? image_2506 : _GEN_21006; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21008 = 12'h9cb == _T_196[11:0] ? image_2507 : _GEN_21007; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21009 = 12'h9cc == _T_196[11:0] ? image_2508 : _GEN_21008; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21010 = 12'h9cd == _T_196[11:0] ? image_2509 : _GEN_21009; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21011 = 12'h9ce == _T_196[11:0] ? image_2510 : _GEN_21010; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21012 = 12'h9cf == _T_196[11:0] ? image_2511 : _GEN_21011; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21013 = 12'h9d0 == _T_196[11:0] ? image_2512 : _GEN_21012; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21014 = 12'h9d1 == _T_196[11:0] ? image_2513 : _GEN_21013; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21015 = 12'h9d2 == _T_196[11:0] ? image_2514 : _GEN_21014; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21016 = 12'h9d3 == _T_196[11:0] ? image_2515 : _GEN_21015; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21017 = 12'h9d4 == _T_196[11:0] ? image_2516 : _GEN_21016; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21018 = 12'h9d5 == _T_196[11:0] ? image_2517 : _GEN_21017; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21019 = 12'h9d6 == _T_196[11:0] ? image_2518 : _GEN_21018; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21020 = 12'h9d7 == _T_196[11:0] ? image_2519 : _GEN_21019; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21021 = 12'h9d8 == _T_196[11:0] ? image_2520 : _GEN_21020; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21022 = 12'h9d9 == _T_196[11:0] ? image_2521 : _GEN_21021; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21023 = 12'h9da == _T_196[11:0] ? image_2522 : _GEN_21022; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21024 = 12'h9db == _T_196[11:0] ? image_2523 : _GEN_21023; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21025 = 12'h9dc == _T_196[11:0] ? image_2524 : _GEN_21024; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21026 = 12'h9dd == _T_196[11:0] ? image_2525 : _GEN_21025; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21027 = 12'h9de == _T_196[11:0] ? image_2526 : _GEN_21026; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21028 = 12'h9df == _T_196[11:0] ? image_2527 : _GEN_21027; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21029 = 12'h9e0 == _T_196[11:0] ? image_2528 : _GEN_21028; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21030 = 12'h9e1 == _T_196[11:0] ? image_2529 : _GEN_21029; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21031 = 12'h9e2 == _T_196[11:0] ? image_2530 : _GEN_21030; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21032 = 12'h9e3 == _T_196[11:0] ? image_2531 : _GEN_21031; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21033 = 12'h9e4 == _T_196[11:0] ? image_2532 : _GEN_21032; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21034 = 12'h9e5 == _T_196[11:0] ? image_2533 : _GEN_21033; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21035 = 12'h9e6 == _T_196[11:0] ? image_2534 : _GEN_21034; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21036 = 12'h9e7 == _T_196[11:0] ? image_2535 : _GEN_21035; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21037 = 12'h9e8 == _T_196[11:0] ? image_2536 : _GEN_21036; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21038 = 12'h9e9 == _T_196[11:0] ? image_2537 : _GEN_21037; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21039 = 12'h9ea == _T_196[11:0] ? image_2538 : _GEN_21038; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21040 = 12'h9eb == _T_196[11:0] ? image_2539 : _GEN_21039; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21041 = 12'h9ec == _T_196[11:0] ? image_2540 : _GEN_21040; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21042 = 12'h9ed == _T_196[11:0] ? image_2541 : _GEN_21041; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21043 = 12'h9ee == _T_196[11:0] ? image_2542 : _GEN_21042; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21044 = 12'h9ef == _T_196[11:0] ? image_2543 : _GEN_21043; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21045 = 12'h9f0 == _T_196[11:0] ? image_2544 : _GEN_21044; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21046 = 12'h9f1 == _T_196[11:0] ? image_2545 : _GEN_21045; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21047 = 12'h9f2 == _T_196[11:0] ? image_2546 : _GEN_21046; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21048 = 12'h9f3 == _T_196[11:0] ? image_2547 : _GEN_21047; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21049 = 12'h9f4 == _T_196[11:0] ? image_2548 : _GEN_21048; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21050 = 12'h9f5 == _T_196[11:0] ? image_2549 : _GEN_21049; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21051 = 12'h9f6 == _T_196[11:0] ? image_2550 : _GEN_21050; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21052 = 12'h9f7 == _T_196[11:0] ? image_2551 : _GEN_21051; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21053 = 12'h9f8 == _T_196[11:0] ? image_2552 : _GEN_21052; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21054 = 12'h9f9 == _T_196[11:0] ? image_2553 : _GEN_21053; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21055 = 12'h9fa == _T_196[11:0] ? image_2554 : _GEN_21054; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21056 = 12'h9fb == _T_196[11:0] ? 4'h0 : _GEN_21055; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21057 = 12'h9fc == _T_196[11:0] ? 4'h0 : _GEN_21056; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21058 = 12'h9fd == _T_196[11:0] ? 4'h0 : _GEN_21057; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21059 = 12'h9fe == _T_196[11:0] ? 4'h0 : _GEN_21058; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21060 = 12'h9ff == _T_196[11:0] ? 4'h0 : _GEN_21059; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21061 = 12'ha00 == _T_196[11:0] ? 4'h0 : _GEN_21060; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21062 = 12'ha01 == _T_196[11:0] ? 4'h0 : _GEN_21061; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21063 = 12'ha02 == _T_196[11:0] ? 4'h0 : _GEN_21062; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21064 = 12'ha03 == _T_196[11:0] ? 4'h0 : _GEN_21063; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21065 = 12'ha04 == _T_196[11:0] ? 4'h0 : _GEN_21064; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21066 = 12'ha05 == _T_196[11:0] ? 4'h0 : _GEN_21065; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21067 = 12'ha06 == _T_196[11:0] ? 4'h0 : _GEN_21066; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21068 = 12'ha07 == _T_196[11:0] ? image_2567 : _GEN_21067; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21069 = 12'ha08 == _T_196[11:0] ? image_2568 : _GEN_21068; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21070 = 12'ha09 == _T_196[11:0] ? image_2569 : _GEN_21069; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21071 = 12'ha0a == _T_196[11:0] ? image_2570 : _GEN_21070; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21072 = 12'ha0b == _T_196[11:0] ? image_2571 : _GEN_21071; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21073 = 12'ha0c == _T_196[11:0] ? image_2572 : _GEN_21072; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21074 = 12'ha0d == _T_196[11:0] ? image_2573 : _GEN_21073; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21075 = 12'ha0e == _T_196[11:0] ? image_2574 : _GEN_21074; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21076 = 12'ha0f == _T_196[11:0] ? image_2575 : _GEN_21075; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21077 = 12'ha10 == _T_196[11:0] ? image_2576 : _GEN_21076; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21078 = 12'ha11 == _T_196[11:0] ? image_2577 : _GEN_21077; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21079 = 12'ha12 == _T_196[11:0] ? image_2578 : _GEN_21078; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21080 = 12'ha13 == _T_196[11:0] ? image_2579 : _GEN_21079; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21081 = 12'ha14 == _T_196[11:0] ? image_2580 : _GEN_21080; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21082 = 12'ha15 == _T_196[11:0] ? image_2581 : _GEN_21081; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21083 = 12'ha16 == _T_196[11:0] ? image_2582 : _GEN_21082; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21084 = 12'ha17 == _T_196[11:0] ? image_2583 : _GEN_21083; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21085 = 12'ha18 == _T_196[11:0] ? image_2584 : _GEN_21084; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21086 = 12'ha19 == _T_196[11:0] ? image_2585 : _GEN_21085; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21087 = 12'ha1a == _T_196[11:0] ? image_2586 : _GEN_21086; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21088 = 12'ha1b == _T_196[11:0] ? image_2587 : _GEN_21087; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21089 = 12'ha1c == _T_196[11:0] ? image_2588 : _GEN_21088; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21090 = 12'ha1d == _T_196[11:0] ? image_2589 : _GEN_21089; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21091 = 12'ha1e == _T_196[11:0] ? image_2590 : _GEN_21090; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21092 = 12'ha1f == _T_196[11:0] ? image_2591 : _GEN_21091; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21093 = 12'ha20 == _T_196[11:0] ? image_2592 : _GEN_21092; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21094 = 12'ha21 == _T_196[11:0] ? image_2593 : _GEN_21093; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21095 = 12'ha22 == _T_196[11:0] ? image_2594 : _GEN_21094; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21096 = 12'ha23 == _T_196[11:0] ? image_2595 : _GEN_21095; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21097 = 12'ha24 == _T_196[11:0] ? image_2596 : _GEN_21096; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21098 = 12'ha25 == _T_196[11:0] ? image_2597 : _GEN_21097; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21099 = 12'ha26 == _T_196[11:0] ? image_2598 : _GEN_21098; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21100 = 12'ha27 == _T_196[11:0] ? image_2599 : _GEN_21099; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21101 = 12'ha28 == _T_196[11:0] ? image_2600 : _GEN_21100; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21102 = 12'ha29 == _T_196[11:0] ? image_2601 : _GEN_21101; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21103 = 12'ha2a == _T_196[11:0] ? image_2602 : _GEN_21102; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21104 = 12'ha2b == _T_196[11:0] ? image_2603 : _GEN_21103; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21105 = 12'ha2c == _T_196[11:0] ? image_2604 : _GEN_21104; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21106 = 12'ha2d == _T_196[11:0] ? image_2605 : _GEN_21105; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21107 = 12'ha2e == _T_196[11:0] ? image_2606 : _GEN_21106; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21108 = 12'ha2f == _T_196[11:0] ? image_2607 : _GEN_21107; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21109 = 12'ha30 == _T_196[11:0] ? image_2608 : _GEN_21108; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21110 = 12'ha31 == _T_196[11:0] ? image_2609 : _GEN_21109; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21111 = 12'ha32 == _T_196[11:0] ? image_2610 : _GEN_21110; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21112 = 12'ha33 == _T_196[11:0] ? image_2611 : _GEN_21111; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21113 = 12'ha34 == _T_196[11:0] ? image_2612 : _GEN_21112; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21114 = 12'ha35 == _T_196[11:0] ? image_2613 : _GEN_21113; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21115 = 12'ha36 == _T_196[11:0] ? image_2614 : _GEN_21114; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21116 = 12'ha37 == _T_196[11:0] ? image_2615 : _GEN_21115; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21117 = 12'ha38 == _T_196[11:0] ? image_2616 : _GEN_21116; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21118 = 12'ha39 == _T_196[11:0] ? image_2617 : _GEN_21117; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21119 = 12'ha3a == _T_196[11:0] ? image_2618 : _GEN_21118; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21120 = 12'ha3b == _T_196[11:0] ? 4'h0 : _GEN_21119; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21121 = 12'ha3c == _T_196[11:0] ? 4'h0 : _GEN_21120; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21122 = 12'ha3d == _T_196[11:0] ? 4'h0 : _GEN_21121; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21123 = 12'ha3e == _T_196[11:0] ? 4'h0 : _GEN_21122; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21124 = 12'ha3f == _T_196[11:0] ? 4'h0 : _GEN_21123; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21125 = 12'ha40 == _T_196[11:0] ? 4'h0 : _GEN_21124; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21126 = 12'ha41 == _T_196[11:0] ? 4'h0 : _GEN_21125; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21127 = 12'ha42 == _T_196[11:0] ? 4'h0 : _GEN_21126; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21128 = 12'ha43 == _T_196[11:0] ? 4'h0 : _GEN_21127; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21129 = 12'ha44 == _T_196[11:0] ? 4'h0 : _GEN_21128; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21130 = 12'ha45 == _T_196[11:0] ? 4'h0 : _GEN_21129; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21131 = 12'ha46 == _T_196[11:0] ? 4'h0 : _GEN_21130; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21132 = 12'ha47 == _T_196[11:0] ? 4'h0 : _GEN_21131; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21133 = 12'ha48 == _T_196[11:0] ? image_2632 : _GEN_21132; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21134 = 12'ha49 == _T_196[11:0] ? image_2633 : _GEN_21133; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21135 = 12'ha4a == _T_196[11:0] ? image_2634 : _GEN_21134; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21136 = 12'ha4b == _T_196[11:0] ? image_2635 : _GEN_21135; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21137 = 12'ha4c == _T_196[11:0] ? image_2636 : _GEN_21136; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21138 = 12'ha4d == _T_196[11:0] ? image_2637 : _GEN_21137; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21139 = 12'ha4e == _T_196[11:0] ? image_2638 : _GEN_21138; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21140 = 12'ha4f == _T_196[11:0] ? image_2639 : _GEN_21139; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21141 = 12'ha50 == _T_196[11:0] ? image_2640 : _GEN_21140; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21142 = 12'ha51 == _T_196[11:0] ? image_2641 : _GEN_21141; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21143 = 12'ha52 == _T_196[11:0] ? image_2642 : _GEN_21142; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21144 = 12'ha53 == _T_196[11:0] ? image_2643 : _GEN_21143; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21145 = 12'ha54 == _T_196[11:0] ? image_2644 : _GEN_21144; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21146 = 12'ha55 == _T_196[11:0] ? image_2645 : _GEN_21145; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21147 = 12'ha56 == _T_196[11:0] ? image_2646 : _GEN_21146; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21148 = 12'ha57 == _T_196[11:0] ? image_2647 : _GEN_21147; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21149 = 12'ha58 == _T_196[11:0] ? image_2648 : _GEN_21148; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21150 = 12'ha59 == _T_196[11:0] ? image_2649 : _GEN_21149; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21151 = 12'ha5a == _T_196[11:0] ? image_2650 : _GEN_21150; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21152 = 12'ha5b == _T_196[11:0] ? image_2651 : _GEN_21151; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21153 = 12'ha5c == _T_196[11:0] ? image_2652 : _GEN_21152; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21154 = 12'ha5d == _T_196[11:0] ? image_2653 : _GEN_21153; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21155 = 12'ha5e == _T_196[11:0] ? image_2654 : _GEN_21154; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21156 = 12'ha5f == _T_196[11:0] ? image_2655 : _GEN_21155; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21157 = 12'ha60 == _T_196[11:0] ? image_2656 : _GEN_21156; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21158 = 12'ha61 == _T_196[11:0] ? image_2657 : _GEN_21157; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21159 = 12'ha62 == _T_196[11:0] ? image_2658 : _GEN_21158; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21160 = 12'ha63 == _T_196[11:0] ? image_2659 : _GEN_21159; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21161 = 12'ha64 == _T_196[11:0] ? image_2660 : _GEN_21160; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21162 = 12'ha65 == _T_196[11:0] ? image_2661 : _GEN_21161; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21163 = 12'ha66 == _T_196[11:0] ? image_2662 : _GEN_21162; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21164 = 12'ha67 == _T_196[11:0] ? image_2663 : _GEN_21163; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21165 = 12'ha68 == _T_196[11:0] ? image_2664 : _GEN_21164; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21166 = 12'ha69 == _T_196[11:0] ? image_2665 : _GEN_21165; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21167 = 12'ha6a == _T_196[11:0] ? image_2666 : _GEN_21166; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21168 = 12'ha6b == _T_196[11:0] ? image_2667 : _GEN_21167; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21169 = 12'ha6c == _T_196[11:0] ? image_2668 : _GEN_21168; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21170 = 12'ha6d == _T_196[11:0] ? image_2669 : _GEN_21169; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21171 = 12'ha6e == _T_196[11:0] ? image_2670 : _GEN_21170; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21172 = 12'ha6f == _T_196[11:0] ? image_2671 : _GEN_21171; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21173 = 12'ha70 == _T_196[11:0] ? image_2672 : _GEN_21172; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21174 = 12'ha71 == _T_196[11:0] ? image_2673 : _GEN_21173; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21175 = 12'ha72 == _T_196[11:0] ? image_2674 : _GEN_21174; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21176 = 12'ha73 == _T_196[11:0] ? image_2675 : _GEN_21175; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21177 = 12'ha74 == _T_196[11:0] ? image_2676 : _GEN_21176; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21178 = 12'ha75 == _T_196[11:0] ? image_2677 : _GEN_21177; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21179 = 12'ha76 == _T_196[11:0] ? image_2678 : _GEN_21178; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21180 = 12'ha77 == _T_196[11:0] ? image_2679 : _GEN_21179; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21181 = 12'ha78 == _T_196[11:0] ? image_2680 : _GEN_21180; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21182 = 12'ha79 == _T_196[11:0] ? image_2681 : _GEN_21181; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21183 = 12'ha7a == _T_196[11:0] ? image_2682 : _GEN_21182; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21184 = 12'ha7b == _T_196[11:0] ? 4'h0 : _GEN_21183; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21185 = 12'ha7c == _T_196[11:0] ? 4'h0 : _GEN_21184; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21186 = 12'ha7d == _T_196[11:0] ? 4'h0 : _GEN_21185; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21187 = 12'ha7e == _T_196[11:0] ? 4'h0 : _GEN_21186; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21188 = 12'ha7f == _T_196[11:0] ? 4'h0 : _GEN_21187; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21189 = 12'ha80 == _T_196[11:0] ? 4'h0 : _GEN_21188; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21190 = 12'ha81 == _T_196[11:0] ? 4'h0 : _GEN_21189; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21191 = 12'ha82 == _T_196[11:0] ? 4'h0 : _GEN_21190; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21192 = 12'ha83 == _T_196[11:0] ? 4'h0 : _GEN_21191; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21193 = 12'ha84 == _T_196[11:0] ? 4'h0 : _GEN_21192; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21194 = 12'ha85 == _T_196[11:0] ? 4'h0 : _GEN_21193; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21195 = 12'ha86 == _T_196[11:0] ? 4'h0 : _GEN_21194; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21196 = 12'ha87 == _T_196[11:0] ? 4'h0 : _GEN_21195; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21197 = 12'ha88 == _T_196[11:0] ? 4'h0 : _GEN_21196; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21198 = 12'ha89 == _T_196[11:0] ? image_2697 : _GEN_21197; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21199 = 12'ha8a == _T_196[11:0] ? image_2698 : _GEN_21198; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21200 = 12'ha8b == _T_196[11:0] ? image_2699 : _GEN_21199; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21201 = 12'ha8c == _T_196[11:0] ? image_2700 : _GEN_21200; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21202 = 12'ha8d == _T_196[11:0] ? image_2701 : _GEN_21201; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21203 = 12'ha8e == _T_196[11:0] ? image_2702 : _GEN_21202; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21204 = 12'ha8f == _T_196[11:0] ? image_2703 : _GEN_21203; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21205 = 12'ha90 == _T_196[11:0] ? image_2704 : _GEN_21204; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21206 = 12'ha91 == _T_196[11:0] ? image_2705 : _GEN_21205; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21207 = 12'ha92 == _T_196[11:0] ? image_2706 : _GEN_21206; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21208 = 12'ha93 == _T_196[11:0] ? image_2707 : _GEN_21207; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21209 = 12'ha94 == _T_196[11:0] ? image_2708 : _GEN_21208; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21210 = 12'ha95 == _T_196[11:0] ? image_2709 : _GEN_21209; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21211 = 12'ha96 == _T_196[11:0] ? image_2710 : _GEN_21210; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21212 = 12'ha97 == _T_196[11:0] ? image_2711 : _GEN_21211; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21213 = 12'ha98 == _T_196[11:0] ? image_2712 : _GEN_21212; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21214 = 12'ha99 == _T_196[11:0] ? image_2713 : _GEN_21213; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21215 = 12'ha9a == _T_196[11:0] ? image_2714 : _GEN_21214; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21216 = 12'ha9b == _T_196[11:0] ? image_2715 : _GEN_21215; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21217 = 12'ha9c == _T_196[11:0] ? image_2716 : _GEN_21216; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21218 = 12'ha9d == _T_196[11:0] ? image_2717 : _GEN_21217; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21219 = 12'ha9e == _T_196[11:0] ? image_2718 : _GEN_21218; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21220 = 12'ha9f == _T_196[11:0] ? image_2719 : _GEN_21219; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21221 = 12'haa0 == _T_196[11:0] ? image_2720 : _GEN_21220; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21222 = 12'haa1 == _T_196[11:0] ? image_2721 : _GEN_21221; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21223 = 12'haa2 == _T_196[11:0] ? image_2722 : _GEN_21222; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21224 = 12'haa3 == _T_196[11:0] ? image_2723 : _GEN_21223; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21225 = 12'haa4 == _T_196[11:0] ? image_2724 : _GEN_21224; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21226 = 12'haa5 == _T_196[11:0] ? image_2725 : _GEN_21225; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21227 = 12'haa6 == _T_196[11:0] ? image_2726 : _GEN_21226; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21228 = 12'haa7 == _T_196[11:0] ? image_2727 : _GEN_21227; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21229 = 12'haa8 == _T_196[11:0] ? image_2728 : _GEN_21228; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21230 = 12'haa9 == _T_196[11:0] ? image_2729 : _GEN_21229; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21231 = 12'haaa == _T_196[11:0] ? image_2730 : _GEN_21230; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21232 = 12'haab == _T_196[11:0] ? image_2731 : _GEN_21231; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21233 = 12'haac == _T_196[11:0] ? image_2732 : _GEN_21232; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21234 = 12'haad == _T_196[11:0] ? image_2733 : _GEN_21233; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21235 = 12'haae == _T_196[11:0] ? image_2734 : _GEN_21234; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21236 = 12'haaf == _T_196[11:0] ? image_2735 : _GEN_21235; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21237 = 12'hab0 == _T_196[11:0] ? image_2736 : _GEN_21236; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21238 = 12'hab1 == _T_196[11:0] ? image_2737 : _GEN_21237; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21239 = 12'hab2 == _T_196[11:0] ? image_2738 : _GEN_21238; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21240 = 12'hab3 == _T_196[11:0] ? image_2739 : _GEN_21239; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21241 = 12'hab4 == _T_196[11:0] ? image_2740 : _GEN_21240; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21242 = 12'hab5 == _T_196[11:0] ? image_2741 : _GEN_21241; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21243 = 12'hab6 == _T_196[11:0] ? image_2742 : _GEN_21242; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21244 = 12'hab7 == _T_196[11:0] ? image_2743 : _GEN_21243; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21245 = 12'hab8 == _T_196[11:0] ? image_2744 : _GEN_21244; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21246 = 12'hab9 == _T_196[11:0] ? image_2745 : _GEN_21245; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21247 = 12'haba == _T_196[11:0] ? 4'h0 : _GEN_21246; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21248 = 12'habb == _T_196[11:0] ? 4'h0 : _GEN_21247; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21249 = 12'habc == _T_196[11:0] ? 4'h0 : _GEN_21248; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21250 = 12'habd == _T_196[11:0] ? 4'h0 : _GEN_21249; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21251 = 12'habe == _T_196[11:0] ? 4'h0 : _GEN_21250; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21252 = 12'habf == _T_196[11:0] ? 4'h0 : _GEN_21251; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21253 = 12'hac0 == _T_196[11:0] ? 4'h0 : _GEN_21252; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21254 = 12'hac1 == _T_196[11:0] ? 4'h0 : _GEN_21253; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21255 = 12'hac2 == _T_196[11:0] ? 4'h0 : _GEN_21254; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21256 = 12'hac3 == _T_196[11:0] ? 4'h0 : _GEN_21255; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21257 = 12'hac4 == _T_196[11:0] ? 4'h0 : _GEN_21256; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21258 = 12'hac5 == _T_196[11:0] ? 4'h0 : _GEN_21257; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21259 = 12'hac6 == _T_196[11:0] ? 4'h0 : _GEN_21258; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21260 = 12'hac7 == _T_196[11:0] ? 4'h0 : _GEN_21259; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21261 = 12'hac8 == _T_196[11:0] ? 4'h0 : _GEN_21260; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21262 = 12'hac9 == _T_196[11:0] ? 4'h0 : _GEN_21261; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21263 = 12'haca == _T_196[11:0] ? 4'h0 : _GEN_21262; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21264 = 12'hacb == _T_196[11:0] ? image_2763 : _GEN_21263; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21265 = 12'hacc == _T_196[11:0] ? image_2764 : _GEN_21264; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21266 = 12'hacd == _T_196[11:0] ? image_2765 : _GEN_21265; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21267 = 12'hace == _T_196[11:0] ? image_2766 : _GEN_21266; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21268 = 12'hacf == _T_196[11:0] ? image_2767 : _GEN_21267; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21269 = 12'had0 == _T_196[11:0] ? image_2768 : _GEN_21268; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21270 = 12'had1 == _T_196[11:0] ? image_2769 : _GEN_21269; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21271 = 12'had2 == _T_196[11:0] ? image_2770 : _GEN_21270; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21272 = 12'had3 == _T_196[11:0] ? image_2771 : _GEN_21271; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21273 = 12'had4 == _T_196[11:0] ? image_2772 : _GEN_21272; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21274 = 12'had5 == _T_196[11:0] ? image_2773 : _GEN_21273; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21275 = 12'had6 == _T_196[11:0] ? image_2774 : _GEN_21274; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21276 = 12'had7 == _T_196[11:0] ? image_2775 : _GEN_21275; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21277 = 12'had8 == _T_196[11:0] ? image_2776 : _GEN_21276; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21278 = 12'had9 == _T_196[11:0] ? image_2777 : _GEN_21277; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21279 = 12'hada == _T_196[11:0] ? image_2778 : _GEN_21278; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21280 = 12'hadb == _T_196[11:0] ? image_2779 : _GEN_21279; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21281 = 12'hadc == _T_196[11:0] ? image_2780 : _GEN_21280; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21282 = 12'hadd == _T_196[11:0] ? image_2781 : _GEN_21281; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21283 = 12'hade == _T_196[11:0] ? image_2782 : _GEN_21282; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21284 = 12'hadf == _T_196[11:0] ? image_2783 : _GEN_21283; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21285 = 12'hae0 == _T_196[11:0] ? image_2784 : _GEN_21284; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21286 = 12'hae1 == _T_196[11:0] ? image_2785 : _GEN_21285; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21287 = 12'hae2 == _T_196[11:0] ? image_2786 : _GEN_21286; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21288 = 12'hae3 == _T_196[11:0] ? image_2787 : _GEN_21287; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21289 = 12'hae4 == _T_196[11:0] ? image_2788 : _GEN_21288; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21290 = 12'hae5 == _T_196[11:0] ? image_2789 : _GEN_21289; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21291 = 12'hae6 == _T_196[11:0] ? image_2790 : _GEN_21290; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21292 = 12'hae7 == _T_196[11:0] ? image_2791 : _GEN_21291; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21293 = 12'hae8 == _T_196[11:0] ? image_2792 : _GEN_21292; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21294 = 12'hae9 == _T_196[11:0] ? image_2793 : _GEN_21293; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21295 = 12'haea == _T_196[11:0] ? image_2794 : _GEN_21294; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21296 = 12'haeb == _T_196[11:0] ? image_2795 : _GEN_21295; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21297 = 12'haec == _T_196[11:0] ? image_2796 : _GEN_21296; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21298 = 12'haed == _T_196[11:0] ? image_2797 : _GEN_21297; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21299 = 12'haee == _T_196[11:0] ? image_2798 : _GEN_21298; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21300 = 12'haef == _T_196[11:0] ? image_2799 : _GEN_21299; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21301 = 12'haf0 == _T_196[11:0] ? image_2800 : _GEN_21300; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21302 = 12'haf1 == _T_196[11:0] ? image_2801 : _GEN_21301; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21303 = 12'haf2 == _T_196[11:0] ? image_2802 : _GEN_21302; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21304 = 12'haf3 == _T_196[11:0] ? image_2803 : _GEN_21303; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21305 = 12'haf4 == _T_196[11:0] ? image_2804 : _GEN_21304; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21306 = 12'haf5 == _T_196[11:0] ? image_2805 : _GEN_21305; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21307 = 12'haf6 == _T_196[11:0] ? image_2806 : _GEN_21306; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21308 = 12'haf7 == _T_196[11:0] ? image_2807 : _GEN_21307; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21309 = 12'haf8 == _T_196[11:0] ? image_2808 : _GEN_21308; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21310 = 12'haf9 == _T_196[11:0] ? 4'h0 : _GEN_21309; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21311 = 12'hafa == _T_196[11:0] ? 4'h0 : _GEN_21310; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21312 = 12'hafb == _T_196[11:0] ? 4'h0 : _GEN_21311; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21313 = 12'hafc == _T_196[11:0] ? 4'h0 : _GEN_21312; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21314 = 12'hafd == _T_196[11:0] ? 4'h0 : _GEN_21313; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21315 = 12'hafe == _T_196[11:0] ? 4'h0 : _GEN_21314; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21316 = 12'haff == _T_196[11:0] ? 4'h0 : _GEN_21315; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21317 = 12'hb00 == _T_196[11:0] ? 4'h0 : _GEN_21316; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21318 = 12'hb01 == _T_196[11:0] ? 4'h0 : _GEN_21317; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21319 = 12'hb02 == _T_196[11:0] ? 4'h0 : _GEN_21318; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21320 = 12'hb03 == _T_196[11:0] ? 4'h0 : _GEN_21319; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21321 = 12'hb04 == _T_196[11:0] ? 4'h0 : _GEN_21320; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21322 = 12'hb05 == _T_196[11:0] ? 4'h0 : _GEN_21321; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21323 = 12'hb06 == _T_196[11:0] ? 4'h0 : _GEN_21322; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21324 = 12'hb07 == _T_196[11:0] ? 4'h0 : _GEN_21323; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21325 = 12'hb08 == _T_196[11:0] ? 4'h0 : _GEN_21324; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21326 = 12'hb09 == _T_196[11:0] ? 4'h0 : _GEN_21325; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21327 = 12'hb0a == _T_196[11:0] ? 4'h0 : _GEN_21326; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21328 = 12'hb0b == _T_196[11:0] ? 4'h0 : _GEN_21327; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21329 = 12'hb0c == _T_196[11:0] ? image_2828 : _GEN_21328; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21330 = 12'hb0d == _T_196[11:0] ? image_2829 : _GEN_21329; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21331 = 12'hb0e == _T_196[11:0] ? image_2830 : _GEN_21330; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21332 = 12'hb0f == _T_196[11:0] ? image_2831 : _GEN_21331; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21333 = 12'hb10 == _T_196[11:0] ? image_2832 : _GEN_21332; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21334 = 12'hb11 == _T_196[11:0] ? image_2833 : _GEN_21333; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21335 = 12'hb12 == _T_196[11:0] ? image_2834 : _GEN_21334; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21336 = 12'hb13 == _T_196[11:0] ? image_2835 : _GEN_21335; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21337 = 12'hb14 == _T_196[11:0] ? image_2836 : _GEN_21336; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21338 = 12'hb15 == _T_196[11:0] ? image_2837 : _GEN_21337; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21339 = 12'hb16 == _T_196[11:0] ? image_2838 : _GEN_21338; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21340 = 12'hb17 == _T_196[11:0] ? image_2839 : _GEN_21339; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21341 = 12'hb18 == _T_196[11:0] ? image_2840 : _GEN_21340; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21342 = 12'hb19 == _T_196[11:0] ? image_2841 : _GEN_21341; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21343 = 12'hb1a == _T_196[11:0] ? image_2842 : _GEN_21342; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21344 = 12'hb1b == _T_196[11:0] ? image_2843 : _GEN_21343; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21345 = 12'hb1c == _T_196[11:0] ? image_2844 : _GEN_21344; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21346 = 12'hb1d == _T_196[11:0] ? image_2845 : _GEN_21345; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21347 = 12'hb1e == _T_196[11:0] ? image_2846 : _GEN_21346; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21348 = 12'hb1f == _T_196[11:0] ? image_2847 : _GEN_21347; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21349 = 12'hb20 == _T_196[11:0] ? image_2848 : _GEN_21348; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21350 = 12'hb21 == _T_196[11:0] ? image_2849 : _GEN_21349; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21351 = 12'hb22 == _T_196[11:0] ? image_2850 : _GEN_21350; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21352 = 12'hb23 == _T_196[11:0] ? image_2851 : _GEN_21351; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21353 = 12'hb24 == _T_196[11:0] ? image_2852 : _GEN_21352; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21354 = 12'hb25 == _T_196[11:0] ? image_2853 : _GEN_21353; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21355 = 12'hb26 == _T_196[11:0] ? image_2854 : _GEN_21354; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21356 = 12'hb27 == _T_196[11:0] ? image_2855 : _GEN_21355; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21357 = 12'hb28 == _T_196[11:0] ? image_2856 : _GEN_21356; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21358 = 12'hb29 == _T_196[11:0] ? image_2857 : _GEN_21357; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21359 = 12'hb2a == _T_196[11:0] ? image_2858 : _GEN_21358; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21360 = 12'hb2b == _T_196[11:0] ? image_2859 : _GEN_21359; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21361 = 12'hb2c == _T_196[11:0] ? image_2860 : _GEN_21360; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21362 = 12'hb2d == _T_196[11:0] ? image_2861 : _GEN_21361; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21363 = 12'hb2e == _T_196[11:0] ? image_2862 : _GEN_21362; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21364 = 12'hb2f == _T_196[11:0] ? image_2863 : _GEN_21363; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21365 = 12'hb30 == _T_196[11:0] ? image_2864 : _GEN_21364; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21366 = 12'hb31 == _T_196[11:0] ? image_2865 : _GEN_21365; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21367 = 12'hb32 == _T_196[11:0] ? image_2866 : _GEN_21366; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21368 = 12'hb33 == _T_196[11:0] ? image_2867 : _GEN_21367; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21369 = 12'hb34 == _T_196[11:0] ? image_2868 : _GEN_21368; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21370 = 12'hb35 == _T_196[11:0] ? image_2869 : _GEN_21369; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21371 = 12'hb36 == _T_196[11:0] ? image_2870 : _GEN_21370; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21372 = 12'hb37 == _T_196[11:0] ? image_2871 : _GEN_21371; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21373 = 12'hb38 == _T_196[11:0] ? 4'h0 : _GEN_21372; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21374 = 12'hb39 == _T_196[11:0] ? 4'h0 : _GEN_21373; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21375 = 12'hb3a == _T_196[11:0] ? 4'h0 : _GEN_21374; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21376 = 12'hb3b == _T_196[11:0] ? 4'h0 : _GEN_21375; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21377 = 12'hb3c == _T_196[11:0] ? 4'h0 : _GEN_21376; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21378 = 12'hb3d == _T_196[11:0] ? 4'h0 : _GEN_21377; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21379 = 12'hb3e == _T_196[11:0] ? 4'h0 : _GEN_21378; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21380 = 12'hb3f == _T_196[11:0] ? 4'h0 : _GEN_21379; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21381 = 12'hb40 == _T_196[11:0] ? 4'h0 : _GEN_21380; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21382 = 12'hb41 == _T_196[11:0] ? 4'h0 : _GEN_21381; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21383 = 12'hb42 == _T_196[11:0] ? 4'h0 : _GEN_21382; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21384 = 12'hb43 == _T_196[11:0] ? 4'h0 : _GEN_21383; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21385 = 12'hb44 == _T_196[11:0] ? 4'h0 : _GEN_21384; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21386 = 12'hb45 == _T_196[11:0] ? 4'h0 : _GEN_21385; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21387 = 12'hb46 == _T_196[11:0] ? 4'h0 : _GEN_21386; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21388 = 12'hb47 == _T_196[11:0] ? 4'h0 : _GEN_21387; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21389 = 12'hb48 == _T_196[11:0] ? 4'h0 : _GEN_21388; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21390 = 12'hb49 == _T_196[11:0] ? 4'h0 : _GEN_21389; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21391 = 12'hb4a == _T_196[11:0] ? 4'h0 : _GEN_21390; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21392 = 12'hb4b == _T_196[11:0] ? 4'h0 : _GEN_21391; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21393 = 12'hb4c == _T_196[11:0] ? 4'h0 : _GEN_21392; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21394 = 12'hb4d == _T_196[11:0] ? 4'h0 : _GEN_21393; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21395 = 12'hb4e == _T_196[11:0] ? 4'h0 : _GEN_21394; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21396 = 12'hb4f == _T_196[11:0] ? image_2895 : _GEN_21395; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21397 = 12'hb50 == _T_196[11:0] ? image_2896 : _GEN_21396; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21398 = 12'hb51 == _T_196[11:0] ? image_2897 : _GEN_21397; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21399 = 12'hb52 == _T_196[11:0] ? image_2898 : _GEN_21398; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21400 = 12'hb53 == _T_196[11:0] ? image_2899 : _GEN_21399; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21401 = 12'hb54 == _T_196[11:0] ? image_2900 : _GEN_21400; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21402 = 12'hb55 == _T_196[11:0] ? image_2901 : _GEN_21401; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21403 = 12'hb56 == _T_196[11:0] ? image_2902 : _GEN_21402; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21404 = 12'hb57 == _T_196[11:0] ? image_2903 : _GEN_21403; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21405 = 12'hb58 == _T_196[11:0] ? image_2904 : _GEN_21404; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21406 = 12'hb59 == _T_196[11:0] ? image_2905 : _GEN_21405; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21407 = 12'hb5a == _T_196[11:0] ? image_2906 : _GEN_21406; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21408 = 12'hb5b == _T_196[11:0] ? image_2907 : _GEN_21407; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21409 = 12'hb5c == _T_196[11:0] ? image_2908 : _GEN_21408; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21410 = 12'hb5d == _T_196[11:0] ? image_2909 : _GEN_21409; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21411 = 12'hb5e == _T_196[11:0] ? image_2910 : _GEN_21410; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21412 = 12'hb5f == _T_196[11:0] ? image_2911 : _GEN_21411; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21413 = 12'hb60 == _T_196[11:0] ? image_2912 : _GEN_21412; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21414 = 12'hb61 == _T_196[11:0] ? image_2913 : _GEN_21413; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21415 = 12'hb62 == _T_196[11:0] ? image_2914 : _GEN_21414; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21416 = 12'hb63 == _T_196[11:0] ? image_2915 : _GEN_21415; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21417 = 12'hb64 == _T_196[11:0] ? image_2916 : _GEN_21416; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21418 = 12'hb65 == _T_196[11:0] ? image_2917 : _GEN_21417; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21419 = 12'hb66 == _T_196[11:0] ? image_2918 : _GEN_21418; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21420 = 12'hb67 == _T_196[11:0] ? image_2919 : _GEN_21419; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21421 = 12'hb68 == _T_196[11:0] ? image_2920 : _GEN_21420; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21422 = 12'hb69 == _T_196[11:0] ? image_2921 : _GEN_21421; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21423 = 12'hb6a == _T_196[11:0] ? image_2922 : _GEN_21422; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21424 = 12'hb6b == _T_196[11:0] ? image_2923 : _GEN_21423; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21425 = 12'hb6c == _T_196[11:0] ? image_2924 : _GEN_21424; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21426 = 12'hb6d == _T_196[11:0] ? image_2925 : _GEN_21425; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21427 = 12'hb6e == _T_196[11:0] ? image_2926 : _GEN_21426; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21428 = 12'hb6f == _T_196[11:0] ? image_2927 : _GEN_21427; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21429 = 12'hb70 == _T_196[11:0] ? image_2928 : _GEN_21428; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21430 = 12'hb71 == _T_196[11:0] ? image_2929 : _GEN_21429; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21431 = 12'hb72 == _T_196[11:0] ? image_2930 : _GEN_21430; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21432 = 12'hb73 == _T_196[11:0] ? image_2931 : _GEN_21431; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21433 = 12'hb74 == _T_196[11:0] ? image_2932 : _GEN_21432; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21434 = 12'hb75 == _T_196[11:0] ? image_2933 : _GEN_21433; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21435 = 12'hb76 == _T_196[11:0] ? image_2934 : _GEN_21434; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21436 = 12'hb77 == _T_196[11:0] ? 4'h0 : _GEN_21435; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21437 = 12'hb78 == _T_196[11:0] ? 4'h0 : _GEN_21436; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21438 = 12'hb79 == _T_196[11:0] ? 4'h0 : _GEN_21437; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21439 = 12'hb7a == _T_196[11:0] ? 4'h0 : _GEN_21438; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21440 = 12'hb7b == _T_196[11:0] ? 4'h0 : _GEN_21439; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21441 = 12'hb7c == _T_196[11:0] ? 4'h0 : _GEN_21440; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21442 = 12'hb7d == _T_196[11:0] ? 4'h0 : _GEN_21441; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21443 = 12'hb7e == _T_196[11:0] ? 4'h0 : _GEN_21442; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21444 = 12'hb7f == _T_196[11:0] ? 4'h0 : _GEN_21443; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21445 = 12'hb80 == _T_196[11:0] ? 4'h0 : _GEN_21444; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21446 = 12'hb81 == _T_196[11:0] ? 4'h0 : _GEN_21445; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21447 = 12'hb82 == _T_196[11:0] ? 4'h0 : _GEN_21446; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21448 = 12'hb83 == _T_196[11:0] ? 4'h0 : _GEN_21447; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21449 = 12'hb84 == _T_196[11:0] ? 4'h0 : _GEN_21448; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21450 = 12'hb85 == _T_196[11:0] ? 4'h0 : _GEN_21449; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21451 = 12'hb86 == _T_196[11:0] ? 4'h0 : _GEN_21450; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21452 = 12'hb87 == _T_196[11:0] ? 4'h0 : _GEN_21451; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21453 = 12'hb88 == _T_196[11:0] ? 4'h0 : _GEN_21452; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21454 = 12'hb89 == _T_196[11:0] ? 4'h0 : _GEN_21453; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21455 = 12'hb8a == _T_196[11:0] ? 4'h0 : _GEN_21454; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21456 = 12'hb8b == _T_196[11:0] ? 4'h0 : _GEN_21455; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21457 = 12'hb8c == _T_196[11:0] ? 4'h0 : _GEN_21456; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21458 = 12'hb8d == _T_196[11:0] ? 4'h0 : _GEN_21457; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21459 = 12'hb8e == _T_196[11:0] ? 4'h0 : _GEN_21458; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21460 = 12'hb8f == _T_196[11:0] ? 4'h0 : _GEN_21459; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21461 = 12'hb90 == _T_196[11:0] ? 4'h0 : _GEN_21460; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21462 = 12'hb91 == _T_196[11:0] ? 4'h0 : _GEN_21461; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21463 = 12'hb92 == _T_196[11:0] ? 4'h0 : _GEN_21462; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21464 = 12'hb93 == _T_196[11:0] ? 4'h0 : _GEN_21463; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21465 = 12'hb94 == _T_196[11:0] ? 4'h0 : _GEN_21464; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21466 = 12'hb95 == _T_196[11:0] ? image_2965 : _GEN_21465; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21467 = 12'hb96 == _T_196[11:0] ? image_2966 : _GEN_21466; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21468 = 12'hb97 == _T_196[11:0] ? image_2967 : _GEN_21467; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21469 = 12'hb98 == _T_196[11:0] ? image_2968 : _GEN_21468; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21470 = 12'hb99 == _T_196[11:0] ? image_2969 : _GEN_21469; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21471 = 12'hb9a == _T_196[11:0] ? image_2970 : _GEN_21470; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21472 = 12'hb9b == _T_196[11:0] ? image_2971 : _GEN_21471; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21473 = 12'hb9c == _T_196[11:0] ? image_2972 : _GEN_21472; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21474 = 12'hb9d == _T_196[11:0] ? image_2973 : _GEN_21473; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21475 = 12'hb9e == _T_196[11:0] ? image_2974 : _GEN_21474; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21476 = 12'hb9f == _T_196[11:0] ? image_2975 : _GEN_21475; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21477 = 12'hba0 == _T_196[11:0] ? image_2976 : _GEN_21476; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21478 = 12'hba1 == _T_196[11:0] ? image_2977 : _GEN_21477; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21479 = 12'hba2 == _T_196[11:0] ? image_2978 : _GEN_21478; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21480 = 12'hba3 == _T_196[11:0] ? image_2979 : _GEN_21479; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21481 = 12'hba4 == _T_196[11:0] ? image_2980 : _GEN_21480; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21482 = 12'hba5 == _T_196[11:0] ? image_2981 : _GEN_21481; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21483 = 12'hba6 == _T_196[11:0] ? image_2982 : _GEN_21482; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21484 = 12'hba7 == _T_196[11:0] ? image_2983 : _GEN_21483; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21485 = 12'hba8 == _T_196[11:0] ? image_2984 : _GEN_21484; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21486 = 12'hba9 == _T_196[11:0] ? image_2985 : _GEN_21485; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21487 = 12'hbaa == _T_196[11:0] ? image_2986 : _GEN_21486; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21488 = 12'hbab == _T_196[11:0] ? image_2987 : _GEN_21487; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21489 = 12'hbac == _T_196[11:0] ? image_2988 : _GEN_21488; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21490 = 12'hbad == _T_196[11:0] ? image_2989 : _GEN_21489; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21491 = 12'hbae == _T_196[11:0] ? image_2990 : _GEN_21490; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21492 = 12'hbaf == _T_196[11:0] ? image_2991 : _GEN_21491; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21493 = 12'hbb0 == _T_196[11:0] ? image_2992 : _GEN_21492; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21494 = 12'hbb1 == _T_196[11:0] ? image_2993 : _GEN_21493; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21495 = 12'hbb2 == _T_196[11:0] ? image_2994 : _GEN_21494; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21496 = 12'hbb3 == _T_196[11:0] ? image_2995 : _GEN_21495; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21497 = 12'hbb4 == _T_196[11:0] ? image_2996 : _GEN_21496; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21498 = 12'hbb5 == _T_196[11:0] ? 4'h0 : _GEN_21497; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21499 = 12'hbb6 == _T_196[11:0] ? 4'h0 : _GEN_21498; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21500 = 12'hbb7 == _T_196[11:0] ? 4'h0 : _GEN_21499; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21501 = 12'hbb8 == _T_196[11:0] ? 4'h0 : _GEN_21500; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21502 = 12'hbb9 == _T_196[11:0] ? 4'h0 : _GEN_21501; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21503 = 12'hbba == _T_196[11:0] ? 4'h0 : _GEN_21502; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21504 = 12'hbbb == _T_196[11:0] ? 4'h0 : _GEN_21503; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21505 = 12'hbbc == _T_196[11:0] ? 4'h0 : _GEN_21504; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21506 = 12'hbbd == _T_196[11:0] ? 4'h0 : _GEN_21505; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21507 = 12'hbbe == _T_196[11:0] ? 4'h0 : _GEN_21506; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21508 = 12'hbbf == _T_196[11:0] ? 4'h0 : _GEN_21507; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21509 = 12'hbc0 == _T_196[11:0] ? 4'h0 : _GEN_21508; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21510 = 12'hbc1 == _T_196[11:0] ? 4'h0 : _GEN_21509; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21511 = 12'hbc2 == _T_196[11:0] ? 4'h0 : _GEN_21510; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21512 = 12'hbc3 == _T_196[11:0] ? 4'h0 : _GEN_21511; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21513 = 12'hbc4 == _T_196[11:0] ? 4'h0 : _GEN_21512; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21514 = 12'hbc5 == _T_196[11:0] ? 4'h0 : _GEN_21513; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21515 = 12'hbc6 == _T_196[11:0] ? 4'h0 : _GEN_21514; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21516 = 12'hbc7 == _T_196[11:0] ? 4'h0 : _GEN_21515; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21517 = 12'hbc8 == _T_196[11:0] ? 4'h0 : _GEN_21516; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21518 = 12'hbc9 == _T_196[11:0] ? 4'h0 : _GEN_21517; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21519 = 12'hbca == _T_196[11:0] ? 4'h0 : _GEN_21518; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21520 = 12'hbcb == _T_196[11:0] ? 4'h0 : _GEN_21519; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21521 = 12'hbcc == _T_196[11:0] ? 4'h0 : _GEN_21520; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21522 = 12'hbcd == _T_196[11:0] ? 4'h0 : _GEN_21521; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21523 = 12'hbce == _T_196[11:0] ? 4'h0 : _GEN_21522; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21524 = 12'hbcf == _T_196[11:0] ? 4'h0 : _GEN_21523; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21525 = 12'hbd0 == _T_196[11:0] ? 4'h0 : _GEN_21524; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21526 = 12'hbd1 == _T_196[11:0] ? 4'h0 : _GEN_21525; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21527 = 12'hbd2 == _T_196[11:0] ? 4'h0 : _GEN_21526; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21528 = 12'hbd3 == _T_196[11:0] ? 4'h0 : _GEN_21527; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21529 = 12'hbd4 == _T_196[11:0] ? 4'h0 : _GEN_21528; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21530 = 12'hbd5 == _T_196[11:0] ? 4'h0 : _GEN_21529; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21531 = 12'hbd6 == _T_196[11:0] ? 4'h0 : _GEN_21530; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21532 = 12'hbd7 == _T_196[11:0] ? 4'h0 : _GEN_21531; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21533 = 12'hbd8 == _T_196[11:0] ? 4'h0 : _GEN_21532; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21534 = 12'hbd9 == _T_196[11:0] ? 4'h0 : _GEN_21533; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21535 = 12'hbda == _T_196[11:0] ? 4'h0 : _GEN_21534; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21536 = 12'hbdb == _T_196[11:0] ? image_3035 : _GEN_21535; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21537 = 12'hbdc == _T_196[11:0] ? image_3036 : _GEN_21536; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21538 = 12'hbdd == _T_196[11:0] ? image_3037 : _GEN_21537; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21539 = 12'hbde == _T_196[11:0] ? image_3038 : _GEN_21538; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21540 = 12'hbdf == _T_196[11:0] ? image_3039 : _GEN_21539; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21541 = 12'hbe0 == _T_196[11:0] ? image_3040 : _GEN_21540; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21542 = 12'hbe1 == _T_196[11:0] ? image_3041 : _GEN_21541; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21543 = 12'hbe2 == _T_196[11:0] ? image_3042 : _GEN_21542; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21544 = 12'hbe3 == _T_196[11:0] ? image_3043 : _GEN_21543; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21545 = 12'hbe4 == _T_196[11:0] ? image_3044 : _GEN_21544; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21546 = 12'hbe5 == _T_196[11:0] ? image_3045 : _GEN_21545; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21547 = 12'hbe6 == _T_196[11:0] ? image_3046 : _GEN_21546; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21548 = 12'hbe7 == _T_196[11:0] ? image_3047 : _GEN_21547; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21549 = 12'hbe8 == _T_196[11:0] ? image_3048 : _GEN_21548; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21550 = 12'hbe9 == _T_196[11:0] ? image_3049 : _GEN_21549; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21551 = 12'hbea == _T_196[11:0] ? image_3050 : _GEN_21550; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21552 = 12'hbeb == _T_196[11:0] ? image_3051 : _GEN_21551; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21553 = 12'hbec == _T_196[11:0] ? image_3052 : _GEN_21552; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21554 = 12'hbed == _T_196[11:0] ? image_3053 : _GEN_21553; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21555 = 12'hbee == _T_196[11:0] ? image_3054 : _GEN_21554; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21556 = 12'hbef == _T_196[11:0] ? image_3055 : _GEN_21555; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21557 = 12'hbf0 == _T_196[11:0] ? image_3056 : _GEN_21556; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21558 = 12'hbf1 == _T_196[11:0] ? 4'h0 : _GEN_21557; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21559 = 12'hbf2 == _T_196[11:0] ? 4'h0 : _GEN_21558; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21560 = 12'hbf3 == _T_196[11:0] ? 4'h0 : _GEN_21559; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21561 = 12'hbf4 == _T_196[11:0] ? 4'h0 : _GEN_21560; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21562 = 12'hbf5 == _T_196[11:0] ? 4'h0 : _GEN_21561; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21563 = 12'hbf6 == _T_196[11:0] ? 4'h0 : _GEN_21562; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21564 = 12'hbf7 == _T_196[11:0] ? 4'h0 : _GEN_21563; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21565 = 12'hbf8 == _T_196[11:0] ? 4'h0 : _GEN_21564; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21566 = 12'hbf9 == _T_196[11:0] ? 4'h0 : _GEN_21565; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21567 = 12'hbfa == _T_196[11:0] ? 4'h0 : _GEN_21566; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21568 = 12'hbfb == _T_196[11:0] ? 4'h0 : _GEN_21567; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21569 = 12'hbfc == _T_196[11:0] ? 4'h0 : _GEN_21568; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21570 = 12'hbfd == _T_196[11:0] ? 4'h0 : _GEN_21569; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21571 = 12'hbfe == _T_196[11:0] ? 4'h0 : _GEN_21570; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21572 = 12'hbff == _T_196[11:0] ? 4'h0 : _GEN_21571; // @[Filter.scala 138:46]
  wire [31:0] _T_199 = pixelIndex + 32'h7; // @[Filter.scala 133:29]
  wire [31:0] _T_200 = _T_199 / 32'h40; // @[Filter.scala 133:36]
  wire [31:0] _T_202 = _T_200 + _GEN_24805; // @[Filter.scala 133:51]
  wire [31:0] _T_204 = _T_202 - 32'h1; // @[Filter.scala 133:67]
  wire [31:0] _GEN_56 = _T_199 % 32'h40; // @[Filter.scala 134:36]
  wire [6:0] _T_207 = _GEN_56[6:0]; // @[Filter.scala 134:36]
  wire [6:0] _T_209 = _T_207 + _GEN_24806; // @[Filter.scala 134:51]
  wire [6:0] _T_211 = _T_209 - 7'h1; // @[Filter.scala 134:67]
  wire  _T_213 = _T_204 >= 32'h40; // @[Filter.scala 135:27]
  wire  _T_217 = _T_211 >= 7'h30; // @[Filter.scala 135:59]
  wire  _T_218 = _T_213 | _T_217; // @[Filter.scala 135:54]
  wire [13:0] _T_219 = _T_211 * 7'h40; // @[Filter.scala 138:57]
  wire [31:0] _GEN_24828 = {{18'd0}, _T_219}; // @[Filter.scala 138:72]
  wire [31:0] _T_221 = _GEN_24828 + _T_204; // @[Filter.scala 138:72]
  wire [3:0] _GEN_21586 = 12'hc == _T_221[11:0] ? image_12 : 4'h0; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21587 = 12'hd == _T_221[11:0] ? 4'h0 : _GEN_21586; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21588 = 12'he == _T_221[11:0] ? image_14 : _GEN_21587; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21589 = 12'hf == _T_221[11:0] ? image_15 : _GEN_21588; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21590 = 12'h10 == _T_221[11:0] ? image_16 : _GEN_21589; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21591 = 12'h11 == _T_221[11:0] ? image_17 : _GEN_21590; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21592 = 12'h12 == _T_221[11:0] ? image_18 : _GEN_21591; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21593 = 12'h13 == _T_221[11:0] ? image_19 : _GEN_21592; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21594 = 12'h14 == _T_221[11:0] ? image_20 : _GEN_21593; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21595 = 12'h15 == _T_221[11:0] ? image_21 : _GEN_21594; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21596 = 12'h16 == _T_221[11:0] ? image_22 : _GEN_21595; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21597 = 12'h17 == _T_221[11:0] ? image_23 : _GEN_21596; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21598 = 12'h18 == _T_221[11:0] ? 4'h0 : _GEN_21597; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21599 = 12'h19 == _T_221[11:0] ? 4'h0 : _GEN_21598; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21600 = 12'h1a == _T_221[11:0] ? 4'h0 : _GEN_21599; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21601 = 12'h1b == _T_221[11:0] ? 4'h0 : _GEN_21600; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21602 = 12'h1c == _T_221[11:0] ? 4'h0 : _GEN_21601; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21603 = 12'h1d == _T_221[11:0] ? 4'h0 : _GEN_21602; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21604 = 12'h1e == _T_221[11:0] ? 4'h0 : _GEN_21603; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21605 = 12'h1f == _T_221[11:0] ? 4'h0 : _GEN_21604; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21606 = 12'h20 == _T_221[11:0] ? 4'h0 : _GEN_21605; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21607 = 12'h21 == _T_221[11:0] ? 4'h0 : _GEN_21606; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21608 = 12'h22 == _T_221[11:0] ? 4'h0 : _GEN_21607; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21609 = 12'h23 == _T_221[11:0] ? image_35 : _GEN_21608; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21610 = 12'h24 == _T_221[11:0] ? image_36 : _GEN_21609; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21611 = 12'h25 == _T_221[11:0] ? image_37 : _GEN_21610; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21612 = 12'h26 == _T_221[11:0] ? image_38 : _GEN_21611; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21613 = 12'h27 == _T_221[11:0] ? image_39 : _GEN_21612; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21614 = 12'h28 == _T_221[11:0] ? image_40 : _GEN_21613; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21615 = 12'h29 == _T_221[11:0] ? image_41 : _GEN_21614; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21616 = 12'h2a == _T_221[11:0] ? image_42 : _GEN_21615; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21617 = 12'h2b == _T_221[11:0] ? 4'h0 : _GEN_21616; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21618 = 12'h2c == _T_221[11:0] ? 4'h0 : _GEN_21617; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21619 = 12'h2d == _T_221[11:0] ? 4'h0 : _GEN_21618; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21620 = 12'h2e == _T_221[11:0] ? 4'h0 : _GEN_21619; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21621 = 12'h2f == _T_221[11:0] ? 4'h0 : _GEN_21620; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21622 = 12'h30 == _T_221[11:0] ? 4'h0 : _GEN_21621; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21623 = 12'h31 == _T_221[11:0] ? 4'h0 : _GEN_21622; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21624 = 12'h32 == _T_221[11:0] ? 4'h0 : _GEN_21623; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21625 = 12'h33 == _T_221[11:0] ? 4'h0 : _GEN_21624; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21626 = 12'h34 == _T_221[11:0] ? 4'h0 : _GEN_21625; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21627 = 12'h35 == _T_221[11:0] ? 4'h0 : _GEN_21626; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21628 = 12'h36 == _T_221[11:0] ? 4'h0 : _GEN_21627; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21629 = 12'h37 == _T_221[11:0] ? 4'h0 : _GEN_21628; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21630 = 12'h38 == _T_221[11:0] ? 4'h0 : _GEN_21629; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21631 = 12'h39 == _T_221[11:0] ? 4'h0 : _GEN_21630; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21632 = 12'h3a == _T_221[11:0] ? 4'h0 : _GEN_21631; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21633 = 12'h3b == _T_221[11:0] ? 4'h0 : _GEN_21632; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21634 = 12'h3c == _T_221[11:0] ? 4'h0 : _GEN_21633; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21635 = 12'h3d == _T_221[11:0] ? 4'h0 : _GEN_21634; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21636 = 12'h3e == _T_221[11:0] ? 4'h0 : _GEN_21635; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21637 = 12'h3f == _T_221[11:0] ? 4'h0 : _GEN_21636; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21638 = 12'h40 == _T_221[11:0] ? 4'h0 : _GEN_21637; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21639 = 12'h41 == _T_221[11:0] ? 4'h0 : _GEN_21638; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21640 = 12'h42 == _T_221[11:0] ? 4'h0 : _GEN_21639; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21641 = 12'h43 == _T_221[11:0] ? 4'h0 : _GEN_21640; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21642 = 12'h44 == _T_221[11:0] ? 4'h0 : _GEN_21641; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21643 = 12'h45 == _T_221[11:0] ? 4'h0 : _GEN_21642; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21644 = 12'h46 == _T_221[11:0] ? 4'h0 : _GEN_21643; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21645 = 12'h47 == _T_221[11:0] ? 4'h0 : _GEN_21644; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21646 = 12'h48 == _T_221[11:0] ? 4'h0 : _GEN_21645; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21647 = 12'h49 == _T_221[11:0] ? 4'h0 : _GEN_21646; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21648 = 12'h4a == _T_221[11:0] ? 4'h0 : _GEN_21647; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21649 = 12'h4b == _T_221[11:0] ? image_75 : _GEN_21648; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21650 = 12'h4c == _T_221[11:0] ? image_76 : _GEN_21649; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21651 = 12'h4d == _T_221[11:0] ? image_77 : _GEN_21650; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21652 = 12'h4e == _T_221[11:0] ? image_78 : _GEN_21651; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21653 = 12'h4f == _T_221[11:0] ? image_79 : _GEN_21652; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21654 = 12'h50 == _T_221[11:0] ? image_80 : _GEN_21653; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21655 = 12'h51 == _T_221[11:0] ? image_81 : _GEN_21654; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21656 = 12'h52 == _T_221[11:0] ? image_82 : _GEN_21655; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21657 = 12'h53 == _T_221[11:0] ? image_83 : _GEN_21656; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21658 = 12'h54 == _T_221[11:0] ? image_84 : _GEN_21657; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21659 = 12'h55 == _T_221[11:0] ? image_85 : _GEN_21658; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21660 = 12'h56 == _T_221[11:0] ? image_86 : _GEN_21659; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21661 = 12'h57 == _T_221[11:0] ? image_87 : _GEN_21660; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21662 = 12'h58 == _T_221[11:0] ? image_88 : _GEN_21661; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21663 = 12'h59 == _T_221[11:0] ? image_89 : _GEN_21662; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21664 = 12'h5a == _T_221[11:0] ? image_90 : _GEN_21663; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21665 = 12'h5b == _T_221[11:0] ? 4'h0 : _GEN_21664; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21666 = 12'h5c == _T_221[11:0] ? 4'h0 : _GEN_21665; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21667 = 12'h5d == _T_221[11:0] ? image_93 : _GEN_21666; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21668 = 12'h5e == _T_221[11:0] ? 4'h0 : _GEN_21667; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21669 = 12'h5f == _T_221[11:0] ? image_95 : _GEN_21668; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21670 = 12'h60 == _T_221[11:0] ? image_96 : _GEN_21669; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21671 = 12'h61 == _T_221[11:0] ? image_97 : _GEN_21670; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21672 = 12'h62 == _T_221[11:0] ? image_98 : _GEN_21671; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21673 = 12'h63 == _T_221[11:0] ? image_99 : _GEN_21672; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21674 = 12'h64 == _T_221[11:0] ? image_100 : _GEN_21673; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21675 = 12'h65 == _T_221[11:0] ? image_101 : _GEN_21674; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21676 = 12'h66 == _T_221[11:0] ? image_102 : _GEN_21675; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21677 = 12'h67 == _T_221[11:0] ? image_103 : _GEN_21676; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21678 = 12'h68 == _T_221[11:0] ? image_104 : _GEN_21677; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21679 = 12'h69 == _T_221[11:0] ? image_105 : _GEN_21678; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21680 = 12'h6a == _T_221[11:0] ? image_106 : _GEN_21679; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21681 = 12'h6b == _T_221[11:0] ? image_107 : _GEN_21680; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21682 = 12'h6c == _T_221[11:0] ? image_108 : _GEN_21681; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21683 = 12'h6d == _T_221[11:0] ? 4'h0 : _GEN_21682; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21684 = 12'h6e == _T_221[11:0] ? 4'h0 : _GEN_21683; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21685 = 12'h6f == _T_221[11:0] ? 4'h0 : _GEN_21684; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21686 = 12'h70 == _T_221[11:0] ? 4'h0 : _GEN_21685; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21687 = 12'h71 == _T_221[11:0] ? 4'h0 : _GEN_21686; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21688 = 12'h72 == _T_221[11:0] ? 4'h0 : _GEN_21687; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21689 = 12'h73 == _T_221[11:0] ? 4'h0 : _GEN_21688; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21690 = 12'h74 == _T_221[11:0] ? 4'h0 : _GEN_21689; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21691 = 12'h75 == _T_221[11:0] ? 4'h0 : _GEN_21690; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21692 = 12'h76 == _T_221[11:0] ? 4'h0 : _GEN_21691; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21693 = 12'h77 == _T_221[11:0] ? 4'h0 : _GEN_21692; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21694 = 12'h78 == _T_221[11:0] ? 4'h0 : _GEN_21693; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21695 = 12'h79 == _T_221[11:0] ? 4'h0 : _GEN_21694; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21696 = 12'h7a == _T_221[11:0] ? 4'h0 : _GEN_21695; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21697 = 12'h7b == _T_221[11:0] ? 4'h0 : _GEN_21696; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21698 = 12'h7c == _T_221[11:0] ? 4'h0 : _GEN_21697; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21699 = 12'h7d == _T_221[11:0] ? 4'h0 : _GEN_21698; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21700 = 12'h7e == _T_221[11:0] ? 4'h0 : _GEN_21699; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21701 = 12'h7f == _T_221[11:0] ? 4'h0 : _GEN_21700; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21702 = 12'h80 == _T_221[11:0] ? 4'h0 : _GEN_21701; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21703 = 12'h81 == _T_221[11:0] ? 4'h0 : _GEN_21702; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21704 = 12'h82 == _T_221[11:0] ? 4'h0 : _GEN_21703; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21705 = 12'h83 == _T_221[11:0] ? 4'h0 : _GEN_21704; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21706 = 12'h84 == _T_221[11:0] ? 4'h0 : _GEN_21705; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21707 = 12'h85 == _T_221[11:0] ? 4'h0 : _GEN_21706; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21708 = 12'h86 == _T_221[11:0] ? 4'h0 : _GEN_21707; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21709 = 12'h87 == _T_221[11:0] ? 4'h0 : _GEN_21708; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21710 = 12'h88 == _T_221[11:0] ? image_136 : _GEN_21709; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21711 = 12'h89 == _T_221[11:0] ? image_137 : _GEN_21710; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21712 = 12'h8a == _T_221[11:0] ? image_138 : _GEN_21711; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21713 = 12'h8b == _T_221[11:0] ? image_139 : _GEN_21712; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21714 = 12'h8c == _T_221[11:0] ? image_140 : _GEN_21713; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21715 = 12'h8d == _T_221[11:0] ? image_141 : _GEN_21714; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21716 = 12'h8e == _T_221[11:0] ? image_142 : _GEN_21715; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21717 = 12'h8f == _T_221[11:0] ? image_143 : _GEN_21716; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21718 = 12'h90 == _T_221[11:0] ? image_144 : _GEN_21717; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21719 = 12'h91 == _T_221[11:0] ? image_145 : _GEN_21718; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21720 = 12'h92 == _T_221[11:0] ? image_146 : _GEN_21719; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21721 = 12'h93 == _T_221[11:0] ? image_147 : _GEN_21720; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21722 = 12'h94 == _T_221[11:0] ? image_148 : _GEN_21721; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21723 = 12'h95 == _T_221[11:0] ? image_149 : _GEN_21722; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21724 = 12'h96 == _T_221[11:0] ? image_150 : _GEN_21723; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21725 = 12'h97 == _T_221[11:0] ? image_151 : _GEN_21724; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21726 = 12'h98 == _T_221[11:0] ? image_152 : _GEN_21725; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21727 = 12'h99 == _T_221[11:0] ? image_153 : _GEN_21726; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21728 = 12'h9a == _T_221[11:0] ? image_154 : _GEN_21727; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21729 = 12'h9b == _T_221[11:0] ? image_155 : _GEN_21728; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21730 = 12'h9c == _T_221[11:0] ? 4'h0 : _GEN_21729; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21731 = 12'h9d == _T_221[11:0] ? image_157 : _GEN_21730; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21732 = 12'h9e == _T_221[11:0] ? image_158 : _GEN_21731; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21733 = 12'h9f == _T_221[11:0] ? image_159 : _GEN_21732; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21734 = 12'ha0 == _T_221[11:0] ? image_160 : _GEN_21733; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21735 = 12'ha1 == _T_221[11:0] ? image_161 : _GEN_21734; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21736 = 12'ha2 == _T_221[11:0] ? image_162 : _GEN_21735; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21737 = 12'ha3 == _T_221[11:0] ? image_163 : _GEN_21736; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21738 = 12'ha4 == _T_221[11:0] ? image_164 : _GEN_21737; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21739 = 12'ha5 == _T_221[11:0] ? image_165 : _GEN_21738; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21740 = 12'ha6 == _T_221[11:0] ? image_166 : _GEN_21739; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21741 = 12'ha7 == _T_221[11:0] ? image_167 : _GEN_21740; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21742 = 12'ha8 == _T_221[11:0] ? image_168 : _GEN_21741; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21743 = 12'ha9 == _T_221[11:0] ? image_169 : _GEN_21742; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21744 = 12'haa == _T_221[11:0] ? image_170 : _GEN_21743; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21745 = 12'hab == _T_221[11:0] ? image_171 : _GEN_21744; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21746 = 12'hac == _T_221[11:0] ? image_172 : _GEN_21745; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21747 = 12'had == _T_221[11:0] ? image_173 : _GEN_21746; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21748 = 12'hae == _T_221[11:0] ? image_174 : _GEN_21747; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21749 = 12'haf == _T_221[11:0] ? image_175 : _GEN_21748; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21750 = 12'hb0 == _T_221[11:0] ? image_176 : _GEN_21749; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21751 = 12'hb1 == _T_221[11:0] ? image_177 : _GEN_21750; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21752 = 12'hb2 == _T_221[11:0] ? image_178 : _GEN_21751; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21753 = 12'hb3 == _T_221[11:0] ? image_179 : _GEN_21752; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21754 = 12'hb4 == _T_221[11:0] ? 4'h0 : _GEN_21753; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21755 = 12'hb5 == _T_221[11:0] ? 4'h0 : _GEN_21754; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21756 = 12'hb6 == _T_221[11:0] ? 4'h0 : _GEN_21755; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21757 = 12'hb7 == _T_221[11:0] ? 4'h0 : _GEN_21756; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21758 = 12'hb8 == _T_221[11:0] ? 4'h0 : _GEN_21757; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21759 = 12'hb9 == _T_221[11:0] ? 4'h0 : _GEN_21758; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21760 = 12'hba == _T_221[11:0] ? 4'h0 : _GEN_21759; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21761 = 12'hbb == _T_221[11:0] ? 4'h0 : _GEN_21760; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21762 = 12'hbc == _T_221[11:0] ? 4'h0 : _GEN_21761; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21763 = 12'hbd == _T_221[11:0] ? 4'h0 : _GEN_21762; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21764 = 12'hbe == _T_221[11:0] ? 4'h0 : _GEN_21763; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21765 = 12'hbf == _T_221[11:0] ? 4'h0 : _GEN_21764; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21766 = 12'hc0 == _T_221[11:0] ? 4'h0 : _GEN_21765; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21767 = 12'hc1 == _T_221[11:0] ? 4'h0 : _GEN_21766; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21768 = 12'hc2 == _T_221[11:0] ? 4'h0 : _GEN_21767; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21769 = 12'hc3 == _T_221[11:0] ? 4'h0 : _GEN_21768; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21770 = 12'hc4 == _T_221[11:0] ? 4'h0 : _GEN_21769; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21771 = 12'hc5 == _T_221[11:0] ? 4'h0 : _GEN_21770; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21772 = 12'hc6 == _T_221[11:0] ? 4'h0 : _GEN_21771; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21773 = 12'hc7 == _T_221[11:0] ? image_199 : _GEN_21772; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21774 = 12'hc8 == _T_221[11:0] ? image_200 : _GEN_21773; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21775 = 12'hc9 == _T_221[11:0] ? image_201 : _GEN_21774; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21776 = 12'hca == _T_221[11:0] ? image_202 : _GEN_21775; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21777 = 12'hcb == _T_221[11:0] ? image_203 : _GEN_21776; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21778 = 12'hcc == _T_221[11:0] ? image_204 : _GEN_21777; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21779 = 12'hcd == _T_221[11:0] ? image_205 : _GEN_21778; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21780 = 12'hce == _T_221[11:0] ? image_206 : _GEN_21779; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21781 = 12'hcf == _T_221[11:0] ? image_207 : _GEN_21780; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21782 = 12'hd0 == _T_221[11:0] ? image_208 : _GEN_21781; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21783 = 12'hd1 == _T_221[11:0] ? image_209 : _GEN_21782; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21784 = 12'hd2 == _T_221[11:0] ? image_210 : _GEN_21783; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21785 = 12'hd3 == _T_221[11:0] ? image_211 : _GEN_21784; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21786 = 12'hd4 == _T_221[11:0] ? image_212 : _GEN_21785; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21787 = 12'hd5 == _T_221[11:0] ? image_213 : _GEN_21786; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21788 = 12'hd6 == _T_221[11:0] ? image_214 : _GEN_21787; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21789 = 12'hd7 == _T_221[11:0] ? image_215 : _GEN_21788; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21790 = 12'hd8 == _T_221[11:0] ? image_216 : _GEN_21789; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21791 = 12'hd9 == _T_221[11:0] ? image_217 : _GEN_21790; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21792 = 12'hda == _T_221[11:0] ? image_218 : _GEN_21791; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21793 = 12'hdb == _T_221[11:0] ? image_219 : _GEN_21792; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21794 = 12'hdc == _T_221[11:0] ? image_220 : _GEN_21793; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21795 = 12'hdd == _T_221[11:0] ? image_221 : _GEN_21794; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21796 = 12'hde == _T_221[11:0] ? image_222 : _GEN_21795; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21797 = 12'hdf == _T_221[11:0] ? image_223 : _GEN_21796; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21798 = 12'he0 == _T_221[11:0] ? image_224 : _GEN_21797; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21799 = 12'he1 == _T_221[11:0] ? image_225 : _GEN_21798; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21800 = 12'he2 == _T_221[11:0] ? image_226 : _GEN_21799; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21801 = 12'he3 == _T_221[11:0] ? image_227 : _GEN_21800; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21802 = 12'he4 == _T_221[11:0] ? image_228 : _GEN_21801; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21803 = 12'he5 == _T_221[11:0] ? image_229 : _GEN_21802; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21804 = 12'he6 == _T_221[11:0] ? image_230 : _GEN_21803; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21805 = 12'he7 == _T_221[11:0] ? image_231 : _GEN_21804; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21806 = 12'he8 == _T_221[11:0] ? image_232 : _GEN_21805; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21807 = 12'he9 == _T_221[11:0] ? image_233 : _GEN_21806; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21808 = 12'hea == _T_221[11:0] ? image_234 : _GEN_21807; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21809 = 12'heb == _T_221[11:0] ? image_235 : _GEN_21808; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21810 = 12'hec == _T_221[11:0] ? image_236 : _GEN_21809; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21811 = 12'hed == _T_221[11:0] ? image_237 : _GEN_21810; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21812 = 12'hee == _T_221[11:0] ? image_238 : _GEN_21811; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21813 = 12'hef == _T_221[11:0] ? image_239 : _GEN_21812; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21814 = 12'hf0 == _T_221[11:0] ? image_240 : _GEN_21813; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21815 = 12'hf1 == _T_221[11:0] ? image_241 : _GEN_21814; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21816 = 12'hf2 == _T_221[11:0] ? image_242 : _GEN_21815; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21817 = 12'hf3 == _T_221[11:0] ? image_243 : _GEN_21816; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21818 = 12'hf4 == _T_221[11:0] ? image_244 : _GEN_21817; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21819 = 12'hf5 == _T_221[11:0] ? image_245 : _GEN_21818; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21820 = 12'hf6 == _T_221[11:0] ? image_246 : _GEN_21819; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21821 = 12'hf7 == _T_221[11:0] ? 4'h0 : _GEN_21820; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21822 = 12'hf8 == _T_221[11:0] ? 4'h0 : _GEN_21821; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21823 = 12'hf9 == _T_221[11:0] ? 4'h0 : _GEN_21822; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21824 = 12'hfa == _T_221[11:0] ? 4'h0 : _GEN_21823; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21825 = 12'hfb == _T_221[11:0] ? 4'h0 : _GEN_21824; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21826 = 12'hfc == _T_221[11:0] ? 4'h0 : _GEN_21825; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21827 = 12'hfd == _T_221[11:0] ? 4'h0 : _GEN_21826; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21828 = 12'hfe == _T_221[11:0] ? 4'h0 : _GEN_21827; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21829 = 12'hff == _T_221[11:0] ? 4'h0 : _GEN_21828; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21830 = 12'h100 == _T_221[11:0] ? 4'h0 : _GEN_21829; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21831 = 12'h101 == _T_221[11:0] ? 4'h0 : _GEN_21830; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21832 = 12'h102 == _T_221[11:0] ? 4'h0 : _GEN_21831; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21833 = 12'h103 == _T_221[11:0] ? 4'h0 : _GEN_21832; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21834 = 12'h104 == _T_221[11:0] ? 4'h0 : _GEN_21833; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21835 = 12'h105 == _T_221[11:0] ? 4'h0 : _GEN_21834; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21836 = 12'h106 == _T_221[11:0] ? image_262 : _GEN_21835; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21837 = 12'h107 == _T_221[11:0] ? image_263 : _GEN_21836; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21838 = 12'h108 == _T_221[11:0] ? image_264 : _GEN_21837; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21839 = 12'h109 == _T_221[11:0] ? image_265 : _GEN_21838; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21840 = 12'h10a == _T_221[11:0] ? image_266 : _GEN_21839; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21841 = 12'h10b == _T_221[11:0] ? image_267 : _GEN_21840; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21842 = 12'h10c == _T_221[11:0] ? image_268 : _GEN_21841; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21843 = 12'h10d == _T_221[11:0] ? image_269 : _GEN_21842; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21844 = 12'h10e == _T_221[11:0] ? image_270 : _GEN_21843; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21845 = 12'h10f == _T_221[11:0] ? image_271 : _GEN_21844; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21846 = 12'h110 == _T_221[11:0] ? image_272 : _GEN_21845; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21847 = 12'h111 == _T_221[11:0] ? image_273 : _GEN_21846; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21848 = 12'h112 == _T_221[11:0] ? image_274 : _GEN_21847; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21849 = 12'h113 == _T_221[11:0] ? image_275 : _GEN_21848; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21850 = 12'h114 == _T_221[11:0] ? image_276 : _GEN_21849; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21851 = 12'h115 == _T_221[11:0] ? image_277 : _GEN_21850; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21852 = 12'h116 == _T_221[11:0] ? image_278 : _GEN_21851; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21853 = 12'h117 == _T_221[11:0] ? image_279 : _GEN_21852; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21854 = 12'h118 == _T_221[11:0] ? image_280 : _GEN_21853; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21855 = 12'h119 == _T_221[11:0] ? image_281 : _GEN_21854; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21856 = 12'h11a == _T_221[11:0] ? image_282 : _GEN_21855; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21857 = 12'h11b == _T_221[11:0] ? image_283 : _GEN_21856; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21858 = 12'h11c == _T_221[11:0] ? image_284 : _GEN_21857; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21859 = 12'h11d == _T_221[11:0] ? image_285 : _GEN_21858; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21860 = 12'h11e == _T_221[11:0] ? image_286 : _GEN_21859; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21861 = 12'h11f == _T_221[11:0] ? image_287 : _GEN_21860; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21862 = 12'h120 == _T_221[11:0] ? image_288 : _GEN_21861; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21863 = 12'h121 == _T_221[11:0] ? image_289 : _GEN_21862; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21864 = 12'h122 == _T_221[11:0] ? image_290 : _GEN_21863; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21865 = 12'h123 == _T_221[11:0] ? image_291 : _GEN_21864; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21866 = 12'h124 == _T_221[11:0] ? image_292 : _GEN_21865; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21867 = 12'h125 == _T_221[11:0] ? image_293 : _GEN_21866; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21868 = 12'h126 == _T_221[11:0] ? image_294 : _GEN_21867; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21869 = 12'h127 == _T_221[11:0] ? image_295 : _GEN_21868; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21870 = 12'h128 == _T_221[11:0] ? image_296 : _GEN_21869; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21871 = 12'h129 == _T_221[11:0] ? image_297 : _GEN_21870; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21872 = 12'h12a == _T_221[11:0] ? image_298 : _GEN_21871; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21873 = 12'h12b == _T_221[11:0] ? image_299 : _GEN_21872; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21874 = 12'h12c == _T_221[11:0] ? image_300 : _GEN_21873; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21875 = 12'h12d == _T_221[11:0] ? image_301 : _GEN_21874; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21876 = 12'h12e == _T_221[11:0] ? image_302 : _GEN_21875; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21877 = 12'h12f == _T_221[11:0] ? image_303 : _GEN_21876; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21878 = 12'h130 == _T_221[11:0] ? image_304 : _GEN_21877; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21879 = 12'h131 == _T_221[11:0] ? image_305 : _GEN_21878; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21880 = 12'h132 == _T_221[11:0] ? image_306 : _GEN_21879; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21881 = 12'h133 == _T_221[11:0] ? image_307 : _GEN_21880; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21882 = 12'h134 == _T_221[11:0] ? image_308 : _GEN_21881; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21883 = 12'h135 == _T_221[11:0] ? image_309 : _GEN_21882; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21884 = 12'h136 == _T_221[11:0] ? image_310 : _GEN_21883; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21885 = 12'h137 == _T_221[11:0] ? image_311 : _GEN_21884; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21886 = 12'h138 == _T_221[11:0] ? image_312 : _GEN_21885; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21887 = 12'h139 == _T_221[11:0] ? image_313 : _GEN_21886; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21888 = 12'h13a == _T_221[11:0] ? image_314 : _GEN_21887; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21889 = 12'h13b == _T_221[11:0] ? image_315 : _GEN_21888; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21890 = 12'h13c == _T_221[11:0] ? 4'h0 : _GEN_21889; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21891 = 12'h13d == _T_221[11:0] ? 4'h0 : _GEN_21890; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21892 = 12'h13e == _T_221[11:0] ? 4'h0 : _GEN_21891; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21893 = 12'h13f == _T_221[11:0] ? 4'h0 : _GEN_21892; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21894 = 12'h140 == _T_221[11:0] ? 4'h0 : _GEN_21893; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21895 = 12'h141 == _T_221[11:0] ? 4'h0 : _GEN_21894; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21896 = 12'h142 == _T_221[11:0] ? 4'h0 : _GEN_21895; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21897 = 12'h143 == _T_221[11:0] ? 4'h0 : _GEN_21896; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21898 = 12'h144 == _T_221[11:0] ? 4'h0 : _GEN_21897; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21899 = 12'h145 == _T_221[11:0] ? image_325 : _GEN_21898; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21900 = 12'h146 == _T_221[11:0] ? image_326 : _GEN_21899; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21901 = 12'h147 == _T_221[11:0] ? image_327 : _GEN_21900; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21902 = 12'h148 == _T_221[11:0] ? image_328 : _GEN_21901; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21903 = 12'h149 == _T_221[11:0] ? image_329 : _GEN_21902; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21904 = 12'h14a == _T_221[11:0] ? image_330 : _GEN_21903; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21905 = 12'h14b == _T_221[11:0] ? image_331 : _GEN_21904; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21906 = 12'h14c == _T_221[11:0] ? image_332 : _GEN_21905; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21907 = 12'h14d == _T_221[11:0] ? image_333 : _GEN_21906; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21908 = 12'h14e == _T_221[11:0] ? image_334 : _GEN_21907; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21909 = 12'h14f == _T_221[11:0] ? image_335 : _GEN_21908; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21910 = 12'h150 == _T_221[11:0] ? image_336 : _GEN_21909; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21911 = 12'h151 == _T_221[11:0] ? image_337 : _GEN_21910; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21912 = 12'h152 == _T_221[11:0] ? image_338 : _GEN_21911; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21913 = 12'h153 == _T_221[11:0] ? image_339 : _GEN_21912; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21914 = 12'h154 == _T_221[11:0] ? image_340 : _GEN_21913; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21915 = 12'h155 == _T_221[11:0] ? image_341 : _GEN_21914; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21916 = 12'h156 == _T_221[11:0] ? image_342 : _GEN_21915; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21917 = 12'h157 == _T_221[11:0] ? image_343 : _GEN_21916; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21918 = 12'h158 == _T_221[11:0] ? image_344 : _GEN_21917; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21919 = 12'h159 == _T_221[11:0] ? image_345 : _GEN_21918; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21920 = 12'h15a == _T_221[11:0] ? image_346 : _GEN_21919; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21921 = 12'h15b == _T_221[11:0] ? image_347 : _GEN_21920; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21922 = 12'h15c == _T_221[11:0] ? image_348 : _GEN_21921; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21923 = 12'h15d == _T_221[11:0] ? image_349 : _GEN_21922; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21924 = 12'h15e == _T_221[11:0] ? image_350 : _GEN_21923; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21925 = 12'h15f == _T_221[11:0] ? image_351 : _GEN_21924; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21926 = 12'h160 == _T_221[11:0] ? image_352 : _GEN_21925; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21927 = 12'h161 == _T_221[11:0] ? image_353 : _GEN_21926; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21928 = 12'h162 == _T_221[11:0] ? image_354 : _GEN_21927; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21929 = 12'h163 == _T_221[11:0] ? image_355 : _GEN_21928; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21930 = 12'h164 == _T_221[11:0] ? image_356 : _GEN_21929; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21931 = 12'h165 == _T_221[11:0] ? image_357 : _GEN_21930; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21932 = 12'h166 == _T_221[11:0] ? image_358 : _GEN_21931; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21933 = 12'h167 == _T_221[11:0] ? image_359 : _GEN_21932; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21934 = 12'h168 == _T_221[11:0] ? image_360 : _GEN_21933; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21935 = 12'h169 == _T_221[11:0] ? image_361 : _GEN_21934; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21936 = 12'h16a == _T_221[11:0] ? image_362 : _GEN_21935; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21937 = 12'h16b == _T_221[11:0] ? image_363 : _GEN_21936; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21938 = 12'h16c == _T_221[11:0] ? image_364 : _GEN_21937; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21939 = 12'h16d == _T_221[11:0] ? image_365 : _GEN_21938; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21940 = 12'h16e == _T_221[11:0] ? image_366 : _GEN_21939; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21941 = 12'h16f == _T_221[11:0] ? image_367 : _GEN_21940; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21942 = 12'h170 == _T_221[11:0] ? image_368 : _GEN_21941; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21943 = 12'h171 == _T_221[11:0] ? image_369 : _GEN_21942; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21944 = 12'h172 == _T_221[11:0] ? image_370 : _GEN_21943; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21945 = 12'h173 == _T_221[11:0] ? image_371 : _GEN_21944; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21946 = 12'h174 == _T_221[11:0] ? image_372 : _GEN_21945; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21947 = 12'h175 == _T_221[11:0] ? image_373 : _GEN_21946; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21948 = 12'h176 == _T_221[11:0] ? image_374 : _GEN_21947; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21949 = 12'h177 == _T_221[11:0] ? image_375 : _GEN_21948; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21950 = 12'h178 == _T_221[11:0] ? image_376 : _GEN_21949; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21951 = 12'h179 == _T_221[11:0] ? image_377 : _GEN_21950; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21952 = 12'h17a == _T_221[11:0] ? image_378 : _GEN_21951; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21953 = 12'h17b == _T_221[11:0] ? image_379 : _GEN_21952; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21954 = 12'h17c == _T_221[11:0] ? 4'h0 : _GEN_21953; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21955 = 12'h17d == _T_221[11:0] ? 4'h0 : _GEN_21954; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21956 = 12'h17e == _T_221[11:0] ? 4'h0 : _GEN_21955; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21957 = 12'h17f == _T_221[11:0] ? 4'h0 : _GEN_21956; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21958 = 12'h180 == _T_221[11:0] ? 4'h0 : _GEN_21957; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21959 = 12'h181 == _T_221[11:0] ? 4'h0 : _GEN_21958; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21960 = 12'h182 == _T_221[11:0] ? 4'h0 : _GEN_21959; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21961 = 12'h183 == _T_221[11:0] ? 4'h0 : _GEN_21960; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21962 = 12'h184 == _T_221[11:0] ? image_388 : _GEN_21961; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21963 = 12'h185 == _T_221[11:0] ? image_389 : _GEN_21962; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21964 = 12'h186 == _T_221[11:0] ? image_390 : _GEN_21963; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21965 = 12'h187 == _T_221[11:0] ? image_391 : _GEN_21964; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21966 = 12'h188 == _T_221[11:0] ? image_392 : _GEN_21965; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21967 = 12'h189 == _T_221[11:0] ? image_393 : _GEN_21966; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21968 = 12'h18a == _T_221[11:0] ? image_394 : _GEN_21967; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21969 = 12'h18b == _T_221[11:0] ? image_395 : _GEN_21968; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21970 = 12'h18c == _T_221[11:0] ? image_396 : _GEN_21969; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21971 = 12'h18d == _T_221[11:0] ? image_397 : _GEN_21970; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21972 = 12'h18e == _T_221[11:0] ? image_398 : _GEN_21971; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21973 = 12'h18f == _T_221[11:0] ? image_399 : _GEN_21972; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21974 = 12'h190 == _T_221[11:0] ? image_400 : _GEN_21973; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21975 = 12'h191 == _T_221[11:0] ? image_401 : _GEN_21974; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21976 = 12'h192 == _T_221[11:0] ? image_402 : _GEN_21975; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21977 = 12'h193 == _T_221[11:0] ? image_403 : _GEN_21976; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21978 = 12'h194 == _T_221[11:0] ? image_404 : _GEN_21977; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21979 = 12'h195 == _T_221[11:0] ? image_405 : _GEN_21978; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21980 = 12'h196 == _T_221[11:0] ? image_406 : _GEN_21979; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21981 = 12'h197 == _T_221[11:0] ? image_407 : _GEN_21980; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21982 = 12'h198 == _T_221[11:0] ? image_408 : _GEN_21981; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21983 = 12'h199 == _T_221[11:0] ? image_409 : _GEN_21982; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21984 = 12'h19a == _T_221[11:0] ? image_410 : _GEN_21983; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21985 = 12'h19b == _T_221[11:0] ? image_411 : _GEN_21984; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21986 = 12'h19c == _T_221[11:0] ? image_412 : _GEN_21985; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21987 = 12'h19d == _T_221[11:0] ? image_413 : _GEN_21986; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21988 = 12'h19e == _T_221[11:0] ? image_414 : _GEN_21987; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21989 = 12'h19f == _T_221[11:0] ? image_415 : _GEN_21988; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21990 = 12'h1a0 == _T_221[11:0] ? image_416 : _GEN_21989; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21991 = 12'h1a1 == _T_221[11:0] ? image_417 : _GEN_21990; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21992 = 12'h1a2 == _T_221[11:0] ? image_418 : _GEN_21991; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21993 = 12'h1a3 == _T_221[11:0] ? image_419 : _GEN_21992; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21994 = 12'h1a4 == _T_221[11:0] ? image_420 : _GEN_21993; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21995 = 12'h1a5 == _T_221[11:0] ? image_421 : _GEN_21994; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21996 = 12'h1a6 == _T_221[11:0] ? image_422 : _GEN_21995; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21997 = 12'h1a7 == _T_221[11:0] ? image_423 : _GEN_21996; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21998 = 12'h1a8 == _T_221[11:0] ? image_424 : _GEN_21997; // @[Filter.scala 138:46]
  wire [3:0] _GEN_21999 = 12'h1a9 == _T_221[11:0] ? image_425 : _GEN_21998; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22000 = 12'h1aa == _T_221[11:0] ? image_426 : _GEN_21999; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22001 = 12'h1ab == _T_221[11:0] ? image_427 : _GEN_22000; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22002 = 12'h1ac == _T_221[11:0] ? image_428 : _GEN_22001; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22003 = 12'h1ad == _T_221[11:0] ? image_429 : _GEN_22002; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22004 = 12'h1ae == _T_221[11:0] ? image_430 : _GEN_22003; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22005 = 12'h1af == _T_221[11:0] ? image_431 : _GEN_22004; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22006 = 12'h1b0 == _T_221[11:0] ? image_432 : _GEN_22005; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22007 = 12'h1b1 == _T_221[11:0] ? image_433 : _GEN_22006; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22008 = 12'h1b2 == _T_221[11:0] ? image_434 : _GEN_22007; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22009 = 12'h1b3 == _T_221[11:0] ? image_435 : _GEN_22008; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22010 = 12'h1b4 == _T_221[11:0] ? image_436 : _GEN_22009; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22011 = 12'h1b5 == _T_221[11:0] ? image_437 : _GEN_22010; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22012 = 12'h1b6 == _T_221[11:0] ? image_438 : _GEN_22011; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22013 = 12'h1b7 == _T_221[11:0] ? image_439 : _GEN_22012; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22014 = 12'h1b8 == _T_221[11:0] ? image_440 : _GEN_22013; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22015 = 12'h1b9 == _T_221[11:0] ? image_441 : _GEN_22014; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22016 = 12'h1ba == _T_221[11:0] ? image_442 : _GEN_22015; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22017 = 12'h1bb == _T_221[11:0] ? image_443 : _GEN_22016; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22018 = 12'h1bc == _T_221[11:0] ? image_444 : _GEN_22017; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22019 = 12'h1bd == _T_221[11:0] ? 4'h0 : _GEN_22018; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22020 = 12'h1be == _T_221[11:0] ? 4'h0 : _GEN_22019; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22021 = 12'h1bf == _T_221[11:0] ? 4'h0 : _GEN_22020; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22022 = 12'h1c0 == _T_221[11:0] ? 4'h0 : _GEN_22021; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22023 = 12'h1c1 == _T_221[11:0] ? 4'h0 : _GEN_22022; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22024 = 12'h1c2 == _T_221[11:0] ? 4'h0 : _GEN_22023; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22025 = 12'h1c3 == _T_221[11:0] ? image_451 : _GEN_22024; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22026 = 12'h1c4 == _T_221[11:0] ? image_452 : _GEN_22025; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22027 = 12'h1c5 == _T_221[11:0] ? image_453 : _GEN_22026; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22028 = 12'h1c6 == _T_221[11:0] ? image_454 : _GEN_22027; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22029 = 12'h1c7 == _T_221[11:0] ? image_455 : _GEN_22028; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22030 = 12'h1c8 == _T_221[11:0] ? image_456 : _GEN_22029; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22031 = 12'h1c9 == _T_221[11:0] ? image_457 : _GEN_22030; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22032 = 12'h1ca == _T_221[11:0] ? image_458 : _GEN_22031; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22033 = 12'h1cb == _T_221[11:0] ? image_459 : _GEN_22032; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22034 = 12'h1cc == _T_221[11:0] ? image_460 : _GEN_22033; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22035 = 12'h1cd == _T_221[11:0] ? image_461 : _GEN_22034; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22036 = 12'h1ce == _T_221[11:0] ? image_462 : _GEN_22035; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22037 = 12'h1cf == _T_221[11:0] ? image_463 : _GEN_22036; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22038 = 12'h1d0 == _T_221[11:0] ? image_464 : _GEN_22037; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22039 = 12'h1d1 == _T_221[11:0] ? image_465 : _GEN_22038; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22040 = 12'h1d2 == _T_221[11:0] ? image_466 : _GEN_22039; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22041 = 12'h1d3 == _T_221[11:0] ? image_467 : _GEN_22040; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22042 = 12'h1d4 == _T_221[11:0] ? image_468 : _GEN_22041; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22043 = 12'h1d5 == _T_221[11:0] ? image_469 : _GEN_22042; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22044 = 12'h1d6 == _T_221[11:0] ? image_470 : _GEN_22043; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22045 = 12'h1d7 == _T_221[11:0] ? image_471 : _GEN_22044; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22046 = 12'h1d8 == _T_221[11:0] ? image_472 : _GEN_22045; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22047 = 12'h1d9 == _T_221[11:0] ? image_473 : _GEN_22046; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22048 = 12'h1da == _T_221[11:0] ? image_474 : _GEN_22047; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22049 = 12'h1db == _T_221[11:0] ? image_475 : _GEN_22048; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22050 = 12'h1dc == _T_221[11:0] ? image_476 : _GEN_22049; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22051 = 12'h1dd == _T_221[11:0] ? image_477 : _GEN_22050; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22052 = 12'h1de == _T_221[11:0] ? image_478 : _GEN_22051; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22053 = 12'h1df == _T_221[11:0] ? image_479 : _GEN_22052; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22054 = 12'h1e0 == _T_221[11:0] ? image_480 : _GEN_22053; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22055 = 12'h1e1 == _T_221[11:0] ? image_481 : _GEN_22054; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22056 = 12'h1e2 == _T_221[11:0] ? image_482 : _GEN_22055; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22057 = 12'h1e3 == _T_221[11:0] ? image_483 : _GEN_22056; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22058 = 12'h1e4 == _T_221[11:0] ? image_484 : _GEN_22057; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22059 = 12'h1e5 == _T_221[11:0] ? image_485 : _GEN_22058; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22060 = 12'h1e6 == _T_221[11:0] ? image_486 : _GEN_22059; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22061 = 12'h1e7 == _T_221[11:0] ? image_487 : _GEN_22060; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22062 = 12'h1e8 == _T_221[11:0] ? image_488 : _GEN_22061; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22063 = 12'h1e9 == _T_221[11:0] ? image_489 : _GEN_22062; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22064 = 12'h1ea == _T_221[11:0] ? image_490 : _GEN_22063; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22065 = 12'h1eb == _T_221[11:0] ? image_491 : _GEN_22064; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22066 = 12'h1ec == _T_221[11:0] ? image_492 : _GEN_22065; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22067 = 12'h1ed == _T_221[11:0] ? image_493 : _GEN_22066; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22068 = 12'h1ee == _T_221[11:0] ? image_494 : _GEN_22067; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22069 = 12'h1ef == _T_221[11:0] ? image_495 : _GEN_22068; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22070 = 12'h1f0 == _T_221[11:0] ? image_496 : _GEN_22069; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22071 = 12'h1f1 == _T_221[11:0] ? image_497 : _GEN_22070; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22072 = 12'h1f2 == _T_221[11:0] ? image_498 : _GEN_22071; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22073 = 12'h1f3 == _T_221[11:0] ? image_499 : _GEN_22072; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22074 = 12'h1f4 == _T_221[11:0] ? image_500 : _GEN_22073; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22075 = 12'h1f5 == _T_221[11:0] ? image_501 : _GEN_22074; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22076 = 12'h1f6 == _T_221[11:0] ? image_502 : _GEN_22075; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22077 = 12'h1f7 == _T_221[11:0] ? image_503 : _GEN_22076; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22078 = 12'h1f8 == _T_221[11:0] ? image_504 : _GEN_22077; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22079 = 12'h1f9 == _T_221[11:0] ? image_505 : _GEN_22078; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22080 = 12'h1fa == _T_221[11:0] ? image_506 : _GEN_22079; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22081 = 12'h1fb == _T_221[11:0] ? image_507 : _GEN_22080; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22082 = 12'h1fc == _T_221[11:0] ? image_508 : _GEN_22081; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22083 = 12'h1fd == _T_221[11:0] ? image_509 : _GEN_22082; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22084 = 12'h1fe == _T_221[11:0] ? 4'h0 : _GEN_22083; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22085 = 12'h1ff == _T_221[11:0] ? 4'h0 : _GEN_22084; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22086 = 12'h200 == _T_221[11:0] ? 4'h0 : _GEN_22085; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22087 = 12'h201 == _T_221[11:0] ? 4'h0 : _GEN_22086; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22088 = 12'h202 == _T_221[11:0] ? 4'h0 : _GEN_22087; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22089 = 12'h203 == _T_221[11:0] ? image_515 : _GEN_22088; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22090 = 12'h204 == _T_221[11:0] ? image_516 : _GEN_22089; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22091 = 12'h205 == _T_221[11:0] ? image_517 : _GEN_22090; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22092 = 12'h206 == _T_221[11:0] ? image_518 : _GEN_22091; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22093 = 12'h207 == _T_221[11:0] ? image_519 : _GEN_22092; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22094 = 12'h208 == _T_221[11:0] ? image_520 : _GEN_22093; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22095 = 12'h209 == _T_221[11:0] ? image_521 : _GEN_22094; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22096 = 12'h20a == _T_221[11:0] ? image_522 : _GEN_22095; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22097 = 12'h20b == _T_221[11:0] ? image_523 : _GEN_22096; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22098 = 12'h20c == _T_221[11:0] ? image_524 : _GEN_22097; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22099 = 12'h20d == _T_221[11:0] ? image_525 : _GEN_22098; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22100 = 12'h20e == _T_221[11:0] ? image_526 : _GEN_22099; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22101 = 12'h20f == _T_221[11:0] ? image_527 : _GEN_22100; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22102 = 12'h210 == _T_221[11:0] ? image_528 : _GEN_22101; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22103 = 12'h211 == _T_221[11:0] ? image_529 : _GEN_22102; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22104 = 12'h212 == _T_221[11:0] ? image_530 : _GEN_22103; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22105 = 12'h213 == _T_221[11:0] ? image_531 : _GEN_22104; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22106 = 12'h214 == _T_221[11:0] ? image_532 : _GEN_22105; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22107 = 12'h215 == _T_221[11:0] ? image_533 : _GEN_22106; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22108 = 12'h216 == _T_221[11:0] ? image_534 : _GEN_22107; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22109 = 12'h217 == _T_221[11:0] ? image_535 : _GEN_22108; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22110 = 12'h218 == _T_221[11:0] ? image_536 : _GEN_22109; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22111 = 12'h219 == _T_221[11:0] ? image_537 : _GEN_22110; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22112 = 12'h21a == _T_221[11:0] ? image_538 : _GEN_22111; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22113 = 12'h21b == _T_221[11:0] ? image_539 : _GEN_22112; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22114 = 12'h21c == _T_221[11:0] ? image_540 : _GEN_22113; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22115 = 12'h21d == _T_221[11:0] ? image_541 : _GEN_22114; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22116 = 12'h21e == _T_221[11:0] ? image_542 : _GEN_22115; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22117 = 12'h21f == _T_221[11:0] ? image_543 : _GEN_22116; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22118 = 12'h220 == _T_221[11:0] ? image_544 : _GEN_22117; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22119 = 12'h221 == _T_221[11:0] ? image_545 : _GEN_22118; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22120 = 12'h222 == _T_221[11:0] ? image_546 : _GEN_22119; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22121 = 12'h223 == _T_221[11:0] ? image_547 : _GEN_22120; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22122 = 12'h224 == _T_221[11:0] ? image_548 : _GEN_22121; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22123 = 12'h225 == _T_221[11:0] ? image_549 : _GEN_22122; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22124 = 12'h226 == _T_221[11:0] ? image_550 : _GEN_22123; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22125 = 12'h227 == _T_221[11:0] ? image_551 : _GEN_22124; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22126 = 12'h228 == _T_221[11:0] ? image_552 : _GEN_22125; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22127 = 12'h229 == _T_221[11:0] ? image_553 : _GEN_22126; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22128 = 12'h22a == _T_221[11:0] ? image_554 : _GEN_22127; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22129 = 12'h22b == _T_221[11:0] ? image_555 : _GEN_22128; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22130 = 12'h22c == _T_221[11:0] ? image_556 : _GEN_22129; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22131 = 12'h22d == _T_221[11:0] ? image_557 : _GEN_22130; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22132 = 12'h22e == _T_221[11:0] ? image_558 : _GEN_22131; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22133 = 12'h22f == _T_221[11:0] ? image_559 : _GEN_22132; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22134 = 12'h230 == _T_221[11:0] ? image_560 : _GEN_22133; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22135 = 12'h231 == _T_221[11:0] ? image_561 : _GEN_22134; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22136 = 12'h232 == _T_221[11:0] ? image_562 : _GEN_22135; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22137 = 12'h233 == _T_221[11:0] ? image_563 : _GEN_22136; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22138 = 12'h234 == _T_221[11:0] ? image_564 : _GEN_22137; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22139 = 12'h235 == _T_221[11:0] ? image_565 : _GEN_22138; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22140 = 12'h236 == _T_221[11:0] ? image_566 : _GEN_22139; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22141 = 12'h237 == _T_221[11:0] ? 4'h0 : _GEN_22140; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22142 = 12'h238 == _T_221[11:0] ? 4'h0 : _GEN_22141; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22143 = 12'h239 == _T_221[11:0] ? 4'h0 : _GEN_22142; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22144 = 12'h23a == _T_221[11:0] ? 4'h0 : _GEN_22143; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22145 = 12'h23b == _T_221[11:0] ? image_571 : _GEN_22144; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22146 = 12'h23c == _T_221[11:0] ? image_572 : _GEN_22145; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22147 = 12'h23d == _T_221[11:0] ? image_573 : _GEN_22146; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22148 = 12'h23e == _T_221[11:0] ? image_574 : _GEN_22147; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22149 = 12'h23f == _T_221[11:0] ? 4'h0 : _GEN_22148; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22150 = 12'h240 == _T_221[11:0] ? 4'h0 : _GEN_22149; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22151 = 12'h241 == _T_221[11:0] ? 4'h0 : _GEN_22150; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22152 = 12'h242 == _T_221[11:0] ? image_578 : _GEN_22151; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22153 = 12'h243 == _T_221[11:0] ? image_579 : _GEN_22152; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22154 = 12'h244 == _T_221[11:0] ? image_580 : _GEN_22153; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22155 = 12'h245 == _T_221[11:0] ? image_581 : _GEN_22154; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22156 = 12'h246 == _T_221[11:0] ? image_582 : _GEN_22155; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22157 = 12'h247 == _T_221[11:0] ? image_583 : _GEN_22156; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22158 = 12'h248 == _T_221[11:0] ? image_584 : _GEN_22157; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22159 = 12'h249 == _T_221[11:0] ? image_585 : _GEN_22158; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22160 = 12'h24a == _T_221[11:0] ? image_586 : _GEN_22159; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22161 = 12'h24b == _T_221[11:0] ? image_587 : _GEN_22160; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22162 = 12'h24c == _T_221[11:0] ? image_588 : _GEN_22161; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22163 = 12'h24d == _T_221[11:0] ? image_589 : _GEN_22162; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22164 = 12'h24e == _T_221[11:0] ? image_590 : _GEN_22163; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22165 = 12'h24f == _T_221[11:0] ? image_591 : _GEN_22164; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22166 = 12'h250 == _T_221[11:0] ? image_592 : _GEN_22165; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22167 = 12'h251 == _T_221[11:0] ? image_593 : _GEN_22166; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22168 = 12'h252 == _T_221[11:0] ? image_594 : _GEN_22167; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22169 = 12'h253 == _T_221[11:0] ? image_595 : _GEN_22168; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22170 = 12'h254 == _T_221[11:0] ? image_596 : _GEN_22169; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22171 = 12'h255 == _T_221[11:0] ? image_597 : _GEN_22170; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22172 = 12'h256 == _T_221[11:0] ? image_598 : _GEN_22171; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22173 = 12'h257 == _T_221[11:0] ? image_599 : _GEN_22172; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22174 = 12'h258 == _T_221[11:0] ? image_600 : _GEN_22173; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22175 = 12'h259 == _T_221[11:0] ? image_601 : _GEN_22174; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22176 = 12'h25a == _T_221[11:0] ? image_602 : _GEN_22175; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22177 = 12'h25b == _T_221[11:0] ? image_603 : _GEN_22176; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22178 = 12'h25c == _T_221[11:0] ? image_604 : _GEN_22177; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22179 = 12'h25d == _T_221[11:0] ? image_605 : _GEN_22178; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22180 = 12'h25e == _T_221[11:0] ? image_606 : _GEN_22179; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22181 = 12'h25f == _T_221[11:0] ? image_607 : _GEN_22180; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22182 = 12'h260 == _T_221[11:0] ? 4'h0 : _GEN_22181; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22183 = 12'h261 == _T_221[11:0] ? 4'h0 : _GEN_22182; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22184 = 12'h262 == _T_221[11:0] ? 4'h0 : _GEN_22183; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22185 = 12'h263 == _T_221[11:0] ? 4'h0 : _GEN_22184; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22186 = 12'h264 == _T_221[11:0] ? 4'h0 : _GEN_22185; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22187 = 12'h265 == _T_221[11:0] ? 4'h0 : _GEN_22186; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22188 = 12'h266 == _T_221[11:0] ? image_614 : _GEN_22187; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22189 = 12'h267 == _T_221[11:0] ? image_615 : _GEN_22188; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22190 = 12'h268 == _T_221[11:0] ? image_616 : _GEN_22189; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22191 = 12'h269 == _T_221[11:0] ? image_617 : _GEN_22190; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22192 = 12'h26a == _T_221[11:0] ? image_618 : _GEN_22191; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22193 = 12'h26b == _T_221[11:0] ? image_619 : _GEN_22192; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22194 = 12'h26c == _T_221[11:0] ? image_620 : _GEN_22193; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22195 = 12'h26d == _T_221[11:0] ? image_621 : _GEN_22194; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22196 = 12'h26e == _T_221[11:0] ? image_622 : _GEN_22195; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22197 = 12'h26f == _T_221[11:0] ? image_623 : _GEN_22196; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22198 = 12'h270 == _T_221[11:0] ? image_624 : _GEN_22197; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22199 = 12'h271 == _T_221[11:0] ? image_625 : _GEN_22198; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22200 = 12'h272 == _T_221[11:0] ? image_626 : _GEN_22199; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22201 = 12'h273 == _T_221[11:0] ? image_627 : _GEN_22200; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22202 = 12'h274 == _T_221[11:0] ? image_628 : _GEN_22201; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22203 = 12'h275 == _T_221[11:0] ? 4'h0 : _GEN_22202; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22204 = 12'h276 == _T_221[11:0] ? 4'h0 : _GEN_22203; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22205 = 12'h277 == _T_221[11:0] ? 4'h0 : _GEN_22204; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22206 = 12'h278 == _T_221[11:0] ? 4'h0 : _GEN_22205; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22207 = 12'h279 == _T_221[11:0] ? 4'h0 : _GEN_22206; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22208 = 12'h27a == _T_221[11:0] ? 4'h0 : _GEN_22207; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22209 = 12'h27b == _T_221[11:0] ? 4'h0 : _GEN_22208; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22210 = 12'h27c == _T_221[11:0] ? image_636 : _GEN_22209; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22211 = 12'h27d == _T_221[11:0] ? image_637 : _GEN_22210; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22212 = 12'h27e == _T_221[11:0] ? image_638 : _GEN_22211; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22213 = 12'h27f == _T_221[11:0] ? image_639 : _GEN_22212; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22214 = 12'h280 == _T_221[11:0] ? 4'h0 : _GEN_22213; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22215 = 12'h281 == _T_221[11:0] ? 4'h0 : _GEN_22214; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22216 = 12'h282 == _T_221[11:0] ? image_642 : _GEN_22215; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22217 = 12'h283 == _T_221[11:0] ? image_643 : _GEN_22216; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22218 = 12'h284 == _T_221[11:0] ? image_644 : _GEN_22217; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22219 = 12'h285 == _T_221[11:0] ? image_645 : _GEN_22218; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22220 = 12'h286 == _T_221[11:0] ? image_646 : _GEN_22219; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22221 = 12'h287 == _T_221[11:0] ? image_647 : _GEN_22220; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22222 = 12'h288 == _T_221[11:0] ? image_648 : _GEN_22221; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22223 = 12'h289 == _T_221[11:0] ? image_649 : _GEN_22222; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22224 = 12'h28a == _T_221[11:0] ? image_650 : _GEN_22223; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22225 = 12'h28b == _T_221[11:0] ? image_651 : _GEN_22224; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22226 = 12'h28c == _T_221[11:0] ? image_652 : _GEN_22225; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22227 = 12'h28d == _T_221[11:0] ? image_653 : _GEN_22226; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22228 = 12'h28e == _T_221[11:0] ? image_654 : _GEN_22227; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22229 = 12'h28f == _T_221[11:0] ? image_655 : _GEN_22228; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22230 = 12'h290 == _T_221[11:0] ? image_656 : _GEN_22229; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22231 = 12'h291 == _T_221[11:0] ? image_657 : _GEN_22230; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22232 = 12'h292 == _T_221[11:0] ? image_658 : _GEN_22231; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22233 = 12'h293 == _T_221[11:0] ? image_659 : _GEN_22232; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22234 = 12'h294 == _T_221[11:0] ? image_660 : _GEN_22233; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22235 = 12'h295 == _T_221[11:0] ? image_661 : _GEN_22234; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22236 = 12'h296 == _T_221[11:0] ? image_662 : _GEN_22235; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22237 = 12'h297 == _T_221[11:0] ? image_663 : _GEN_22236; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22238 = 12'h298 == _T_221[11:0] ? image_664 : _GEN_22237; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22239 = 12'h299 == _T_221[11:0] ? image_665 : _GEN_22238; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22240 = 12'h29a == _T_221[11:0] ? image_666 : _GEN_22239; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22241 = 12'h29b == _T_221[11:0] ? image_667 : _GEN_22240; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22242 = 12'h29c == _T_221[11:0] ? image_668 : _GEN_22241; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22243 = 12'h29d == _T_221[11:0] ? image_669 : _GEN_22242; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22244 = 12'h29e == _T_221[11:0] ? image_670 : _GEN_22243; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22245 = 12'h29f == _T_221[11:0] ? 4'h0 : _GEN_22244; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22246 = 12'h2a0 == _T_221[11:0] ? 4'h0 : _GEN_22245; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22247 = 12'h2a1 == _T_221[11:0] ? 4'h0 : _GEN_22246; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22248 = 12'h2a2 == _T_221[11:0] ? 4'h0 : _GEN_22247; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22249 = 12'h2a3 == _T_221[11:0] ? 4'h0 : _GEN_22248; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22250 = 12'h2a4 == _T_221[11:0] ? 4'h0 : _GEN_22249; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22251 = 12'h2a5 == _T_221[11:0] ? 4'h0 : _GEN_22250; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22252 = 12'h2a6 == _T_221[11:0] ? 4'h0 : _GEN_22251; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22253 = 12'h2a7 == _T_221[11:0] ? image_679 : _GEN_22252; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22254 = 12'h2a8 == _T_221[11:0] ? image_680 : _GEN_22253; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22255 = 12'h2a9 == _T_221[11:0] ? image_681 : _GEN_22254; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22256 = 12'h2aa == _T_221[11:0] ? image_682 : _GEN_22255; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22257 = 12'h2ab == _T_221[11:0] ? image_683 : _GEN_22256; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22258 = 12'h2ac == _T_221[11:0] ? image_684 : _GEN_22257; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22259 = 12'h2ad == _T_221[11:0] ? image_685 : _GEN_22258; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22260 = 12'h2ae == _T_221[11:0] ? image_686 : _GEN_22259; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22261 = 12'h2af == _T_221[11:0] ? image_687 : _GEN_22260; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22262 = 12'h2b0 == _T_221[11:0] ? image_688 : _GEN_22261; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22263 = 12'h2b1 == _T_221[11:0] ? image_689 : _GEN_22262; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22264 = 12'h2b2 == _T_221[11:0] ? image_690 : _GEN_22263; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22265 = 12'h2b3 == _T_221[11:0] ? image_691 : _GEN_22264; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22266 = 12'h2b4 == _T_221[11:0] ? image_692 : _GEN_22265; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22267 = 12'h2b5 == _T_221[11:0] ? image_693 : _GEN_22266; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22268 = 12'h2b6 == _T_221[11:0] ? image_694 : _GEN_22267; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22269 = 12'h2b7 == _T_221[11:0] ? image_695 : _GEN_22268; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22270 = 12'h2b8 == _T_221[11:0] ? image_696 : _GEN_22269; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22271 = 12'h2b9 == _T_221[11:0] ? image_697 : _GEN_22270; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22272 = 12'h2ba == _T_221[11:0] ? image_698 : _GEN_22271; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22273 = 12'h2bb == _T_221[11:0] ? 4'h0 : _GEN_22272; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22274 = 12'h2bc == _T_221[11:0] ? 4'h0 : _GEN_22273; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22275 = 12'h2bd == _T_221[11:0] ? image_701 : _GEN_22274; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22276 = 12'h2be == _T_221[11:0] ? image_702 : _GEN_22275; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22277 = 12'h2bf == _T_221[11:0] ? image_703 : _GEN_22276; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22278 = 12'h2c0 == _T_221[11:0] ? 4'h0 : _GEN_22277; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22279 = 12'h2c1 == _T_221[11:0] ? image_705 : _GEN_22278; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22280 = 12'h2c2 == _T_221[11:0] ? image_706 : _GEN_22279; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22281 = 12'h2c3 == _T_221[11:0] ? image_707 : _GEN_22280; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22282 = 12'h2c4 == _T_221[11:0] ? image_708 : _GEN_22281; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22283 = 12'h2c5 == _T_221[11:0] ? image_709 : _GEN_22282; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22284 = 12'h2c6 == _T_221[11:0] ? image_710 : _GEN_22283; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22285 = 12'h2c7 == _T_221[11:0] ? image_711 : _GEN_22284; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22286 = 12'h2c8 == _T_221[11:0] ? image_712 : _GEN_22285; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22287 = 12'h2c9 == _T_221[11:0] ? image_713 : _GEN_22286; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22288 = 12'h2ca == _T_221[11:0] ? image_714 : _GEN_22287; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22289 = 12'h2cb == _T_221[11:0] ? image_715 : _GEN_22288; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22290 = 12'h2cc == _T_221[11:0] ? image_716 : _GEN_22289; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22291 = 12'h2cd == _T_221[11:0] ? image_717 : _GEN_22290; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22292 = 12'h2ce == _T_221[11:0] ? image_718 : _GEN_22291; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22293 = 12'h2cf == _T_221[11:0] ? image_719 : _GEN_22292; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22294 = 12'h2d0 == _T_221[11:0] ? image_720 : _GEN_22293; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22295 = 12'h2d1 == _T_221[11:0] ? image_721 : _GEN_22294; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22296 = 12'h2d2 == _T_221[11:0] ? image_722 : _GEN_22295; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22297 = 12'h2d3 == _T_221[11:0] ? image_723 : _GEN_22296; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22298 = 12'h2d4 == _T_221[11:0] ? image_724 : _GEN_22297; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22299 = 12'h2d5 == _T_221[11:0] ? image_725 : _GEN_22298; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22300 = 12'h2d6 == _T_221[11:0] ? image_726 : _GEN_22299; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22301 = 12'h2d7 == _T_221[11:0] ? image_727 : _GEN_22300; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22302 = 12'h2d8 == _T_221[11:0] ? image_728 : _GEN_22301; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22303 = 12'h2d9 == _T_221[11:0] ? image_729 : _GEN_22302; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22304 = 12'h2da == _T_221[11:0] ? image_730 : _GEN_22303; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22305 = 12'h2db == _T_221[11:0] ? image_731 : _GEN_22304; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22306 = 12'h2dc == _T_221[11:0] ? image_732 : _GEN_22305; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22307 = 12'h2dd == _T_221[11:0] ? image_733 : _GEN_22306; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22308 = 12'h2de == _T_221[11:0] ? image_734 : _GEN_22307; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22309 = 12'h2df == _T_221[11:0] ? 4'h0 : _GEN_22308; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22310 = 12'h2e0 == _T_221[11:0] ? image_736 : _GEN_22309; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22311 = 12'h2e1 == _T_221[11:0] ? image_737 : _GEN_22310; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22312 = 12'h2e2 == _T_221[11:0] ? 4'h0 : _GEN_22311; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22313 = 12'h2e3 == _T_221[11:0] ? image_739 : _GEN_22312; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22314 = 12'h2e4 == _T_221[11:0] ? image_740 : _GEN_22313; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22315 = 12'h2e5 == _T_221[11:0] ? image_741 : _GEN_22314; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22316 = 12'h2e6 == _T_221[11:0] ? 4'h0 : _GEN_22315; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22317 = 12'h2e7 == _T_221[11:0] ? 4'h0 : _GEN_22316; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22318 = 12'h2e8 == _T_221[11:0] ? image_744 : _GEN_22317; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22319 = 12'h2e9 == _T_221[11:0] ? image_745 : _GEN_22318; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22320 = 12'h2ea == _T_221[11:0] ? image_746 : _GEN_22319; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22321 = 12'h2eb == _T_221[11:0] ? image_747 : _GEN_22320; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22322 = 12'h2ec == _T_221[11:0] ? image_748 : _GEN_22321; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22323 = 12'h2ed == _T_221[11:0] ? image_749 : _GEN_22322; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22324 = 12'h2ee == _T_221[11:0] ? image_750 : _GEN_22323; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22325 = 12'h2ef == _T_221[11:0] ? image_751 : _GEN_22324; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22326 = 12'h2f0 == _T_221[11:0] ? image_752 : _GEN_22325; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22327 = 12'h2f1 == _T_221[11:0] ? image_753 : _GEN_22326; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22328 = 12'h2f2 == _T_221[11:0] ? image_754 : _GEN_22327; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22329 = 12'h2f3 == _T_221[11:0] ? image_755 : _GEN_22328; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22330 = 12'h2f4 == _T_221[11:0] ? image_756 : _GEN_22329; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22331 = 12'h2f5 == _T_221[11:0] ? 4'h0 : _GEN_22330; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22332 = 12'h2f6 == _T_221[11:0] ? image_758 : _GEN_22331; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22333 = 12'h2f7 == _T_221[11:0] ? 4'h0 : _GEN_22332; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22334 = 12'h2f8 == _T_221[11:0] ? image_760 : _GEN_22333; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22335 = 12'h2f9 == _T_221[11:0] ? image_761 : _GEN_22334; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22336 = 12'h2fa == _T_221[11:0] ? image_762 : _GEN_22335; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22337 = 12'h2fb == _T_221[11:0] ? image_763 : _GEN_22336; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22338 = 12'h2fc == _T_221[11:0] ? 4'h0 : _GEN_22337; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22339 = 12'h2fd == _T_221[11:0] ? image_765 : _GEN_22338; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22340 = 12'h2fe == _T_221[11:0] ? image_766 : _GEN_22339; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22341 = 12'h2ff == _T_221[11:0] ? image_767 : _GEN_22340; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22342 = 12'h300 == _T_221[11:0] ? image_768 : _GEN_22341; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22343 = 12'h301 == _T_221[11:0] ? image_769 : _GEN_22342; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22344 = 12'h302 == _T_221[11:0] ? image_770 : _GEN_22343; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22345 = 12'h303 == _T_221[11:0] ? image_771 : _GEN_22344; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22346 = 12'h304 == _T_221[11:0] ? image_772 : _GEN_22345; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22347 = 12'h305 == _T_221[11:0] ? image_773 : _GEN_22346; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22348 = 12'h306 == _T_221[11:0] ? image_774 : _GEN_22347; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22349 = 12'h307 == _T_221[11:0] ? image_775 : _GEN_22348; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22350 = 12'h308 == _T_221[11:0] ? image_776 : _GEN_22349; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22351 = 12'h309 == _T_221[11:0] ? image_777 : _GEN_22350; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22352 = 12'h30a == _T_221[11:0] ? image_778 : _GEN_22351; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22353 = 12'h30b == _T_221[11:0] ? image_779 : _GEN_22352; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22354 = 12'h30c == _T_221[11:0] ? image_780 : _GEN_22353; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22355 = 12'h30d == _T_221[11:0] ? image_781 : _GEN_22354; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22356 = 12'h30e == _T_221[11:0] ? image_782 : _GEN_22355; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22357 = 12'h30f == _T_221[11:0] ? image_783 : _GEN_22356; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22358 = 12'h310 == _T_221[11:0] ? image_784 : _GEN_22357; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22359 = 12'h311 == _T_221[11:0] ? image_785 : _GEN_22358; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22360 = 12'h312 == _T_221[11:0] ? image_786 : _GEN_22359; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22361 = 12'h313 == _T_221[11:0] ? image_787 : _GEN_22360; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22362 = 12'h314 == _T_221[11:0] ? image_788 : _GEN_22361; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22363 = 12'h315 == _T_221[11:0] ? image_789 : _GEN_22362; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22364 = 12'h316 == _T_221[11:0] ? image_790 : _GEN_22363; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22365 = 12'h317 == _T_221[11:0] ? image_791 : _GEN_22364; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22366 = 12'h318 == _T_221[11:0] ? image_792 : _GEN_22365; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22367 = 12'h319 == _T_221[11:0] ? image_793 : _GEN_22366; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22368 = 12'h31a == _T_221[11:0] ? image_794 : _GEN_22367; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22369 = 12'h31b == _T_221[11:0] ? image_795 : _GEN_22368; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22370 = 12'h31c == _T_221[11:0] ? image_796 : _GEN_22369; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22371 = 12'h31d == _T_221[11:0] ? image_797 : _GEN_22370; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22372 = 12'h31e == _T_221[11:0] ? 4'h0 : _GEN_22371; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22373 = 12'h31f == _T_221[11:0] ? 4'h0 : _GEN_22372; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22374 = 12'h320 == _T_221[11:0] ? image_800 : _GEN_22373; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22375 = 12'h321 == _T_221[11:0] ? image_801 : _GEN_22374; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22376 = 12'h322 == _T_221[11:0] ? image_802 : _GEN_22375; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22377 = 12'h323 == _T_221[11:0] ? image_803 : _GEN_22376; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22378 = 12'h324 == _T_221[11:0] ? image_804 : _GEN_22377; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22379 = 12'h325 == _T_221[11:0] ? image_805 : _GEN_22378; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22380 = 12'h326 == _T_221[11:0] ? image_806 : _GEN_22379; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22381 = 12'h327 == _T_221[11:0] ? 4'h0 : _GEN_22380; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22382 = 12'h328 == _T_221[11:0] ? image_808 : _GEN_22381; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22383 = 12'h329 == _T_221[11:0] ? image_809 : _GEN_22382; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22384 = 12'h32a == _T_221[11:0] ? image_810 : _GEN_22383; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22385 = 12'h32b == _T_221[11:0] ? image_811 : _GEN_22384; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22386 = 12'h32c == _T_221[11:0] ? image_812 : _GEN_22385; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22387 = 12'h32d == _T_221[11:0] ? image_813 : _GEN_22386; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22388 = 12'h32e == _T_221[11:0] ? image_814 : _GEN_22387; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22389 = 12'h32f == _T_221[11:0] ? image_815 : _GEN_22388; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22390 = 12'h330 == _T_221[11:0] ? image_816 : _GEN_22389; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22391 = 12'h331 == _T_221[11:0] ? image_817 : _GEN_22390; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22392 = 12'h332 == _T_221[11:0] ? image_818 : _GEN_22391; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22393 = 12'h333 == _T_221[11:0] ? image_819 : _GEN_22392; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22394 = 12'h334 == _T_221[11:0] ? image_820 : _GEN_22393; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22395 = 12'h335 == _T_221[11:0] ? 4'h0 : _GEN_22394; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22396 = 12'h336 == _T_221[11:0] ? image_822 : _GEN_22395; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22397 = 12'h337 == _T_221[11:0] ? image_823 : _GEN_22396; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22398 = 12'h338 == _T_221[11:0] ? image_824 : _GEN_22397; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22399 = 12'h339 == _T_221[11:0] ? image_825 : _GEN_22398; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22400 = 12'h33a == _T_221[11:0] ? image_826 : _GEN_22399; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22401 = 12'h33b == _T_221[11:0] ? 4'h0 : _GEN_22400; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22402 = 12'h33c == _T_221[11:0] ? image_828 : _GEN_22401; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22403 = 12'h33d == _T_221[11:0] ? image_829 : _GEN_22402; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22404 = 12'h33e == _T_221[11:0] ? image_830 : _GEN_22403; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22405 = 12'h33f == _T_221[11:0] ? image_831 : _GEN_22404; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22406 = 12'h340 == _T_221[11:0] ? 4'h0 : _GEN_22405; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22407 = 12'h341 == _T_221[11:0] ? image_833 : _GEN_22406; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22408 = 12'h342 == _T_221[11:0] ? image_834 : _GEN_22407; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22409 = 12'h343 == _T_221[11:0] ? image_835 : _GEN_22408; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22410 = 12'h344 == _T_221[11:0] ? image_836 : _GEN_22409; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22411 = 12'h345 == _T_221[11:0] ? image_837 : _GEN_22410; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22412 = 12'h346 == _T_221[11:0] ? image_838 : _GEN_22411; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22413 = 12'h347 == _T_221[11:0] ? image_839 : _GEN_22412; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22414 = 12'h348 == _T_221[11:0] ? image_840 : _GEN_22413; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22415 = 12'h349 == _T_221[11:0] ? image_841 : _GEN_22414; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22416 = 12'h34a == _T_221[11:0] ? image_842 : _GEN_22415; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22417 = 12'h34b == _T_221[11:0] ? image_843 : _GEN_22416; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22418 = 12'h34c == _T_221[11:0] ? image_844 : _GEN_22417; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22419 = 12'h34d == _T_221[11:0] ? image_845 : _GEN_22418; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22420 = 12'h34e == _T_221[11:0] ? image_846 : _GEN_22419; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22421 = 12'h34f == _T_221[11:0] ? image_847 : _GEN_22420; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22422 = 12'h350 == _T_221[11:0] ? image_848 : _GEN_22421; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22423 = 12'h351 == _T_221[11:0] ? image_849 : _GEN_22422; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22424 = 12'h352 == _T_221[11:0] ? image_850 : _GEN_22423; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22425 = 12'h353 == _T_221[11:0] ? image_851 : _GEN_22424; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22426 = 12'h354 == _T_221[11:0] ? image_852 : _GEN_22425; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22427 = 12'h355 == _T_221[11:0] ? image_853 : _GEN_22426; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22428 = 12'h356 == _T_221[11:0] ? image_854 : _GEN_22427; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22429 = 12'h357 == _T_221[11:0] ? image_855 : _GEN_22428; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22430 = 12'h358 == _T_221[11:0] ? image_856 : _GEN_22429; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22431 = 12'h359 == _T_221[11:0] ? image_857 : _GEN_22430; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22432 = 12'h35a == _T_221[11:0] ? image_858 : _GEN_22431; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22433 = 12'h35b == _T_221[11:0] ? image_859 : _GEN_22432; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22434 = 12'h35c == _T_221[11:0] ? image_860 : _GEN_22433; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22435 = 12'h35d == _T_221[11:0] ? image_861 : _GEN_22434; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22436 = 12'h35e == _T_221[11:0] ? image_862 : _GEN_22435; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22437 = 12'h35f == _T_221[11:0] ? 4'h0 : _GEN_22436; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22438 = 12'h360 == _T_221[11:0] ? 4'h0 : _GEN_22437; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22439 = 12'h361 == _T_221[11:0] ? image_865 : _GEN_22438; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22440 = 12'h362 == _T_221[11:0] ? image_866 : _GEN_22439; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22441 = 12'h363 == _T_221[11:0] ? image_867 : _GEN_22440; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22442 = 12'h364 == _T_221[11:0] ? image_868 : _GEN_22441; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22443 = 12'h365 == _T_221[11:0] ? image_869 : _GEN_22442; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22444 = 12'h366 == _T_221[11:0] ? 4'h0 : _GEN_22443; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22445 = 12'h367 == _T_221[11:0] ? 4'h0 : _GEN_22444; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22446 = 12'h368 == _T_221[11:0] ? image_872 : _GEN_22445; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22447 = 12'h369 == _T_221[11:0] ? image_873 : _GEN_22446; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22448 = 12'h36a == _T_221[11:0] ? image_874 : _GEN_22447; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22449 = 12'h36b == _T_221[11:0] ? image_875 : _GEN_22448; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22450 = 12'h36c == _T_221[11:0] ? image_876 : _GEN_22449; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22451 = 12'h36d == _T_221[11:0] ? image_877 : _GEN_22450; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22452 = 12'h36e == _T_221[11:0] ? image_878 : _GEN_22451; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22453 = 12'h36f == _T_221[11:0] ? image_879 : _GEN_22452; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22454 = 12'h370 == _T_221[11:0] ? image_880 : _GEN_22453; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22455 = 12'h371 == _T_221[11:0] ? image_881 : _GEN_22454; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22456 = 12'h372 == _T_221[11:0] ? image_882 : _GEN_22455; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22457 = 12'h373 == _T_221[11:0] ? image_883 : _GEN_22456; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22458 = 12'h374 == _T_221[11:0] ? image_884 : _GEN_22457; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22459 = 12'h375 == _T_221[11:0] ? image_885 : _GEN_22458; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22460 = 12'h376 == _T_221[11:0] ? 4'h0 : _GEN_22459; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22461 = 12'h377 == _T_221[11:0] ? 4'h0 : _GEN_22460; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22462 = 12'h378 == _T_221[11:0] ? 4'h0 : _GEN_22461; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22463 = 12'h379 == _T_221[11:0] ? 4'h0 : _GEN_22462; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22464 = 12'h37a == _T_221[11:0] ? 4'h0 : _GEN_22463; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22465 = 12'h37b == _T_221[11:0] ? image_891 : _GEN_22464; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22466 = 12'h37c == _T_221[11:0] ? image_892 : _GEN_22465; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22467 = 12'h37d == _T_221[11:0] ? image_893 : _GEN_22466; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22468 = 12'h37e == _T_221[11:0] ? image_894 : _GEN_22467; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22469 = 12'h37f == _T_221[11:0] ? image_895 : _GEN_22468; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22470 = 12'h380 == _T_221[11:0] ? 4'h0 : _GEN_22469; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22471 = 12'h381 == _T_221[11:0] ? image_897 : _GEN_22470; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22472 = 12'h382 == _T_221[11:0] ? image_898 : _GEN_22471; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22473 = 12'h383 == _T_221[11:0] ? image_899 : _GEN_22472; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22474 = 12'h384 == _T_221[11:0] ? image_900 : _GEN_22473; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22475 = 12'h385 == _T_221[11:0] ? image_901 : _GEN_22474; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22476 = 12'h386 == _T_221[11:0] ? image_902 : _GEN_22475; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22477 = 12'h387 == _T_221[11:0] ? image_903 : _GEN_22476; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22478 = 12'h388 == _T_221[11:0] ? image_904 : _GEN_22477; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22479 = 12'h389 == _T_221[11:0] ? image_905 : _GEN_22478; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22480 = 12'h38a == _T_221[11:0] ? image_906 : _GEN_22479; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22481 = 12'h38b == _T_221[11:0] ? image_907 : _GEN_22480; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22482 = 12'h38c == _T_221[11:0] ? image_908 : _GEN_22481; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22483 = 12'h38d == _T_221[11:0] ? image_909 : _GEN_22482; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22484 = 12'h38e == _T_221[11:0] ? image_910 : _GEN_22483; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22485 = 12'h38f == _T_221[11:0] ? image_911 : _GEN_22484; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22486 = 12'h390 == _T_221[11:0] ? image_912 : _GEN_22485; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22487 = 12'h391 == _T_221[11:0] ? image_913 : _GEN_22486; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22488 = 12'h392 == _T_221[11:0] ? image_914 : _GEN_22487; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22489 = 12'h393 == _T_221[11:0] ? image_915 : _GEN_22488; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22490 = 12'h394 == _T_221[11:0] ? image_916 : _GEN_22489; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22491 = 12'h395 == _T_221[11:0] ? image_917 : _GEN_22490; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22492 = 12'h396 == _T_221[11:0] ? image_918 : _GEN_22491; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22493 = 12'h397 == _T_221[11:0] ? image_919 : _GEN_22492; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22494 = 12'h398 == _T_221[11:0] ? image_920 : _GEN_22493; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22495 = 12'h399 == _T_221[11:0] ? image_921 : _GEN_22494; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22496 = 12'h39a == _T_221[11:0] ? image_922 : _GEN_22495; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22497 = 12'h39b == _T_221[11:0] ? image_923 : _GEN_22496; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22498 = 12'h39c == _T_221[11:0] ? image_924 : _GEN_22497; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22499 = 12'h39d == _T_221[11:0] ? image_925 : _GEN_22498; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22500 = 12'h39e == _T_221[11:0] ? image_926 : _GEN_22499; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22501 = 12'h39f == _T_221[11:0] ? image_927 : _GEN_22500; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22502 = 12'h3a0 == _T_221[11:0] ? 4'h0 : _GEN_22501; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22503 = 12'h3a1 == _T_221[11:0] ? image_929 : _GEN_22502; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22504 = 12'h3a2 == _T_221[11:0] ? image_930 : _GEN_22503; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22505 = 12'h3a3 == _T_221[11:0] ? 4'h0 : _GEN_22504; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22506 = 12'h3a4 == _T_221[11:0] ? 4'h0 : _GEN_22505; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22507 = 12'h3a5 == _T_221[11:0] ? 4'h0 : _GEN_22506; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22508 = 12'h3a6 == _T_221[11:0] ? 4'h0 : _GEN_22507; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22509 = 12'h3a7 == _T_221[11:0] ? image_935 : _GEN_22508; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22510 = 12'h3a8 == _T_221[11:0] ? image_936 : _GEN_22509; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22511 = 12'h3a9 == _T_221[11:0] ? image_937 : _GEN_22510; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22512 = 12'h3aa == _T_221[11:0] ? image_938 : _GEN_22511; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22513 = 12'h3ab == _T_221[11:0] ? image_939 : _GEN_22512; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22514 = 12'h3ac == _T_221[11:0] ? image_940 : _GEN_22513; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22515 = 12'h3ad == _T_221[11:0] ? image_941 : _GEN_22514; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22516 = 12'h3ae == _T_221[11:0] ? image_942 : _GEN_22515; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22517 = 12'h3af == _T_221[11:0] ? image_943 : _GEN_22516; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22518 = 12'h3b0 == _T_221[11:0] ? image_944 : _GEN_22517; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22519 = 12'h3b1 == _T_221[11:0] ? image_945 : _GEN_22518; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22520 = 12'h3b2 == _T_221[11:0] ? image_946 : _GEN_22519; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22521 = 12'h3b3 == _T_221[11:0] ? image_947 : _GEN_22520; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22522 = 12'h3b4 == _T_221[11:0] ? image_948 : _GEN_22521; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22523 = 12'h3b5 == _T_221[11:0] ? image_949 : _GEN_22522; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22524 = 12'h3b6 == _T_221[11:0] ? image_950 : _GEN_22523; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22525 = 12'h3b7 == _T_221[11:0] ? image_951 : _GEN_22524; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22526 = 12'h3b8 == _T_221[11:0] ? image_952 : _GEN_22525; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22527 = 12'h3b9 == _T_221[11:0] ? image_953 : _GEN_22526; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22528 = 12'h3ba == _T_221[11:0] ? image_954 : _GEN_22527; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22529 = 12'h3bb == _T_221[11:0] ? image_955 : _GEN_22528; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22530 = 12'h3bc == _T_221[11:0] ? image_956 : _GEN_22529; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22531 = 12'h3bd == _T_221[11:0] ? image_957 : _GEN_22530; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22532 = 12'h3be == _T_221[11:0] ? image_958 : _GEN_22531; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22533 = 12'h3bf == _T_221[11:0] ? image_959 : _GEN_22532; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22534 = 12'h3c0 == _T_221[11:0] ? 4'h0 : _GEN_22533; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22535 = 12'h3c1 == _T_221[11:0] ? image_961 : _GEN_22534; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22536 = 12'h3c2 == _T_221[11:0] ? image_962 : _GEN_22535; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22537 = 12'h3c3 == _T_221[11:0] ? image_963 : _GEN_22536; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22538 = 12'h3c4 == _T_221[11:0] ? image_964 : _GEN_22537; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22539 = 12'h3c5 == _T_221[11:0] ? image_965 : _GEN_22538; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22540 = 12'h3c6 == _T_221[11:0] ? image_966 : _GEN_22539; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22541 = 12'h3c7 == _T_221[11:0] ? image_967 : _GEN_22540; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22542 = 12'h3c8 == _T_221[11:0] ? image_968 : _GEN_22541; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22543 = 12'h3c9 == _T_221[11:0] ? image_969 : _GEN_22542; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22544 = 12'h3ca == _T_221[11:0] ? image_970 : _GEN_22543; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22545 = 12'h3cb == _T_221[11:0] ? image_971 : _GEN_22544; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22546 = 12'h3cc == _T_221[11:0] ? image_972 : _GEN_22545; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22547 = 12'h3cd == _T_221[11:0] ? image_973 : _GEN_22546; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22548 = 12'h3ce == _T_221[11:0] ? image_974 : _GEN_22547; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22549 = 12'h3cf == _T_221[11:0] ? image_975 : _GEN_22548; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22550 = 12'h3d0 == _T_221[11:0] ? image_976 : _GEN_22549; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22551 = 12'h3d1 == _T_221[11:0] ? image_977 : _GEN_22550; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22552 = 12'h3d2 == _T_221[11:0] ? image_978 : _GEN_22551; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22553 = 12'h3d3 == _T_221[11:0] ? image_979 : _GEN_22552; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22554 = 12'h3d4 == _T_221[11:0] ? image_980 : _GEN_22553; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22555 = 12'h3d5 == _T_221[11:0] ? image_981 : _GEN_22554; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22556 = 12'h3d6 == _T_221[11:0] ? image_982 : _GEN_22555; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22557 = 12'h3d7 == _T_221[11:0] ? image_983 : _GEN_22556; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22558 = 12'h3d8 == _T_221[11:0] ? image_984 : _GEN_22557; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22559 = 12'h3d9 == _T_221[11:0] ? image_985 : _GEN_22558; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22560 = 12'h3da == _T_221[11:0] ? image_986 : _GEN_22559; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22561 = 12'h3db == _T_221[11:0] ? image_987 : _GEN_22560; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22562 = 12'h3dc == _T_221[11:0] ? image_988 : _GEN_22561; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22563 = 12'h3dd == _T_221[11:0] ? image_989 : _GEN_22562; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22564 = 12'h3de == _T_221[11:0] ? image_990 : _GEN_22563; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22565 = 12'h3df == _T_221[11:0] ? image_991 : _GEN_22564; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22566 = 12'h3e0 == _T_221[11:0] ? image_992 : _GEN_22565; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22567 = 12'h3e1 == _T_221[11:0] ? 4'h0 : _GEN_22566; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22568 = 12'h3e2 == _T_221[11:0] ? 4'h0 : _GEN_22567; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22569 = 12'h3e3 == _T_221[11:0] ? 4'h0 : _GEN_22568; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22570 = 12'h3e4 == _T_221[11:0] ? 4'h0 : _GEN_22569; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22571 = 12'h3e5 == _T_221[11:0] ? image_997 : _GEN_22570; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22572 = 12'h3e6 == _T_221[11:0] ? image_998 : _GEN_22571; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22573 = 12'h3e7 == _T_221[11:0] ? image_999 : _GEN_22572; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22574 = 12'h3e8 == _T_221[11:0] ? image_1000 : _GEN_22573; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22575 = 12'h3e9 == _T_221[11:0] ? image_1001 : _GEN_22574; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22576 = 12'h3ea == _T_221[11:0] ? image_1002 : _GEN_22575; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22577 = 12'h3eb == _T_221[11:0] ? image_1003 : _GEN_22576; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22578 = 12'h3ec == _T_221[11:0] ? image_1004 : _GEN_22577; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22579 = 12'h3ed == _T_221[11:0] ? image_1005 : _GEN_22578; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22580 = 12'h3ee == _T_221[11:0] ? image_1006 : _GEN_22579; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22581 = 12'h3ef == _T_221[11:0] ? image_1007 : _GEN_22580; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22582 = 12'h3f0 == _T_221[11:0] ? image_1008 : _GEN_22581; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22583 = 12'h3f1 == _T_221[11:0] ? image_1009 : _GEN_22582; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22584 = 12'h3f2 == _T_221[11:0] ? image_1010 : _GEN_22583; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22585 = 12'h3f3 == _T_221[11:0] ? image_1011 : _GEN_22584; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22586 = 12'h3f4 == _T_221[11:0] ? image_1012 : _GEN_22585; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22587 = 12'h3f5 == _T_221[11:0] ? image_1013 : _GEN_22586; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22588 = 12'h3f6 == _T_221[11:0] ? image_1014 : _GEN_22587; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22589 = 12'h3f7 == _T_221[11:0] ? image_1015 : _GEN_22588; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22590 = 12'h3f8 == _T_221[11:0] ? image_1016 : _GEN_22589; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22591 = 12'h3f9 == _T_221[11:0] ? image_1017 : _GEN_22590; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22592 = 12'h3fa == _T_221[11:0] ? image_1018 : _GEN_22591; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22593 = 12'h3fb == _T_221[11:0] ? image_1019 : _GEN_22592; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22594 = 12'h3fc == _T_221[11:0] ? image_1020 : _GEN_22593; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22595 = 12'h3fd == _T_221[11:0] ? 4'h0 : _GEN_22594; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22596 = 12'h3fe == _T_221[11:0] ? 4'h0 : _GEN_22595; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22597 = 12'h3ff == _T_221[11:0] ? 4'h0 : _GEN_22596; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22598 = 12'h400 == _T_221[11:0] ? image_1024 : _GEN_22597; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22599 = 12'h401 == _T_221[11:0] ? image_1025 : _GEN_22598; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22600 = 12'h402 == _T_221[11:0] ? image_1026 : _GEN_22599; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22601 = 12'h403 == _T_221[11:0] ? image_1027 : _GEN_22600; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22602 = 12'h404 == _T_221[11:0] ? image_1028 : _GEN_22601; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22603 = 12'h405 == _T_221[11:0] ? image_1029 : _GEN_22602; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22604 = 12'h406 == _T_221[11:0] ? image_1030 : _GEN_22603; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22605 = 12'h407 == _T_221[11:0] ? image_1031 : _GEN_22604; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22606 = 12'h408 == _T_221[11:0] ? image_1032 : _GEN_22605; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22607 = 12'h409 == _T_221[11:0] ? image_1033 : _GEN_22606; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22608 = 12'h40a == _T_221[11:0] ? image_1034 : _GEN_22607; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22609 = 12'h40b == _T_221[11:0] ? image_1035 : _GEN_22608; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22610 = 12'h40c == _T_221[11:0] ? image_1036 : _GEN_22609; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22611 = 12'h40d == _T_221[11:0] ? image_1037 : _GEN_22610; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22612 = 12'h40e == _T_221[11:0] ? image_1038 : _GEN_22611; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22613 = 12'h40f == _T_221[11:0] ? image_1039 : _GEN_22612; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22614 = 12'h410 == _T_221[11:0] ? image_1040 : _GEN_22613; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22615 = 12'h411 == _T_221[11:0] ? image_1041 : _GEN_22614; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22616 = 12'h412 == _T_221[11:0] ? image_1042 : _GEN_22615; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22617 = 12'h413 == _T_221[11:0] ? image_1043 : _GEN_22616; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22618 = 12'h414 == _T_221[11:0] ? image_1044 : _GEN_22617; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22619 = 12'h415 == _T_221[11:0] ? image_1045 : _GEN_22618; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22620 = 12'h416 == _T_221[11:0] ? image_1046 : _GEN_22619; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22621 = 12'h417 == _T_221[11:0] ? image_1047 : _GEN_22620; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22622 = 12'h418 == _T_221[11:0] ? image_1048 : _GEN_22621; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22623 = 12'h419 == _T_221[11:0] ? image_1049 : _GEN_22622; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22624 = 12'h41a == _T_221[11:0] ? image_1050 : _GEN_22623; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22625 = 12'h41b == _T_221[11:0] ? image_1051 : _GEN_22624; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22626 = 12'h41c == _T_221[11:0] ? image_1052 : _GEN_22625; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22627 = 12'h41d == _T_221[11:0] ? image_1053 : _GEN_22626; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22628 = 12'h41e == _T_221[11:0] ? image_1054 : _GEN_22627; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22629 = 12'h41f == _T_221[11:0] ? image_1055 : _GEN_22628; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22630 = 12'h420 == _T_221[11:0] ? image_1056 : _GEN_22629; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22631 = 12'h421 == _T_221[11:0] ? image_1057 : _GEN_22630; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22632 = 12'h422 == _T_221[11:0] ? image_1058 : _GEN_22631; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22633 = 12'h423 == _T_221[11:0] ? image_1059 : _GEN_22632; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22634 = 12'h424 == _T_221[11:0] ? image_1060 : _GEN_22633; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22635 = 12'h425 == _T_221[11:0] ? image_1061 : _GEN_22634; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22636 = 12'h426 == _T_221[11:0] ? image_1062 : _GEN_22635; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22637 = 12'h427 == _T_221[11:0] ? image_1063 : _GEN_22636; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22638 = 12'h428 == _T_221[11:0] ? image_1064 : _GEN_22637; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22639 = 12'h429 == _T_221[11:0] ? image_1065 : _GEN_22638; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22640 = 12'h42a == _T_221[11:0] ? image_1066 : _GEN_22639; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22641 = 12'h42b == _T_221[11:0] ? image_1067 : _GEN_22640; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22642 = 12'h42c == _T_221[11:0] ? image_1068 : _GEN_22641; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22643 = 12'h42d == _T_221[11:0] ? image_1069 : _GEN_22642; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22644 = 12'h42e == _T_221[11:0] ? image_1070 : _GEN_22643; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22645 = 12'h42f == _T_221[11:0] ? image_1071 : _GEN_22644; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22646 = 12'h430 == _T_221[11:0] ? image_1072 : _GEN_22645; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22647 = 12'h431 == _T_221[11:0] ? image_1073 : _GEN_22646; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22648 = 12'h432 == _T_221[11:0] ? image_1074 : _GEN_22647; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22649 = 12'h433 == _T_221[11:0] ? image_1075 : _GEN_22648; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22650 = 12'h434 == _T_221[11:0] ? image_1076 : _GEN_22649; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22651 = 12'h435 == _T_221[11:0] ? image_1077 : _GEN_22650; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22652 = 12'h436 == _T_221[11:0] ? image_1078 : _GEN_22651; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22653 = 12'h437 == _T_221[11:0] ? image_1079 : _GEN_22652; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22654 = 12'h438 == _T_221[11:0] ? image_1080 : _GEN_22653; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22655 = 12'h439 == _T_221[11:0] ? image_1081 : _GEN_22654; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22656 = 12'h43a == _T_221[11:0] ? image_1082 : _GEN_22655; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22657 = 12'h43b == _T_221[11:0] ? image_1083 : _GEN_22656; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22658 = 12'h43c == _T_221[11:0] ? image_1084 : _GEN_22657; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22659 = 12'h43d == _T_221[11:0] ? image_1085 : _GEN_22658; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22660 = 12'h43e == _T_221[11:0] ? 4'h0 : _GEN_22659; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22661 = 12'h43f == _T_221[11:0] ? 4'h0 : _GEN_22660; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22662 = 12'h440 == _T_221[11:0] ? image_1088 : _GEN_22661; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22663 = 12'h441 == _T_221[11:0] ? image_1089 : _GEN_22662; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22664 = 12'h442 == _T_221[11:0] ? image_1090 : _GEN_22663; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22665 = 12'h443 == _T_221[11:0] ? image_1091 : _GEN_22664; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22666 = 12'h444 == _T_221[11:0] ? image_1092 : _GEN_22665; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22667 = 12'h445 == _T_221[11:0] ? image_1093 : _GEN_22666; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22668 = 12'h446 == _T_221[11:0] ? image_1094 : _GEN_22667; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22669 = 12'h447 == _T_221[11:0] ? image_1095 : _GEN_22668; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22670 = 12'h448 == _T_221[11:0] ? image_1096 : _GEN_22669; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22671 = 12'h449 == _T_221[11:0] ? image_1097 : _GEN_22670; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22672 = 12'h44a == _T_221[11:0] ? image_1098 : _GEN_22671; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22673 = 12'h44b == _T_221[11:0] ? image_1099 : _GEN_22672; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22674 = 12'h44c == _T_221[11:0] ? image_1100 : _GEN_22673; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22675 = 12'h44d == _T_221[11:0] ? image_1101 : _GEN_22674; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22676 = 12'h44e == _T_221[11:0] ? image_1102 : _GEN_22675; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22677 = 12'h44f == _T_221[11:0] ? image_1103 : _GEN_22676; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22678 = 12'h450 == _T_221[11:0] ? image_1104 : _GEN_22677; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22679 = 12'h451 == _T_221[11:0] ? image_1105 : _GEN_22678; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22680 = 12'h452 == _T_221[11:0] ? image_1106 : _GEN_22679; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22681 = 12'h453 == _T_221[11:0] ? image_1107 : _GEN_22680; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22682 = 12'h454 == _T_221[11:0] ? image_1108 : _GEN_22681; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22683 = 12'h455 == _T_221[11:0] ? image_1109 : _GEN_22682; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22684 = 12'h456 == _T_221[11:0] ? image_1110 : _GEN_22683; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22685 = 12'h457 == _T_221[11:0] ? image_1111 : _GEN_22684; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22686 = 12'h458 == _T_221[11:0] ? image_1112 : _GEN_22685; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22687 = 12'h459 == _T_221[11:0] ? image_1113 : _GEN_22686; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22688 = 12'h45a == _T_221[11:0] ? image_1114 : _GEN_22687; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22689 = 12'h45b == _T_221[11:0] ? image_1115 : _GEN_22688; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22690 = 12'h45c == _T_221[11:0] ? image_1116 : _GEN_22689; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22691 = 12'h45d == _T_221[11:0] ? image_1117 : _GEN_22690; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22692 = 12'h45e == _T_221[11:0] ? image_1118 : _GEN_22691; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22693 = 12'h45f == _T_221[11:0] ? image_1119 : _GEN_22692; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22694 = 12'h460 == _T_221[11:0] ? image_1120 : _GEN_22693; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22695 = 12'h461 == _T_221[11:0] ? image_1121 : _GEN_22694; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22696 = 12'h462 == _T_221[11:0] ? image_1122 : _GEN_22695; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22697 = 12'h463 == _T_221[11:0] ? image_1123 : _GEN_22696; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22698 = 12'h464 == _T_221[11:0] ? image_1124 : _GEN_22697; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22699 = 12'h465 == _T_221[11:0] ? image_1125 : _GEN_22698; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22700 = 12'h466 == _T_221[11:0] ? image_1126 : _GEN_22699; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22701 = 12'h467 == _T_221[11:0] ? image_1127 : _GEN_22700; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22702 = 12'h468 == _T_221[11:0] ? image_1128 : _GEN_22701; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22703 = 12'h469 == _T_221[11:0] ? image_1129 : _GEN_22702; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22704 = 12'h46a == _T_221[11:0] ? image_1130 : _GEN_22703; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22705 = 12'h46b == _T_221[11:0] ? image_1131 : _GEN_22704; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22706 = 12'h46c == _T_221[11:0] ? image_1132 : _GEN_22705; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22707 = 12'h46d == _T_221[11:0] ? image_1133 : _GEN_22706; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22708 = 12'h46e == _T_221[11:0] ? image_1134 : _GEN_22707; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22709 = 12'h46f == _T_221[11:0] ? image_1135 : _GEN_22708; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22710 = 12'h470 == _T_221[11:0] ? image_1136 : _GEN_22709; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22711 = 12'h471 == _T_221[11:0] ? image_1137 : _GEN_22710; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22712 = 12'h472 == _T_221[11:0] ? image_1138 : _GEN_22711; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22713 = 12'h473 == _T_221[11:0] ? image_1139 : _GEN_22712; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22714 = 12'h474 == _T_221[11:0] ? image_1140 : _GEN_22713; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22715 = 12'h475 == _T_221[11:0] ? image_1141 : _GEN_22714; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22716 = 12'h476 == _T_221[11:0] ? image_1142 : _GEN_22715; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22717 = 12'h477 == _T_221[11:0] ? image_1143 : _GEN_22716; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22718 = 12'h478 == _T_221[11:0] ? image_1144 : _GEN_22717; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22719 = 12'h479 == _T_221[11:0] ? image_1145 : _GEN_22718; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22720 = 12'h47a == _T_221[11:0] ? image_1146 : _GEN_22719; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22721 = 12'h47b == _T_221[11:0] ? image_1147 : _GEN_22720; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22722 = 12'h47c == _T_221[11:0] ? image_1148 : _GEN_22721; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22723 = 12'h47d == _T_221[11:0] ? 4'h0 : _GEN_22722; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22724 = 12'h47e == _T_221[11:0] ? 4'h0 : _GEN_22723; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22725 = 12'h47f == _T_221[11:0] ? 4'h0 : _GEN_22724; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22726 = 12'h480 == _T_221[11:0] ? image_1152 : _GEN_22725; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22727 = 12'h481 == _T_221[11:0] ? image_1153 : _GEN_22726; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22728 = 12'h482 == _T_221[11:0] ? image_1154 : _GEN_22727; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22729 = 12'h483 == _T_221[11:0] ? image_1155 : _GEN_22728; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22730 = 12'h484 == _T_221[11:0] ? image_1156 : _GEN_22729; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22731 = 12'h485 == _T_221[11:0] ? image_1157 : _GEN_22730; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22732 = 12'h486 == _T_221[11:0] ? image_1158 : _GEN_22731; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22733 = 12'h487 == _T_221[11:0] ? image_1159 : _GEN_22732; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22734 = 12'h488 == _T_221[11:0] ? image_1160 : _GEN_22733; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22735 = 12'h489 == _T_221[11:0] ? image_1161 : _GEN_22734; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22736 = 12'h48a == _T_221[11:0] ? image_1162 : _GEN_22735; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22737 = 12'h48b == _T_221[11:0] ? image_1163 : _GEN_22736; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22738 = 12'h48c == _T_221[11:0] ? image_1164 : _GEN_22737; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22739 = 12'h48d == _T_221[11:0] ? image_1165 : _GEN_22738; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22740 = 12'h48e == _T_221[11:0] ? image_1166 : _GEN_22739; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22741 = 12'h48f == _T_221[11:0] ? image_1167 : _GEN_22740; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22742 = 12'h490 == _T_221[11:0] ? image_1168 : _GEN_22741; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22743 = 12'h491 == _T_221[11:0] ? image_1169 : _GEN_22742; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22744 = 12'h492 == _T_221[11:0] ? image_1170 : _GEN_22743; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22745 = 12'h493 == _T_221[11:0] ? image_1171 : _GEN_22744; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22746 = 12'h494 == _T_221[11:0] ? image_1172 : _GEN_22745; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22747 = 12'h495 == _T_221[11:0] ? image_1173 : _GEN_22746; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22748 = 12'h496 == _T_221[11:0] ? image_1174 : _GEN_22747; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22749 = 12'h497 == _T_221[11:0] ? image_1175 : _GEN_22748; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22750 = 12'h498 == _T_221[11:0] ? image_1176 : _GEN_22749; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22751 = 12'h499 == _T_221[11:0] ? image_1177 : _GEN_22750; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22752 = 12'h49a == _T_221[11:0] ? image_1178 : _GEN_22751; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22753 = 12'h49b == _T_221[11:0] ? image_1179 : _GEN_22752; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22754 = 12'h49c == _T_221[11:0] ? image_1180 : _GEN_22753; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22755 = 12'h49d == _T_221[11:0] ? image_1181 : _GEN_22754; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22756 = 12'h49e == _T_221[11:0] ? image_1182 : _GEN_22755; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22757 = 12'h49f == _T_221[11:0] ? image_1183 : _GEN_22756; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22758 = 12'h4a0 == _T_221[11:0] ? image_1184 : _GEN_22757; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22759 = 12'h4a1 == _T_221[11:0] ? image_1185 : _GEN_22758; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22760 = 12'h4a2 == _T_221[11:0] ? image_1186 : _GEN_22759; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22761 = 12'h4a3 == _T_221[11:0] ? image_1187 : _GEN_22760; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22762 = 12'h4a4 == _T_221[11:0] ? image_1188 : _GEN_22761; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22763 = 12'h4a5 == _T_221[11:0] ? image_1189 : _GEN_22762; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22764 = 12'h4a6 == _T_221[11:0] ? image_1190 : _GEN_22763; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22765 = 12'h4a7 == _T_221[11:0] ? image_1191 : _GEN_22764; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22766 = 12'h4a8 == _T_221[11:0] ? image_1192 : _GEN_22765; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22767 = 12'h4a9 == _T_221[11:0] ? image_1193 : _GEN_22766; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22768 = 12'h4aa == _T_221[11:0] ? image_1194 : _GEN_22767; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22769 = 12'h4ab == _T_221[11:0] ? image_1195 : _GEN_22768; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22770 = 12'h4ac == _T_221[11:0] ? image_1196 : _GEN_22769; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22771 = 12'h4ad == _T_221[11:0] ? image_1197 : _GEN_22770; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22772 = 12'h4ae == _T_221[11:0] ? image_1198 : _GEN_22771; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22773 = 12'h4af == _T_221[11:0] ? image_1199 : _GEN_22772; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22774 = 12'h4b0 == _T_221[11:0] ? image_1200 : _GEN_22773; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22775 = 12'h4b1 == _T_221[11:0] ? image_1201 : _GEN_22774; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22776 = 12'h4b2 == _T_221[11:0] ? image_1202 : _GEN_22775; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22777 = 12'h4b3 == _T_221[11:0] ? image_1203 : _GEN_22776; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22778 = 12'h4b4 == _T_221[11:0] ? image_1204 : _GEN_22777; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22779 = 12'h4b5 == _T_221[11:0] ? image_1205 : _GEN_22778; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22780 = 12'h4b6 == _T_221[11:0] ? image_1206 : _GEN_22779; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22781 = 12'h4b7 == _T_221[11:0] ? image_1207 : _GEN_22780; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22782 = 12'h4b8 == _T_221[11:0] ? image_1208 : _GEN_22781; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22783 = 12'h4b9 == _T_221[11:0] ? 4'h0 : _GEN_22782; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22784 = 12'h4ba == _T_221[11:0] ? 4'h0 : _GEN_22783; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22785 = 12'h4bb == _T_221[11:0] ? 4'h0 : _GEN_22784; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22786 = 12'h4bc == _T_221[11:0] ? 4'h0 : _GEN_22785; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22787 = 12'h4bd == _T_221[11:0] ? 4'h0 : _GEN_22786; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22788 = 12'h4be == _T_221[11:0] ? 4'h0 : _GEN_22787; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22789 = 12'h4bf == _T_221[11:0] ? 4'h0 : _GEN_22788; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22790 = 12'h4c0 == _T_221[11:0] ? image_1216 : _GEN_22789; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22791 = 12'h4c1 == _T_221[11:0] ? image_1217 : _GEN_22790; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22792 = 12'h4c2 == _T_221[11:0] ? image_1218 : _GEN_22791; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22793 = 12'h4c3 == _T_221[11:0] ? image_1219 : _GEN_22792; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22794 = 12'h4c4 == _T_221[11:0] ? image_1220 : _GEN_22793; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22795 = 12'h4c5 == _T_221[11:0] ? image_1221 : _GEN_22794; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22796 = 12'h4c6 == _T_221[11:0] ? image_1222 : _GEN_22795; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22797 = 12'h4c7 == _T_221[11:0] ? image_1223 : _GEN_22796; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22798 = 12'h4c8 == _T_221[11:0] ? image_1224 : _GEN_22797; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22799 = 12'h4c9 == _T_221[11:0] ? image_1225 : _GEN_22798; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22800 = 12'h4ca == _T_221[11:0] ? image_1226 : _GEN_22799; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22801 = 12'h4cb == _T_221[11:0] ? image_1227 : _GEN_22800; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22802 = 12'h4cc == _T_221[11:0] ? image_1228 : _GEN_22801; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22803 = 12'h4cd == _T_221[11:0] ? image_1229 : _GEN_22802; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22804 = 12'h4ce == _T_221[11:0] ? image_1230 : _GEN_22803; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22805 = 12'h4cf == _T_221[11:0] ? image_1231 : _GEN_22804; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22806 = 12'h4d0 == _T_221[11:0] ? image_1232 : _GEN_22805; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22807 = 12'h4d1 == _T_221[11:0] ? image_1233 : _GEN_22806; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22808 = 12'h4d2 == _T_221[11:0] ? image_1234 : _GEN_22807; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22809 = 12'h4d3 == _T_221[11:0] ? image_1235 : _GEN_22808; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22810 = 12'h4d4 == _T_221[11:0] ? image_1236 : _GEN_22809; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22811 = 12'h4d5 == _T_221[11:0] ? image_1237 : _GEN_22810; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22812 = 12'h4d6 == _T_221[11:0] ? image_1238 : _GEN_22811; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22813 = 12'h4d7 == _T_221[11:0] ? image_1239 : _GEN_22812; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22814 = 12'h4d8 == _T_221[11:0] ? image_1240 : _GEN_22813; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22815 = 12'h4d9 == _T_221[11:0] ? image_1241 : _GEN_22814; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22816 = 12'h4da == _T_221[11:0] ? image_1242 : _GEN_22815; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22817 = 12'h4db == _T_221[11:0] ? image_1243 : _GEN_22816; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22818 = 12'h4dc == _T_221[11:0] ? image_1244 : _GEN_22817; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22819 = 12'h4dd == _T_221[11:0] ? image_1245 : _GEN_22818; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22820 = 12'h4de == _T_221[11:0] ? image_1246 : _GEN_22819; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22821 = 12'h4df == _T_221[11:0] ? image_1247 : _GEN_22820; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22822 = 12'h4e0 == _T_221[11:0] ? image_1248 : _GEN_22821; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22823 = 12'h4e1 == _T_221[11:0] ? image_1249 : _GEN_22822; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22824 = 12'h4e2 == _T_221[11:0] ? image_1250 : _GEN_22823; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22825 = 12'h4e3 == _T_221[11:0] ? image_1251 : _GEN_22824; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22826 = 12'h4e4 == _T_221[11:0] ? image_1252 : _GEN_22825; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22827 = 12'h4e5 == _T_221[11:0] ? image_1253 : _GEN_22826; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22828 = 12'h4e6 == _T_221[11:0] ? image_1254 : _GEN_22827; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22829 = 12'h4e7 == _T_221[11:0] ? image_1255 : _GEN_22828; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22830 = 12'h4e8 == _T_221[11:0] ? image_1256 : _GEN_22829; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22831 = 12'h4e9 == _T_221[11:0] ? image_1257 : _GEN_22830; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22832 = 12'h4ea == _T_221[11:0] ? image_1258 : _GEN_22831; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22833 = 12'h4eb == _T_221[11:0] ? image_1259 : _GEN_22832; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22834 = 12'h4ec == _T_221[11:0] ? image_1260 : _GEN_22833; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22835 = 12'h4ed == _T_221[11:0] ? image_1261 : _GEN_22834; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22836 = 12'h4ee == _T_221[11:0] ? image_1262 : _GEN_22835; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22837 = 12'h4ef == _T_221[11:0] ? image_1263 : _GEN_22836; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22838 = 12'h4f0 == _T_221[11:0] ? image_1264 : _GEN_22837; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22839 = 12'h4f1 == _T_221[11:0] ? image_1265 : _GEN_22838; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22840 = 12'h4f2 == _T_221[11:0] ? image_1266 : _GEN_22839; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22841 = 12'h4f3 == _T_221[11:0] ? image_1267 : _GEN_22840; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22842 = 12'h4f4 == _T_221[11:0] ? image_1268 : _GEN_22841; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22843 = 12'h4f5 == _T_221[11:0] ? image_1269 : _GEN_22842; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22844 = 12'h4f6 == _T_221[11:0] ? image_1270 : _GEN_22843; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22845 = 12'h4f7 == _T_221[11:0] ? image_1271 : _GEN_22844; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22846 = 12'h4f8 == _T_221[11:0] ? image_1272 : _GEN_22845; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22847 = 12'h4f9 == _T_221[11:0] ? image_1273 : _GEN_22846; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22848 = 12'h4fa == _T_221[11:0] ? image_1274 : _GEN_22847; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22849 = 12'h4fb == _T_221[11:0] ? image_1275 : _GEN_22848; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22850 = 12'h4fc == _T_221[11:0] ? 4'h0 : _GEN_22849; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22851 = 12'h4fd == _T_221[11:0] ? 4'h0 : _GEN_22850; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22852 = 12'h4fe == _T_221[11:0] ? 4'h0 : _GEN_22851; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22853 = 12'h4ff == _T_221[11:0] ? 4'h0 : _GEN_22852; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22854 = 12'h500 == _T_221[11:0] ? image_1280 : _GEN_22853; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22855 = 12'h501 == _T_221[11:0] ? image_1281 : _GEN_22854; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22856 = 12'h502 == _T_221[11:0] ? image_1282 : _GEN_22855; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22857 = 12'h503 == _T_221[11:0] ? image_1283 : _GEN_22856; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22858 = 12'h504 == _T_221[11:0] ? image_1284 : _GEN_22857; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22859 = 12'h505 == _T_221[11:0] ? image_1285 : _GEN_22858; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22860 = 12'h506 == _T_221[11:0] ? image_1286 : _GEN_22859; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22861 = 12'h507 == _T_221[11:0] ? image_1287 : _GEN_22860; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22862 = 12'h508 == _T_221[11:0] ? image_1288 : _GEN_22861; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22863 = 12'h509 == _T_221[11:0] ? image_1289 : _GEN_22862; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22864 = 12'h50a == _T_221[11:0] ? image_1290 : _GEN_22863; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22865 = 12'h50b == _T_221[11:0] ? image_1291 : _GEN_22864; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22866 = 12'h50c == _T_221[11:0] ? image_1292 : _GEN_22865; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22867 = 12'h50d == _T_221[11:0] ? image_1293 : _GEN_22866; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22868 = 12'h50e == _T_221[11:0] ? image_1294 : _GEN_22867; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22869 = 12'h50f == _T_221[11:0] ? image_1295 : _GEN_22868; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22870 = 12'h510 == _T_221[11:0] ? image_1296 : _GEN_22869; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22871 = 12'h511 == _T_221[11:0] ? image_1297 : _GEN_22870; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22872 = 12'h512 == _T_221[11:0] ? image_1298 : _GEN_22871; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22873 = 12'h513 == _T_221[11:0] ? image_1299 : _GEN_22872; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22874 = 12'h514 == _T_221[11:0] ? image_1300 : _GEN_22873; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22875 = 12'h515 == _T_221[11:0] ? image_1301 : _GEN_22874; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22876 = 12'h516 == _T_221[11:0] ? image_1302 : _GEN_22875; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22877 = 12'h517 == _T_221[11:0] ? image_1303 : _GEN_22876; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22878 = 12'h518 == _T_221[11:0] ? image_1304 : _GEN_22877; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22879 = 12'h519 == _T_221[11:0] ? image_1305 : _GEN_22878; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22880 = 12'h51a == _T_221[11:0] ? image_1306 : _GEN_22879; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22881 = 12'h51b == _T_221[11:0] ? image_1307 : _GEN_22880; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22882 = 12'h51c == _T_221[11:0] ? image_1308 : _GEN_22881; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22883 = 12'h51d == _T_221[11:0] ? image_1309 : _GEN_22882; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22884 = 12'h51e == _T_221[11:0] ? image_1310 : _GEN_22883; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22885 = 12'h51f == _T_221[11:0] ? image_1311 : _GEN_22884; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22886 = 12'h520 == _T_221[11:0] ? image_1312 : _GEN_22885; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22887 = 12'h521 == _T_221[11:0] ? image_1313 : _GEN_22886; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22888 = 12'h522 == _T_221[11:0] ? image_1314 : _GEN_22887; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22889 = 12'h523 == _T_221[11:0] ? image_1315 : _GEN_22888; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22890 = 12'h524 == _T_221[11:0] ? image_1316 : _GEN_22889; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22891 = 12'h525 == _T_221[11:0] ? image_1317 : _GEN_22890; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22892 = 12'h526 == _T_221[11:0] ? image_1318 : _GEN_22891; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22893 = 12'h527 == _T_221[11:0] ? image_1319 : _GEN_22892; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22894 = 12'h528 == _T_221[11:0] ? image_1320 : _GEN_22893; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22895 = 12'h529 == _T_221[11:0] ? image_1321 : _GEN_22894; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22896 = 12'h52a == _T_221[11:0] ? image_1322 : _GEN_22895; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22897 = 12'h52b == _T_221[11:0] ? image_1323 : _GEN_22896; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22898 = 12'h52c == _T_221[11:0] ? image_1324 : _GEN_22897; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22899 = 12'h52d == _T_221[11:0] ? image_1325 : _GEN_22898; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22900 = 12'h52e == _T_221[11:0] ? image_1326 : _GEN_22899; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22901 = 12'h52f == _T_221[11:0] ? image_1327 : _GEN_22900; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22902 = 12'h530 == _T_221[11:0] ? image_1328 : _GEN_22901; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22903 = 12'h531 == _T_221[11:0] ? image_1329 : _GEN_22902; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22904 = 12'h532 == _T_221[11:0] ? image_1330 : _GEN_22903; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22905 = 12'h533 == _T_221[11:0] ? image_1331 : _GEN_22904; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22906 = 12'h534 == _T_221[11:0] ? image_1332 : _GEN_22905; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22907 = 12'h535 == _T_221[11:0] ? image_1333 : _GEN_22906; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22908 = 12'h536 == _T_221[11:0] ? image_1334 : _GEN_22907; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22909 = 12'h537 == _T_221[11:0] ? image_1335 : _GEN_22908; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22910 = 12'h538 == _T_221[11:0] ? image_1336 : _GEN_22909; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22911 = 12'h539 == _T_221[11:0] ? image_1337 : _GEN_22910; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22912 = 12'h53a == _T_221[11:0] ? image_1338 : _GEN_22911; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22913 = 12'h53b == _T_221[11:0] ? image_1339 : _GEN_22912; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22914 = 12'h53c == _T_221[11:0] ? image_1340 : _GEN_22913; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22915 = 12'h53d == _T_221[11:0] ? image_1341 : _GEN_22914; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22916 = 12'h53e == _T_221[11:0] ? 4'h0 : _GEN_22915; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22917 = 12'h53f == _T_221[11:0] ? 4'h0 : _GEN_22916; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22918 = 12'h540 == _T_221[11:0] ? image_1344 : _GEN_22917; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22919 = 12'h541 == _T_221[11:0] ? image_1345 : _GEN_22918; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22920 = 12'h542 == _T_221[11:0] ? image_1346 : _GEN_22919; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22921 = 12'h543 == _T_221[11:0] ? image_1347 : _GEN_22920; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22922 = 12'h544 == _T_221[11:0] ? image_1348 : _GEN_22921; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22923 = 12'h545 == _T_221[11:0] ? image_1349 : _GEN_22922; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22924 = 12'h546 == _T_221[11:0] ? image_1350 : _GEN_22923; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22925 = 12'h547 == _T_221[11:0] ? image_1351 : _GEN_22924; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22926 = 12'h548 == _T_221[11:0] ? image_1352 : _GEN_22925; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22927 = 12'h549 == _T_221[11:0] ? image_1353 : _GEN_22926; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22928 = 12'h54a == _T_221[11:0] ? image_1354 : _GEN_22927; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22929 = 12'h54b == _T_221[11:0] ? image_1355 : _GEN_22928; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22930 = 12'h54c == _T_221[11:0] ? image_1356 : _GEN_22929; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22931 = 12'h54d == _T_221[11:0] ? image_1357 : _GEN_22930; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22932 = 12'h54e == _T_221[11:0] ? image_1358 : _GEN_22931; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22933 = 12'h54f == _T_221[11:0] ? image_1359 : _GEN_22932; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22934 = 12'h550 == _T_221[11:0] ? image_1360 : _GEN_22933; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22935 = 12'h551 == _T_221[11:0] ? image_1361 : _GEN_22934; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22936 = 12'h552 == _T_221[11:0] ? image_1362 : _GEN_22935; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22937 = 12'h553 == _T_221[11:0] ? image_1363 : _GEN_22936; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22938 = 12'h554 == _T_221[11:0] ? image_1364 : _GEN_22937; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22939 = 12'h555 == _T_221[11:0] ? image_1365 : _GEN_22938; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22940 = 12'h556 == _T_221[11:0] ? image_1366 : _GEN_22939; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22941 = 12'h557 == _T_221[11:0] ? image_1367 : _GEN_22940; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22942 = 12'h558 == _T_221[11:0] ? image_1368 : _GEN_22941; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22943 = 12'h559 == _T_221[11:0] ? image_1369 : _GEN_22942; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22944 = 12'h55a == _T_221[11:0] ? image_1370 : _GEN_22943; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22945 = 12'h55b == _T_221[11:0] ? image_1371 : _GEN_22944; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22946 = 12'h55c == _T_221[11:0] ? image_1372 : _GEN_22945; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22947 = 12'h55d == _T_221[11:0] ? image_1373 : _GEN_22946; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22948 = 12'h55e == _T_221[11:0] ? image_1374 : _GEN_22947; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22949 = 12'h55f == _T_221[11:0] ? image_1375 : _GEN_22948; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22950 = 12'h560 == _T_221[11:0] ? image_1376 : _GEN_22949; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22951 = 12'h561 == _T_221[11:0] ? image_1377 : _GEN_22950; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22952 = 12'h562 == _T_221[11:0] ? image_1378 : _GEN_22951; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22953 = 12'h563 == _T_221[11:0] ? image_1379 : _GEN_22952; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22954 = 12'h564 == _T_221[11:0] ? image_1380 : _GEN_22953; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22955 = 12'h565 == _T_221[11:0] ? image_1381 : _GEN_22954; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22956 = 12'h566 == _T_221[11:0] ? image_1382 : _GEN_22955; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22957 = 12'h567 == _T_221[11:0] ? image_1383 : _GEN_22956; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22958 = 12'h568 == _T_221[11:0] ? image_1384 : _GEN_22957; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22959 = 12'h569 == _T_221[11:0] ? image_1385 : _GEN_22958; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22960 = 12'h56a == _T_221[11:0] ? image_1386 : _GEN_22959; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22961 = 12'h56b == _T_221[11:0] ? image_1387 : _GEN_22960; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22962 = 12'h56c == _T_221[11:0] ? image_1388 : _GEN_22961; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22963 = 12'h56d == _T_221[11:0] ? image_1389 : _GEN_22962; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22964 = 12'h56e == _T_221[11:0] ? image_1390 : _GEN_22963; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22965 = 12'h56f == _T_221[11:0] ? image_1391 : _GEN_22964; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22966 = 12'h570 == _T_221[11:0] ? image_1392 : _GEN_22965; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22967 = 12'h571 == _T_221[11:0] ? image_1393 : _GEN_22966; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22968 = 12'h572 == _T_221[11:0] ? image_1394 : _GEN_22967; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22969 = 12'h573 == _T_221[11:0] ? image_1395 : _GEN_22968; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22970 = 12'h574 == _T_221[11:0] ? image_1396 : _GEN_22969; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22971 = 12'h575 == _T_221[11:0] ? image_1397 : _GEN_22970; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22972 = 12'h576 == _T_221[11:0] ? image_1398 : _GEN_22971; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22973 = 12'h577 == _T_221[11:0] ? image_1399 : _GEN_22972; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22974 = 12'h578 == _T_221[11:0] ? image_1400 : _GEN_22973; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22975 = 12'h579 == _T_221[11:0] ? image_1401 : _GEN_22974; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22976 = 12'h57a == _T_221[11:0] ? image_1402 : _GEN_22975; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22977 = 12'h57b == _T_221[11:0] ? image_1403 : _GEN_22976; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22978 = 12'h57c == _T_221[11:0] ? image_1404 : _GEN_22977; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22979 = 12'h57d == _T_221[11:0] ? image_1405 : _GEN_22978; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22980 = 12'h57e == _T_221[11:0] ? 4'h0 : _GEN_22979; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22981 = 12'h57f == _T_221[11:0] ? 4'h0 : _GEN_22980; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22982 = 12'h580 == _T_221[11:0] ? image_1408 : _GEN_22981; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22983 = 12'h581 == _T_221[11:0] ? image_1409 : _GEN_22982; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22984 = 12'h582 == _T_221[11:0] ? image_1410 : _GEN_22983; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22985 = 12'h583 == _T_221[11:0] ? image_1411 : _GEN_22984; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22986 = 12'h584 == _T_221[11:0] ? image_1412 : _GEN_22985; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22987 = 12'h585 == _T_221[11:0] ? image_1413 : _GEN_22986; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22988 = 12'h586 == _T_221[11:0] ? image_1414 : _GEN_22987; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22989 = 12'h587 == _T_221[11:0] ? image_1415 : _GEN_22988; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22990 = 12'h588 == _T_221[11:0] ? image_1416 : _GEN_22989; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22991 = 12'h589 == _T_221[11:0] ? image_1417 : _GEN_22990; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22992 = 12'h58a == _T_221[11:0] ? image_1418 : _GEN_22991; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22993 = 12'h58b == _T_221[11:0] ? image_1419 : _GEN_22992; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22994 = 12'h58c == _T_221[11:0] ? image_1420 : _GEN_22993; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22995 = 12'h58d == _T_221[11:0] ? image_1421 : _GEN_22994; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22996 = 12'h58e == _T_221[11:0] ? image_1422 : _GEN_22995; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22997 = 12'h58f == _T_221[11:0] ? image_1423 : _GEN_22996; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22998 = 12'h590 == _T_221[11:0] ? image_1424 : _GEN_22997; // @[Filter.scala 138:46]
  wire [3:0] _GEN_22999 = 12'h591 == _T_221[11:0] ? image_1425 : _GEN_22998; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23000 = 12'h592 == _T_221[11:0] ? image_1426 : _GEN_22999; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23001 = 12'h593 == _T_221[11:0] ? image_1427 : _GEN_23000; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23002 = 12'h594 == _T_221[11:0] ? image_1428 : _GEN_23001; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23003 = 12'h595 == _T_221[11:0] ? image_1429 : _GEN_23002; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23004 = 12'h596 == _T_221[11:0] ? image_1430 : _GEN_23003; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23005 = 12'h597 == _T_221[11:0] ? image_1431 : _GEN_23004; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23006 = 12'h598 == _T_221[11:0] ? image_1432 : _GEN_23005; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23007 = 12'h599 == _T_221[11:0] ? image_1433 : _GEN_23006; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23008 = 12'h59a == _T_221[11:0] ? image_1434 : _GEN_23007; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23009 = 12'h59b == _T_221[11:0] ? image_1435 : _GEN_23008; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23010 = 12'h59c == _T_221[11:0] ? image_1436 : _GEN_23009; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23011 = 12'h59d == _T_221[11:0] ? image_1437 : _GEN_23010; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23012 = 12'h59e == _T_221[11:0] ? image_1438 : _GEN_23011; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23013 = 12'h59f == _T_221[11:0] ? image_1439 : _GEN_23012; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23014 = 12'h5a0 == _T_221[11:0] ? image_1440 : _GEN_23013; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23015 = 12'h5a1 == _T_221[11:0] ? image_1441 : _GEN_23014; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23016 = 12'h5a2 == _T_221[11:0] ? image_1442 : _GEN_23015; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23017 = 12'h5a3 == _T_221[11:0] ? image_1443 : _GEN_23016; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23018 = 12'h5a4 == _T_221[11:0] ? image_1444 : _GEN_23017; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23019 = 12'h5a5 == _T_221[11:0] ? image_1445 : _GEN_23018; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23020 = 12'h5a6 == _T_221[11:0] ? image_1446 : _GEN_23019; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23021 = 12'h5a7 == _T_221[11:0] ? image_1447 : _GEN_23020; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23022 = 12'h5a8 == _T_221[11:0] ? image_1448 : _GEN_23021; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23023 = 12'h5a9 == _T_221[11:0] ? image_1449 : _GEN_23022; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23024 = 12'h5aa == _T_221[11:0] ? image_1450 : _GEN_23023; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23025 = 12'h5ab == _T_221[11:0] ? image_1451 : _GEN_23024; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23026 = 12'h5ac == _T_221[11:0] ? image_1452 : _GEN_23025; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23027 = 12'h5ad == _T_221[11:0] ? image_1453 : _GEN_23026; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23028 = 12'h5ae == _T_221[11:0] ? image_1454 : _GEN_23027; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23029 = 12'h5af == _T_221[11:0] ? image_1455 : _GEN_23028; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23030 = 12'h5b0 == _T_221[11:0] ? image_1456 : _GEN_23029; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23031 = 12'h5b1 == _T_221[11:0] ? image_1457 : _GEN_23030; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23032 = 12'h5b2 == _T_221[11:0] ? image_1458 : _GEN_23031; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23033 = 12'h5b3 == _T_221[11:0] ? image_1459 : _GEN_23032; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23034 = 12'h5b4 == _T_221[11:0] ? image_1460 : _GEN_23033; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23035 = 12'h5b5 == _T_221[11:0] ? image_1461 : _GEN_23034; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23036 = 12'h5b6 == _T_221[11:0] ? image_1462 : _GEN_23035; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23037 = 12'h5b7 == _T_221[11:0] ? image_1463 : _GEN_23036; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23038 = 12'h5b8 == _T_221[11:0] ? image_1464 : _GEN_23037; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23039 = 12'h5b9 == _T_221[11:0] ? image_1465 : _GEN_23038; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23040 = 12'h5ba == _T_221[11:0] ? image_1466 : _GEN_23039; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23041 = 12'h5bb == _T_221[11:0] ? image_1467 : _GEN_23040; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23042 = 12'h5bc == _T_221[11:0] ? image_1468 : _GEN_23041; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23043 = 12'h5bd == _T_221[11:0] ? image_1469 : _GEN_23042; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23044 = 12'h5be == _T_221[11:0] ? 4'h0 : _GEN_23043; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23045 = 12'h5bf == _T_221[11:0] ? 4'h0 : _GEN_23044; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23046 = 12'h5c0 == _T_221[11:0] ? image_1472 : _GEN_23045; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23047 = 12'h5c1 == _T_221[11:0] ? image_1473 : _GEN_23046; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23048 = 12'h5c2 == _T_221[11:0] ? image_1474 : _GEN_23047; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23049 = 12'h5c3 == _T_221[11:0] ? image_1475 : _GEN_23048; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23050 = 12'h5c4 == _T_221[11:0] ? image_1476 : _GEN_23049; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23051 = 12'h5c5 == _T_221[11:0] ? image_1477 : _GEN_23050; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23052 = 12'h5c6 == _T_221[11:0] ? image_1478 : _GEN_23051; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23053 = 12'h5c7 == _T_221[11:0] ? image_1479 : _GEN_23052; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23054 = 12'h5c8 == _T_221[11:0] ? image_1480 : _GEN_23053; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23055 = 12'h5c9 == _T_221[11:0] ? image_1481 : _GEN_23054; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23056 = 12'h5ca == _T_221[11:0] ? image_1482 : _GEN_23055; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23057 = 12'h5cb == _T_221[11:0] ? image_1483 : _GEN_23056; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23058 = 12'h5cc == _T_221[11:0] ? image_1484 : _GEN_23057; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23059 = 12'h5cd == _T_221[11:0] ? image_1485 : _GEN_23058; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23060 = 12'h5ce == _T_221[11:0] ? image_1486 : _GEN_23059; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23061 = 12'h5cf == _T_221[11:0] ? image_1487 : _GEN_23060; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23062 = 12'h5d0 == _T_221[11:0] ? image_1488 : _GEN_23061; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23063 = 12'h5d1 == _T_221[11:0] ? image_1489 : _GEN_23062; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23064 = 12'h5d2 == _T_221[11:0] ? image_1490 : _GEN_23063; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23065 = 12'h5d3 == _T_221[11:0] ? image_1491 : _GEN_23064; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23066 = 12'h5d4 == _T_221[11:0] ? image_1492 : _GEN_23065; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23067 = 12'h5d5 == _T_221[11:0] ? image_1493 : _GEN_23066; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23068 = 12'h5d6 == _T_221[11:0] ? image_1494 : _GEN_23067; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23069 = 12'h5d7 == _T_221[11:0] ? image_1495 : _GEN_23068; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23070 = 12'h5d8 == _T_221[11:0] ? image_1496 : _GEN_23069; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23071 = 12'h5d9 == _T_221[11:0] ? image_1497 : _GEN_23070; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23072 = 12'h5da == _T_221[11:0] ? image_1498 : _GEN_23071; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23073 = 12'h5db == _T_221[11:0] ? image_1499 : _GEN_23072; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23074 = 12'h5dc == _T_221[11:0] ? image_1500 : _GEN_23073; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23075 = 12'h5dd == _T_221[11:0] ? image_1501 : _GEN_23074; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23076 = 12'h5de == _T_221[11:0] ? image_1502 : _GEN_23075; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23077 = 12'h5df == _T_221[11:0] ? image_1503 : _GEN_23076; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23078 = 12'h5e0 == _T_221[11:0] ? image_1504 : _GEN_23077; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23079 = 12'h5e1 == _T_221[11:0] ? image_1505 : _GEN_23078; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23080 = 12'h5e2 == _T_221[11:0] ? image_1506 : _GEN_23079; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23081 = 12'h5e3 == _T_221[11:0] ? image_1507 : _GEN_23080; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23082 = 12'h5e4 == _T_221[11:0] ? image_1508 : _GEN_23081; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23083 = 12'h5e5 == _T_221[11:0] ? image_1509 : _GEN_23082; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23084 = 12'h5e6 == _T_221[11:0] ? image_1510 : _GEN_23083; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23085 = 12'h5e7 == _T_221[11:0] ? image_1511 : _GEN_23084; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23086 = 12'h5e8 == _T_221[11:0] ? image_1512 : _GEN_23085; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23087 = 12'h5e9 == _T_221[11:0] ? image_1513 : _GEN_23086; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23088 = 12'h5ea == _T_221[11:0] ? image_1514 : _GEN_23087; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23089 = 12'h5eb == _T_221[11:0] ? image_1515 : _GEN_23088; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23090 = 12'h5ec == _T_221[11:0] ? image_1516 : _GEN_23089; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23091 = 12'h5ed == _T_221[11:0] ? image_1517 : _GEN_23090; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23092 = 12'h5ee == _T_221[11:0] ? image_1518 : _GEN_23091; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23093 = 12'h5ef == _T_221[11:0] ? image_1519 : _GEN_23092; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23094 = 12'h5f0 == _T_221[11:0] ? image_1520 : _GEN_23093; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23095 = 12'h5f1 == _T_221[11:0] ? image_1521 : _GEN_23094; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23096 = 12'h5f2 == _T_221[11:0] ? image_1522 : _GEN_23095; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23097 = 12'h5f3 == _T_221[11:0] ? image_1523 : _GEN_23096; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23098 = 12'h5f4 == _T_221[11:0] ? image_1524 : _GEN_23097; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23099 = 12'h5f5 == _T_221[11:0] ? image_1525 : _GEN_23098; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23100 = 12'h5f6 == _T_221[11:0] ? image_1526 : _GEN_23099; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23101 = 12'h5f7 == _T_221[11:0] ? image_1527 : _GEN_23100; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23102 = 12'h5f8 == _T_221[11:0] ? image_1528 : _GEN_23101; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23103 = 12'h5f9 == _T_221[11:0] ? image_1529 : _GEN_23102; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23104 = 12'h5fa == _T_221[11:0] ? image_1530 : _GEN_23103; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23105 = 12'h5fb == _T_221[11:0] ? image_1531 : _GEN_23104; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23106 = 12'h5fc == _T_221[11:0] ? image_1532 : _GEN_23105; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23107 = 12'h5fd == _T_221[11:0] ? image_1533 : _GEN_23106; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23108 = 12'h5fe == _T_221[11:0] ? 4'h0 : _GEN_23107; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23109 = 12'h5ff == _T_221[11:0] ? 4'h0 : _GEN_23108; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23110 = 12'h600 == _T_221[11:0] ? image_1536 : _GEN_23109; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23111 = 12'h601 == _T_221[11:0] ? image_1537 : _GEN_23110; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23112 = 12'h602 == _T_221[11:0] ? image_1538 : _GEN_23111; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23113 = 12'h603 == _T_221[11:0] ? image_1539 : _GEN_23112; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23114 = 12'h604 == _T_221[11:0] ? image_1540 : _GEN_23113; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23115 = 12'h605 == _T_221[11:0] ? image_1541 : _GEN_23114; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23116 = 12'h606 == _T_221[11:0] ? image_1542 : _GEN_23115; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23117 = 12'h607 == _T_221[11:0] ? image_1543 : _GEN_23116; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23118 = 12'h608 == _T_221[11:0] ? image_1544 : _GEN_23117; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23119 = 12'h609 == _T_221[11:0] ? image_1545 : _GEN_23118; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23120 = 12'h60a == _T_221[11:0] ? image_1546 : _GEN_23119; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23121 = 12'h60b == _T_221[11:0] ? image_1547 : _GEN_23120; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23122 = 12'h60c == _T_221[11:0] ? image_1548 : _GEN_23121; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23123 = 12'h60d == _T_221[11:0] ? image_1549 : _GEN_23122; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23124 = 12'h60e == _T_221[11:0] ? image_1550 : _GEN_23123; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23125 = 12'h60f == _T_221[11:0] ? image_1551 : _GEN_23124; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23126 = 12'h610 == _T_221[11:0] ? image_1552 : _GEN_23125; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23127 = 12'h611 == _T_221[11:0] ? image_1553 : _GEN_23126; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23128 = 12'h612 == _T_221[11:0] ? image_1554 : _GEN_23127; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23129 = 12'h613 == _T_221[11:0] ? image_1555 : _GEN_23128; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23130 = 12'h614 == _T_221[11:0] ? image_1556 : _GEN_23129; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23131 = 12'h615 == _T_221[11:0] ? image_1557 : _GEN_23130; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23132 = 12'h616 == _T_221[11:0] ? image_1558 : _GEN_23131; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23133 = 12'h617 == _T_221[11:0] ? image_1559 : _GEN_23132; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23134 = 12'h618 == _T_221[11:0] ? image_1560 : _GEN_23133; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23135 = 12'h619 == _T_221[11:0] ? image_1561 : _GEN_23134; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23136 = 12'h61a == _T_221[11:0] ? image_1562 : _GEN_23135; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23137 = 12'h61b == _T_221[11:0] ? image_1563 : _GEN_23136; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23138 = 12'h61c == _T_221[11:0] ? image_1564 : _GEN_23137; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23139 = 12'h61d == _T_221[11:0] ? image_1565 : _GEN_23138; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23140 = 12'h61e == _T_221[11:0] ? image_1566 : _GEN_23139; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23141 = 12'h61f == _T_221[11:0] ? image_1567 : _GEN_23140; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23142 = 12'h620 == _T_221[11:0] ? image_1568 : _GEN_23141; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23143 = 12'h621 == _T_221[11:0] ? image_1569 : _GEN_23142; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23144 = 12'h622 == _T_221[11:0] ? image_1570 : _GEN_23143; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23145 = 12'h623 == _T_221[11:0] ? image_1571 : _GEN_23144; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23146 = 12'h624 == _T_221[11:0] ? image_1572 : _GEN_23145; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23147 = 12'h625 == _T_221[11:0] ? image_1573 : _GEN_23146; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23148 = 12'h626 == _T_221[11:0] ? image_1574 : _GEN_23147; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23149 = 12'h627 == _T_221[11:0] ? image_1575 : _GEN_23148; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23150 = 12'h628 == _T_221[11:0] ? image_1576 : _GEN_23149; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23151 = 12'h629 == _T_221[11:0] ? image_1577 : _GEN_23150; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23152 = 12'h62a == _T_221[11:0] ? image_1578 : _GEN_23151; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23153 = 12'h62b == _T_221[11:0] ? image_1579 : _GEN_23152; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23154 = 12'h62c == _T_221[11:0] ? image_1580 : _GEN_23153; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23155 = 12'h62d == _T_221[11:0] ? image_1581 : _GEN_23154; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23156 = 12'h62e == _T_221[11:0] ? image_1582 : _GEN_23155; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23157 = 12'h62f == _T_221[11:0] ? image_1583 : _GEN_23156; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23158 = 12'h630 == _T_221[11:0] ? image_1584 : _GEN_23157; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23159 = 12'h631 == _T_221[11:0] ? image_1585 : _GEN_23158; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23160 = 12'h632 == _T_221[11:0] ? image_1586 : _GEN_23159; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23161 = 12'h633 == _T_221[11:0] ? image_1587 : _GEN_23160; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23162 = 12'h634 == _T_221[11:0] ? image_1588 : _GEN_23161; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23163 = 12'h635 == _T_221[11:0] ? image_1589 : _GEN_23162; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23164 = 12'h636 == _T_221[11:0] ? image_1590 : _GEN_23163; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23165 = 12'h637 == _T_221[11:0] ? image_1591 : _GEN_23164; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23166 = 12'h638 == _T_221[11:0] ? image_1592 : _GEN_23165; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23167 = 12'h639 == _T_221[11:0] ? image_1593 : _GEN_23166; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23168 = 12'h63a == _T_221[11:0] ? image_1594 : _GEN_23167; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23169 = 12'h63b == _T_221[11:0] ? image_1595 : _GEN_23168; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23170 = 12'h63c == _T_221[11:0] ? image_1596 : _GEN_23169; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23171 = 12'h63d == _T_221[11:0] ? image_1597 : _GEN_23170; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23172 = 12'h63e == _T_221[11:0] ? 4'h0 : _GEN_23171; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23173 = 12'h63f == _T_221[11:0] ? 4'h0 : _GEN_23172; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23174 = 12'h640 == _T_221[11:0] ? image_1600 : _GEN_23173; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23175 = 12'h641 == _T_221[11:0] ? image_1601 : _GEN_23174; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23176 = 12'h642 == _T_221[11:0] ? image_1602 : _GEN_23175; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23177 = 12'h643 == _T_221[11:0] ? image_1603 : _GEN_23176; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23178 = 12'h644 == _T_221[11:0] ? image_1604 : _GEN_23177; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23179 = 12'h645 == _T_221[11:0] ? image_1605 : _GEN_23178; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23180 = 12'h646 == _T_221[11:0] ? image_1606 : _GEN_23179; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23181 = 12'h647 == _T_221[11:0] ? image_1607 : _GEN_23180; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23182 = 12'h648 == _T_221[11:0] ? image_1608 : _GEN_23181; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23183 = 12'h649 == _T_221[11:0] ? image_1609 : _GEN_23182; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23184 = 12'h64a == _T_221[11:0] ? image_1610 : _GEN_23183; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23185 = 12'h64b == _T_221[11:0] ? image_1611 : _GEN_23184; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23186 = 12'h64c == _T_221[11:0] ? image_1612 : _GEN_23185; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23187 = 12'h64d == _T_221[11:0] ? image_1613 : _GEN_23186; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23188 = 12'h64e == _T_221[11:0] ? image_1614 : _GEN_23187; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23189 = 12'h64f == _T_221[11:0] ? image_1615 : _GEN_23188; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23190 = 12'h650 == _T_221[11:0] ? image_1616 : _GEN_23189; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23191 = 12'h651 == _T_221[11:0] ? image_1617 : _GEN_23190; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23192 = 12'h652 == _T_221[11:0] ? image_1618 : _GEN_23191; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23193 = 12'h653 == _T_221[11:0] ? image_1619 : _GEN_23192; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23194 = 12'h654 == _T_221[11:0] ? image_1620 : _GEN_23193; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23195 = 12'h655 == _T_221[11:0] ? image_1621 : _GEN_23194; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23196 = 12'h656 == _T_221[11:0] ? image_1622 : _GEN_23195; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23197 = 12'h657 == _T_221[11:0] ? image_1623 : _GEN_23196; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23198 = 12'h658 == _T_221[11:0] ? image_1624 : _GEN_23197; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23199 = 12'h659 == _T_221[11:0] ? image_1625 : _GEN_23198; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23200 = 12'h65a == _T_221[11:0] ? image_1626 : _GEN_23199; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23201 = 12'h65b == _T_221[11:0] ? image_1627 : _GEN_23200; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23202 = 12'h65c == _T_221[11:0] ? image_1628 : _GEN_23201; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23203 = 12'h65d == _T_221[11:0] ? image_1629 : _GEN_23202; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23204 = 12'h65e == _T_221[11:0] ? image_1630 : _GEN_23203; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23205 = 12'h65f == _T_221[11:0] ? image_1631 : _GEN_23204; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23206 = 12'h660 == _T_221[11:0] ? image_1632 : _GEN_23205; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23207 = 12'h661 == _T_221[11:0] ? image_1633 : _GEN_23206; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23208 = 12'h662 == _T_221[11:0] ? image_1634 : _GEN_23207; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23209 = 12'h663 == _T_221[11:0] ? image_1635 : _GEN_23208; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23210 = 12'h664 == _T_221[11:0] ? image_1636 : _GEN_23209; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23211 = 12'h665 == _T_221[11:0] ? image_1637 : _GEN_23210; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23212 = 12'h666 == _T_221[11:0] ? image_1638 : _GEN_23211; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23213 = 12'h667 == _T_221[11:0] ? image_1639 : _GEN_23212; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23214 = 12'h668 == _T_221[11:0] ? image_1640 : _GEN_23213; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23215 = 12'h669 == _T_221[11:0] ? image_1641 : _GEN_23214; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23216 = 12'h66a == _T_221[11:0] ? image_1642 : _GEN_23215; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23217 = 12'h66b == _T_221[11:0] ? image_1643 : _GEN_23216; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23218 = 12'h66c == _T_221[11:0] ? image_1644 : _GEN_23217; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23219 = 12'h66d == _T_221[11:0] ? image_1645 : _GEN_23218; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23220 = 12'h66e == _T_221[11:0] ? image_1646 : _GEN_23219; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23221 = 12'h66f == _T_221[11:0] ? image_1647 : _GEN_23220; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23222 = 12'h670 == _T_221[11:0] ? image_1648 : _GEN_23221; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23223 = 12'h671 == _T_221[11:0] ? image_1649 : _GEN_23222; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23224 = 12'h672 == _T_221[11:0] ? image_1650 : _GEN_23223; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23225 = 12'h673 == _T_221[11:0] ? image_1651 : _GEN_23224; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23226 = 12'h674 == _T_221[11:0] ? image_1652 : _GEN_23225; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23227 = 12'h675 == _T_221[11:0] ? image_1653 : _GEN_23226; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23228 = 12'h676 == _T_221[11:0] ? image_1654 : _GEN_23227; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23229 = 12'h677 == _T_221[11:0] ? image_1655 : _GEN_23228; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23230 = 12'h678 == _T_221[11:0] ? image_1656 : _GEN_23229; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23231 = 12'h679 == _T_221[11:0] ? image_1657 : _GEN_23230; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23232 = 12'h67a == _T_221[11:0] ? image_1658 : _GEN_23231; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23233 = 12'h67b == _T_221[11:0] ? image_1659 : _GEN_23232; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23234 = 12'h67c == _T_221[11:0] ? image_1660 : _GEN_23233; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23235 = 12'h67d == _T_221[11:0] ? 4'h0 : _GEN_23234; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23236 = 12'h67e == _T_221[11:0] ? 4'h0 : _GEN_23235; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23237 = 12'h67f == _T_221[11:0] ? 4'h0 : _GEN_23236; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23238 = 12'h680 == _T_221[11:0] ? image_1664 : _GEN_23237; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23239 = 12'h681 == _T_221[11:0] ? image_1665 : _GEN_23238; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23240 = 12'h682 == _T_221[11:0] ? image_1666 : _GEN_23239; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23241 = 12'h683 == _T_221[11:0] ? image_1667 : _GEN_23240; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23242 = 12'h684 == _T_221[11:0] ? image_1668 : _GEN_23241; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23243 = 12'h685 == _T_221[11:0] ? image_1669 : _GEN_23242; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23244 = 12'h686 == _T_221[11:0] ? image_1670 : _GEN_23243; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23245 = 12'h687 == _T_221[11:0] ? image_1671 : _GEN_23244; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23246 = 12'h688 == _T_221[11:0] ? image_1672 : _GEN_23245; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23247 = 12'h689 == _T_221[11:0] ? image_1673 : _GEN_23246; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23248 = 12'h68a == _T_221[11:0] ? image_1674 : _GEN_23247; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23249 = 12'h68b == _T_221[11:0] ? image_1675 : _GEN_23248; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23250 = 12'h68c == _T_221[11:0] ? image_1676 : _GEN_23249; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23251 = 12'h68d == _T_221[11:0] ? image_1677 : _GEN_23250; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23252 = 12'h68e == _T_221[11:0] ? image_1678 : _GEN_23251; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23253 = 12'h68f == _T_221[11:0] ? image_1679 : _GEN_23252; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23254 = 12'h690 == _T_221[11:0] ? image_1680 : _GEN_23253; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23255 = 12'h691 == _T_221[11:0] ? image_1681 : _GEN_23254; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23256 = 12'h692 == _T_221[11:0] ? image_1682 : _GEN_23255; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23257 = 12'h693 == _T_221[11:0] ? image_1683 : _GEN_23256; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23258 = 12'h694 == _T_221[11:0] ? image_1684 : _GEN_23257; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23259 = 12'h695 == _T_221[11:0] ? image_1685 : _GEN_23258; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23260 = 12'h696 == _T_221[11:0] ? image_1686 : _GEN_23259; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23261 = 12'h697 == _T_221[11:0] ? image_1687 : _GEN_23260; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23262 = 12'h698 == _T_221[11:0] ? image_1688 : _GEN_23261; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23263 = 12'h699 == _T_221[11:0] ? image_1689 : _GEN_23262; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23264 = 12'h69a == _T_221[11:0] ? image_1690 : _GEN_23263; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23265 = 12'h69b == _T_221[11:0] ? image_1691 : _GEN_23264; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23266 = 12'h69c == _T_221[11:0] ? image_1692 : _GEN_23265; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23267 = 12'h69d == _T_221[11:0] ? image_1693 : _GEN_23266; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23268 = 12'h69e == _T_221[11:0] ? image_1694 : _GEN_23267; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23269 = 12'h69f == _T_221[11:0] ? image_1695 : _GEN_23268; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23270 = 12'h6a0 == _T_221[11:0] ? image_1696 : _GEN_23269; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23271 = 12'h6a1 == _T_221[11:0] ? image_1697 : _GEN_23270; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23272 = 12'h6a2 == _T_221[11:0] ? image_1698 : _GEN_23271; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23273 = 12'h6a3 == _T_221[11:0] ? image_1699 : _GEN_23272; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23274 = 12'h6a4 == _T_221[11:0] ? image_1700 : _GEN_23273; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23275 = 12'h6a5 == _T_221[11:0] ? image_1701 : _GEN_23274; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23276 = 12'h6a6 == _T_221[11:0] ? image_1702 : _GEN_23275; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23277 = 12'h6a7 == _T_221[11:0] ? image_1703 : _GEN_23276; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23278 = 12'h6a8 == _T_221[11:0] ? image_1704 : _GEN_23277; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23279 = 12'h6a9 == _T_221[11:0] ? image_1705 : _GEN_23278; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23280 = 12'h6aa == _T_221[11:0] ? image_1706 : _GEN_23279; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23281 = 12'h6ab == _T_221[11:0] ? image_1707 : _GEN_23280; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23282 = 12'h6ac == _T_221[11:0] ? image_1708 : _GEN_23281; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23283 = 12'h6ad == _T_221[11:0] ? image_1709 : _GEN_23282; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23284 = 12'h6ae == _T_221[11:0] ? image_1710 : _GEN_23283; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23285 = 12'h6af == _T_221[11:0] ? image_1711 : _GEN_23284; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23286 = 12'h6b0 == _T_221[11:0] ? image_1712 : _GEN_23285; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23287 = 12'h6b1 == _T_221[11:0] ? image_1713 : _GEN_23286; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23288 = 12'h6b2 == _T_221[11:0] ? image_1714 : _GEN_23287; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23289 = 12'h6b3 == _T_221[11:0] ? image_1715 : _GEN_23288; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23290 = 12'h6b4 == _T_221[11:0] ? image_1716 : _GEN_23289; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23291 = 12'h6b5 == _T_221[11:0] ? image_1717 : _GEN_23290; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23292 = 12'h6b6 == _T_221[11:0] ? image_1718 : _GEN_23291; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23293 = 12'h6b7 == _T_221[11:0] ? image_1719 : _GEN_23292; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23294 = 12'h6b8 == _T_221[11:0] ? image_1720 : _GEN_23293; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23295 = 12'h6b9 == _T_221[11:0] ? image_1721 : _GEN_23294; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23296 = 12'h6ba == _T_221[11:0] ? image_1722 : _GEN_23295; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23297 = 12'h6bb == _T_221[11:0] ? image_1723 : _GEN_23296; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23298 = 12'h6bc == _T_221[11:0] ? 4'h0 : _GEN_23297; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23299 = 12'h6bd == _T_221[11:0] ? 4'h0 : _GEN_23298; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23300 = 12'h6be == _T_221[11:0] ? 4'h0 : _GEN_23299; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23301 = 12'h6bf == _T_221[11:0] ? 4'h0 : _GEN_23300; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23302 = 12'h6c0 == _T_221[11:0] ? image_1728 : _GEN_23301; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23303 = 12'h6c1 == _T_221[11:0] ? image_1729 : _GEN_23302; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23304 = 12'h6c2 == _T_221[11:0] ? image_1730 : _GEN_23303; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23305 = 12'h6c3 == _T_221[11:0] ? image_1731 : _GEN_23304; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23306 = 12'h6c4 == _T_221[11:0] ? image_1732 : _GEN_23305; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23307 = 12'h6c5 == _T_221[11:0] ? image_1733 : _GEN_23306; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23308 = 12'h6c6 == _T_221[11:0] ? image_1734 : _GEN_23307; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23309 = 12'h6c7 == _T_221[11:0] ? image_1735 : _GEN_23308; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23310 = 12'h6c8 == _T_221[11:0] ? image_1736 : _GEN_23309; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23311 = 12'h6c9 == _T_221[11:0] ? image_1737 : _GEN_23310; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23312 = 12'h6ca == _T_221[11:0] ? image_1738 : _GEN_23311; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23313 = 12'h6cb == _T_221[11:0] ? image_1739 : _GEN_23312; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23314 = 12'h6cc == _T_221[11:0] ? image_1740 : _GEN_23313; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23315 = 12'h6cd == _T_221[11:0] ? image_1741 : _GEN_23314; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23316 = 12'h6ce == _T_221[11:0] ? image_1742 : _GEN_23315; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23317 = 12'h6cf == _T_221[11:0] ? image_1743 : _GEN_23316; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23318 = 12'h6d0 == _T_221[11:0] ? image_1744 : _GEN_23317; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23319 = 12'h6d1 == _T_221[11:0] ? image_1745 : _GEN_23318; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23320 = 12'h6d2 == _T_221[11:0] ? image_1746 : _GEN_23319; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23321 = 12'h6d3 == _T_221[11:0] ? image_1747 : _GEN_23320; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23322 = 12'h6d4 == _T_221[11:0] ? image_1748 : _GEN_23321; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23323 = 12'h6d5 == _T_221[11:0] ? image_1749 : _GEN_23322; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23324 = 12'h6d6 == _T_221[11:0] ? image_1750 : _GEN_23323; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23325 = 12'h6d7 == _T_221[11:0] ? image_1751 : _GEN_23324; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23326 = 12'h6d8 == _T_221[11:0] ? image_1752 : _GEN_23325; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23327 = 12'h6d9 == _T_221[11:0] ? image_1753 : _GEN_23326; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23328 = 12'h6da == _T_221[11:0] ? image_1754 : _GEN_23327; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23329 = 12'h6db == _T_221[11:0] ? image_1755 : _GEN_23328; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23330 = 12'h6dc == _T_221[11:0] ? image_1756 : _GEN_23329; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23331 = 12'h6dd == _T_221[11:0] ? image_1757 : _GEN_23330; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23332 = 12'h6de == _T_221[11:0] ? image_1758 : _GEN_23331; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23333 = 12'h6df == _T_221[11:0] ? image_1759 : _GEN_23332; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23334 = 12'h6e0 == _T_221[11:0] ? image_1760 : _GEN_23333; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23335 = 12'h6e1 == _T_221[11:0] ? image_1761 : _GEN_23334; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23336 = 12'h6e2 == _T_221[11:0] ? image_1762 : _GEN_23335; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23337 = 12'h6e3 == _T_221[11:0] ? image_1763 : _GEN_23336; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23338 = 12'h6e4 == _T_221[11:0] ? image_1764 : _GEN_23337; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23339 = 12'h6e5 == _T_221[11:0] ? image_1765 : _GEN_23338; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23340 = 12'h6e6 == _T_221[11:0] ? image_1766 : _GEN_23339; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23341 = 12'h6e7 == _T_221[11:0] ? image_1767 : _GEN_23340; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23342 = 12'h6e8 == _T_221[11:0] ? image_1768 : _GEN_23341; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23343 = 12'h6e9 == _T_221[11:0] ? image_1769 : _GEN_23342; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23344 = 12'h6ea == _T_221[11:0] ? image_1770 : _GEN_23343; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23345 = 12'h6eb == _T_221[11:0] ? image_1771 : _GEN_23344; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23346 = 12'h6ec == _T_221[11:0] ? image_1772 : _GEN_23345; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23347 = 12'h6ed == _T_221[11:0] ? image_1773 : _GEN_23346; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23348 = 12'h6ee == _T_221[11:0] ? image_1774 : _GEN_23347; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23349 = 12'h6ef == _T_221[11:0] ? image_1775 : _GEN_23348; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23350 = 12'h6f0 == _T_221[11:0] ? image_1776 : _GEN_23349; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23351 = 12'h6f1 == _T_221[11:0] ? image_1777 : _GEN_23350; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23352 = 12'h6f2 == _T_221[11:0] ? image_1778 : _GEN_23351; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23353 = 12'h6f3 == _T_221[11:0] ? image_1779 : _GEN_23352; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23354 = 12'h6f4 == _T_221[11:0] ? image_1780 : _GEN_23353; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23355 = 12'h6f5 == _T_221[11:0] ? image_1781 : _GEN_23354; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23356 = 12'h6f6 == _T_221[11:0] ? image_1782 : _GEN_23355; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23357 = 12'h6f7 == _T_221[11:0] ? image_1783 : _GEN_23356; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23358 = 12'h6f8 == _T_221[11:0] ? image_1784 : _GEN_23357; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23359 = 12'h6f9 == _T_221[11:0] ? image_1785 : _GEN_23358; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23360 = 12'h6fa == _T_221[11:0] ? image_1786 : _GEN_23359; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23361 = 12'h6fb == _T_221[11:0] ? 4'h0 : _GEN_23360; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23362 = 12'h6fc == _T_221[11:0] ? 4'h0 : _GEN_23361; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23363 = 12'h6fd == _T_221[11:0] ? 4'h0 : _GEN_23362; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23364 = 12'h6fe == _T_221[11:0] ? 4'h0 : _GEN_23363; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23365 = 12'h6ff == _T_221[11:0] ? 4'h0 : _GEN_23364; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23366 = 12'h700 == _T_221[11:0] ? 4'h0 : _GEN_23365; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23367 = 12'h701 == _T_221[11:0] ? image_1793 : _GEN_23366; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23368 = 12'h702 == _T_221[11:0] ? image_1794 : _GEN_23367; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23369 = 12'h703 == _T_221[11:0] ? image_1795 : _GEN_23368; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23370 = 12'h704 == _T_221[11:0] ? image_1796 : _GEN_23369; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23371 = 12'h705 == _T_221[11:0] ? image_1797 : _GEN_23370; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23372 = 12'h706 == _T_221[11:0] ? image_1798 : _GEN_23371; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23373 = 12'h707 == _T_221[11:0] ? image_1799 : _GEN_23372; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23374 = 12'h708 == _T_221[11:0] ? image_1800 : _GEN_23373; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23375 = 12'h709 == _T_221[11:0] ? image_1801 : _GEN_23374; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23376 = 12'h70a == _T_221[11:0] ? image_1802 : _GEN_23375; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23377 = 12'h70b == _T_221[11:0] ? image_1803 : _GEN_23376; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23378 = 12'h70c == _T_221[11:0] ? image_1804 : _GEN_23377; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23379 = 12'h70d == _T_221[11:0] ? image_1805 : _GEN_23378; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23380 = 12'h70e == _T_221[11:0] ? image_1806 : _GEN_23379; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23381 = 12'h70f == _T_221[11:0] ? image_1807 : _GEN_23380; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23382 = 12'h710 == _T_221[11:0] ? image_1808 : _GEN_23381; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23383 = 12'h711 == _T_221[11:0] ? image_1809 : _GEN_23382; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23384 = 12'h712 == _T_221[11:0] ? image_1810 : _GEN_23383; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23385 = 12'h713 == _T_221[11:0] ? image_1811 : _GEN_23384; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23386 = 12'h714 == _T_221[11:0] ? image_1812 : _GEN_23385; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23387 = 12'h715 == _T_221[11:0] ? image_1813 : _GEN_23386; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23388 = 12'h716 == _T_221[11:0] ? image_1814 : _GEN_23387; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23389 = 12'h717 == _T_221[11:0] ? image_1815 : _GEN_23388; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23390 = 12'h718 == _T_221[11:0] ? image_1816 : _GEN_23389; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23391 = 12'h719 == _T_221[11:0] ? image_1817 : _GEN_23390; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23392 = 12'h71a == _T_221[11:0] ? image_1818 : _GEN_23391; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23393 = 12'h71b == _T_221[11:0] ? image_1819 : _GEN_23392; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23394 = 12'h71c == _T_221[11:0] ? image_1820 : _GEN_23393; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23395 = 12'h71d == _T_221[11:0] ? image_1821 : _GEN_23394; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23396 = 12'h71e == _T_221[11:0] ? image_1822 : _GEN_23395; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23397 = 12'h71f == _T_221[11:0] ? image_1823 : _GEN_23396; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23398 = 12'h720 == _T_221[11:0] ? image_1824 : _GEN_23397; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23399 = 12'h721 == _T_221[11:0] ? image_1825 : _GEN_23398; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23400 = 12'h722 == _T_221[11:0] ? image_1826 : _GEN_23399; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23401 = 12'h723 == _T_221[11:0] ? image_1827 : _GEN_23400; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23402 = 12'h724 == _T_221[11:0] ? image_1828 : _GEN_23401; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23403 = 12'h725 == _T_221[11:0] ? image_1829 : _GEN_23402; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23404 = 12'h726 == _T_221[11:0] ? image_1830 : _GEN_23403; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23405 = 12'h727 == _T_221[11:0] ? image_1831 : _GEN_23404; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23406 = 12'h728 == _T_221[11:0] ? image_1832 : _GEN_23405; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23407 = 12'h729 == _T_221[11:0] ? image_1833 : _GEN_23406; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23408 = 12'h72a == _T_221[11:0] ? image_1834 : _GEN_23407; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23409 = 12'h72b == _T_221[11:0] ? image_1835 : _GEN_23408; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23410 = 12'h72c == _T_221[11:0] ? image_1836 : _GEN_23409; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23411 = 12'h72d == _T_221[11:0] ? image_1837 : _GEN_23410; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23412 = 12'h72e == _T_221[11:0] ? image_1838 : _GEN_23411; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23413 = 12'h72f == _T_221[11:0] ? image_1839 : _GEN_23412; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23414 = 12'h730 == _T_221[11:0] ? image_1840 : _GEN_23413; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23415 = 12'h731 == _T_221[11:0] ? image_1841 : _GEN_23414; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23416 = 12'h732 == _T_221[11:0] ? image_1842 : _GEN_23415; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23417 = 12'h733 == _T_221[11:0] ? image_1843 : _GEN_23416; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23418 = 12'h734 == _T_221[11:0] ? image_1844 : _GEN_23417; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23419 = 12'h735 == _T_221[11:0] ? image_1845 : _GEN_23418; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23420 = 12'h736 == _T_221[11:0] ? image_1846 : _GEN_23419; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23421 = 12'h737 == _T_221[11:0] ? image_1847 : _GEN_23420; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23422 = 12'h738 == _T_221[11:0] ? image_1848 : _GEN_23421; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23423 = 12'h739 == _T_221[11:0] ? image_1849 : _GEN_23422; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23424 = 12'h73a == _T_221[11:0] ? 4'h0 : _GEN_23423; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23425 = 12'h73b == _T_221[11:0] ? 4'h0 : _GEN_23424; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23426 = 12'h73c == _T_221[11:0] ? 4'h0 : _GEN_23425; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23427 = 12'h73d == _T_221[11:0] ? 4'h0 : _GEN_23426; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23428 = 12'h73e == _T_221[11:0] ? 4'h0 : _GEN_23427; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23429 = 12'h73f == _T_221[11:0] ? 4'h0 : _GEN_23428; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23430 = 12'h740 == _T_221[11:0] ? 4'h0 : _GEN_23429; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23431 = 12'h741 == _T_221[11:0] ? image_1857 : _GEN_23430; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23432 = 12'h742 == _T_221[11:0] ? image_1858 : _GEN_23431; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23433 = 12'h743 == _T_221[11:0] ? image_1859 : _GEN_23432; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23434 = 12'h744 == _T_221[11:0] ? image_1860 : _GEN_23433; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23435 = 12'h745 == _T_221[11:0] ? image_1861 : _GEN_23434; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23436 = 12'h746 == _T_221[11:0] ? image_1862 : _GEN_23435; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23437 = 12'h747 == _T_221[11:0] ? image_1863 : _GEN_23436; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23438 = 12'h748 == _T_221[11:0] ? image_1864 : _GEN_23437; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23439 = 12'h749 == _T_221[11:0] ? image_1865 : _GEN_23438; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23440 = 12'h74a == _T_221[11:0] ? image_1866 : _GEN_23439; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23441 = 12'h74b == _T_221[11:0] ? image_1867 : _GEN_23440; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23442 = 12'h74c == _T_221[11:0] ? image_1868 : _GEN_23441; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23443 = 12'h74d == _T_221[11:0] ? image_1869 : _GEN_23442; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23444 = 12'h74e == _T_221[11:0] ? image_1870 : _GEN_23443; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23445 = 12'h74f == _T_221[11:0] ? image_1871 : _GEN_23444; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23446 = 12'h750 == _T_221[11:0] ? image_1872 : _GEN_23445; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23447 = 12'h751 == _T_221[11:0] ? image_1873 : _GEN_23446; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23448 = 12'h752 == _T_221[11:0] ? image_1874 : _GEN_23447; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23449 = 12'h753 == _T_221[11:0] ? image_1875 : _GEN_23448; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23450 = 12'h754 == _T_221[11:0] ? image_1876 : _GEN_23449; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23451 = 12'h755 == _T_221[11:0] ? image_1877 : _GEN_23450; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23452 = 12'h756 == _T_221[11:0] ? image_1878 : _GEN_23451; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23453 = 12'h757 == _T_221[11:0] ? image_1879 : _GEN_23452; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23454 = 12'h758 == _T_221[11:0] ? image_1880 : _GEN_23453; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23455 = 12'h759 == _T_221[11:0] ? image_1881 : _GEN_23454; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23456 = 12'h75a == _T_221[11:0] ? image_1882 : _GEN_23455; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23457 = 12'h75b == _T_221[11:0] ? image_1883 : _GEN_23456; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23458 = 12'h75c == _T_221[11:0] ? image_1884 : _GEN_23457; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23459 = 12'h75d == _T_221[11:0] ? image_1885 : _GEN_23458; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23460 = 12'h75e == _T_221[11:0] ? image_1886 : _GEN_23459; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23461 = 12'h75f == _T_221[11:0] ? image_1887 : _GEN_23460; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23462 = 12'h760 == _T_221[11:0] ? image_1888 : _GEN_23461; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23463 = 12'h761 == _T_221[11:0] ? image_1889 : _GEN_23462; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23464 = 12'h762 == _T_221[11:0] ? image_1890 : _GEN_23463; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23465 = 12'h763 == _T_221[11:0] ? image_1891 : _GEN_23464; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23466 = 12'h764 == _T_221[11:0] ? image_1892 : _GEN_23465; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23467 = 12'h765 == _T_221[11:0] ? image_1893 : _GEN_23466; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23468 = 12'h766 == _T_221[11:0] ? image_1894 : _GEN_23467; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23469 = 12'h767 == _T_221[11:0] ? image_1895 : _GEN_23468; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23470 = 12'h768 == _T_221[11:0] ? image_1896 : _GEN_23469; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23471 = 12'h769 == _T_221[11:0] ? image_1897 : _GEN_23470; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23472 = 12'h76a == _T_221[11:0] ? image_1898 : _GEN_23471; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23473 = 12'h76b == _T_221[11:0] ? image_1899 : _GEN_23472; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23474 = 12'h76c == _T_221[11:0] ? image_1900 : _GEN_23473; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23475 = 12'h76d == _T_221[11:0] ? image_1901 : _GEN_23474; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23476 = 12'h76e == _T_221[11:0] ? image_1902 : _GEN_23475; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23477 = 12'h76f == _T_221[11:0] ? image_1903 : _GEN_23476; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23478 = 12'h770 == _T_221[11:0] ? image_1904 : _GEN_23477; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23479 = 12'h771 == _T_221[11:0] ? image_1905 : _GEN_23478; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23480 = 12'h772 == _T_221[11:0] ? image_1906 : _GEN_23479; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23481 = 12'h773 == _T_221[11:0] ? image_1907 : _GEN_23480; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23482 = 12'h774 == _T_221[11:0] ? image_1908 : _GEN_23481; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23483 = 12'h775 == _T_221[11:0] ? image_1909 : _GEN_23482; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23484 = 12'h776 == _T_221[11:0] ? image_1910 : _GEN_23483; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23485 = 12'h777 == _T_221[11:0] ? image_1911 : _GEN_23484; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23486 = 12'h778 == _T_221[11:0] ? image_1912 : _GEN_23485; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23487 = 12'h779 == _T_221[11:0] ? image_1913 : _GEN_23486; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23488 = 12'h77a == _T_221[11:0] ? 4'h0 : _GEN_23487; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23489 = 12'h77b == _T_221[11:0] ? 4'h0 : _GEN_23488; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23490 = 12'h77c == _T_221[11:0] ? 4'h0 : _GEN_23489; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23491 = 12'h77d == _T_221[11:0] ? 4'h0 : _GEN_23490; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23492 = 12'h77e == _T_221[11:0] ? 4'h0 : _GEN_23491; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23493 = 12'h77f == _T_221[11:0] ? 4'h0 : _GEN_23492; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23494 = 12'h780 == _T_221[11:0] ? 4'h0 : _GEN_23493; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23495 = 12'h781 == _T_221[11:0] ? image_1921 : _GEN_23494; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23496 = 12'h782 == _T_221[11:0] ? image_1922 : _GEN_23495; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23497 = 12'h783 == _T_221[11:0] ? image_1923 : _GEN_23496; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23498 = 12'h784 == _T_221[11:0] ? image_1924 : _GEN_23497; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23499 = 12'h785 == _T_221[11:0] ? image_1925 : _GEN_23498; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23500 = 12'h786 == _T_221[11:0] ? image_1926 : _GEN_23499; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23501 = 12'h787 == _T_221[11:0] ? image_1927 : _GEN_23500; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23502 = 12'h788 == _T_221[11:0] ? image_1928 : _GEN_23501; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23503 = 12'h789 == _T_221[11:0] ? image_1929 : _GEN_23502; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23504 = 12'h78a == _T_221[11:0] ? image_1930 : _GEN_23503; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23505 = 12'h78b == _T_221[11:0] ? image_1931 : _GEN_23504; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23506 = 12'h78c == _T_221[11:0] ? image_1932 : _GEN_23505; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23507 = 12'h78d == _T_221[11:0] ? image_1933 : _GEN_23506; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23508 = 12'h78e == _T_221[11:0] ? image_1934 : _GEN_23507; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23509 = 12'h78f == _T_221[11:0] ? image_1935 : _GEN_23508; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23510 = 12'h790 == _T_221[11:0] ? image_1936 : _GEN_23509; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23511 = 12'h791 == _T_221[11:0] ? image_1937 : _GEN_23510; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23512 = 12'h792 == _T_221[11:0] ? image_1938 : _GEN_23511; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23513 = 12'h793 == _T_221[11:0] ? image_1939 : _GEN_23512; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23514 = 12'h794 == _T_221[11:0] ? image_1940 : _GEN_23513; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23515 = 12'h795 == _T_221[11:0] ? image_1941 : _GEN_23514; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23516 = 12'h796 == _T_221[11:0] ? image_1942 : _GEN_23515; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23517 = 12'h797 == _T_221[11:0] ? image_1943 : _GEN_23516; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23518 = 12'h798 == _T_221[11:0] ? image_1944 : _GEN_23517; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23519 = 12'h799 == _T_221[11:0] ? image_1945 : _GEN_23518; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23520 = 12'h79a == _T_221[11:0] ? image_1946 : _GEN_23519; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23521 = 12'h79b == _T_221[11:0] ? image_1947 : _GEN_23520; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23522 = 12'h79c == _T_221[11:0] ? image_1948 : _GEN_23521; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23523 = 12'h79d == _T_221[11:0] ? image_1949 : _GEN_23522; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23524 = 12'h79e == _T_221[11:0] ? image_1950 : _GEN_23523; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23525 = 12'h79f == _T_221[11:0] ? image_1951 : _GEN_23524; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23526 = 12'h7a0 == _T_221[11:0] ? image_1952 : _GEN_23525; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23527 = 12'h7a1 == _T_221[11:0] ? image_1953 : _GEN_23526; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23528 = 12'h7a2 == _T_221[11:0] ? image_1954 : _GEN_23527; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23529 = 12'h7a3 == _T_221[11:0] ? image_1955 : _GEN_23528; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23530 = 12'h7a4 == _T_221[11:0] ? image_1956 : _GEN_23529; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23531 = 12'h7a5 == _T_221[11:0] ? image_1957 : _GEN_23530; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23532 = 12'h7a6 == _T_221[11:0] ? image_1958 : _GEN_23531; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23533 = 12'h7a7 == _T_221[11:0] ? image_1959 : _GEN_23532; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23534 = 12'h7a8 == _T_221[11:0] ? image_1960 : _GEN_23533; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23535 = 12'h7a9 == _T_221[11:0] ? image_1961 : _GEN_23534; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23536 = 12'h7aa == _T_221[11:0] ? image_1962 : _GEN_23535; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23537 = 12'h7ab == _T_221[11:0] ? image_1963 : _GEN_23536; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23538 = 12'h7ac == _T_221[11:0] ? image_1964 : _GEN_23537; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23539 = 12'h7ad == _T_221[11:0] ? image_1965 : _GEN_23538; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23540 = 12'h7ae == _T_221[11:0] ? image_1966 : _GEN_23539; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23541 = 12'h7af == _T_221[11:0] ? image_1967 : _GEN_23540; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23542 = 12'h7b0 == _T_221[11:0] ? image_1968 : _GEN_23541; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23543 = 12'h7b1 == _T_221[11:0] ? image_1969 : _GEN_23542; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23544 = 12'h7b2 == _T_221[11:0] ? image_1970 : _GEN_23543; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23545 = 12'h7b3 == _T_221[11:0] ? image_1971 : _GEN_23544; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23546 = 12'h7b4 == _T_221[11:0] ? image_1972 : _GEN_23545; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23547 = 12'h7b5 == _T_221[11:0] ? image_1973 : _GEN_23546; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23548 = 12'h7b6 == _T_221[11:0] ? image_1974 : _GEN_23547; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23549 = 12'h7b7 == _T_221[11:0] ? image_1975 : _GEN_23548; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23550 = 12'h7b8 == _T_221[11:0] ? image_1976 : _GEN_23549; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23551 = 12'h7b9 == _T_221[11:0] ? image_1977 : _GEN_23550; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23552 = 12'h7ba == _T_221[11:0] ? 4'h0 : _GEN_23551; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23553 = 12'h7bb == _T_221[11:0] ? 4'h0 : _GEN_23552; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23554 = 12'h7bc == _T_221[11:0] ? 4'h0 : _GEN_23553; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23555 = 12'h7bd == _T_221[11:0] ? 4'h0 : _GEN_23554; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23556 = 12'h7be == _T_221[11:0] ? 4'h0 : _GEN_23555; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23557 = 12'h7bf == _T_221[11:0] ? 4'h0 : _GEN_23556; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23558 = 12'h7c0 == _T_221[11:0] ? 4'h0 : _GEN_23557; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23559 = 12'h7c1 == _T_221[11:0] ? image_1985 : _GEN_23558; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23560 = 12'h7c2 == _T_221[11:0] ? image_1986 : _GEN_23559; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23561 = 12'h7c3 == _T_221[11:0] ? image_1987 : _GEN_23560; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23562 = 12'h7c4 == _T_221[11:0] ? image_1988 : _GEN_23561; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23563 = 12'h7c5 == _T_221[11:0] ? image_1989 : _GEN_23562; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23564 = 12'h7c6 == _T_221[11:0] ? image_1990 : _GEN_23563; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23565 = 12'h7c7 == _T_221[11:0] ? image_1991 : _GEN_23564; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23566 = 12'h7c8 == _T_221[11:0] ? image_1992 : _GEN_23565; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23567 = 12'h7c9 == _T_221[11:0] ? image_1993 : _GEN_23566; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23568 = 12'h7ca == _T_221[11:0] ? image_1994 : _GEN_23567; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23569 = 12'h7cb == _T_221[11:0] ? image_1995 : _GEN_23568; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23570 = 12'h7cc == _T_221[11:0] ? image_1996 : _GEN_23569; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23571 = 12'h7cd == _T_221[11:0] ? image_1997 : _GEN_23570; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23572 = 12'h7ce == _T_221[11:0] ? image_1998 : _GEN_23571; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23573 = 12'h7cf == _T_221[11:0] ? image_1999 : _GEN_23572; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23574 = 12'h7d0 == _T_221[11:0] ? image_2000 : _GEN_23573; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23575 = 12'h7d1 == _T_221[11:0] ? image_2001 : _GEN_23574; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23576 = 12'h7d2 == _T_221[11:0] ? image_2002 : _GEN_23575; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23577 = 12'h7d3 == _T_221[11:0] ? image_2003 : _GEN_23576; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23578 = 12'h7d4 == _T_221[11:0] ? image_2004 : _GEN_23577; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23579 = 12'h7d5 == _T_221[11:0] ? image_2005 : _GEN_23578; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23580 = 12'h7d6 == _T_221[11:0] ? image_2006 : _GEN_23579; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23581 = 12'h7d7 == _T_221[11:0] ? image_2007 : _GEN_23580; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23582 = 12'h7d8 == _T_221[11:0] ? image_2008 : _GEN_23581; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23583 = 12'h7d9 == _T_221[11:0] ? image_2009 : _GEN_23582; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23584 = 12'h7da == _T_221[11:0] ? image_2010 : _GEN_23583; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23585 = 12'h7db == _T_221[11:0] ? image_2011 : _GEN_23584; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23586 = 12'h7dc == _T_221[11:0] ? image_2012 : _GEN_23585; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23587 = 12'h7dd == _T_221[11:0] ? image_2013 : _GEN_23586; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23588 = 12'h7de == _T_221[11:0] ? image_2014 : _GEN_23587; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23589 = 12'h7df == _T_221[11:0] ? image_2015 : _GEN_23588; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23590 = 12'h7e0 == _T_221[11:0] ? image_2016 : _GEN_23589; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23591 = 12'h7e1 == _T_221[11:0] ? image_2017 : _GEN_23590; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23592 = 12'h7e2 == _T_221[11:0] ? image_2018 : _GEN_23591; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23593 = 12'h7e3 == _T_221[11:0] ? image_2019 : _GEN_23592; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23594 = 12'h7e4 == _T_221[11:0] ? image_2020 : _GEN_23593; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23595 = 12'h7e5 == _T_221[11:0] ? image_2021 : _GEN_23594; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23596 = 12'h7e6 == _T_221[11:0] ? image_2022 : _GEN_23595; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23597 = 12'h7e7 == _T_221[11:0] ? image_2023 : _GEN_23596; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23598 = 12'h7e8 == _T_221[11:0] ? image_2024 : _GEN_23597; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23599 = 12'h7e9 == _T_221[11:0] ? image_2025 : _GEN_23598; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23600 = 12'h7ea == _T_221[11:0] ? image_2026 : _GEN_23599; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23601 = 12'h7eb == _T_221[11:0] ? image_2027 : _GEN_23600; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23602 = 12'h7ec == _T_221[11:0] ? image_2028 : _GEN_23601; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23603 = 12'h7ed == _T_221[11:0] ? image_2029 : _GEN_23602; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23604 = 12'h7ee == _T_221[11:0] ? image_2030 : _GEN_23603; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23605 = 12'h7ef == _T_221[11:0] ? image_2031 : _GEN_23604; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23606 = 12'h7f0 == _T_221[11:0] ? image_2032 : _GEN_23605; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23607 = 12'h7f1 == _T_221[11:0] ? image_2033 : _GEN_23606; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23608 = 12'h7f2 == _T_221[11:0] ? image_2034 : _GEN_23607; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23609 = 12'h7f3 == _T_221[11:0] ? image_2035 : _GEN_23608; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23610 = 12'h7f4 == _T_221[11:0] ? image_2036 : _GEN_23609; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23611 = 12'h7f5 == _T_221[11:0] ? image_2037 : _GEN_23610; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23612 = 12'h7f6 == _T_221[11:0] ? image_2038 : _GEN_23611; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23613 = 12'h7f7 == _T_221[11:0] ? image_2039 : _GEN_23612; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23614 = 12'h7f8 == _T_221[11:0] ? image_2040 : _GEN_23613; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23615 = 12'h7f9 == _T_221[11:0] ? image_2041 : _GEN_23614; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23616 = 12'h7fa == _T_221[11:0] ? 4'h0 : _GEN_23615; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23617 = 12'h7fb == _T_221[11:0] ? 4'h0 : _GEN_23616; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23618 = 12'h7fc == _T_221[11:0] ? 4'h0 : _GEN_23617; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23619 = 12'h7fd == _T_221[11:0] ? 4'h0 : _GEN_23618; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23620 = 12'h7fe == _T_221[11:0] ? 4'h0 : _GEN_23619; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23621 = 12'h7ff == _T_221[11:0] ? 4'h0 : _GEN_23620; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23622 = 12'h800 == _T_221[11:0] ? 4'h0 : _GEN_23621; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23623 = 12'h801 == _T_221[11:0] ? image_2049 : _GEN_23622; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23624 = 12'h802 == _T_221[11:0] ? image_2050 : _GEN_23623; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23625 = 12'h803 == _T_221[11:0] ? image_2051 : _GEN_23624; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23626 = 12'h804 == _T_221[11:0] ? image_2052 : _GEN_23625; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23627 = 12'h805 == _T_221[11:0] ? image_2053 : _GEN_23626; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23628 = 12'h806 == _T_221[11:0] ? image_2054 : _GEN_23627; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23629 = 12'h807 == _T_221[11:0] ? image_2055 : _GEN_23628; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23630 = 12'h808 == _T_221[11:0] ? image_2056 : _GEN_23629; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23631 = 12'h809 == _T_221[11:0] ? image_2057 : _GEN_23630; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23632 = 12'h80a == _T_221[11:0] ? image_2058 : _GEN_23631; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23633 = 12'h80b == _T_221[11:0] ? image_2059 : _GEN_23632; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23634 = 12'h80c == _T_221[11:0] ? image_2060 : _GEN_23633; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23635 = 12'h80d == _T_221[11:0] ? image_2061 : _GEN_23634; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23636 = 12'h80e == _T_221[11:0] ? image_2062 : _GEN_23635; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23637 = 12'h80f == _T_221[11:0] ? image_2063 : _GEN_23636; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23638 = 12'h810 == _T_221[11:0] ? image_2064 : _GEN_23637; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23639 = 12'h811 == _T_221[11:0] ? image_2065 : _GEN_23638; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23640 = 12'h812 == _T_221[11:0] ? image_2066 : _GEN_23639; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23641 = 12'h813 == _T_221[11:0] ? image_2067 : _GEN_23640; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23642 = 12'h814 == _T_221[11:0] ? image_2068 : _GEN_23641; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23643 = 12'h815 == _T_221[11:0] ? image_2069 : _GEN_23642; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23644 = 12'h816 == _T_221[11:0] ? image_2070 : _GEN_23643; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23645 = 12'h817 == _T_221[11:0] ? image_2071 : _GEN_23644; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23646 = 12'h818 == _T_221[11:0] ? image_2072 : _GEN_23645; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23647 = 12'h819 == _T_221[11:0] ? image_2073 : _GEN_23646; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23648 = 12'h81a == _T_221[11:0] ? image_2074 : _GEN_23647; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23649 = 12'h81b == _T_221[11:0] ? image_2075 : _GEN_23648; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23650 = 12'h81c == _T_221[11:0] ? image_2076 : _GEN_23649; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23651 = 12'h81d == _T_221[11:0] ? image_2077 : _GEN_23650; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23652 = 12'h81e == _T_221[11:0] ? image_2078 : _GEN_23651; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23653 = 12'h81f == _T_221[11:0] ? image_2079 : _GEN_23652; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23654 = 12'h820 == _T_221[11:0] ? image_2080 : _GEN_23653; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23655 = 12'h821 == _T_221[11:0] ? image_2081 : _GEN_23654; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23656 = 12'h822 == _T_221[11:0] ? image_2082 : _GEN_23655; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23657 = 12'h823 == _T_221[11:0] ? image_2083 : _GEN_23656; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23658 = 12'h824 == _T_221[11:0] ? image_2084 : _GEN_23657; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23659 = 12'h825 == _T_221[11:0] ? image_2085 : _GEN_23658; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23660 = 12'h826 == _T_221[11:0] ? image_2086 : _GEN_23659; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23661 = 12'h827 == _T_221[11:0] ? image_2087 : _GEN_23660; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23662 = 12'h828 == _T_221[11:0] ? image_2088 : _GEN_23661; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23663 = 12'h829 == _T_221[11:0] ? image_2089 : _GEN_23662; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23664 = 12'h82a == _T_221[11:0] ? image_2090 : _GEN_23663; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23665 = 12'h82b == _T_221[11:0] ? image_2091 : _GEN_23664; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23666 = 12'h82c == _T_221[11:0] ? image_2092 : _GEN_23665; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23667 = 12'h82d == _T_221[11:0] ? image_2093 : _GEN_23666; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23668 = 12'h82e == _T_221[11:0] ? image_2094 : _GEN_23667; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23669 = 12'h82f == _T_221[11:0] ? image_2095 : _GEN_23668; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23670 = 12'h830 == _T_221[11:0] ? image_2096 : _GEN_23669; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23671 = 12'h831 == _T_221[11:0] ? image_2097 : _GEN_23670; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23672 = 12'h832 == _T_221[11:0] ? image_2098 : _GEN_23671; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23673 = 12'h833 == _T_221[11:0] ? image_2099 : _GEN_23672; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23674 = 12'h834 == _T_221[11:0] ? image_2100 : _GEN_23673; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23675 = 12'h835 == _T_221[11:0] ? image_2101 : _GEN_23674; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23676 = 12'h836 == _T_221[11:0] ? image_2102 : _GEN_23675; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23677 = 12'h837 == _T_221[11:0] ? image_2103 : _GEN_23676; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23678 = 12'h838 == _T_221[11:0] ? image_2104 : _GEN_23677; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23679 = 12'h839 == _T_221[11:0] ? image_2105 : _GEN_23678; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23680 = 12'h83a == _T_221[11:0] ? image_2106 : _GEN_23679; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23681 = 12'h83b == _T_221[11:0] ? 4'h0 : _GEN_23680; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23682 = 12'h83c == _T_221[11:0] ? 4'h0 : _GEN_23681; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23683 = 12'h83d == _T_221[11:0] ? 4'h0 : _GEN_23682; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23684 = 12'h83e == _T_221[11:0] ? 4'h0 : _GEN_23683; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23685 = 12'h83f == _T_221[11:0] ? 4'h0 : _GEN_23684; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23686 = 12'h840 == _T_221[11:0] ? 4'h0 : _GEN_23685; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23687 = 12'h841 == _T_221[11:0] ? 4'h0 : _GEN_23686; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23688 = 12'h842 == _T_221[11:0] ? image_2114 : _GEN_23687; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23689 = 12'h843 == _T_221[11:0] ? image_2115 : _GEN_23688; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23690 = 12'h844 == _T_221[11:0] ? image_2116 : _GEN_23689; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23691 = 12'h845 == _T_221[11:0] ? image_2117 : _GEN_23690; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23692 = 12'h846 == _T_221[11:0] ? image_2118 : _GEN_23691; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23693 = 12'h847 == _T_221[11:0] ? image_2119 : _GEN_23692; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23694 = 12'h848 == _T_221[11:0] ? image_2120 : _GEN_23693; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23695 = 12'h849 == _T_221[11:0] ? image_2121 : _GEN_23694; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23696 = 12'h84a == _T_221[11:0] ? image_2122 : _GEN_23695; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23697 = 12'h84b == _T_221[11:0] ? image_2123 : _GEN_23696; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23698 = 12'h84c == _T_221[11:0] ? image_2124 : _GEN_23697; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23699 = 12'h84d == _T_221[11:0] ? image_2125 : _GEN_23698; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23700 = 12'h84e == _T_221[11:0] ? image_2126 : _GEN_23699; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23701 = 12'h84f == _T_221[11:0] ? image_2127 : _GEN_23700; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23702 = 12'h850 == _T_221[11:0] ? image_2128 : _GEN_23701; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23703 = 12'h851 == _T_221[11:0] ? image_2129 : _GEN_23702; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23704 = 12'h852 == _T_221[11:0] ? image_2130 : _GEN_23703; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23705 = 12'h853 == _T_221[11:0] ? image_2131 : _GEN_23704; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23706 = 12'h854 == _T_221[11:0] ? image_2132 : _GEN_23705; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23707 = 12'h855 == _T_221[11:0] ? image_2133 : _GEN_23706; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23708 = 12'h856 == _T_221[11:0] ? image_2134 : _GEN_23707; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23709 = 12'h857 == _T_221[11:0] ? image_2135 : _GEN_23708; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23710 = 12'h858 == _T_221[11:0] ? image_2136 : _GEN_23709; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23711 = 12'h859 == _T_221[11:0] ? image_2137 : _GEN_23710; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23712 = 12'h85a == _T_221[11:0] ? image_2138 : _GEN_23711; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23713 = 12'h85b == _T_221[11:0] ? image_2139 : _GEN_23712; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23714 = 12'h85c == _T_221[11:0] ? image_2140 : _GEN_23713; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23715 = 12'h85d == _T_221[11:0] ? image_2141 : _GEN_23714; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23716 = 12'h85e == _T_221[11:0] ? image_2142 : _GEN_23715; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23717 = 12'h85f == _T_221[11:0] ? image_2143 : _GEN_23716; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23718 = 12'h860 == _T_221[11:0] ? image_2144 : _GEN_23717; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23719 = 12'h861 == _T_221[11:0] ? image_2145 : _GEN_23718; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23720 = 12'h862 == _T_221[11:0] ? image_2146 : _GEN_23719; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23721 = 12'h863 == _T_221[11:0] ? image_2147 : _GEN_23720; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23722 = 12'h864 == _T_221[11:0] ? image_2148 : _GEN_23721; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23723 = 12'h865 == _T_221[11:0] ? image_2149 : _GEN_23722; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23724 = 12'h866 == _T_221[11:0] ? image_2150 : _GEN_23723; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23725 = 12'h867 == _T_221[11:0] ? image_2151 : _GEN_23724; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23726 = 12'h868 == _T_221[11:0] ? image_2152 : _GEN_23725; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23727 = 12'h869 == _T_221[11:0] ? image_2153 : _GEN_23726; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23728 = 12'h86a == _T_221[11:0] ? image_2154 : _GEN_23727; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23729 = 12'h86b == _T_221[11:0] ? image_2155 : _GEN_23728; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23730 = 12'h86c == _T_221[11:0] ? image_2156 : _GEN_23729; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23731 = 12'h86d == _T_221[11:0] ? image_2157 : _GEN_23730; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23732 = 12'h86e == _T_221[11:0] ? image_2158 : _GEN_23731; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23733 = 12'h86f == _T_221[11:0] ? image_2159 : _GEN_23732; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23734 = 12'h870 == _T_221[11:0] ? image_2160 : _GEN_23733; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23735 = 12'h871 == _T_221[11:0] ? image_2161 : _GEN_23734; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23736 = 12'h872 == _T_221[11:0] ? image_2162 : _GEN_23735; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23737 = 12'h873 == _T_221[11:0] ? image_2163 : _GEN_23736; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23738 = 12'h874 == _T_221[11:0] ? image_2164 : _GEN_23737; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23739 = 12'h875 == _T_221[11:0] ? image_2165 : _GEN_23738; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23740 = 12'h876 == _T_221[11:0] ? image_2166 : _GEN_23739; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23741 = 12'h877 == _T_221[11:0] ? image_2167 : _GEN_23740; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23742 = 12'h878 == _T_221[11:0] ? image_2168 : _GEN_23741; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23743 = 12'h879 == _T_221[11:0] ? image_2169 : _GEN_23742; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23744 = 12'h87a == _T_221[11:0] ? image_2170 : _GEN_23743; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23745 = 12'h87b == _T_221[11:0] ? 4'h0 : _GEN_23744; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23746 = 12'h87c == _T_221[11:0] ? 4'h0 : _GEN_23745; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23747 = 12'h87d == _T_221[11:0] ? 4'h0 : _GEN_23746; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23748 = 12'h87e == _T_221[11:0] ? 4'h0 : _GEN_23747; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23749 = 12'h87f == _T_221[11:0] ? 4'h0 : _GEN_23748; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23750 = 12'h880 == _T_221[11:0] ? 4'h0 : _GEN_23749; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23751 = 12'h881 == _T_221[11:0] ? image_2177 : _GEN_23750; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23752 = 12'h882 == _T_221[11:0] ? image_2178 : _GEN_23751; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23753 = 12'h883 == _T_221[11:0] ? image_2179 : _GEN_23752; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23754 = 12'h884 == _T_221[11:0] ? image_2180 : _GEN_23753; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23755 = 12'h885 == _T_221[11:0] ? image_2181 : _GEN_23754; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23756 = 12'h886 == _T_221[11:0] ? image_2182 : _GEN_23755; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23757 = 12'h887 == _T_221[11:0] ? image_2183 : _GEN_23756; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23758 = 12'h888 == _T_221[11:0] ? image_2184 : _GEN_23757; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23759 = 12'h889 == _T_221[11:0] ? image_2185 : _GEN_23758; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23760 = 12'h88a == _T_221[11:0] ? image_2186 : _GEN_23759; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23761 = 12'h88b == _T_221[11:0] ? image_2187 : _GEN_23760; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23762 = 12'h88c == _T_221[11:0] ? image_2188 : _GEN_23761; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23763 = 12'h88d == _T_221[11:0] ? image_2189 : _GEN_23762; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23764 = 12'h88e == _T_221[11:0] ? image_2190 : _GEN_23763; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23765 = 12'h88f == _T_221[11:0] ? image_2191 : _GEN_23764; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23766 = 12'h890 == _T_221[11:0] ? image_2192 : _GEN_23765; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23767 = 12'h891 == _T_221[11:0] ? image_2193 : _GEN_23766; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23768 = 12'h892 == _T_221[11:0] ? image_2194 : _GEN_23767; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23769 = 12'h893 == _T_221[11:0] ? image_2195 : _GEN_23768; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23770 = 12'h894 == _T_221[11:0] ? image_2196 : _GEN_23769; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23771 = 12'h895 == _T_221[11:0] ? image_2197 : _GEN_23770; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23772 = 12'h896 == _T_221[11:0] ? image_2198 : _GEN_23771; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23773 = 12'h897 == _T_221[11:0] ? image_2199 : _GEN_23772; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23774 = 12'h898 == _T_221[11:0] ? image_2200 : _GEN_23773; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23775 = 12'h899 == _T_221[11:0] ? image_2201 : _GEN_23774; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23776 = 12'h89a == _T_221[11:0] ? image_2202 : _GEN_23775; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23777 = 12'h89b == _T_221[11:0] ? image_2203 : _GEN_23776; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23778 = 12'h89c == _T_221[11:0] ? image_2204 : _GEN_23777; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23779 = 12'h89d == _T_221[11:0] ? image_2205 : _GEN_23778; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23780 = 12'h89e == _T_221[11:0] ? image_2206 : _GEN_23779; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23781 = 12'h89f == _T_221[11:0] ? image_2207 : _GEN_23780; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23782 = 12'h8a0 == _T_221[11:0] ? image_2208 : _GEN_23781; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23783 = 12'h8a1 == _T_221[11:0] ? image_2209 : _GEN_23782; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23784 = 12'h8a2 == _T_221[11:0] ? image_2210 : _GEN_23783; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23785 = 12'h8a3 == _T_221[11:0] ? image_2211 : _GEN_23784; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23786 = 12'h8a4 == _T_221[11:0] ? image_2212 : _GEN_23785; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23787 = 12'h8a5 == _T_221[11:0] ? image_2213 : _GEN_23786; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23788 = 12'h8a6 == _T_221[11:0] ? image_2214 : _GEN_23787; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23789 = 12'h8a7 == _T_221[11:0] ? image_2215 : _GEN_23788; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23790 = 12'h8a8 == _T_221[11:0] ? image_2216 : _GEN_23789; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23791 = 12'h8a9 == _T_221[11:0] ? image_2217 : _GEN_23790; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23792 = 12'h8aa == _T_221[11:0] ? image_2218 : _GEN_23791; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23793 = 12'h8ab == _T_221[11:0] ? image_2219 : _GEN_23792; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23794 = 12'h8ac == _T_221[11:0] ? image_2220 : _GEN_23793; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23795 = 12'h8ad == _T_221[11:0] ? image_2221 : _GEN_23794; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23796 = 12'h8ae == _T_221[11:0] ? image_2222 : _GEN_23795; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23797 = 12'h8af == _T_221[11:0] ? image_2223 : _GEN_23796; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23798 = 12'h8b0 == _T_221[11:0] ? image_2224 : _GEN_23797; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23799 = 12'h8b1 == _T_221[11:0] ? image_2225 : _GEN_23798; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23800 = 12'h8b2 == _T_221[11:0] ? image_2226 : _GEN_23799; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23801 = 12'h8b3 == _T_221[11:0] ? image_2227 : _GEN_23800; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23802 = 12'h8b4 == _T_221[11:0] ? image_2228 : _GEN_23801; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23803 = 12'h8b5 == _T_221[11:0] ? image_2229 : _GEN_23802; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23804 = 12'h8b6 == _T_221[11:0] ? image_2230 : _GEN_23803; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23805 = 12'h8b7 == _T_221[11:0] ? image_2231 : _GEN_23804; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23806 = 12'h8b8 == _T_221[11:0] ? image_2232 : _GEN_23805; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23807 = 12'h8b9 == _T_221[11:0] ? image_2233 : _GEN_23806; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23808 = 12'h8ba == _T_221[11:0] ? image_2234 : _GEN_23807; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23809 = 12'h8bb == _T_221[11:0] ? 4'h0 : _GEN_23808; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23810 = 12'h8bc == _T_221[11:0] ? 4'h0 : _GEN_23809; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23811 = 12'h8bd == _T_221[11:0] ? 4'h0 : _GEN_23810; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23812 = 12'h8be == _T_221[11:0] ? 4'h0 : _GEN_23811; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23813 = 12'h8bf == _T_221[11:0] ? 4'h0 : _GEN_23812; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23814 = 12'h8c0 == _T_221[11:0] ? 4'h0 : _GEN_23813; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23815 = 12'h8c1 == _T_221[11:0] ? 4'h0 : _GEN_23814; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23816 = 12'h8c2 == _T_221[11:0] ? 4'h0 : _GEN_23815; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23817 = 12'h8c3 == _T_221[11:0] ? image_2243 : _GEN_23816; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23818 = 12'h8c4 == _T_221[11:0] ? image_2244 : _GEN_23817; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23819 = 12'h8c5 == _T_221[11:0] ? image_2245 : _GEN_23818; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23820 = 12'h8c6 == _T_221[11:0] ? image_2246 : _GEN_23819; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23821 = 12'h8c7 == _T_221[11:0] ? image_2247 : _GEN_23820; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23822 = 12'h8c8 == _T_221[11:0] ? image_2248 : _GEN_23821; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23823 = 12'h8c9 == _T_221[11:0] ? image_2249 : _GEN_23822; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23824 = 12'h8ca == _T_221[11:0] ? image_2250 : _GEN_23823; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23825 = 12'h8cb == _T_221[11:0] ? image_2251 : _GEN_23824; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23826 = 12'h8cc == _T_221[11:0] ? image_2252 : _GEN_23825; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23827 = 12'h8cd == _T_221[11:0] ? image_2253 : _GEN_23826; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23828 = 12'h8ce == _T_221[11:0] ? image_2254 : _GEN_23827; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23829 = 12'h8cf == _T_221[11:0] ? image_2255 : _GEN_23828; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23830 = 12'h8d0 == _T_221[11:0] ? image_2256 : _GEN_23829; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23831 = 12'h8d1 == _T_221[11:0] ? image_2257 : _GEN_23830; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23832 = 12'h8d2 == _T_221[11:0] ? image_2258 : _GEN_23831; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23833 = 12'h8d3 == _T_221[11:0] ? image_2259 : _GEN_23832; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23834 = 12'h8d4 == _T_221[11:0] ? image_2260 : _GEN_23833; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23835 = 12'h8d5 == _T_221[11:0] ? image_2261 : _GEN_23834; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23836 = 12'h8d6 == _T_221[11:0] ? image_2262 : _GEN_23835; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23837 = 12'h8d7 == _T_221[11:0] ? image_2263 : _GEN_23836; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23838 = 12'h8d8 == _T_221[11:0] ? image_2264 : _GEN_23837; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23839 = 12'h8d9 == _T_221[11:0] ? image_2265 : _GEN_23838; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23840 = 12'h8da == _T_221[11:0] ? image_2266 : _GEN_23839; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23841 = 12'h8db == _T_221[11:0] ? image_2267 : _GEN_23840; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23842 = 12'h8dc == _T_221[11:0] ? image_2268 : _GEN_23841; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23843 = 12'h8dd == _T_221[11:0] ? image_2269 : _GEN_23842; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23844 = 12'h8de == _T_221[11:0] ? image_2270 : _GEN_23843; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23845 = 12'h8df == _T_221[11:0] ? image_2271 : _GEN_23844; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23846 = 12'h8e0 == _T_221[11:0] ? image_2272 : _GEN_23845; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23847 = 12'h8e1 == _T_221[11:0] ? image_2273 : _GEN_23846; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23848 = 12'h8e2 == _T_221[11:0] ? image_2274 : _GEN_23847; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23849 = 12'h8e3 == _T_221[11:0] ? image_2275 : _GEN_23848; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23850 = 12'h8e4 == _T_221[11:0] ? image_2276 : _GEN_23849; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23851 = 12'h8e5 == _T_221[11:0] ? image_2277 : _GEN_23850; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23852 = 12'h8e6 == _T_221[11:0] ? image_2278 : _GEN_23851; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23853 = 12'h8e7 == _T_221[11:0] ? image_2279 : _GEN_23852; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23854 = 12'h8e8 == _T_221[11:0] ? image_2280 : _GEN_23853; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23855 = 12'h8e9 == _T_221[11:0] ? image_2281 : _GEN_23854; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23856 = 12'h8ea == _T_221[11:0] ? image_2282 : _GEN_23855; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23857 = 12'h8eb == _T_221[11:0] ? image_2283 : _GEN_23856; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23858 = 12'h8ec == _T_221[11:0] ? image_2284 : _GEN_23857; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23859 = 12'h8ed == _T_221[11:0] ? image_2285 : _GEN_23858; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23860 = 12'h8ee == _T_221[11:0] ? image_2286 : _GEN_23859; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23861 = 12'h8ef == _T_221[11:0] ? image_2287 : _GEN_23860; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23862 = 12'h8f0 == _T_221[11:0] ? image_2288 : _GEN_23861; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23863 = 12'h8f1 == _T_221[11:0] ? image_2289 : _GEN_23862; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23864 = 12'h8f2 == _T_221[11:0] ? image_2290 : _GEN_23863; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23865 = 12'h8f3 == _T_221[11:0] ? image_2291 : _GEN_23864; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23866 = 12'h8f4 == _T_221[11:0] ? image_2292 : _GEN_23865; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23867 = 12'h8f5 == _T_221[11:0] ? image_2293 : _GEN_23866; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23868 = 12'h8f6 == _T_221[11:0] ? image_2294 : _GEN_23867; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23869 = 12'h8f7 == _T_221[11:0] ? image_2295 : _GEN_23868; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23870 = 12'h8f8 == _T_221[11:0] ? image_2296 : _GEN_23869; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23871 = 12'h8f9 == _T_221[11:0] ? image_2297 : _GEN_23870; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23872 = 12'h8fa == _T_221[11:0] ? image_2298 : _GEN_23871; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23873 = 12'h8fb == _T_221[11:0] ? 4'h0 : _GEN_23872; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23874 = 12'h8fc == _T_221[11:0] ? 4'h0 : _GEN_23873; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23875 = 12'h8fd == _T_221[11:0] ? 4'h0 : _GEN_23874; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23876 = 12'h8fe == _T_221[11:0] ? 4'h0 : _GEN_23875; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23877 = 12'h8ff == _T_221[11:0] ? 4'h0 : _GEN_23876; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23878 = 12'h900 == _T_221[11:0] ? 4'h0 : _GEN_23877; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23879 = 12'h901 == _T_221[11:0] ? 4'h0 : _GEN_23878; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23880 = 12'h902 == _T_221[11:0] ? 4'h0 : _GEN_23879; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23881 = 12'h903 == _T_221[11:0] ? image_2307 : _GEN_23880; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23882 = 12'h904 == _T_221[11:0] ? image_2308 : _GEN_23881; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23883 = 12'h905 == _T_221[11:0] ? image_2309 : _GEN_23882; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23884 = 12'h906 == _T_221[11:0] ? image_2310 : _GEN_23883; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23885 = 12'h907 == _T_221[11:0] ? image_2311 : _GEN_23884; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23886 = 12'h908 == _T_221[11:0] ? image_2312 : _GEN_23885; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23887 = 12'h909 == _T_221[11:0] ? image_2313 : _GEN_23886; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23888 = 12'h90a == _T_221[11:0] ? image_2314 : _GEN_23887; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23889 = 12'h90b == _T_221[11:0] ? image_2315 : _GEN_23888; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23890 = 12'h90c == _T_221[11:0] ? image_2316 : _GEN_23889; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23891 = 12'h90d == _T_221[11:0] ? image_2317 : _GEN_23890; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23892 = 12'h90e == _T_221[11:0] ? image_2318 : _GEN_23891; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23893 = 12'h90f == _T_221[11:0] ? image_2319 : _GEN_23892; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23894 = 12'h910 == _T_221[11:0] ? image_2320 : _GEN_23893; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23895 = 12'h911 == _T_221[11:0] ? image_2321 : _GEN_23894; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23896 = 12'h912 == _T_221[11:0] ? image_2322 : _GEN_23895; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23897 = 12'h913 == _T_221[11:0] ? image_2323 : _GEN_23896; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23898 = 12'h914 == _T_221[11:0] ? image_2324 : _GEN_23897; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23899 = 12'h915 == _T_221[11:0] ? image_2325 : _GEN_23898; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23900 = 12'h916 == _T_221[11:0] ? image_2326 : _GEN_23899; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23901 = 12'h917 == _T_221[11:0] ? image_2327 : _GEN_23900; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23902 = 12'h918 == _T_221[11:0] ? image_2328 : _GEN_23901; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23903 = 12'h919 == _T_221[11:0] ? image_2329 : _GEN_23902; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23904 = 12'h91a == _T_221[11:0] ? image_2330 : _GEN_23903; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23905 = 12'h91b == _T_221[11:0] ? image_2331 : _GEN_23904; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23906 = 12'h91c == _T_221[11:0] ? image_2332 : _GEN_23905; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23907 = 12'h91d == _T_221[11:0] ? image_2333 : _GEN_23906; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23908 = 12'h91e == _T_221[11:0] ? image_2334 : _GEN_23907; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23909 = 12'h91f == _T_221[11:0] ? image_2335 : _GEN_23908; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23910 = 12'h920 == _T_221[11:0] ? image_2336 : _GEN_23909; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23911 = 12'h921 == _T_221[11:0] ? image_2337 : _GEN_23910; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23912 = 12'h922 == _T_221[11:0] ? image_2338 : _GEN_23911; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23913 = 12'h923 == _T_221[11:0] ? image_2339 : _GEN_23912; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23914 = 12'h924 == _T_221[11:0] ? image_2340 : _GEN_23913; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23915 = 12'h925 == _T_221[11:0] ? image_2341 : _GEN_23914; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23916 = 12'h926 == _T_221[11:0] ? image_2342 : _GEN_23915; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23917 = 12'h927 == _T_221[11:0] ? image_2343 : _GEN_23916; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23918 = 12'h928 == _T_221[11:0] ? image_2344 : _GEN_23917; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23919 = 12'h929 == _T_221[11:0] ? image_2345 : _GEN_23918; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23920 = 12'h92a == _T_221[11:0] ? image_2346 : _GEN_23919; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23921 = 12'h92b == _T_221[11:0] ? image_2347 : _GEN_23920; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23922 = 12'h92c == _T_221[11:0] ? image_2348 : _GEN_23921; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23923 = 12'h92d == _T_221[11:0] ? image_2349 : _GEN_23922; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23924 = 12'h92e == _T_221[11:0] ? image_2350 : _GEN_23923; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23925 = 12'h92f == _T_221[11:0] ? image_2351 : _GEN_23924; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23926 = 12'h930 == _T_221[11:0] ? image_2352 : _GEN_23925; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23927 = 12'h931 == _T_221[11:0] ? image_2353 : _GEN_23926; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23928 = 12'h932 == _T_221[11:0] ? image_2354 : _GEN_23927; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23929 = 12'h933 == _T_221[11:0] ? image_2355 : _GEN_23928; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23930 = 12'h934 == _T_221[11:0] ? image_2356 : _GEN_23929; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23931 = 12'h935 == _T_221[11:0] ? image_2357 : _GEN_23930; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23932 = 12'h936 == _T_221[11:0] ? image_2358 : _GEN_23931; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23933 = 12'h937 == _T_221[11:0] ? image_2359 : _GEN_23932; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23934 = 12'h938 == _T_221[11:0] ? image_2360 : _GEN_23933; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23935 = 12'h939 == _T_221[11:0] ? image_2361 : _GEN_23934; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23936 = 12'h93a == _T_221[11:0] ? image_2362 : _GEN_23935; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23937 = 12'h93b == _T_221[11:0] ? 4'h0 : _GEN_23936; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23938 = 12'h93c == _T_221[11:0] ? 4'h0 : _GEN_23937; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23939 = 12'h93d == _T_221[11:0] ? 4'h0 : _GEN_23938; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23940 = 12'h93e == _T_221[11:0] ? 4'h0 : _GEN_23939; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23941 = 12'h93f == _T_221[11:0] ? 4'h0 : _GEN_23940; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23942 = 12'h940 == _T_221[11:0] ? 4'h0 : _GEN_23941; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23943 = 12'h941 == _T_221[11:0] ? 4'h0 : _GEN_23942; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23944 = 12'h942 == _T_221[11:0] ? 4'h0 : _GEN_23943; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23945 = 12'h943 == _T_221[11:0] ? 4'h0 : _GEN_23944; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23946 = 12'h944 == _T_221[11:0] ? image_2372 : _GEN_23945; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23947 = 12'h945 == _T_221[11:0] ? image_2373 : _GEN_23946; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23948 = 12'h946 == _T_221[11:0] ? image_2374 : _GEN_23947; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23949 = 12'h947 == _T_221[11:0] ? image_2375 : _GEN_23948; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23950 = 12'h948 == _T_221[11:0] ? image_2376 : _GEN_23949; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23951 = 12'h949 == _T_221[11:0] ? image_2377 : _GEN_23950; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23952 = 12'h94a == _T_221[11:0] ? image_2378 : _GEN_23951; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23953 = 12'h94b == _T_221[11:0] ? image_2379 : _GEN_23952; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23954 = 12'h94c == _T_221[11:0] ? image_2380 : _GEN_23953; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23955 = 12'h94d == _T_221[11:0] ? image_2381 : _GEN_23954; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23956 = 12'h94e == _T_221[11:0] ? image_2382 : _GEN_23955; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23957 = 12'h94f == _T_221[11:0] ? image_2383 : _GEN_23956; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23958 = 12'h950 == _T_221[11:0] ? image_2384 : _GEN_23957; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23959 = 12'h951 == _T_221[11:0] ? image_2385 : _GEN_23958; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23960 = 12'h952 == _T_221[11:0] ? image_2386 : _GEN_23959; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23961 = 12'h953 == _T_221[11:0] ? image_2387 : _GEN_23960; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23962 = 12'h954 == _T_221[11:0] ? image_2388 : _GEN_23961; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23963 = 12'h955 == _T_221[11:0] ? image_2389 : _GEN_23962; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23964 = 12'h956 == _T_221[11:0] ? image_2390 : _GEN_23963; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23965 = 12'h957 == _T_221[11:0] ? image_2391 : _GEN_23964; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23966 = 12'h958 == _T_221[11:0] ? image_2392 : _GEN_23965; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23967 = 12'h959 == _T_221[11:0] ? image_2393 : _GEN_23966; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23968 = 12'h95a == _T_221[11:0] ? image_2394 : _GEN_23967; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23969 = 12'h95b == _T_221[11:0] ? image_2395 : _GEN_23968; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23970 = 12'h95c == _T_221[11:0] ? image_2396 : _GEN_23969; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23971 = 12'h95d == _T_221[11:0] ? image_2397 : _GEN_23970; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23972 = 12'h95e == _T_221[11:0] ? image_2398 : _GEN_23971; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23973 = 12'h95f == _T_221[11:0] ? image_2399 : _GEN_23972; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23974 = 12'h960 == _T_221[11:0] ? image_2400 : _GEN_23973; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23975 = 12'h961 == _T_221[11:0] ? image_2401 : _GEN_23974; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23976 = 12'h962 == _T_221[11:0] ? image_2402 : _GEN_23975; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23977 = 12'h963 == _T_221[11:0] ? image_2403 : _GEN_23976; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23978 = 12'h964 == _T_221[11:0] ? image_2404 : _GEN_23977; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23979 = 12'h965 == _T_221[11:0] ? image_2405 : _GEN_23978; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23980 = 12'h966 == _T_221[11:0] ? image_2406 : _GEN_23979; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23981 = 12'h967 == _T_221[11:0] ? image_2407 : _GEN_23980; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23982 = 12'h968 == _T_221[11:0] ? image_2408 : _GEN_23981; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23983 = 12'h969 == _T_221[11:0] ? image_2409 : _GEN_23982; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23984 = 12'h96a == _T_221[11:0] ? image_2410 : _GEN_23983; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23985 = 12'h96b == _T_221[11:0] ? image_2411 : _GEN_23984; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23986 = 12'h96c == _T_221[11:0] ? image_2412 : _GEN_23985; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23987 = 12'h96d == _T_221[11:0] ? image_2413 : _GEN_23986; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23988 = 12'h96e == _T_221[11:0] ? image_2414 : _GEN_23987; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23989 = 12'h96f == _T_221[11:0] ? image_2415 : _GEN_23988; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23990 = 12'h970 == _T_221[11:0] ? image_2416 : _GEN_23989; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23991 = 12'h971 == _T_221[11:0] ? image_2417 : _GEN_23990; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23992 = 12'h972 == _T_221[11:0] ? image_2418 : _GEN_23991; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23993 = 12'h973 == _T_221[11:0] ? image_2419 : _GEN_23992; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23994 = 12'h974 == _T_221[11:0] ? image_2420 : _GEN_23993; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23995 = 12'h975 == _T_221[11:0] ? image_2421 : _GEN_23994; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23996 = 12'h976 == _T_221[11:0] ? image_2422 : _GEN_23995; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23997 = 12'h977 == _T_221[11:0] ? image_2423 : _GEN_23996; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23998 = 12'h978 == _T_221[11:0] ? image_2424 : _GEN_23997; // @[Filter.scala 138:46]
  wire [3:0] _GEN_23999 = 12'h979 == _T_221[11:0] ? image_2425 : _GEN_23998; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24000 = 12'h97a == _T_221[11:0] ? image_2426 : _GEN_23999; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24001 = 12'h97b == _T_221[11:0] ? 4'h0 : _GEN_24000; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24002 = 12'h97c == _T_221[11:0] ? 4'h0 : _GEN_24001; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24003 = 12'h97d == _T_221[11:0] ? 4'h0 : _GEN_24002; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24004 = 12'h97e == _T_221[11:0] ? 4'h0 : _GEN_24003; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24005 = 12'h97f == _T_221[11:0] ? 4'h0 : _GEN_24004; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24006 = 12'h980 == _T_221[11:0] ? 4'h0 : _GEN_24005; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24007 = 12'h981 == _T_221[11:0] ? 4'h0 : _GEN_24006; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24008 = 12'h982 == _T_221[11:0] ? 4'h0 : _GEN_24007; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24009 = 12'h983 == _T_221[11:0] ? 4'h0 : _GEN_24008; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24010 = 12'h984 == _T_221[11:0] ? 4'h0 : _GEN_24009; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24011 = 12'h985 == _T_221[11:0] ? image_2437 : _GEN_24010; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24012 = 12'h986 == _T_221[11:0] ? image_2438 : _GEN_24011; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24013 = 12'h987 == _T_221[11:0] ? image_2439 : _GEN_24012; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24014 = 12'h988 == _T_221[11:0] ? image_2440 : _GEN_24013; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24015 = 12'h989 == _T_221[11:0] ? image_2441 : _GEN_24014; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24016 = 12'h98a == _T_221[11:0] ? image_2442 : _GEN_24015; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24017 = 12'h98b == _T_221[11:0] ? image_2443 : _GEN_24016; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24018 = 12'h98c == _T_221[11:0] ? image_2444 : _GEN_24017; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24019 = 12'h98d == _T_221[11:0] ? image_2445 : _GEN_24018; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24020 = 12'h98e == _T_221[11:0] ? image_2446 : _GEN_24019; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24021 = 12'h98f == _T_221[11:0] ? image_2447 : _GEN_24020; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24022 = 12'h990 == _T_221[11:0] ? image_2448 : _GEN_24021; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24023 = 12'h991 == _T_221[11:0] ? image_2449 : _GEN_24022; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24024 = 12'h992 == _T_221[11:0] ? image_2450 : _GEN_24023; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24025 = 12'h993 == _T_221[11:0] ? image_2451 : _GEN_24024; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24026 = 12'h994 == _T_221[11:0] ? image_2452 : _GEN_24025; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24027 = 12'h995 == _T_221[11:0] ? image_2453 : _GEN_24026; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24028 = 12'h996 == _T_221[11:0] ? image_2454 : _GEN_24027; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24029 = 12'h997 == _T_221[11:0] ? image_2455 : _GEN_24028; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24030 = 12'h998 == _T_221[11:0] ? image_2456 : _GEN_24029; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24031 = 12'h999 == _T_221[11:0] ? image_2457 : _GEN_24030; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24032 = 12'h99a == _T_221[11:0] ? image_2458 : _GEN_24031; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24033 = 12'h99b == _T_221[11:0] ? image_2459 : _GEN_24032; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24034 = 12'h99c == _T_221[11:0] ? image_2460 : _GEN_24033; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24035 = 12'h99d == _T_221[11:0] ? image_2461 : _GEN_24034; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24036 = 12'h99e == _T_221[11:0] ? image_2462 : _GEN_24035; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24037 = 12'h99f == _T_221[11:0] ? image_2463 : _GEN_24036; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24038 = 12'h9a0 == _T_221[11:0] ? image_2464 : _GEN_24037; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24039 = 12'h9a1 == _T_221[11:0] ? image_2465 : _GEN_24038; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24040 = 12'h9a2 == _T_221[11:0] ? image_2466 : _GEN_24039; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24041 = 12'h9a3 == _T_221[11:0] ? image_2467 : _GEN_24040; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24042 = 12'h9a4 == _T_221[11:0] ? image_2468 : _GEN_24041; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24043 = 12'h9a5 == _T_221[11:0] ? image_2469 : _GEN_24042; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24044 = 12'h9a6 == _T_221[11:0] ? image_2470 : _GEN_24043; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24045 = 12'h9a7 == _T_221[11:0] ? image_2471 : _GEN_24044; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24046 = 12'h9a8 == _T_221[11:0] ? image_2472 : _GEN_24045; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24047 = 12'h9a9 == _T_221[11:0] ? image_2473 : _GEN_24046; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24048 = 12'h9aa == _T_221[11:0] ? image_2474 : _GEN_24047; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24049 = 12'h9ab == _T_221[11:0] ? image_2475 : _GEN_24048; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24050 = 12'h9ac == _T_221[11:0] ? image_2476 : _GEN_24049; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24051 = 12'h9ad == _T_221[11:0] ? image_2477 : _GEN_24050; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24052 = 12'h9ae == _T_221[11:0] ? image_2478 : _GEN_24051; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24053 = 12'h9af == _T_221[11:0] ? image_2479 : _GEN_24052; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24054 = 12'h9b0 == _T_221[11:0] ? image_2480 : _GEN_24053; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24055 = 12'h9b1 == _T_221[11:0] ? image_2481 : _GEN_24054; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24056 = 12'h9b2 == _T_221[11:0] ? image_2482 : _GEN_24055; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24057 = 12'h9b3 == _T_221[11:0] ? image_2483 : _GEN_24056; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24058 = 12'h9b4 == _T_221[11:0] ? image_2484 : _GEN_24057; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24059 = 12'h9b5 == _T_221[11:0] ? image_2485 : _GEN_24058; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24060 = 12'h9b6 == _T_221[11:0] ? image_2486 : _GEN_24059; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24061 = 12'h9b7 == _T_221[11:0] ? image_2487 : _GEN_24060; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24062 = 12'h9b8 == _T_221[11:0] ? image_2488 : _GEN_24061; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24063 = 12'h9b9 == _T_221[11:0] ? image_2489 : _GEN_24062; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24064 = 12'h9ba == _T_221[11:0] ? image_2490 : _GEN_24063; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24065 = 12'h9bb == _T_221[11:0] ? 4'h0 : _GEN_24064; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24066 = 12'h9bc == _T_221[11:0] ? 4'h0 : _GEN_24065; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24067 = 12'h9bd == _T_221[11:0] ? 4'h0 : _GEN_24066; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24068 = 12'h9be == _T_221[11:0] ? 4'h0 : _GEN_24067; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24069 = 12'h9bf == _T_221[11:0] ? 4'h0 : _GEN_24068; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24070 = 12'h9c0 == _T_221[11:0] ? 4'h0 : _GEN_24069; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24071 = 12'h9c1 == _T_221[11:0] ? 4'h0 : _GEN_24070; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24072 = 12'h9c2 == _T_221[11:0] ? 4'h0 : _GEN_24071; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24073 = 12'h9c3 == _T_221[11:0] ? 4'h0 : _GEN_24072; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24074 = 12'h9c4 == _T_221[11:0] ? 4'h0 : _GEN_24073; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24075 = 12'h9c5 == _T_221[11:0] ? 4'h0 : _GEN_24074; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24076 = 12'h9c6 == _T_221[11:0] ? image_2502 : _GEN_24075; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24077 = 12'h9c7 == _T_221[11:0] ? image_2503 : _GEN_24076; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24078 = 12'h9c8 == _T_221[11:0] ? image_2504 : _GEN_24077; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24079 = 12'h9c9 == _T_221[11:0] ? image_2505 : _GEN_24078; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24080 = 12'h9ca == _T_221[11:0] ? image_2506 : _GEN_24079; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24081 = 12'h9cb == _T_221[11:0] ? image_2507 : _GEN_24080; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24082 = 12'h9cc == _T_221[11:0] ? image_2508 : _GEN_24081; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24083 = 12'h9cd == _T_221[11:0] ? image_2509 : _GEN_24082; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24084 = 12'h9ce == _T_221[11:0] ? image_2510 : _GEN_24083; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24085 = 12'h9cf == _T_221[11:0] ? image_2511 : _GEN_24084; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24086 = 12'h9d0 == _T_221[11:0] ? image_2512 : _GEN_24085; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24087 = 12'h9d1 == _T_221[11:0] ? image_2513 : _GEN_24086; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24088 = 12'h9d2 == _T_221[11:0] ? image_2514 : _GEN_24087; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24089 = 12'h9d3 == _T_221[11:0] ? image_2515 : _GEN_24088; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24090 = 12'h9d4 == _T_221[11:0] ? image_2516 : _GEN_24089; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24091 = 12'h9d5 == _T_221[11:0] ? image_2517 : _GEN_24090; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24092 = 12'h9d6 == _T_221[11:0] ? image_2518 : _GEN_24091; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24093 = 12'h9d7 == _T_221[11:0] ? image_2519 : _GEN_24092; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24094 = 12'h9d8 == _T_221[11:0] ? image_2520 : _GEN_24093; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24095 = 12'h9d9 == _T_221[11:0] ? image_2521 : _GEN_24094; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24096 = 12'h9da == _T_221[11:0] ? image_2522 : _GEN_24095; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24097 = 12'h9db == _T_221[11:0] ? image_2523 : _GEN_24096; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24098 = 12'h9dc == _T_221[11:0] ? image_2524 : _GEN_24097; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24099 = 12'h9dd == _T_221[11:0] ? image_2525 : _GEN_24098; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24100 = 12'h9de == _T_221[11:0] ? image_2526 : _GEN_24099; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24101 = 12'h9df == _T_221[11:0] ? image_2527 : _GEN_24100; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24102 = 12'h9e0 == _T_221[11:0] ? image_2528 : _GEN_24101; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24103 = 12'h9e1 == _T_221[11:0] ? image_2529 : _GEN_24102; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24104 = 12'h9e2 == _T_221[11:0] ? image_2530 : _GEN_24103; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24105 = 12'h9e3 == _T_221[11:0] ? image_2531 : _GEN_24104; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24106 = 12'h9e4 == _T_221[11:0] ? image_2532 : _GEN_24105; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24107 = 12'h9e5 == _T_221[11:0] ? image_2533 : _GEN_24106; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24108 = 12'h9e6 == _T_221[11:0] ? image_2534 : _GEN_24107; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24109 = 12'h9e7 == _T_221[11:0] ? image_2535 : _GEN_24108; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24110 = 12'h9e8 == _T_221[11:0] ? image_2536 : _GEN_24109; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24111 = 12'h9e9 == _T_221[11:0] ? image_2537 : _GEN_24110; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24112 = 12'h9ea == _T_221[11:0] ? image_2538 : _GEN_24111; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24113 = 12'h9eb == _T_221[11:0] ? image_2539 : _GEN_24112; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24114 = 12'h9ec == _T_221[11:0] ? image_2540 : _GEN_24113; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24115 = 12'h9ed == _T_221[11:0] ? image_2541 : _GEN_24114; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24116 = 12'h9ee == _T_221[11:0] ? image_2542 : _GEN_24115; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24117 = 12'h9ef == _T_221[11:0] ? image_2543 : _GEN_24116; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24118 = 12'h9f0 == _T_221[11:0] ? image_2544 : _GEN_24117; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24119 = 12'h9f1 == _T_221[11:0] ? image_2545 : _GEN_24118; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24120 = 12'h9f2 == _T_221[11:0] ? image_2546 : _GEN_24119; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24121 = 12'h9f3 == _T_221[11:0] ? image_2547 : _GEN_24120; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24122 = 12'h9f4 == _T_221[11:0] ? image_2548 : _GEN_24121; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24123 = 12'h9f5 == _T_221[11:0] ? image_2549 : _GEN_24122; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24124 = 12'h9f6 == _T_221[11:0] ? image_2550 : _GEN_24123; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24125 = 12'h9f7 == _T_221[11:0] ? image_2551 : _GEN_24124; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24126 = 12'h9f8 == _T_221[11:0] ? image_2552 : _GEN_24125; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24127 = 12'h9f9 == _T_221[11:0] ? image_2553 : _GEN_24126; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24128 = 12'h9fa == _T_221[11:0] ? image_2554 : _GEN_24127; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24129 = 12'h9fb == _T_221[11:0] ? 4'h0 : _GEN_24128; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24130 = 12'h9fc == _T_221[11:0] ? 4'h0 : _GEN_24129; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24131 = 12'h9fd == _T_221[11:0] ? 4'h0 : _GEN_24130; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24132 = 12'h9fe == _T_221[11:0] ? 4'h0 : _GEN_24131; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24133 = 12'h9ff == _T_221[11:0] ? 4'h0 : _GEN_24132; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24134 = 12'ha00 == _T_221[11:0] ? 4'h0 : _GEN_24133; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24135 = 12'ha01 == _T_221[11:0] ? 4'h0 : _GEN_24134; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24136 = 12'ha02 == _T_221[11:0] ? 4'h0 : _GEN_24135; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24137 = 12'ha03 == _T_221[11:0] ? 4'h0 : _GEN_24136; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24138 = 12'ha04 == _T_221[11:0] ? 4'h0 : _GEN_24137; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24139 = 12'ha05 == _T_221[11:0] ? 4'h0 : _GEN_24138; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24140 = 12'ha06 == _T_221[11:0] ? 4'h0 : _GEN_24139; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24141 = 12'ha07 == _T_221[11:0] ? image_2567 : _GEN_24140; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24142 = 12'ha08 == _T_221[11:0] ? image_2568 : _GEN_24141; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24143 = 12'ha09 == _T_221[11:0] ? image_2569 : _GEN_24142; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24144 = 12'ha0a == _T_221[11:0] ? image_2570 : _GEN_24143; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24145 = 12'ha0b == _T_221[11:0] ? image_2571 : _GEN_24144; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24146 = 12'ha0c == _T_221[11:0] ? image_2572 : _GEN_24145; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24147 = 12'ha0d == _T_221[11:0] ? image_2573 : _GEN_24146; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24148 = 12'ha0e == _T_221[11:0] ? image_2574 : _GEN_24147; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24149 = 12'ha0f == _T_221[11:0] ? image_2575 : _GEN_24148; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24150 = 12'ha10 == _T_221[11:0] ? image_2576 : _GEN_24149; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24151 = 12'ha11 == _T_221[11:0] ? image_2577 : _GEN_24150; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24152 = 12'ha12 == _T_221[11:0] ? image_2578 : _GEN_24151; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24153 = 12'ha13 == _T_221[11:0] ? image_2579 : _GEN_24152; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24154 = 12'ha14 == _T_221[11:0] ? image_2580 : _GEN_24153; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24155 = 12'ha15 == _T_221[11:0] ? image_2581 : _GEN_24154; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24156 = 12'ha16 == _T_221[11:0] ? image_2582 : _GEN_24155; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24157 = 12'ha17 == _T_221[11:0] ? image_2583 : _GEN_24156; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24158 = 12'ha18 == _T_221[11:0] ? image_2584 : _GEN_24157; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24159 = 12'ha19 == _T_221[11:0] ? image_2585 : _GEN_24158; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24160 = 12'ha1a == _T_221[11:0] ? image_2586 : _GEN_24159; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24161 = 12'ha1b == _T_221[11:0] ? image_2587 : _GEN_24160; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24162 = 12'ha1c == _T_221[11:0] ? image_2588 : _GEN_24161; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24163 = 12'ha1d == _T_221[11:0] ? image_2589 : _GEN_24162; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24164 = 12'ha1e == _T_221[11:0] ? image_2590 : _GEN_24163; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24165 = 12'ha1f == _T_221[11:0] ? image_2591 : _GEN_24164; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24166 = 12'ha20 == _T_221[11:0] ? image_2592 : _GEN_24165; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24167 = 12'ha21 == _T_221[11:0] ? image_2593 : _GEN_24166; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24168 = 12'ha22 == _T_221[11:0] ? image_2594 : _GEN_24167; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24169 = 12'ha23 == _T_221[11:0] ? image_2595 : _GEN_24168; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24170 = 12'ha24 == _T_221[11:0] ? image_2596 : _GEN_24169; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24171 = 12'ha25 == _T_221[11:0] ? image_2597 : _GEN_24170; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24172 = 12'ha26 == _T_221[11:0] ? image_2598 : _GEN_24171; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24173 = 12'ha27 == _T_221[11:0] ? image_2599 : _GEN_24172; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24174 = 12'ha28 == _T_221[11:0] ? image_2600 : _GEN_24173; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24175 = 12'ha29 == _T_221[11:0] ? image_2601 : _GEN_24174; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24176 = 12'ha2a == _T_221[11:0] ? image_2602 : _GEN_24175; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24177 = 12'ha2b == _T_221[11:0] ? image_2603 : _GEN_24176; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24178 = 12'ha2c == _T_221[11:0] ? image_2604 : _GEN_24177; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24179 = 12'ha2d == _T_221[11:0] ? image_2605 : _GEN_24178; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24180 = 12'ha2e == _T_221[11:0] ? image_2606 : _GEN_24179; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24181 = 12'ha2f == _T_221[11:0] ? image_2607 : _GEN_24180; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24182 = 12'ha30 == _T_221[11:0] ? image_2608 : _GEN_24181; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24183 = 12'ha31 == _T_221[11:0] ? image_2609 : _GEN_24182; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24184 = 12'ha32 == _T_221[11:0] ? image_2610 : _GEN_24183; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24185 = 12'ha33 == _T_221[11:0] ? image_2611 : _GEN_24184; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24186 = 12'ha34 == _T_221[11:0] ? image_2612 : _GEN_24185; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24187 = 12'ha35 == _T_221[11:0] ? image_2613 : _GEN_24186; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24188 = 12'ha36 == _T_221[11:0] ? image_2614 : _GEN_24187; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24189 = 12'ha37 == _T_221[11:0] ? image_2615 : _GEN_24188; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24190 = 12'ha38 == _T_221[11:0] ? image_2616 : _GEN_24189; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24191 = 12'ha39 == _T_221[11:0] ? image_2617 : _GEN_24190; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24192 = 12'ha3a == _T_221[11:0] ? image_2618 : _GEN_24191; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24193 = 12'ha3b == _T_221[11:0] ? 4'h0 : _GEN_24192; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24194 = 12'ha3c == _T_221[11:0] ? 4'h0 : _GEN_24193; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24195 = 12'ha3d == _T_221[11:0] ? 4'h0 : _GEN_24194; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24196 = 12'ha3e == _T_221[11:0] ? 4'h0 : _GEN_24195; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24197 = 12'ha3f == _T_221[11:0] ? 4'h0 : _GEN_24196; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24198 = 12'ha40 == _T_221[11:0] ? 4'h0 : _GEN_24197; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24199 = 12'ha41 == _T_221[11:0] ? 4'h0 : _GEN_24198; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24200 = 12'ha42 == _T_221[11:0] ? 4'h0 : _GEN_24199; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24201 = 12'ha43 == _T_221[11:0] ? 4'h0 : _GEN_24200; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24202 = 12'ha44 == _T_221[11:0] ? 4'h0 : _GEN_24201; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24203 = 12'ha45 == _T_221[11:0] ? 4'h0 : _GEN_24202; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24204 = 12'ha46 == _T_221[11:0] ? 4'h0 : _GEN_24203; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24205 = 12'ha47 == _T_221[11:0] ? 4'h0 : _GEN_24204; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24206 = 12'ha48 == _T_221[11:0] ? image_2632 : _GEN_24205; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24207 = 12'ha49 == _T_221[11:0] ? image_2633 : _GEN_24206; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24208 = 12'ha4a == _T_221[11:0] ? image_2634 : _GEN_24207; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24209 = 12'ha4b == _T_221[11:0] ? image_2635 : _GEN_24208; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24210 = 12'ha4c == _T_221[11:0] ? image_2636 : _GEN_24209; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24211 = 12'ha4d == _T_221[11:0] ? image_2637 : _GEN_24210; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24212 = 12'ha4e == _T_221[11:0] ? image_2638 : _GEN_24211; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24213 = 12'ha4f == _T_221[11:0] ? image_2639 : _GEN_24212; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24214 = 12'ha50 == _T_221[11:0] ? image_2640 : _GEN_24213; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24215 = 12'ha51 == _T_221[11:0] ? image_2641 : _GEN_24214; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24216 = 12'ha52 == _T_221[11:0] ? image_2642 : _GEN_24215; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24217 = 12'ha53 == _T_221[11:0] ? image_2643 : _GEN_24216; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24218 = 12'ha54 == _T_221[11:0] ? image_2644 : _GEN_24217; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24219 = 12'ha55 == _T_221[11:0] ? image_2645 : _GEN_24218; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24220 = 12'ha56 == _T_221[11:0] ? image_2646 : _GEN_24219; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24221 = 12'ha57 == _T_221[11:0] ? image_2647 : _GEN_24220; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24222 = 12'ha58 == _T_221[11:0] ? image_2648 : _GEN_24221; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24223 = 12'ha59 == _T_221[11:0] ? image_2649 : _GEN_24222; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24224 = 12'ha5a == _T_221[11:0] ? image_2650 : _GEN_24223; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24225 = 12'ha5b == _T_221[11:0] ? image_2651 : _GEN_24224; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24226 = 12'ha5c == _T_221[11:0] ? image_2652 : _GEN_24225; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24227 = 12'ha5d == _T_221[11:0] ? image_2653 : _GEN_24226; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24228 = 12'ha5e == _T_221[11:0] ? image_2654 : _GEN_24227; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24229 = 12'ha5f == _T_221[11:0] ? image_2655 : _GEN_24228; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24230 = 12'ha60 == _T_221[11:0] ? image_2656 : _GEN_24229; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24231 = 12'ha61 == _T_221[11:0] ? image_2657 : _GEN_24230; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24232 = 12'ha62 == _T_221[11:0] ? image_2658 : _GEN_24231; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24233 = 12'ha63 == _T_221[11:0] ? image_2659 : _GEN_24232; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24234 = 12'ha64 == _T_221[11:0] ? image_2660 : _GEN_24233; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24235 = 12'ha65 == _T_221[11:0] ? image_2661 : _GEN_24234; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24236 = 12'ha66 == _T_221[11:0] ? image_2662 : _GEN_24235; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24237 = 12'ha67 == _T_221[11:0] ? image_2663 : _GEN_24236; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24238 = 12'ha68 == _T_221[11:0] ? image_2664 : _GEN_24237; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24239 = 12'ha69 == _T_221[11:0] ? image_2665 : _GEN_24238; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24240 = 12'ha6a == _T_221[11:0] ? image_2666 : _GEN_24239; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24241 = 12'ha6b == _T_221[11:0] ? image_2667 : _GEN_24240; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24242 = 12'ha6c == _T_221[11:0] ? image_2668 : _GEN_24241; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24243 = 12'ha6d == _T_221[11:0] ? image_2669 : _GEN_24242; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24244 = 12'ha6e == _T_221[11:0] ? image_2670 : _GEN_24243; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24245 = 12'ha6f == _T_221[11:0] ? image_2671 : _GEN_24244; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24246 = 12'ha70 == _T_221[11:0] ? image_2672 : _GEN_24245; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24247 = 12'ha71 == _T_221[11:0] ? image_2673 : _GEN_24246; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24248 = 12'ha72 == _T_221[11:0] ? image_2674 : _GEN_24247; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24249 = 12'ha73 == _T_221[11:0] ? image_2675 : _GEN_24248; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24250 = 12'ha74 == _T_221[11:0] ? image_2676 : _GEN_24249; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24251 = 12'ha75 == _T_221[11:0] ? image_2677 : _GEN_24250; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24252 = 12'ha76 == _T_221[11:0] ? image_2678 : _GEN_24251; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24253 = 12'ha77 == _T_221[11:0] ? image_2679 : _GEN_24252; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24254 = 12'ha78 == _T_221[11:0] ? image_2680 : _GEN_24253; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24255 = 12'ha79 == _T_221[11:0] ? image_2681 : _GEN_24254; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24256 = 12'ha7a == _T_221[11:0] ? image_2682 : _GEN_24255; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24257 = 12'ha7b == _T_221[11:0] ? 4'h0 : _GEN_24256; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24258 = 12'ha7c == _T_221[11:0] ? 4'h0 : _GEN_24257; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24259 = 12'ha7d == _T_221[11:0] ? 4'h0 : _GEN_24258; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24260 = 12'ha7e == _T_221[11:0] ? 4'h0 : _GEN_24259; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24261 = 12'ha7f == _T_221[11:0] ? 4'h0 : _GEN_24260; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24262 = 12'ha80 == _T_221[11:0] ? 4'h0 : _GEN_24261; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24263 = 12'ha81 == _T_221[11:0] ? 4'h0 : _GEN_24262; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24264 = 12'ha82 == _T_221[11:0] ? 4'h0 : _GEN_24263; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24265 = 12'ha83 == _T_221[11:0] ? 4'h0 : _GEN_24264; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24266 = 12'ha84 == _T_221[11:0] ? 4'h0 : _GEN_24265; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24267 = 12'ha85 == _T_221[11:0] ? 4'h0 : _GEN_24266; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24268 = 12'ha86 == _T_221[11:0] ? 4'h0 : _GEN_24267; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24269 = 12'ha87 == _T_221[11:0] ? 4'h0 : _GEN_24268; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24270 = 12'ha88 == _T_221[11:0] ? 4'h0 : _GEN_24269; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24271 = 12'ha89 == _T_221[11:0] ? image_2697 : _GEN_24270; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24272 = 12'ha8a == _T_221[11:0] ? image_2698 : _GEN_24271; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24273 = 12'ha8b == _T_221[11:0] ? image_2699 : _GEN_24272; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24274 = 12'ha8c == _T_221[11:0] ? image_2700 : _GEN_24273; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24275 = 12'ha8d == _T_221[11:0] ? image_2701 : _GEN_24274; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24276 = 12'ha8e == _T_221[11:0] ? image_2702 : _GEN_24275; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24277 = 12'ha8f == _T_221[11:0] ? image_2703 : _GEN_24276; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24278 = 12'ha90 == _T_221[11:0] ? image_2704 : _GEN_24277; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24279 = 12'ha91 == _T_221[11:0] ? image_2705 : _GEN_24278; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24280 = 12'ha92 == _T_221[11:0] ? image_2706 : _GEN_24279; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24281 = 12'ha93 == _T_221[11:0] ? image_2707 : _GEN_24280; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24282 = 12'ha94 == _T_221[11:0] ? image_2708 : _GEN_24281; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24283 = 12'ha95 == _T_221[11:0] ? image_2709 : _GEN_24282; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24284 = 12'ha96 == _T_221[11:0] ? image_2710 : _GEN_24283; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24285 = 12'ha97 == _T_221[11:0] ? image_2711 : _GEN_24284; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24286 = 12'ha98 == _T_221[11:0] ? image_2712 : _GEN_24285; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24287 = 12'ha99 == _T_221[11:0] ? image_2713 : _GEN_24286; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24288 = 12'ha9a == _T_221[11:0] ? image_2714 : _GEN_24287; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24289 = 12'ha9b == _T_221[11:0] ? image_2715 : _GEN_24288; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24290 = 12'ha9c == _T_221[11:0] ? image_2716 : _GEN_24289; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24291 = 12'ha9d == _T_221[11:0] ? image_2717 : _GEN_24290; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24292 = 12'ha9e == _T_221[11:0] ? image_2718 : _GEN_24291; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24293 = 12'ha9f == _T_221[11:0] ? image_2719 : _GEN_24292; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24294 = 12'haa0 == _T_221[11:0] ? image_2720 : _GEN_24293; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24295 = 12'haa1 == _T_221[11:0] ? image_2721 : _GEN_24294; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24296 = 12'haa2 == _T_221[11:0] ? image_2722 : _GEN_24295; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24297 = 12'haa3 == _T_221[11:0] ? image_2723 : _GEN_24296; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24298 = 12'haa4 == _T_221[11:0] ? image_2724 : _GEN_24297; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24299 = 12'haa5 == _T_221[11:0] ? image_2725 : _GEN_24298; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24300 = 12'haa6 == _T_221[11:0] ? image_2726 : _GEN_24299; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24301 = 12'haa7 == _T_221[11:0] ? image_2727 : _GEN_24300; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24302 = 12'haa8 == _T_221[11:0] ? image_2728 : _GEN_24301; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24303 = 12'haa9 == _T_221[11:0] ? image_2729 : _GEN_24302; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24304 = 12'haaa == _T_221[11:0] ? image_2730 : _GEN_24303; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24305 = 12'haab == _T_221[11:0] ? image_2731 : _GEN_24304; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24306 = 12'haac == _T_221[11:0] ? image_2732 : _GEN_24305; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24307 = 12'haad == _T_221[11:0] ? image_2733 : _GEN_24306; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24308 = 12'haae == _T_221[11:0] ? image_2734 : _GEN_24307; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24309 = 12'haaf == _T_221[11:0] ? image_2735 : _GEN_24308; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24310 = 12'hab0 == _T_221[11:0] ? image_2736 : _GEN_24309; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24311 = 12'hab1 == _T_221[11:0] ? image_2737 : _GEN_24310; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24312 = 12'hab2 == _T_221[11:0] ? image_2738 : _GEN_24311; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24313 = 12'hab3 == _T_221[11:0] ? image_2739 : _GEN_24312; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24314 = 12'hab4 == _T_221[11:0] ? image_2740 : _GEN_24313; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24315 = 12'hab5 == _T_221[11:0] ? image_2741 : _GEN_24314; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24316 = 12'hab6 == _T_221[11:0] ? image_2742 : _GEN_24315; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24317 = 12'hab7 == _T_221[11:0] ? image_2743 : _GEN_24316; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24318 = 12'hab8 == _T_221[11:0] ? image_2744 : _GEN_24317; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24319 = 12'hab9 == _T_221[11:0] ? image_2745 : _GEN_24318; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24320 = 12'haba == _T_221[11:0] ? 4'h0 : _GEN_24319; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24321 = 12'habb == _T_221[11:0] ? 4'h0 : _GEN_24320; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24322 = 12'habc == _T_221[11:0] ? 4'h0 : _GEN_24321; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24323 = 12'habd == _T_221[11:0] ? 4'h0 : _GEN_24322; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24324 = 12'habe == _T_221[11:0] ? 4'h0 : _GEN_24323; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24325 = 12'habf == _T_221[11:0] ? 4'h0 : _GEN_24324; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24326 = 12'hac0 == _T_221[11:0] ? 4'h0 : _GEN_24325; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24327 = 12'hac1 == _T_221[11:0] ? 4'h0 : _GEN_24326; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24328 = 12'hac2 == _T_221[11:0] ? 4'h0 : _GEN_24327; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24329 = 12'hac3 == _T_221[11:0] ? 4'h0 : _GEN_24328; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24330 = 12'hac4 == _T_221[11:0] ? 4'h0 : _GEN_24329; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24331 = 12'hac5 == _T_221[11:0] ? 4'h0 : _GEN_24330; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24332 = 12'hac6 == _T_221[11:0] ? 4'h0 : _GEN_24331; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24333 = 12'hac7 == _T_221[11:0] ? 4'h0 : _GEN_24332; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24334 = 12'hac8 == _T_221[11:0] ? 4'h0 : _GEN_24333; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24335 = 12'hac9 == _T_221[11:0] ? 4'h0 : _GEN_24334; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24336 = 12'haca == _T_221[11:0] ? 4'h0 : _GEN_24335; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24337 = 12'hacb == _T_221[11:0] ? image_2763 : _GEN_24336; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24338 = 12'hacc == _T_221[11:0] ? image_2764 : _GEN_24337; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24339 = 12'hacd == _T_221[11:0] ? image_2765 : _GEN_24338; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24340 = 12'hace == _T_221[11:0] ? image_2766 : _GEN_24339; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24341 = 12'hacf == _T_221[11:0] ? image_2767 : _GEN_24340; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24342 = 12'had0 == _T_221[11:0] ? image_2768 : _GEN_24341; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24343 = 12'had1 == _T_221[11:0] ? image_2769 : _GEN_24342; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24344 = 12'had2 == _T_221[11:0] ? image_2770 : _GEN_24343; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24345 = 12'had3 == _T_221[11:0] ? image_2771 : _GEN_24344; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24346 = 12'had4 == _T_221[11:0] ? image_2772 : _GEN_24345; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24347 = 12'had5 == _T_221[11:0] ? image_2773 : _GEN_24346; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24348 = 12'had6 == _T_221[11:0] ? image_2774 : _GEN_24347; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24349 = 12'had7 == _T_221[11:0] ? image_2775 : _GEN_24348; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24350 = 12'had8 == _T_221[11:0] ? image_2776 : _GEN_24349; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24351 = 12'had9 == _T_221[11:0] ? image_2777 : _GEN_24350; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24352 = 12'hada == _T_221[11:0] ? image_2778 : _GEN_24351; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24353 = 12'hadb == _T_221[11:0] ? image_2779 : _GEN_24352; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24354 = 12'hadc == _T_221[11:0] ? image_2780 : _GEN_24353; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24355 = 12'hadd == _T_221[11:0] ? image_2781 : _GEN_24354; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24356 = 12'hade == _T_221[11:0] ? image_2782 : _GEN_24355; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24357 = 12'hadf == _T_221[11:0] ? image_2783 : _GEN_24356; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24358 = 12'hae0 == _T_221[11:0] ? image_2784 : _GEN_24357; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24359 = 12'hae1 == _T_221[11:0] ? image_2785 : _GEN_24358; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24360 = 12'hae2 == _T_221[11:0] ? image_2786 : _GEN_24359; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24361 = 12'hae3 == _T_221[11:0] ? image_2787 : _GEN_24360; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24362 = 12'hae4 == _T_221[11:0] ? image_2788 : _GEN_24361; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24363 = 12'hae5 == _T_221[11:0] ? image_2789 : _GEN_24362; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24364 = 12'hae6 == _T_221[11:0] ? image_2790 : _GEN_24363; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24365 = 12'hae7 == _T_221[11:0] ? image_2791 : _GEN_24364; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24366 = 12'hae8 == _T_221[11:0] ? image_2792 : _GEN_24365; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24367 = 12'hae9 == _T_221[11:0] ? image_2793 : _GEN_24366; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24368 = 12'haea == _T_221[11:0] ? image_2794 : _GEN_24367; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24369 = 12'haeb == _T_221[11:0] ? image_2795 : _GEN_24368; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24370 = 12'haec == _T_221[11:0] ? image_2796 : _GEN_24369; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24371 = 12'haed == _T_221[11:0] ? image_2797 : _GEN_24370; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24372 = 12'haee == _T_221[11:0] ? image_2798 : _GEN_24371; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24373 = 12'haef == _T_221[11:0] ? image_2799 : _GEN_24372; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24374 = 12'haf0 == _T_221[11:0] ? image_2800 : _GEN_24373; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24375 = 12'haf1 == _T_221[11:0] ? image_2801 : _GEN_24374; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24376 = 12'haf2 == _T_221[11:0] ? image_2802 : _GEN_24375; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24377 = 12'haf3 == _T_221[11:0] ? image_2803 : _GEN_24376; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24378 = 12'haf4 == _T_221[11:0] ? image_2804 : _GEN_24377; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24379 = 12'haf5 == _T_221[11:0] ? image_2805 : _GEN_24378; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24380 = 12'haf6 == _T_221[11:0] ? image_2806 : _GEN_24379; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24381 = 12'haf7 == _T_221[11:0] ? image_2807 : _GEN_24380; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24382 = 12'haf8 == _T_221[11:0] ? image_2808 : _GEN_24381; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24383 = 12'haf9 == _T_221[11:0] ? 4'h0 : _GEN_24382; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24384 = 12'hafa == _T_221[11:0] ? 4'h0 : _GEN_24383; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24385 = 12'hafb == _T_221[11:0] ? 4'h0 : _GEN_24384; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24386 = 12'hafc == _T_221[11:0] ? 4'h0 : _GEN_24385; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24387 = 12'hafd == _T_221[11:0] ? 4'h0 : _GEN_24386; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24388 = 12'hafe == _T_221[11:0] ? 4'h0 : _GEN_24387; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24389 = 12'haff == _T_221[11:0] ? 4'h0 : _GEN_24388; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24390 = 12'hb00 == _T_221[11:0] ? 4'h0 : _GEN_24389; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24391 = 12'hb01 == _T_221[11:0] ? 4'h0 : _GEN_24390; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24392 = 12'hb02 == _T_221[11:0] ? 4'h0 : _GEN_24391; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24393 = 12'hb03 == _T_221[11:0] ? 4'h0 : _GEN_24392; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24394 = 12'hb04 == _T_221[11:0] ? 4'h0 : _GEN_24393; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24395 = 12'hb05 == _T_221[11:0] ? 4'h0 : _GEN_24394; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24396 = 12'hb06 == _T_221[11:0] ? 4'h0 : _GEN_24395; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24397 = 12'hb07 == _T_221[11:0] ? 4'h0 : _GEN_24396; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24398 = 12'hb08 == _T_221[11:0] ? 4'h0 : _GEN_24397; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24399 = 12'hb09 == _T_221[11:0] ? 4'h0 : _GEN_24398; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24400 = 12'hb0a == _T_221[11:0] ? 4'h0 : _GEN_24399; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24401 = 12'hb0b == _T_221[11:0] ? 4'h0 : _GEN_24400; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24402 = 12'hb0c == _T_221[11:0] ? image_2828 : _GEN_24401; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24403 = 12'hb0d == _T_221[11:0] ? image_2829 : _GEN_24402; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24404 = 12'hb0e == _T_221[11:0] ? image_2830 : _GEN_24403; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24405 = 12'hb0f == _T_221[11:0] ? image_2831 : _GEN_24404; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24406 = 12'hb10 == _T_221[11:0] ? image_2832 : _GEN_24405; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24407 = 12'hb11 == _T_221[11:0] ? image_2833 : _GEN_24406; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24408 = 12'hb12 == _T_221[11:0] ? image_2834 : _GEN_24407; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24409 = 12'hb13 == _T_221[11:0] ? image_2835 : _GEN_24408; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24410 = 12'hb14 == _T_221[11:0] ? image_2836 : _GEN_24409; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24411 = 12'hb15 == _T_221[11:0] ? image_2837 : _GEN_24410; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24412 = 12'hb16 == _T_221[11:0] ? image_2838 : _GEN_24411; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24413 = 12'hb17 == _T_221[11:0] ? image_2839 : _GEN_24412; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24414 = 12'hb18 == _T_221[11:0] ? image_2840 : _GEN_24413; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24415 = 12'hb19 == _T_221[11:0] ? image_2841 : _GEN_24414; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24416 = 12'hb1a == _T_221[11:0] ? image_2842 : _GEN_24415; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24417 = 12'hb1b == _T_221[11:0] ? image_2843 : _GEN_24416; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24418 = 12'hb1c == _T_221[11:0] ? image_2844 : _GEN_24417; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24419 = 12'hb1d == _T_221[11:0] ? image_2845 : _GEN_24418; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24420 = 12'hb1e == _T_221[11:0] ? image_2846 : _GEN_24419; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24421 = 12'hb1f == _T_221[11:0] ? image_2847 : _GEN_24420; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24422 = 12'hb20 == _T_221[11:0] ? image_2848 : _GEN_24421; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24423 = 12'hb21 == _T_221[11:0] ? image_2849 : _GEN_24422; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24424 = 12'hb22 == _T_221[11:0] ? image_2850 : _GEN_24423; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24425 = 12'hb23 == _T_221[11:0] ? image_2851 : _GEN_24424; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24426 = 12'hb24 == _T_221[11:0] ? image_2852 : _GEN_24425; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24427 = 12'hb25 == _T_221[11:0] ? image_2853 : _GEN_24426; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24428 = 12'hb26 == _T_221[11:0] ? image_2854 : _GEN_24427; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24429 = 12'hb27 == _T_221[11:0] ? image_2855 : _GEN_24428; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24430 = 12'hb28 == _T_221[11:0] ? image_2856 : _GEN_24429; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24431 = 12'hb29 == _T_221[11:0] ? image_2857 : _GEN_24430; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24432 = 12'hb2a == _T_221[11:0] ? image_2858 : _GEN_24431; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24433 = 12'hb2b == _T_221[11:0] ? image_2859 : _GEN_24432; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24434 = 12'hb2c == _T_221[11:0] ? image_2860 : _GEN_24433; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24435 = 12'hb2d == _T_221[11:0] ? image_2861 : _GEN_24434; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24436 = 12'hb2e == _T_221[11:0] ? image_2862 : _GEN_24435; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24437 = 12'hb2f == _T_221[11:0] ? image_2863 : _GEN_24436; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24438 = 12'hb30 == _T_221[11:0] ? image_2864 : _GEN_24437; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24439 = 12'hb31 == _T_221[11:0] ? image_2865 : _GEN_24438; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24440 = 12'hb32 == _T_221[11:0] ? image_2866 : _GEN_24439; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24441 = 12'hb33 == _T_221[11:0] ? image_2867 : _GEN_24440; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24442 = 12'hb34 == _T_221[11:0] ? image_2868 : _GEN_24441; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24443 = 12'hb35 == _T_221[11:0] ? image_2869 : _GEN_24442; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24444 = 12'hb36 == _T_221[11:0] ? image_2870 : _GEN_24443; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24445 = 12'hb37 == _T_221[11:0] ? image_2871 : _GEN_24444; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24446 = 12'hb38 == _T_221[11:0] ? 4'h0 : _GEN_24445; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24447 = 12'hb39 == _T_221[11:0] ? 4'h0 : _GEN_24446; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24448 = 12'hb3a == _T_221[11:0] ? 4'h0 : _GEN_24447; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24449 = 12'hb3b == _T_221[11:0] ? 4'h0 : _GEN_24448; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24450 = 12'hb3c == _T_221[11:0] ? 4'h0 : _GEN_24449; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24451 = 12'hb3d == _T_221[11:0] ? 4'h0 : _GEN_24450; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24452 = 12'hb3e == _T_221[11:0] ? 4'h0 : _GEN_24451; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24453 = 12'hb3f == _T_221[11:0] ? 4'h0 : _GEN_24452; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24454 = 12'hb40 == _T_221[11:0] ? 4'h0 : _GEN_24453; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24455 = 12'hb41 == _T_221[11:0] ? 4'h0 : _GEN_24454; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24456 = 12'hb42 == _T_221[11:0] ? 4'h0 : _GEN_24455; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24457 = 12'hb43 == _T_221[11:0] ? 4'h0 : _GEN_24456; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24458 = 12'hb44 == _T_221[11:0] ? 4'h0 : _GEN_24457; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24459 = 12'hb45 == _T_221[11:0] ? 4'h0 : _GEN_24458; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24460 = 12'hb46 == _T_221[11:0] ? 4'h0 : _GEN_24459; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24461 = 12'hb47 == _T_221[11:0] ? 4'h0 : _GEN_24460; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24462 = 12'hb48 == _T_221[11:0] ? 4'h0 : _GEN_24461; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24463 = 12'hb49 == _T_221[11:0] ? 4'h0 : _GEN_24462; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24464 = 12'hb4a == _T_221[11:0] ? 4'h0 : _GEN_24463; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24465 = 12'hb4b == _T_221[11:0] ? 4'h0 : _GEN_24464; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24466 = 12'hb4c == _T_221[11:0] ? 4'h0 : _GEN_24465; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24467 = 12'hb4d == _T_221[11:0] ? 4'h0 : _GEN_24466; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24468 = 12'hb4e == _T_221[11:0] ? 4'h0 : _GEN_24467; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24469 = 12'hb4f == _T_221[11:0] ? image_2895 : _GEN_24468; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24470 = 12'hb50 == _T_221[11:0] ? image_2896 : _GEN_24469; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24471 = 12'hb51 == _T_221[11:0] ? image_2897 : _GEN_24470; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24472 = 12'hb52 == _T_221[11:0] ? image_2898 : _GEN_24471; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24473 = 12'hb53 == _T_221[11:0] ? image_2899 : _GEN_24472; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24474 = 12'hb54 == _T_221[11:0] ? image_2900 : _GEN_24473; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24475 = 12'hb55 == _T_221[11:0] ? image_2901 : _GEN_24474; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24476 = 12'hb56 == _T_221[11:0] ? image_2902 : _GEN_24475; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24477 = 12'hb57 == _T_221[11:0] ? image_2903 : _GEN_24476; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24478 = 12'hb58 == _T_221[11:0] ? image_2904 : _GEN_24477; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24479 = 12'hb59 == _T_221[11:0] ? image_2905 : _GEN_24478; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24480 = 12'hb5a == _T_221[11:0] ? image_2906 : _GEN_24479; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24481 = 12'hb5b == _T_221[11:0] ? image_2907 : _GEN_24480; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24482 = 12'hb5c == _T_221[11:0] ? image_2908 : _GEN_24481; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24483 = 12'hb5d == _T_221[11:0] ? image_2909 : _GEN_24482; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24484 = 12'hb5e == _T_221[11:0] ? image_2910 : _GEN_24483; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24485 = 12'hb5f == _T_221[11:0] ? image_2911 : _GEN_24484; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24486 = 12'hb60 == _T_221[11:0] ? image_2912 : _GEN_24485; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24487 = 12'hb61 == _T_221[11:0] ? image_2913 : _GEN_24486; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24488 = 12'hb62 == _T_221[11:0] ? image_2914 : _GEN_24487; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24489 = 12'hb63 == _T_221[11:0] ? image_2915 : _GEN_24488; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24490 = 12'hb64 == _T_221[11:0] ? image_2916 : _GEN_24489; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24491 = 12'hb65 == _T_221[11:0] ? image_2917 : _GEN_24490; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24492 = 12'hb66 == _T_221[11:0] ? image_2918 : _GEN_24491; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24493 = 12'hb67 == _T_221[11:0] ? image_2919 : _GEN_24492; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24494 = 12'hb68 == _T_221[11:0] ? image_2920 : _GEN_24493; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24495 = 12'hb69 == _T_221[11:0] ? image_2921 : _GEN_24494; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24496 = 12'hb6a == _T_221[11:0] ? image_2922 : _GEN_24495; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24497 = 12'hb6b == _T_221[11:0] ? image_2923 : _GEN_24496; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24498 = 12'hb6c == _T_221[11:0] ? image_2924 : _GEN_24497; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24499 = 12'hb6d == _T_221[11:0] ? image_2925 : _GEN_24498; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24500 = 12'hb6e == _T_221[11:0] ? image_2926 : _GEN_24499; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24501 = 12'hb6f == _T_221[11:0] ? image_2927 : _GEN_24500; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24502 = 12'hb70 == _T_221[11:0] ? image_2928 : _GEN_24501; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24503 = 12'hb71 == _T_221[11:0] ? image_2929 : _GEN_24502; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24504 = 12'hb72 == _T_221[11:0] ? image_2930 : _GEN_24503; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24505 = 12'hb73 == _T_221[11:0] ? image_2931 : _GEN_24504; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24506 = 12'hb74 == _T_221[11:0] ? image_2932 : _GEN_24505; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24507 = 12'hb75 == _T_221[11:0] ? image_2933 : _GEN_24506; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24508 = 12'hb76 == _T_221[11:0] ? image_2934 : _GEN_24507; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24509 = 12'hb77 == _T_221[11:0] ? 4'h0 : _GEN_24508; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24510 = 12'hb78 == _T_221[11:0] ? 4'h0 : _GEN_24509; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24511 = 12'hb79 == _T_221[11:0] ? 4'h0 : _GEN_24510; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24512 = 12'hb7a == _T_221[11:0] ? 4'h0 : _GEN_24511; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24513 = 12'hb7b == _T_221[11:0] ? 4'h0 : _GEN_24512; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24514 = 12'hb7c == _T_221[11:0] ? 4'h0 : _GEN_24513; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24515 = 12'hb7d == _T_221[11:0] ? 4'h0 : _GEN_24514; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24516 = 12'hb7e == _T_221[11:0] ? 4'h0 : _GEN_24515; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24517 = 12'hb7f == _T_221[11:0] ? 4'h0 : _GEN_24516; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24518 = 12'hb80 == _T_221[11:0] ? 4'h0 : _GEN_24517; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24519 = 12'hb81 == _T_221[11:0] ? 4'h0 : _GEN_24518; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24520 = 12'hb82 == _T_221[11:0] ? 4'h0 : _GEN_24519; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24521 = 12'hb83 == _T_221[11:0] ? 4'h0 : _GEN_24520; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24522 = 12'hb84 == _T_221[11:0] ? 4'h0 : _GEN_24521; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24523 = 12'hb85 == _T_221[11:0] ? 4'h0 : _GEN_24522; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24524 = 12'hb86 == _T_221[11:0] ? 4'h0 : _GEN_24523; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24525 = 12'hb87 == _T_221[11:0] ? 4'h0 : _GEN_24524; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24526 = 12'hb88 == _T_221[11:0] ? 4'h0 : _GEN_24525; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24527 = 12'hb89 == _T_221[11:0] ? 4'h0 : _GEN_24526; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24528 = 12'hb8a == _T_221[11:0] ? 4'h0 : _GEN_24527; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24529 = 12'hb8b == _T_221[11:0] ? 4'h0 : _GEN_24528; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24530 = 12'hb8c == _T_221[11:0] ? 4'h0 : _GEN_24529; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24531 = 12'hb8d == _T_221[11:0] ? 4'h0 : _GEN_24530; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24532 = 12'hb8e == _T_221[11:0] ? 4'h0 : _GEN_24531; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24533 = 12'hb8f == _T_221[11:0] ? 4'h0 : _GEN_24532; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24534 = 12'hb90 == _T_221[11:0] ? 4'h0 : _GEN_24533; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24535 = 12'hb91 == _T_221[11:0] ? 4'h0 : _GEN_24534; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24536 = 12'hb92 == _T_221[11:0] ? 4'h0 : _GEN_24535; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24537 = 12'hb93 == _T_221[11:0] ? 4'h0 : _GEN_24536; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24538 = 12'hb94 == _T_221[11:0] ? 4'h0 : _GEN_24537; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24539 = 12'hb95 == _T_221[11:0] ? image_2965 : _GEN_24538; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24540 = 12'hb96 == _T_221[11:0] ? image_2966 : _GEN_24539; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24541 = 12'hb97 == _T_221[11:0] ? image_2967 : _GEN_24540; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24542 = 12'hb98 == _T_221[11:0] ? image_2968 : _GEN_24541; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24543 = 12'hb99 == _T_221[11:0] ? image_2969 : _GEN_24542; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24544 = 12'hb9a == _T_221[11:0] ? image_2970 : _GEN_24543; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24545 = 12'hb9b == _T_221[11:0] ? image_2971 : _GEN_24544; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24546 = 12'hb9c == _T_221[11:0] ? image_2972 : _GEN_24545; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24547 = 12'hb9d == _T_221[11:0] ? image_2973 : _GEN_24546; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24548 = 12'hb9e == _T_221[11:0] ? image_2974 : _GEN_24547; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24549 = 12'hb9f == _T_221[11:0] ? image_2975 : _GEN_24548; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24550 = 12'hba0 == _T_221[11:0] ? image_2976 : _GEN_24549; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24551 = 12'hba1 == _T_221[11:0] ? image_2977 : _GEN_24550; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24552 = 12'hba2 == _T_221[11:0] ? image_2978 : _GEN_24551; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24553 = 12'hba3 == _T_221[11:0] ? image_2979 : _GEN_24552; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24554 = 12'hba4 == _T_221[11:0] ? image_2980 : _GEN_24553; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24555 = 12'hba5 == _T_221[11:0] ? image_2981 : _GEN_24554; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24556 = 12'hba6 == _T_221[11:0] ? image_2982 : _GEN_24555; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24557 = 12'hba7 == _T_221[11:0] ? image_2983 : _GEN_24556; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24558 = 12'hba8 == _T_221[11:0] ? image_2984 : _GEN_24557; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24559 = 12'hba9 == _T_221[11:0] ? image_2985 : _GEN_24558; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24560 = 12'hbaa == _T_221[11:0] ? image_2986 : _GEN_24559; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24561 = 12'hbab == _T_221[11:0] ? image_2987 : _GEN_24560; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24562 = 12'hbac == _T_221[11:0] ? image_2988 : _GEN_24561; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24563 = 12'hbad == _T_221[11:0] ? image_2989 : _GEN_24562; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24564 = 12'hbae == _T_221[11:0] ? image_2990 : _GEN_24563; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24565 = 12'hbaf == _T_221[11:0] ? image_2991 : _GEN_24564; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24566 = 12'hbb0 == _T_221[11:0] ? image_2992 : _GEN_24565; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24567 = 12'hbb1 == _T_221[11:0] ? image_2993 : _GEN_24566; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24568 = 12'hbb2 == _T_221[11:0] ? image_2994 : _GEN_24567; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24569 = 12'hbb3 == _T_221[11:0] ? image_2995 : _GEN_24568; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24570 = 12'hbb4 == _T_221[11:0] ? image_2996 : _GEN_24569; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24571 = 12'hbb5 == _T_221[11:0] ? 4'h0 : _GEN_24570; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24572 = 12'hbb6 == _T_221[11:0] ? 4'h0 : _GEN_24571; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24573 = 12'hbb7 == _T_221[11:0] ? 4'h0 : _GEN_24572; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24574 = 12'hbb8 == _T_221[11:0] ? 4'h0 : _GEN_24573; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24575 = 12'hbb9 == _T_221[11:0] ? 4'h0 : _GEN_24574; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24576 = 12'hbba == _T_221[11:0] ? 4'h0 : _GEN_24575; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24577 = 12'hbbb == _T_221[11:0] ? 4'h0 : _GEN_24576; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24578 = 12'hbbc == _T_221[11:0] ? 4'h0 : _GEN_24577; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24579 = 12'hbbd == _T_221[11:0] ? 4'h0 : _GEN_24578; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24580 = 12'hbbe == _T_221[11:0] ? 4'h0 : _GEN_24579; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24581 = 12'hbbf == _T_221[11:0] ? 4'h0 : _GEN_24580; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24582 = 12'hbc0 == _T_221[11:0] ? 4'h0 : _GEN_24581; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24583 = 12'hbc1 == _T_221[11:0] ? 4'h0 : _GEN_24582; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24584 = 12'hbc2 == _T_221[11:0] ? 4'h0 : _GEN_24583; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24585 = 12'hbc3 == _T_221[11:0] ? 4'h0 : _GEN_24584; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24586 = 12'hbc4 == _T_221[11:0] ? 4'h0 : _GEN_24585; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24587 = 12'hbc5 == _T_221[11:0] ? 4'h0 : _GEN_24586; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24588 = 12'hbc6 == _T_221[11:0] ? 4'h0 : _GEN_24587; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24589 = 12'hbc7 == _T_221[11:0] ? 4'h0 : _GEN_24588; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24590 = 12'hbc8 == _T_221[11:0] ? 4'h0 : _GEN_24589; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24591 = 12'hbc9 == _T_221[11:0] ? 4'h0 : _GEN_24590; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24592 = 12'hbca == _T_221[11:0] ? 4'h0 : _GEN_24591; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24593 = 12'hbcb == _T_221[11:0] ? 4'h0 : _GEN_24592; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24594 = 12'hbcc == _T_221[11:0] ? 4'h0 : _GEN_24593; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24595 = 12'hbcd == _T_221[11:0] ? 4'h0 : _GEN_24594; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24596 = 12'hbce == _T_221[11:0] ? 4'h0 : _GEN_24595; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24597 = 12'hbcf == _T_221[11:0] ? 4'h0 : _GEN_24596; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24598 = 12'hbd0 == _T_221[11:0] ? 4'h0 : _GEN_24597; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24599 = 12'hbd1 == _T_221[11:0] ? 4'h0 : _GEN_24598; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24600 = 12'hbd2 == _T_221[11:0] ? 4'h0 : _GEN_24599; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24601 = 12'hbd3 == _T_221[11:0] ? 4'h0 : _GEN_24600; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24602 = 12'hbd4 == _T_221[11:0] ? 4'h0 : _GEN_24601; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24603 = 12'hbd5 == _T_221[11:0] ? 4'h0 : _GEN_24602; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24604 = 12'hbd6 == _T_221[11:0] ? 4'h0 : _GEN_24603; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24605 = 12'hbd7 == _T_221[11:0] ? 4'h0 : _GEN_24604; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24606 = 12'hbd8 == _T_221[11:0] ? 4'h0 : _GEN_24605; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24607 = 12'hbd9 == _T_221[11:0] ? 4'h0 : _GEN_24606; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24608 = 12'hbda == _T_221[11:0] ? 4'h0 : _GEN_24607; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24609 = 12'hbdb == _T_221[11:0] ? image_3035 : _GEN_24608; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24610 = 12'hbdc == _T_221[11:0] ? image_3036 : _GEN_24609; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24611 = 12'hbdd == _T_221[11:0] ? image_3037 : _GEN_24610; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24612 = 12'hbde == _T_221[11:0] ? image_3038 : _GEN_24611; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24613 = 12'hbdf == _T_221[11:0] ? image_3039 : _GEN_24612; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24614 = 12'hbe0 == _T_221[11:0] ? image_3040 : _GEN_24613; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24615 = 12'hbe1 == _T_221[11:0] ? image_3041 : _GEN_24614; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24616 = 12'hbe2 == _T_221[11:0] ? image_3042 : _GEN_24615; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24617 = 12'hbe3 == _T_221[11:0] ? image_3043 : _GEN_24616; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24618 = 12'hbe4 == _T_221[11:0] ? image_3044 : _GEN_24617; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24619 = 12'hbe5 == _T_221[11:0] ? image_3045 : _GEN_24618; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24620 = 12'hbe6 == _T_221[11:0] ? image_3046 : _GEN_24619; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24621 = 12'hbe7 == _T_221[11:0] ? image_3047 : _GEN_24620; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24622 = 12'hbe8 == _T_221[11:0] ? image_3048 : _GEN_24621; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24623 = 12'hbe9 == _T_221[11:0] ? image_3049 : _GEN_24622; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24624 = 12'hbea == _T_221[11:0] ? image_3050 : _GEN_24623; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24625 = 12'hbeb == _T_221[11:0] ? image_3051 : _GEN_24624; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24626 = 12'hbec == _T_221[11:0] ? image_3052 : _GEN_24625; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24627 = 12'hbed == _T_221[11:0] ? image_3053 : _GEN_24626; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24628 = 12'hbee == _T_221[11:0] ? image_3054 : _GEN_24627; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24629 = 12'hbef == _T_221[11:0] ? image_3055 : _GEN_24628; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24630 = 12'hbf0 == _T_221[11:0] ? image_3056 : _GEN_24629; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24631 = 12'hbf1 == _T_221[11:0] ? 4'h0 : _GEN_24630; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24632 = 12'hbf2 == _T_221[11:0] ? 4'h0 : _GEN_24631; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24633 = 12'hbf3 == _T_221[11:0] ? 4'h0 : _GEN_24632; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24634 = 12'hbf4 == _T_221[11:0] ? 4'h0 : _GEN_24633; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24635 = 12'hbf5 == _T_221[11:0] ? 4'h0 : _GEN_24634; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24636 = 12'hbf6 == _T_221[11:0] ? 4'h0 : _GEN_24635; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24637 = 12'hbf7 == _T_221[11:0] ? 4'h0 : _GEN_24636; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24638 = 12'hbf8 == _T_221[11:0] ? 4'h0 : _GEN_24637; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24639 = 12'hbf9 == _T_221[11:0] ? 4'h0 : _GEN_24638; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24640 = 12'hbfa == _T_221[11:0] ? 4'h0 : _GEN_24639; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24641 = 12'hbfb == _T_221[11:0] ? 4'h0 : _GEN_24640; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24642 = 12'hbfc == _T_221[11:0] ? 4'h0 : _GEN_24641; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24643 = 12'hbfd == _T_221[11:0] ? 4'h0 : _GEN_24642; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24644 = 12'hbfe == _T_221[11:0] ? 4'h0 : _GEN_24643; // @[Filter.scala 138:46]
  wire [3:0] _GEN_24645 = 12'hbff == _T_221[11:0] ? 4'h0 : _GEN_24644; // @[Filter.scala 138:46]
  wire [7:0] _GEN_24648 = 3'h1 == io_SPI_filterIndex[2:0] ? $signed(8'sh9) : $signed(8'sh1); // @[Filter.scala 154:53]
  wire [7:0] _GEN_24649 = 3'h2 == io_SPI_filterIndex[2:0] ? $signed(8'sh10) : $signed(_GEN_24648); // @[Filter.scala 154:53]
  wire [7:0] _GEN_24650 = 3'h3 == io_SPI_filterIndex[2:0] ? $signed(8'sh1) : $signed(_GEN_24649); // @[Filter.scala 154:53]
  wire [7:0] _GEN_24651 = 3'h4 == io_SPI_filterIndex[2:0] ? $signed(8'sh1) : $signed(_GEN_24650); // @[Filter.scala 154:53]
  wire [7:0] _GEN_24652 = 3'h5 == io_SPI_filterIndex[2:0] ? $signed(8'sh1) : $signed(_GEN_24651); // @[Filter.scala 154:53]
  wire [8:0] _GEN_24829 = {{1{_GEN_24652[7]}},_GEN_24652}; // @[Filter.scala 154:53]
  wire [9:0] _T_225 = $signed(KernelConvolution_io_pixelVal_out_0) / $signed(_GEN_24829); // @[Filter.scala 154:64]
  wire [9:0] _T_232 = $signed(KernelConvolution_io_pixelVal_out_1) / $signed(_GEN_24829); // @[Filter.scala 154:64]
  wire [9:0] _T_239 = $signed(KernelConvolution_io_pixelVal_out_2) / $signed(_GEN_24829); // @[Filter.scala 154:64]
  wire [9:0] _T_246 = $signed(KernelConvolution_io_pixelVal_out_3) / $signed(_GEN_24829); // @[Filter.scala 154:64]
  wire [9:0] _T_253 = $signed(KernelConvolution_io_pixelVal_out_4) / $signed(_GEN_24829); // @[Filter.scala 154:64]
  wire [9:0] _T_260 = $signed(KernelConvolution_io_pixelVal_out_5) / $signed(_GEN_24829); // @[Filter.scala 154:64]
  wire [9:0] _T_267 = $signed(KernelConvolution_io_pixelVal_out_6) / $signed(_GEN_24829); // @[Filter.scala 154:64]
  wire [9:0] _T_274 = $signed(KernelConvolution_io_pixelVal_out_7) / $signed(_GEN_24829); // @[Filter.scala 154:64]
  wire [31:0] _T_280 = pixelIndex + 32'h8; // @[Filter.scala 163:34]
  wire [12:0] _T_281 = 7'h40 * 7'h30; // @[Filter.scala 164:42]
  wire [31:0] _GEN_24845 = {{19'd0}, _T_281}; // @[Filter.scala 164:25]
  wire  _T_282 = pixelIndex == _GEN_24845; // @[Filter.scala 164:25]
  KernelConvolution KernelConvolution ( // @[Filter.scala 122:35]
    .clock(KernelConvolution_clock),
    .reset(KernelConvolution_reset),
    .io_kernelVal_in(KernelConvolution_io_kernelVal_in),
    .io_pixelVal_in_0(KernelConvolution_io_pixelVal_in_0),
    .io_pixelVal_in_1(KernelConvolution_io_pixelVal_in_1),
    .io_pixelVal_in_2(KernelConvolution_io_pixelVal_in_2),
    .io_pixelVal_in_3(KernelConvolution_io_pixelVal_in_3),
    .io_pixelVal_in_4(KernelConvolution_io_pixelVal_in_4),
    .io_pixelVal_in_5(KernelConvolution_io_pixelVal_in_5),
    .io_pixelVal_in_6(KernelConvolution_io_pixelVal_in_6),
    .io_pixelVal_in_7(KernelConvolution_io_pixelVal_in_7),
    .io_pixelVal_out_0(KernelConvolution_io_pixelVal_out_0),
    .io_pixelVal_out_1(KernelConvolution_io_pixelVal_out_1),
    .io_pixelVal_out_2(KernelConvolution_io_pixelVal_out_2),
    .io_pixelVal_out_3(KernelConvolution_io_pixelVal_out_3),
    .io_pixelVal_out_4(KernelConvolution_io_pixelVal_out_4),
    .io_pixelVal_out_5(KernelConvolution_io_pixelVal_out_5),
    .io_pixelVal_out_6(KernelConvolution_io_pixelVal_out_6),
    .io_pixelVal_out_7(KernelConvolution_io_pixelVal_out_7),
    .io_valid_out(KernelConvolution_io_valid_out)
  );
  assign io_pixelVal_out_0 = _T_225[3:0]; // @[Filter.scala 154:32 Filter.scala 156:32]
  assign io_pixelVal_out_1 = _T_232[3:0]; // @[Filter.scala 154:32 Filter.scala 156:32]
  assign io_pixelVal_out_2 = _T_239[3:0]; // @[Filter.scala 154:32 Filter.scala 156:32]
  assign io_pixelVal_out_3 = _T_246[3:0]; // @[Filter.scala 154:32 Filter.scala 156:32]
  assign io_pixelVal_out_4 = _T_253[3:0]; // @[Filter.scala 154:32 Filter.scala 156:32]
  assign io_pixelVal_out_5 = _T_260[3:0]; // @[Filter.scala 154:32 Filter.scala 156:32]
  assign io_pixelVal_out_6 = _T_267[3:0]; // @[Filter.scala 154:32 Filter.scala 156:32]
  assign io_pixelVal_out_7 = _T_274[3:0]; // @[Filter.scala 154:32 Filter.scala 156:32]
  assign io_valid_out = KernelConvolution_io_valid_out; // @[Filter.scala 160:18]
  assign KernelConvolution_clock = clock;
  assign KernelConvolution_reset = reset;
  assign KernelConvolution_io_kernelVal_in = _GEN_24787 & _GEN_24714 ? $signed(5'sh0) : $signed(_GEN_55); // @[Filter.scala 125:36]
  assign KernelConvolution_io_pixelVal_in_0 = _T_43 ? 4'h0 : _GEN_3134; // @[Filter.scala 136:46 Filter.scala 138:46]
  assign KernelConvolution_io_pixelVal_in_1 = _T_68 ? 4'h0 : _GEN_6207; // @[Filter.scala 136:46 Filter.scala 138:46]
  assign KernelConvolution_io_pixelVal_in_2 = _T_93 ? 4'h0 : _GEN_9280; // @[Filter.scala 136:46 Filter.scala 138:46]
  assign KernelConvolution_io_pixelVal_in_3 = _T_118 ? 4'h0 : _GEN_12353; // @[Filter.scala 136:46 Filter.scala 138:46]
  assign KernelConvolution_io_pixelVal_in_4 = _T_143 ? 4'h0 : _GEN_15426; // @[Filter.scala 136:46 Filter.scala 138:46]
  assign KernelConvolution_io_pixelVal_in_5 = _T_168 ? 4'h0 : _GEN_18499; // @[Filter.scala 136:46 Filter.scala 138:46]
  assign KernelConvolution_io_pixelVal_in_6 = _T_193 ? 4'h0 : _GEN_21572; // @[Filter.scala 136:46 Filter.scala 138:46]
  assign KernelConvolution_io_pixelVal_in_7 = _T_218 ? 4'h0 : _GEN_24645; // @[Filter.scala 136:46 Filter.scala 138:46]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  image_12 = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  image_14 = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  image_15 = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  image_16 = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  image_17 = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  image_18 = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  image_19 = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  image_20 = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  image_21 = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  image_22 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  image_23 = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  image_35 = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  image_36 = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  image_37 = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  image_38 = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  image_39 = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  image_40 = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  image_41 = _RAND_17[3:0];
  _RAND_18 = {1{`RANDOM}};
  image_42 = _RAND_18[3:0];
  _RAND_19 = {1{`RANDOM}};
  image_75 = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  image_76 = _RAND_20[3:0];
  _RAND_21 = {1{`RANDOM}};
  image_77 = _RAND_21[3:0];
  _RAND_22 = {1{`RANDOM}};
  image_78 = _RAND_22[3:0];
  _RAND_23 = {1{`RANDOM}};
  image_79 = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
  image_80 = _RAND_24[3:0];
  _RAND_25 = {1{`RANDOM}};
  image_81 = _RAND_25[3:0];
  _RAND_26 = {1{`RANDOM}};
  image_82 = _RAND_26[3:0];
  _RAND_27 = {1{`RANDOM}};
  image_83 = _RAND_27[3:0];
  _RAND_28 = {1{`RANDOM}};
  image_84 = _RAND_28[3:0];
  _RAND_29 = {1{`RANDOM}};
  image_85 = _RAND_29[3:0];
  _RAND_30 = {1{`RANDOM}};
  image_86 = _RAND_30[3:0];
  _RAND_31 = {1{`RANDOM}};
  image_87 = _RAND_31[3:0];
  _RAND_32 = {1{`RANDOM}};
  image_88 = _RAND_32[3:0];
  _RAND_33 = {1{`RANDOM}};
  image_89 = _RAND_33[3:0];
  _RAND_34 = {1{`RANDOM}};
  image_90 = _RAND_34[3:0];
  _RAND_35 = {1{`RANDOM}};
  image_93 = _RAND_35[3:0];
  _RAND_36 = {1{`RANDOM}};
  image_95 = _RAND_36[3:0];
  _RAND_37 = {1{`RANDOM}};
  image_96 = _RAND_37[3:0];
  _RAND_38 = {1{`RANDOM}};
  image_97 = _RAND_38[3:0];
  _RAND_39 = {1{`RANDOM}};
  image_98 = _RAND_39[3:0];
  _RAND_40 = {1{`RANDOM}};
  image_99 = _RAND_40[3:0];
  _RAND_41 = {1{`RANDOM}};
  image_100 = _RAND_41[3:0];
  _RAND_42 = {1{`RANDOM}};
  image_101 = _RAND_42[3:0];
  _RAND_43 = {1{`RANDOM}};
  image_102 = _RAND_43[3:0];
  _RAND_44 = {1{`RANDOM}};
  image_103 = _RAND_44[3:0];
  _RAND_45 = {1{`RANDOM}};
  image_104 = _RAND_45[3:0];
  _RAND_46 = {1{`RANDOM}};
  image_105 = _RAND_46[3:0];
  _RAND_47 = {1{`RANDOM}};
  image_106 = _RAND_47[3:0];
  _RAND_48 = {1{`RANDOM}};
  image_107 = _RAND_48[3:0];
  _RAND_49 = {1{`RANDOM}};
  image_108 = _RAND_49[3:0];
  _RAND_50 = {1{`RANDOM}};
  image_136 = _RAND_50[3:0];
  _RAND_51 = {1{`RANDOM}};
  image_137 = _RAND_51[3:0];
  _RAND_52 = {1{`RANDOM}};
  image_138 = _RAND_52[3:0];
  _RAND_53 = {1{`RANDOM}};
  image_139 = _RAND_53[3:0];
  _RAND_54 = {1{`RANDOM}};
  image_140 = _RAND_54[3:0];
  _RAND_55 = {1{`RANDOM}};
  image_141 = _RAND_55[3:0];
  _RAND_56 = {1{`RANDOM}};
  image_142 = _RAND_56[3:0];
  _RAND_57 = {1{`RANDOM}};
  image_143 = _RAND_57[3:0];
  _RAND_58 = {1{`RANDOM}};
  image_144 = _RAND_58[3:0];
  _RAND_59 = {1{`RANDOM}};
  image_145 = _RAND_59[3:0];
  _RAND_60 = {1{`RANDOM}};
  image_146 = _RAND_60[3:0];
  _RAND_61 = {1{`RANDOM}};
  image_147 = _RAND_61[3:0];
  _RAND_62 = {1{`RANDOM}};
  image_148 = _RAND_62[3:0];
  _RAND_63 = {1{`RANDOM}};
  image_149 = _RAND_63[3:0];
  _RAND_64 = {1{`RANDOM}};
  image_150 = _RAND_64[3:0];
  _RAND_65 = {1{`RANDOM}};
  image_151 = _RAND_65[3:0];
  _RAND_66 = {1{`RANDOM}};
  image_152 = _RAND_66[3:0];
  _RAND_67 = {1{`RANDOM}};
  image_153 = _RAND_67[3:0];
  _RAND_68 = {1{`RANDOM}};
  image_154 = _RAND_68[3:0];
  _RAND_69 = {1{`RANDOM}};
  image_155 = _RAND_69[3:0];
  _RAND_70 = {1{`RANDOM}};
  image_157 = _RAND_70[3:0];
  _RAND_71 = {1{`RANDOM}};
  image_158 = _RAND_71[3:0];
  _RAND_72 = {1{`RANDOM}};
  image_159 = _RAND_72[3:0];
  _RAND_73 = {1{`RANDOM}};
  image_160 = _RAND_73[3:0];
  _RAND_74 = {1{`RANDOM}};
  image_161 = _RAND_74[3:0];
  _RAND_75 = {1{`RANDOM}};
  image_162 = _RAND_75[3:0];
  _RAND_76 = {1{`RANDOM}};
  image_163 = _RAND_76[3:0];
  _RAND_77 = {1{`RANDOM}};
  image_164 = _RAND_77[3:0];
  _RAND_78 = {1{`RANDOM}};
  image_165 = _RAND_78[3:0];
  _RAND_79 = {1{`RANDOM}};
  image_166 = _RAND_79[3:0];
  _RAND_80 = {1{`RANDOM}};
  image_167 = _RAND_80[3:0];
  _RAND_81 = {1{`RANDOM}};
  image_168 = _RAND_81[3:0];
  _RAND_82 = {1{`RANDOM}};
  image_169 = _RAND_82[3:0];
  _RAND_83 = {1{`RANDOM}};
  image_170 = _RAND_83[3:0];
  _RAND_84 = {1{`RANDOM}};
  image_171 = _RAND_84[3:0];
  _RAND_85 = {1{`RANDOM}};
  image_172 = _RAND_85[3:0];
  _RAND_86 = {1{`RANDOM}};
  image_173 = _RAND_86[3:0];
  _RAND_87 = {1{`RANDOM}};
  image_174 = _RAND_87[3:0];
  _RAND_88 = {1{`RANDOM}};
  image_175 = _RAND_88[3:0];
  _RAND_89 = {1{`RANDOM}};
  image_176 = _RAND_89[3:0];
  _RAND_90 = {1{`RANDOM}};
  image_177 = _RAND_90[3:0];
  _RAND_91 = {1{`RANDOM}};
  image_178 = _RAND_91[3:0];
  _RAND_92 = {1{`RANDOM}};
  image_179 = _RAND_92[3:0];
  _RAND_93 = {1{`RANDOM}};
  image_199 = _RAND_93[3:0];
  _RAND_94 = {1{`RANDOM}};
  image_200 = _RAND_94[3:0];
  _RAND_95 = {1{`RANDOM}};
  image_201 = _RAND_95[3:0];
  _RAND_96 = {1{`RANDOM}};
  image_202 = _RAND_96[3:0];
  _RAND_97 = {1{`RANDOM}};
  image_203 = _RAND_97[3:0];
  _RAND_98 = {1{`RANDOM}};
  image_204 = _RAND_98[3:0];
  _RAND_99 = {1{`RANDOM}};
  image_205 = _RAND_99[3:0];
  _RAND_100 = {1{`RANDOM}};
  image_206 = _RAND_100[3:0];
  _RAND_101 = {1{`RANDOM}};
  image_207 = _RAND_101[3:0];
  _RAND_102 = {1{`RANDOM}};
  image_208 = _RAND_102[3:0];
  _RAND_103 = {1{`RANDOM}};
  image_209 = _RAND_103[3:0];
  _RAND_104 = {1{`RANDOM}};
  image_210 = _RAND_104[3:0];
  _RAND_105 = {1{`RANDOM}};
  image_211 = _RAND_105[3:0];
  _RAND_106 = {1{`RANDOM}};
  image_212 = _RAND_106[3:0];
  _RAND_107 = {1{`RANDOM}};
  image_213 = _RAND_107[3:0];
  _RAND_108 = {1{`RANDOM}};
  image_214 = _RAND_108[3:0];
  _RAND_109 = {1{`RANDOM}};
  image_215 = _RAND_109[3:0];
  _RAND_110 = {1{`RANDOM}};
  image_216 = _RAND_110[3:0];
  _RAND_111 = {1{`RANDOM}};
  image_217 = _RAND_111[3:0];
  _RAND_112 = {1{`RANDOM}};
  image_218 = _RAND_112[3:0];
  _RAND_113 = {1{`RANDOM}};
  image_219 = _RAND_113[3:0];
  _RAND_114 = {1{`RANDOM}};
  image_220 = _RAND_114[3:0];
  _RAND_115 = {1{`RANDOM}};
  image_221 = _RAND_115[3:0];
  _RAND_116 = {1{`RANDOM}};
  image_222 = _RAND_116[3:0];
  _RAND_117 = {1{`RANDOM}};
  image_223 = _RAND_117[3:0];
  _RAND_118 = {1{`RANDOM}};
  image_224 = _RAND_118[3:0];
  _RAND_119 = {1{`RANDOM}};
  image_225 = _RAND_119[3:0];
  _RAND_120 = {1{`RANDOM}};
  image_226 = _RAND_120[3:0];
  _RAND_121 = {1{`RANDOM}};
  image_227 = _RAND_121[3:0];
  _RAND_122 = {1{`RANDOM}};
  image_228 = _RAND_122[3:0];
  _RAND_123 = {1{`RANDOM}};
  image_229 = _RAND_123[3:0];
  _RAND_124 = {1{`RANDOM}};
  image_230 = _RAND_124[3:0];
  _RAND_125 = {1{`RANDOM}};
  image_231 = _RAND_125[3:0];
  _RAND_126 = {1{`RANDOM}};
  image_232 = _RAND_126[3:0];
  _RAND_127 = {1{`RANDOM}};
  image_233 = _RAND_127[3:0];
  _RAND_128 = {1{`RANDOM}};
  image_234 = _RAND_128[3:0];
  _RAND_129 = {1{`RANDOM}};
  image_235 = _RAND_129[3:0];
  _RAND_130 = {1{`RANDOM}};
  image_236 = _RAND_130[3:0];
  _RAND_131 = {1{`RANDOM}};
  image_237 = _RAND_131[3:0];
  _RAND_132 = {1{`RANDOM}};
  image_238 = _RAND_132[3:0];
  _RAND_133 = {1{`RANDOM}};
  image_239 = _RAND_133[3:0];
  _RAND_134 = {1{`RANDOM}};
  image_240 = _RAND_134[3:0];
  _RAND_135 = {1{`RANDOM}};
  image_241 = _RAND_135[3:0];
  _RAND_136 = {1{`RANDOM}};
  image_242 = _RAND_136[3:0];
  _RAND_137 = {1{`RANDOM}};
  image_243 = _RAND_137[3:0];
  _RAND_138 = {1{`RANDOM}};
  image_244 = _RAND_138[3:0];
  _RAND_139 = {1{`RANDOM}};
  image_245 = _RAND_139[3:0];
  _RAND_140 = {1{`RANDOM}};
  image_246 = _RAND_140[3:0];
  _RAND_141 = {1{`RANDOM}};
  image_262 = _RAND_141[3:0];
  _RAND_142 = {1{`RANDOM}};
  image_263 = _RAND_142[3:0];
  _RAND_143 = {1{`RANDOM}};
  image_264 = _RAND_143[3:0];
  _RAND_144 = {1{`RANDOM}};
  image_265 = _RAND_144[3:0];
  _RAND_145 = {1{`RANDOM}};
  image_266 = _RAND_145[3:0];
  _RAND_146 = {1{`RANDOM}};
  image_267 = _RAND_146[3:0];
  _RAND_147 = {1{`RANDOM}};
  image_268 = _RAND_147[3:0];
  _RAND_148 = {1{`RANDOM}};
  image_269 = _RAND_148[3:0];
  _RAND_149 = {1{`RANDOM}};
  image_270 = _RAND_149[3:0];
  _RAND_150 = {1{`RANDOM}};
  image_271 = _RAND_150[3:0];
  _RAND_151 = {1{`RANDOM}};
  image_272 = _RAND_151[3:0];
  _RAND_152 = {1{`RANDOM}};
  image_273 = _RAND_152[3:0];
  _RAND_153 = {1{`RANDOM}};
  image_274 = _RAND_153[3:0];
  _RAND_154 = {1{`RANDOM}};
  image_275 = _RAND_154[3:0];
  _RAND_155 = {1{`RANDOM}};
  image_276 = _RAND_155[3:0];
  _RAND_156 = {1{`RANDOM}};
  image_277 = _RAND_156[3:0];
  _RAND_157 = {1{`RANDOM}};
  image_278 = _RAND_157[3:0];
  _RAND_158 = {1{`RANDOM}};
  image_279 = _RAND_158[3:0];
  _RAND_159 = {1{`RANDOM}};
  image_280 = _RAND_159[3:0];
  _RAND_160 = {1{`RANDOM}};
  image_281 = _RAND_160[3:0];
  _RAND_161 = {1{`RANDOM}};
  image_282 = _RAND_161[3:0];
  _RAND_162 = {1{`RANDOM}};
  image_283 = _RAND_162[3:0];
  _RAND_163 = {1{`RANDOM}};
  image_284 = _RAND_163[3:0];
  _RAND_164 = {1{`RANDOM}};
  image_285 = _RAND_164[3:0];
  _RAND_165 = {1{`RANDOM}};
  image_286 = _RAND_165[3:0];
  _RAND_166 = {1{`RANDOM}};
  image_287 = _RAND_166[3:0];
  _RAND_167 = {1{`RANDOM}};
  image_288 = _RAND_167[3:0];
  _RAND_168 = {1{`RANDOM}};
  image_289 = _RAND_168[3:0];
  _RAND_169 = {1{`RANDOM}};
  image_290 = _RAND_169[3:0];
  _RAND_170 = {1{`RANDOM}};
  image_291 = _RAND_170[3:0];
  _RAND_171 = {1{`RANDOM}};
  image_292 = _RAND_171[3:0];
  _RAND_172 = {1{`RANDOM}};
  image_293 = _RAND_172[3:0];
  _RAND_173 = {1{`RANDOM}};
  image_294 = _RAND_173[3:0];
  _RAND_174 = {1{`RANDOM}};
  image_295 = _RAND_174[3:0];
  _RAND_175 = {1{`RANDOM}};
  image_296 = _RAND_175[3:0];
  _RAND_176 = {1{`RANDOM}};
  image_297 = _RAND_176[3:0];
  _RAND_177 = {1{`RANDOM}};
  image_298 = _RAND_177[3:0];
  _RAND_178 = {1{`RANDOM}};
  image_299 = _RAND_178[3:0];
  _RAND_179 = {1{`RANDOM}};
  image_300 = _RAND_179[3:0];
  _RAND_180 = {1{`RANDOM}};
  image_301 = _RAND_180[3:0];
  _RAND_181 = {1{`RANDOM}};
  image_302 = _RAND_181[3:0];
  _RAND_182 = {1{`RANDOM}};
  image_303 = _RAND_182[3:0];
  _RAND_183 = {1{`RANDOM}};
  image_304 = _RAND_183[3:0];
  _RAND_184 = {1{`RANDOM}};
  image_305 = _RAND_184[3:0];
  _RAND_185 = {1{`RANDOM}};
  image_306 = _RAND_185[3:0];
  _RAND_186 = {1{`RANDOM}};
  image_307 = _RAND_186[3:0];
  _RAND_187 = {1{`RANDOM}};
  image_308 = _RAND_187[3:0];
  _RAND_188 = {1{`RANDOM}};
  image_309 = _RAND_188[3:0];
  _RAND_189 = {1{`RANDOM}};
  image_310 = _RAND_189[3:0];
  _RAND_190 = {1{`RANDOM}};
  image_311 = _RAND_190[3:0];
  _RAND_191 = {1{`RANDOM}};
  image_312 = _RAND_191[3:0];
  _RAND_192 = {1{`RANDOM}};
  image_313 = _RAND_192[3:0];
  _RAND_193 = {1{`RANDOM}};
  image_314 = _RAND_193[3:0];
  _RAND_194 = {1{`RANDOM}};
  image_315 = _RAND_194[3:0];
  _RAND_195 = {1{`RANDOM}};
  image_325 = _RAND_195[3:0];
  _RAND_196 = {1{`RANDOM}};
  image_326 = _RAND_196[3:0];
  _RAND_197 = {1{`RANDOM}};
  image_327 = _RAND_197[3:0];
  _RAND_198 = {1{`RANDOM}};
  image_328 = _RAND_198[3:0];
  _RAND_199 = {1{`RANDOM}};
  image_329 = _RAND_199[3:0];
  _RAND_200 = {1{`RANDOM}};
  image_330 = _RAND_200[3:0];
  _RAND_201 = {1{`RANDOM}};
  image_331 = _RAND_201[3:0];
  _RAND_202 = {1{`RANDOM}};
  image_332 = _RAND_202[3:0];
  _RAND_203 = {1{`RANDOM}};
  image_333 = _RAND_203[3:0];
  _RAND_204 = {1{`RANDOM}};
  image_334 = _RAND_204[3:0];
  _RAND_205 = {1{`RANDOM}};
  image_335 = _RAND_205[3:0];
  _RAND_206 = {1{`RANDOM}};
  image_336 = _RAND_206[3:0];
  _RAND_207 = {1{`RANDOM}};
  image_337 = _RAND_207[3:0];
  _RAND_208 = {1{`RANDOM}};
  image_338 = _RAND_208[3:0];
  _RAND_209 = {1{`RANDOM}};
  image_339 = _RAND_209[3:0];
  _RAND_210 = {1{`RANDOM}};
  image_340 = _RAND_210[3:0];
  _RAND_211 = {1{`RANDOM}};
  image_341 = _RAND_211[3:0];
  _RAND_212 = {1{`RANDOM}};
  image_342 = _RAND_212[3:0];
  _RAND_213 = {1{`RANDOM}};
  image_343 = _RAND_213[3:0];
  _RAND_214 = {1{`RANDOM}};
  image_344 = _RAND_214[3:0];
  _RAND_215 = {1{`RANDOM}};
  image_345 = _RAND_215[3:0];
  _RAND_216 = {1{`RANDOM}};
  image_346 = _RAND_216[3:0];
  _RAND_217 = {1{`RANDOM}};
  image_347 = _RAND_217[3:0];
  _RAND_218 = {1{`RANDOM}};
  image_348 = _RAND_218[3:0];
  _RAND_219 = {1{`RANDOM}};
  image_349 = _RAND_219[3:0];
  _RAND_220 = {1{`RANDOM}};
  image_350 = _RAND_220[3:0];
  _RAND_221 = {1{`RANDOM}};
  image_351 = _RAND_221[3:0];
  _RAND_222 = {1{`RANDOM}};
  image_352 = _RAND_222[3:0];
  _RAND_223 = {1{`RANDOM}};
  image_353 = _RAND_223[3:0];
  _RAND_224 = {1{`RANDOM}};
  image_354 = _RAND_224[3:0];
  _RAND_225 = {1{`RANDOM}};
  image_355 = _RAND_225[3:0];
  _RAND_226 = {1{`RANDOM}};
  image_356 = _RAND_226[3:0];
  _RAND_227 = {1{`RANDOM}};
  image_357 = _RAND_227[3:0];
  _RAND_228 = {1{`RANDOM}};
  image_358 = _RAND_228[3:0];
  _RAND_229 = {1{`RANDOM}};
  image_359 = _RAND_229[3:0];
  _RAND_230 = {1{`RANDOM}};
  image_360 = _RAND_230[3:0];
  _RAND_231 = {1{`RANDOM}};
  image_361 = _RAND_231[3:0];
  _RAND_232 = {1{`RANDOM}};
  image_362 = _RAND_232[3:0];
  _RAND_233 = {1{`RANDOM}};
  image_363 = _RAND_233[3:0];
  _RAND_234 = {1{`RANDOM}};
  image_364 = _RAND_234[3:0];
  _RAND_235 = {1{`RANDOM}};
  image_365 = _RAND_235[3:0];
  _RAND_236 = {1{`RANDOM}};
  image_366 = _RAND_236[3:0];
  _RAND_237 = {1{`RANDOM}};
  image_367 = _RAND_237[3:0];
  _RAND_238 = {1{`RANDOM}};
  image_368 = _RAND_238[3:0];
  _RAND_239 = {1{`RANDOM}};
  image_369 = _RAND_239[3:0];
  _RAND_240 = {1{`RANDOM}};
  image_370 = _RAND_240[3:0];
  _RAND_241 = {1{`RANDOM}};
  image_371 = _RAND_241[3:0];
  _RAND_242 = {1{`RANDOM}};
  image_372 = _RAND_242[3:0];
  _RAND_243 = {1{`RANDOM}};
  image_373 = _RAND_243[3:0];
  _RAND_244 = {1{`RANDOM}};
  image_374 = _RAND_244[3:0];
  _RAND_245 = {1{`RANDOM}};
  image_375 = _RAND_245[3:0];
  _RAND_246 = {1{`RANDOM}};
  image_376 = _RAND_246[3:0];
  _RAND_247 = {1{`RANDOM}};
  image_377 = _RAND_247[3:0];
  _RAND_248 = {1{`RANDOM}};
  image_378 = _RAND_248[3:0];
  _RAND_249 = {1{`RANDOM}};
  image_379 = _RAND_249[3:0];
  _RAND_250 = {1{`RANDOM}};
  image_388 = _RAND_250[3:0];
  _RAND_251 = {1{`RANDOM}};
  image_389 = _RAND_251[3:0];
  _RAND_252 = {1{`RANDOM}};
  image_390 = _RAND_252[3:0];
  _RAND_253 = {1{`RANDOM}};
  image_391 = _RAND_253[3:0];
  _RAND_254 = {1{`RANDOM}};
  image_392 = _RAND_254[3:0];
  _RAND_255 = {1{`RANDOM}};
  image_393 = _RAND_255[3:0];
  _RAND_256 = {1{`RANDOM}};
  image_394 = _RAND_256[3:0];
  _RAND_257 = {1{`RANDOM}};
  image_395 = _RAND_257[3:0];
  _RAND_258 = {1{`RANDOM}};
  image_396 = _RAND_258[3:0];
  _RAND_259 = {1{`RANDOM}};
  image_397 = _RAND_259[3:0];
  _RAND_260 = {1{`RANDOM}};
  image_398 = _RAND_260[3:0];
  _RAND_261 = {1{`RANDOM}};
  image_399 = _RAND_261[3:0];
  _RAND_262 = {1{`RANDOM}};
  image_400 = _RAND_262[3:0];
  _RAND_263 = {1{`RANDOM}};
  image_401 = _RAND_263[3:0];
  _RAND_264 = {1{`RANDOM}};
  image_402 = _RAND_264[3:0];
  _RAND_265 = {1{`RANDOM}};
  image_403 = _RAND_265[3:0];
  _RAND_266 = {1{`RANDOM}};
  image_404 = _RAND_266[3:0];
  _RAND_267 = {1{`RANDOM}};
  image_405 = _RAND_267[3:0];
  _RAND_268 = {1{`RANDOM}};
  image_406 = _RAND_268[3:0];
  _RAND_269 = {1{`RANDOM}};
  image_407 = _RAND_269[3:0];
  _RAND_270 = {1{`RANDOM}};
  image_408 = _RAND_270[3:0];
  _RAND_271 = {1{`RANDOM}};
  image_409 = _RAND_271[3:0];
  _RAND_272 = {1{`RANDOM}};
  image_410 = _RAND_272[3:0];
  _RAND_273 = {1{`RANDOM}};
  image_411 = _RAND_273[3:0];
  _RAND_274 = {1{`RANDOM}};
  image_412 = _RAND_274[3:0];
  _RAND_275 = {1{`RANDOM}};
  image_413 = _RAND_275[3:0];
  _RAND_276 = {1{`RANDOM}};
  image_414 = _RAND_276[3:0];
  _RAND_277 = {1{`RANDOM}};
  image_415 = _RAND_277[3:0];
  _RAND_278 = {1{`RANDOM}};
  image_416 = _RAND_278[3:0];
  _RAND_279 = {1{`RANDOM}};
  image_417 = _RAND_279[3:0];
  _RAND_280 = {1{`RANDOM}};
  image_418 = _RAND_280[3:0];
  _RAND_281 = {1{`RANDOM}};
  image_419 = _RAND_281[3:0];
  _RAND_282 = {1{`RANDOM}};
  image_420 = _RAND_282[3:0];
  _RAND_283 = {1{`RANDOM}};
  image_421 = _RAND_283[3:0];
  _RAND_284 = {1{`RANDOM}};
  image_422 = _RAND_284[3:0];
  _RAND_285 = {1{`RANDOM}};
  image_423 = _RAND_285[3:0];
  _RAND_286 = {1{`RANDOM}};
  image_424 = _RAND_286[3:0];
  _RAND_287 = {1{`RANDOM}};
  image_425 = _RAND_287[3:0];
  _RAND_288 = {1{`RANDOM}};
  image_426 = _RAND_288[3:0];
  _RAND_289 = {1{`RANDOM}};
  image_427 = _RAND_289[3:0];
  _RAND_290 = {1{`RANDOM}};
  image_428 = _RAND_290[3:0];
  _RAND_291 = {1{`RANDOM}};
  image_429 = _RAND_291[3:0];
  _RAND_292 = {1{`RANDOM}};
  image_430 = _RAND_292[3:0];
  _RAND_293 = {1{`RANDOM}};
  image_431 = _RAND_293[3:0];
  _RAND_294 = {1{`RANDOM}};
  image_432 = _RAND_294[3:0];
  _RAND_295 = {1{`RANDOM}};
  image_433 = _RAND_295[3:0];
  _RAND_296 = {1{`RANDOM}};
  image_434 = _RAND_296[3:0];
  _RAND_297 = {1{`RANDOM}};
  image_435 = _RAND_297[3:0];
  _RAND_298 = {1{`RANDOM}};
  image_436 = _RAND_298[3:0];
  _RAND_299 = {1{`RANDOM}};
  image_437 = _RAND_299[3:0];
  _RAND_300 = {1{`RANDOM}};
  image_438 = _RAND_300[3:0];
  _RAND_301 = {1{`RANDOM}};
  image_439 = _RAND_301[3:0];
  _RAND_302 = {1{`RANDOM}};
  image_440 = _RAND_302[3:0];
  _RAND_303 = {1{`RANDOM}};
  image_441 = _RAND_303[3:0];
  _RAND_304 = {1{`RANDOM}};
  image_442 = _RAND_304[3:0];
  _RAND_305 = {1{`RANDOM}};
  image_443 = _RAND_305[3:0];
  _RAND_306 = {1{`RANDOM}};
  image_444 = _RAND_306[3:0];
  _RAND_307 = {1{`RANDOM}};
  image_451 = _RAND_307[3:0];
  _RAND_308 = {1{`RANDOM}};
  image_452 = _RAND_308[3:0];
  _RAND_309 = {1{`RANDOM}};
  image_453 = _RAND_309[3:0];
  _RAND_310 = {1{`RANDOM}};
  image_454 = _RAND_310[3:0];
  _RAND_311 = {1{`RANDOM}};
  image_455 = _RAND_311[3:0];
  _RAND_312 = {1{`RANDOM}};
  image_456 = _RAND_312[3:0];
  _RAND_313 = {1{`RANDOM}};
  image_457 = _RAND_313[3:0];
  _RAND_314 = {1{`RANDOM}};
  image_458 = _RAND_314[3:0];
  _RAND_315 = {1{`RANDOM}};
  image_459 = _RAND_315[3:0];
  _RAND_316 = {1{`RANDOM}};
  image_460 = _RAND_316[3:0];
  _RAND_317 = {1{`RANDOM}};
  image_461 = _RAND_317[3:0];
  _RAND_318 = {1{`RANDOM}};
  image_462 = _RAND_318[3:0];
  _RAND_319 = {1{`RANDOM}};
  image_463 = _RAND_319[3:0];
  _RAND_320 = {1{`RANDOM}};
  image_464 = _RAND_320[3:0];
  _RAND_321 = {1{`RANDOM}};
  image_465 = _RAND_321[3:0];
  _RAND_322 = {1{`RANDOM}};
  image_466 = _RAND_322[3:0];
  _RAND_323 = {1{`RANDOM}};
  image_467 = _RAND_323[3:0];
  _RAND_324 = {1{`RANDOM}};
  image_468 = _RAND_324[3:0];
  _RAND_325 = {1{`RANDOM}};
  image_469 = _RAND_325[3:0];
  _RAND_326 = {1{`RANDOM}};
  image_470 = _RAND_326[3:0];
  _RAND_327 = {1{`RANDOM}};
  image_471 = _RAND_327[3:0];
  _RAND_328 = {1{`RANDOM}};
  image_472 = _RAND_328[3:0];
  _RAND_329 = {1{`RANDOM}};
  image_473 = _RAND_329[3:0];
  _RAND_330 = {1{`RANDOM}};
  image_474 = _RAND_330[3:0];
  _RAND_331 = {1{`RANDOM}};
  image_475 = _RAND_331[3:0];
  _RAND_332 = {1{`RANDOM}};
  image_476 = _RAND_332[3:0];
  _RAND_333 = {1{`RANDOM}};
  image_477 = _RAND_333[3:0];
  _RAND_334 = {1{`RANDOM}};
  image_478 = _RAND_334[3:0];
  _RAND_335 = {1{`RANDOM}};
  image_479 = _RAND_335[3:0];
  _RAND_336 = {1{`RANDOM}};
  image_480 = _RAND_336[3:0];
  _RAND_337 = {1{`RANDOM}};
  image_481 = _RAND_337[3:0];
  _RAND_338 = {1{`RANDOM}};
  image_482 = _RAND_338[3:0];
  _RAND_339 = {1{`RANDOM}};
  image_483 = _RAND_339[3:0];
  _RAND_340 = {1{`RANDOM}};
  image_484 = _RAND_340[3:0];
  _RAND_341 = {1{`RANDOM}};
  image_485 = _RAND_341[3:0];
  _RAND_342 = {1{`RANDOM}};
  image_486 = _RAND_342[3:0];
  _RAND_343 = {1{`RANDOM}};
  image_487 = _RAND_343[3:0];
  _RAND_344 = {1{`RANDOM}};
  image_488 = _RAND_344[3:0];
  _RAND_345 = {1{`RANDOM}};
  image_489 = _RAND_345[3:0];
  _RAND_346 = {1{`RANDOM}};
  image_490 = _RAND_346[3:0];
  _RAND_347 = {1{`RANDOM}};
  image_491 = _RAND_347[3:0];
  _RAND_348 = {1{`RANDOM}};
  image_492 = _RAND_348[3:0];
  _RAND_349 = {1{`RANDOM}};
  image_493 = _RAND_349[3:0];
  _RAND_350 = {1{`RANDOM}};
  image_494 = _RAND_350[3:0];
  _RAND_351 = {1{`RANDOM}};
  image_495 = _RAND_351[3:0];
  _RAND_352 = {1{`RANDOM}};
  image_496 = _RAND_352[3:0];
  _RAND_353 = {1{`RANDOM}};
  image_497 = _RAND_353[3:0];
  _RAND_354 = {1{`RANDOM}};
  image_498 = _RAND_354[3:0];
  _RAND_355 = {1{`RANDOM}};
  image_499 = _RAND_355[3:0];
  _RAND_356 = {1{`RANDOM}};
  image_500 = _RAND_356[3:0];
  _RAND_357 = {1{`RANDOM}};
  image_501 = _RAND_357[3:0];
  _RAND_358 = {1{`RANDOM}};
  image_502 = _RAND_358[3:0];
  _RAND_359 = {1{`RANDOM}};
  image_503 = _RAND_359[3:0];
  _RAND_360 = {1{`RANDOM}};
  image_504 = _RAND_360[3:0];
  _RAND_361 = {1{`RANDOM}};
  image_505 = _RAND_361[3:0];
  _RAND_362 = {1{`RANDOM}};
  image_506 = _RAND_362[3:0];
  _RAND_363 = {1{`RANDOM}};
  image_507 = _RAND_363[3:0];
  _RAND_364 = {1{`RANDOM}};
  image_508 = _RAND_364[3:0];
  _RAND_365 = {1{`RANDOM}};
  image_509 = _RAND_365[3:0];
  _RAND_366 = {1{`RANDOM}};
  image_515 = _RAND_366[3:0];
  _RAND_367 = {1{`RANDOM}};
  image_516 = _RAND_367[3:0];
  _RAND_368 = {1{`RANDOM}};
  image_517 = _RAND_368[3:0];
  _RAND_369 = {1{`RANDOM}};
  image_518 = _RAND_369[3:0];
  _RAND_370 = {1{`RANDOM}};
  image_519 = _RAND_370[3:0];
  _RAND_371 = {1{`RANDOM}};
  image_520 = _RAND_371[3:0];
  _RAND_372 = {1{`RANDOM}};
  image_521 = _RAND_372[3:0];
  _RAND_373 = {1{`RANDOM}};
  image_522 = _RAND_373[3:0];
  _RAND_374 = {1{`RANDOM}};
  image_523 = _RAND_374[3:0];
  _RAND_375 = {1{`RANDOM}};
  image_524 = _RAND_375[3:0];
  _RAND_376 = {1{`RANDOM}};
  image_525 = _RAND_376[3:0];
  _RAND_377 = {1{`RANDOM}};
  image_526 = _RAND_377[3:0];
  _RAND_378 = {1{`RANDOM}};
  image_527 = _RAND_378[3:0];
  _RAND_379 = {1{`RANDOM}};
  image_528 = _RAND_379[3:0];
  _RAND_380 = {1{`RANDOM}};
  image_529 = _RAND_380[3:0];
  _RAND_381 = {1{`RANDOM}};
  image_530 = _RAND_381[3:0];
  _RAND_382 = {1{`RANDOM}};
  image_531 = _RAND_382[3:0];
  _RAND_383 = {1{`RANDOM}};
  image_532 = _RAND_383[3:0];
  _RAND_384 = {1{`RANDOM}};
  image_533 = _RAND_384[3:0];
  _RAND_385 = {1{`RANDOM}};
  image_534 = _RAND_385[3:0];
  _RAND_386 = {1{`RANDOM}};
  image_535 = _RAND_386[3:0];
  _RAND_387 = {1{`RANDOM}};
  image_536 = _RAND_387[3:0];
  _RAND_388 = {1{`RANDOM}};
  image_537 = _RAND_388[3:0];
  _RAND_389 = {1{`RANDOM}};
  image_538 = _RAND_389[3:0];
  _RAND_390 = {1{`RANDOM}};
  image_539 = _RAND_390[3:0];
  _RAND_391 = {1{`RANDOM}};
  image_540 = _RAND_391[3:0];
  _RAND_392 = {1{`RANDOM}};
  image_541 = _RAND_392[3:0];
  _RAND_393 = {1{`RANDOM}};
  image_542 = _RAND_393[3:0];
  _RAND_394 = {1{`RANDOM}};
  image_543 = _RAND_394[3:0];
  _RAND_395 = {1{`RANDOM}};
  image_544 = _RAND_395[3:0];
  _RAND_396 = {1{`RANDOM}};
  image_545 = _RAND_396[3:0];
  _RAND_397 = {1{`RANDOM}};
  image_546 = _RAND_397[3:0];
  _RAND_398 = {1{`RANDOM}};
  image_547 = _RAND_398[3:0];
  _RAND_399 = {1{`RANDOM}};
  image_548 = _RAND_399[3:0];
  _RAND_400 = {1{`RANDOM}};
  image_549 = _RAND_400[3:0];
  _RAND_401 = {1{`RANDOM}};
  image_550 = _RAND_401[3:0];
  _RAND_402 = {1{`RANDOM}};
  image_551 = _RAND_402[3:0];
  _RAND_403 = {1{`RANDOM}};
  image_552 = _RAND_403[3:0];
  _RAND_404 = {1{`RANDOM}};
  image_553 = _RAND_404[3:0];
  _RAND_405 = {1{`RANDOM}};
  image_554 = _RAND_405[3:0];
  _RAND_406 = {1{`RANDOM}};
  image_555 = _RAND_406[3:0];
  _RAND_407 = {1{`RANDOM}};
  image_556 = _RAND_407[3:0];
  _RAND_408 = {1{`RANDOM}};
  image_557 = _RAND_408[3:0];
  _RAND_409 = {1{`RANDOM}};
  image_558 = _RAND_409[3:0];
  _RAND_410 = {1{`RANDOM}};
  image_559 = _RAND_410[3:0];
  _RAND_411 = {1{`RANDOM}};
  image_560 = _RAND_411[3:0];
  _RAND_412 = {1{`RANDOM}};
  image_561 = _RAND_412[3:0];
  _RAND_413 = {1{`RANDOM}};
  image_562 = _RAND_413[3:0];
  _RAND_414 = {1{`RANDOM}};
  image_563 = _RAND_414[3:0];
  _RAND_415 = {1{`RANDOM}};
  image_564 = _RAND_415[3:0];
  _RAND_416 = {1{`RANDOM}};
  image_565 = _RAND_416[3:0];
  _RAND_417 = {1{`RANDOM}};
  image_566 = _RAND_417[3:0];
  _RAND_418 = {1{`RANDOM}};
  image_571 = _RAND_418[3:0];
  _RAND_419 = {1{`RANDOM}};
  image_572 = _RAND_419[3:0];
  _RAND_420 = {1{`RANDOM}};
  image_573 = _RAND_420[3:0];
  _RAND_421 = {1{`RANDOM}};
  image_574 = _RAND_421[3:0];
  _RAND_422 = {1{`RANDOM}};
  image_578 = _RAND_422[3:0];
  _RAND_423 = {1{`RANDOM}};
  image_579 = _RAND_423[3:0];
  _RAND_424 = {1{`RANDOM}};
  image_580 = _RAND_424[3:0];
  _RAND_425 = {1{`RANDOM}};
  image_581 = _RAND_425[3:0];
  _RAND_426 = {1{`RANDOM}};
  image_582 = _RAND_426[3:0];
  _RAND_427 = {1{`RANDOM}};
  image_583 = _RAND_427[3:0];
  _RAND_428 = {1{`RANDOM}};
  image_584 = _RAND_428[3:0];
  _RAND_429 = {1{`RANDOM}};
  image_585 = _RAND_429[3:0];
  _RAND_430 = {1{`RANDOM}};
  image_586 = _RAND_430[3:0];
  _RAND_431 = {1{`RANDOM}};
  image_587 = _RAND_431[3:0];
  _RAND_432 = {1{`RANDOM}};
  image_588 = _RAND_432[3:0];
  _RAND_433 = {1{`RANDOM}};
  image_589 = _RAND_433[3:0];
  _RAND_434 = {1{`RANDOM}};
  image_590 = _RAND_434[3:0];
  _RAND_435 = {1{`RANDOM}};
  image_591 = _RAND_435[3:0];
  _RAND_436 = {1{`RANDOM}};
  image_592 = _RAND_436[3:0];
  _RAND_437 = {1{`RANDOM}};
  image_593 = _RAND_437[3:0];
  _RAND_438 = {1{`RANDOM}};
  image_594 = _RAND_438[3:0];
  _RAND_439 = {1{`RANDOM}};
  image_595 = _RAND_439[3:0];
  _RAND_440 = {1{`RANDOM}};
  image_596 = _RAND_440[3:0];
  _RAND_441 = {1{`RANDOM}};
  image_597 = _RAND_441[3:0];
  _RAND_442 = {1{`RANDOM}};
  image_598 = _RAND_442[3:0];
  _RAND_443 = {1{`RANDOM}};
  image_599 = _RAND_443[3:0];
  _RAND_444 = {1{`RANDOM}};
  image_600 = _RAND_444[3:0];
  _RAND_445 = {1{`RANDOM}};
  image_601 = _RAND_445[3:0];
  _RAND_446 = {1{`RANDOM}};
  image_602 = _RAND_446[3:0];
  _RAND_447 = {1{`RANDOM}};
  image_603 = _RAND_447[3:0];
  _RAND_448 = {1{`RANDOM}};
  image_604 = _RAND_448[3:0];
  _RAND_449 = {1{`RANDOM}};
  image_605 = _RAND_449[3:0];
  _RAND_450 = {1{`RANDOM}};
  image_606 = _RAND_450[3:0];
  _RAND_451 = {1{`RANDOM}};
  image_607 = _RAND_451[3:0];
  _RAND_452 = {1{`RANDOM}};
  image_614 = _RAND_452[3:0];
  _RAND_453 = {1{`RANDOM}};
  image_615 = _RAND_453[3:0];
  _RAND_454 = {1{`RANDOM}};
  image_616 = _RAND_454[3:0];
  _RAND_455 = {1{`RANDOM}};
  image_617 = _RAND_455[3:0];
  _RAND_456 = {1{`RANDOM}};
  image_618 = _RAND_456[3:0];
  _RAND_457 = {1{`RANDOM}};
  image_619 = _RAND_457[3:0];
  _RAND_458 = {1{`RANDOM}};
  image_620 = _RAND_458[3:0];
  _RAND_459 = {1{`RANDOM}};
  image_621 = _RAND_459[3:0];
  _RAND_460 = {1{`RANDOM}};
  image_622 = _RAND_460[3:0];
  _RAND_461 = {1{`RANDOM}};
  image_623 = _RAND_461[3:0];
  _RAND_462 = {1{`RANDOM}};
  image_624 = _RAND_462[3:0];
  _RAND_463 = {1{`RANDOM}};
  image_625 = _RAND_463[3:0];
  _RAND_464 = {1{`RANDOM}};
  image_626 = _RAND_464[3:0];
  _RAND_465 = {1{`RANDOM}};
  image_627 = _RAND_465[3:0];
  _RAND_466 = {1{`RANDOM}};
  image_628 = _RAND_466[3:0];
  _RAND_467 = {1{`RANDOM}};
  image_636 = _RAND_467[3:0];
  _RAND_468 = {1{`RANDOM}};
  image_637 = _RAND_468[3:0];
  _RAND_469 = {1{`RANDOM}};
  image_638 = _RAND_469[3:0];
  _RAND_470 = {1{`RANDOM}};
  image_639 = _RAND_470[3:0];
  _RAND_471 = {1{`RANDOM}};
  image_642 = _RAND_471[3:0];
  _RAND_472 = {1{`RANDOM}};
  image_643 = _RAND_472[3:0];
  _RAND_473 = {1{`RANDOM}};
  image_644 = _RAND_473[3:0];
  _RAND_474 = {1{`RANDOM}};
  image_645 = _RAND_474[3:0];
  _RAND_475 = {1{`RANDOM}};
  image_646 = _RAND_475[3:0];
  _RAND_476 = {1{`RANDOM}};
  image_647 = _RAND_476[3:0];
  _RAND_477 = {1{`RANDOM}};
  image_648 = _RAND_477[3:0];
  _RAND_478 = {1{`RANDOM}};
  image_649 = _RAND_478[3:0];
  _RAND_479 = {1{`RANDOM}};
  image_650 = _RAND_479[3:0];
  _RAND_480 = {1{`RANDOM}};
  image_651 = _RAND_480[3:0];
  _RAND_481 = {1{`RANDOM}};
  image_652 = _RAND_481[3:0];
  _RAND_482 = {1{`RANDOM}};
  image_653 = _RAND_482[3:0];
  _RAND_483 = {1{`RANDOM}};
  image_654 = _RAND_483[3:0];
  _RAND_484 = {1{`RANDOM}};
  image_655 = _RAND_484[3:0];
  _RAND_485 = {1{`RANDOM}};
  image_656 = _RAND_485[3:0];
  _RAND_486 = {1{`RANDOM}};
  image_657 = _RAND_486[3:0];
  _RAND_487 = {1{`RANDOM}};
  image_658 = _RAND_487[3:0];
  _RAND_488 = {1{`RANDOM}};
  image_659 = _RAND_488[3:0];
  _RAND_489 = {1{`RANDOM}};
  image_660 = _RAND_489[3:0];
  _RAND_490 = {1{`RANDOM}};
  image_661 = _RAND_490[3:0];
  _RAND_491 = {1{`RANDOM}};
  image_662 = _RAND_491[3:0];
  _RAND_492 = {1{`RANDOM}};
  image_663 = _RAND_492[3:0];
  _RAND_493 = {1{`RANDOM}};
  image_664 = _RAND_493[3:0];
  _RAND_494 = {1{`RANDOM}};
  image_665 = _RAND_494[3:0];
  _RAND_495 = {1{`RANDOM}};
  image_666 = _RAND_495[3:0];
  _RAND_496 = {1{`RANDOM}};
  image_667 = _RAND_496[3:0];
  _RAND_497 = {1{`RANDOM}};
  image_668 = _RAND_497[3:0];
  _RAND_498 = {1{`RANDOM}};
  image_669 = _RAND_498[3:0];
  _RAND_499 = {1{`RANDOM}};
  image_670 = _RAND_499[3:0];
  _RAND_500 = {1{`RANDOM}};
  image_679 = _RAND_500[3:0];
  _RAND_501 = {1{`RANDOM}};
  image_680 = _RAND_501[3:0];
  _RAND_502 = {1{`RANDOM}};
  image_681 = _RAND_502[3:0];
  _RAND_503 = {1{`RANDOM}};
  image_682 = _RAND_503[3:0];
  _RAND_504 = {1{`RANDOM}};
  image_683 = _RAND_504[3:0];
  _RAND_505 = {1{`RANDOM}};
  image_684 = _RAND_505[3:0];
  _RAND_506 = {1{`RANDOM}};
  image_685 = _RAND_506[3:0];
  _RAND_507 = {1{`RANDOM}};
  image_686 = _RAND_507[3:0];
  _RAND_508 = {1{`RANDOM}};
  image_687 = _RAND_508[3:0];
  _RAND_509 = {1{`RANDOM}};
  image_688 = _RAND_509[3:0];
  _RAND_510 = {1{`RANDOM}};
  image_689 = _RAND_510[3:0];
  _RAND_511 = {1{`RANDOM}};
  image_690 = _RAND_511[3:0];
  _RAND_512 = {1{`RANDOM}};
  image_691 = _RAND_512[3:0];
  _RAND_513 = {1{`RANDOM}};
  image_692 = _RAND_513[3:0];
  _RAND_514 = {1{`RANDOM}};
  image_693 = _RAND_514[3:0];
  _RAND_515 = {1{`RANDOM}};
  image_694 = _RAND_515[3:0];
  _RAND_516 = {1{`RANDOM}};
  image_695 = _RAND_516[3:0];
  _RAND_517 = {1{`RANDOM}};
  image_696 = _RAND_517[3:0];
  _RAND_518 = {1{`RANDOM}};
  image_697 = _RAND_518[3:0];
  _RAND_519 = {1{`RANDOM}};
  image_698 = _RAND_519[3:0];
  _RAND_520 = {1{`RANDOM}};
  image_701 = _RAND_520[3:0];
  _RAND_521 = {1{`RANDOM}};
  image_702 = _RAND_521[3:0];
  _RAND_522 = {1{`RANDOM}};
  image_703 = _RAND_522[3:0];
  _RAND_523 = {1{`RANDOM}};
  image_705 = _RAND_523[3:0];
  _RAND_524 = {1{`RANDOM}};
  image_706 = _RAND_524[3:0];
  _RAND_525 = {1{`RANDOM}};
  image_707 = _RAND_525[3:0];
  _RAND_526 = {1{`RANDOM}};
  image_708 = _RAND_526[3:0];
  _RAND_527 = {1{`RANDOM}};
  image_709 = _RAND_527[3:0];
  _RAND_528 = {1{`RANDOM}};
  image_710 = _RAND_528[3:0];
  _RAND_529 = {1{`RANDOM}};
  image_711 = _RAND_529[3:0];
  _RAND_530 = {1{`RANDOM}};
  image_712 = _RAND_530[3:0];
  _RAND_531 = {1{`RANDOM}};
  image_713 = _RAND_531[3:0];
  _RAND_532 = {1{`RANDOM}};
  image_714 = _RAND_532[3:0];
  _RAND_533 = {1{`RANDOM}};
  image_715 = _RAND_533[3:0];
  _RAND_534 = {1{`RANDOM}};
  image_716 = _RAND_534[3:0];
  _RAND_535 = {1{`RANDOM}};
  image_717 = _RAND_535[3:0];
  _RAND_536 = {1{`RANDOM}};
  image_718 = _RAND_536[3:0];
  _RAND_537 = {1{`RANDOM}};
  image_719 = _RAND_537[3:0];
  _RAND_538 = {1{`RANDOM}};
  image_720 = _RAND_538[3:0];
  _RAND_539 = {1{`RANDOM}};
  image_721 = _RAND_539[3:0];
  _RAND_540 = {1{`RANDOM}};
  image_722 = _RAND_540[3:0];
  _RAND_541 = {1{`RANDOM}};
  image_723 = _RAND_541[3:0];
  _RAND_542 = {1{`RANDOM}};
  image_724 = _RAND_542[3:0];
  _RAND_543 = {1{`RANDOM}};
  image_725 = _RAND_543[3:0];
  _RAND_544 = {1{`RANDOM}};
  image_726 = _RAND_544[3:0];
  _RAND_545 = {1{`RANDOM}};
  image_727 = _RAND_545[3:0];
  _RAND_546 = {1{`RANDOM}};
  image_728 = _RAND_546[3:0];
  _RAND_547 = {1{`RANDOM}};
  image_729 = _RAND_547[3:0];
  _RAND_548 = {1{`RANDOM}};
  image_730 = _RAND_548[3:0];
  _RAND_549 = {1{`RANDOM}};
  image_731 = _RAND_549[3:0];
  _RAND_550 = {1{`RANDOM}};
  image_732 = _RAND_550[3:0];
  _RAND_551 = {1{`RANDOM}};
  image_733 = _RAND_551[3:0];
  _RAND_552 = {1{`RANDOM}};
  image_734 = _RAND_552[3:0];
  _RAND_553 = {1{`RANDOM}};
  image_736 = _RAND_553[3:0];
  _RAND_554 = {1{`RANDOM}};
  image_737 = _RAND_554[3:0];
  _RAND_555 = {1{`RANDOM}};
  image_739 = _RAND_555[3:0];
  _RAND_556 = {1{`RANDOM}};
  image_740 = _RAND_556[3:0];
  _RAND_557 = {1{`RANDOM}};
  image_741 = _RAND_557[3:0];
  _RAND_558 = {1{`RANDOM}};
  image_744 = _RAND_558[3:0];
  _RAND_559 = {1{`RANDOM}};
  image_745 = _RAND_559[3:0];
  _RAND_560 = {1{`RANDOM}};
  image_746 = _RAND_560[3:0];
  _RAND_561 = {1{`RANDOM}};
  image_747 = _RAND_561[3:0];
  _RAND_562 = {1{`RANDOM}};
  image_748 = _RAND_562[3:0];
  _RAND_563 = {1{`RANDOM}};
  image_749 = _RAND_563[3:0];
  _RAND_564 = {1{`RANDOM}};
  image_750 = _RAND_564[3:0];
  _RAND_565 = {1{`RANDOM}};
  image_751 = _RAND_565[3:0];
  _RAND_566 = {1{`RANDOM}};
  image_752 = _RAND_566[3:0];
  _RAND_567 = {1{`RANDOM}};
  image_753 = _RAND_567[3:0];
  _RAND_568 = {1{`RANDOM}};
  image_754 = _RAND_568[3:0];
  _RAND_569 = {1{`RANDOM}};
  image_755 = _RAND_569[3:0];
  _RAND_570 = {1{`RANDOM}};
  image_756 = _RAND_570[3:0];
  _RAND_571 = {1{`RANDOM}};
  image_758 = _RAND_571[3:0];
  _RAND_572 = {1{`RANDOM}};
  image_760 = _RAND_572[3:0];
  _RAND_573 = {1{`RANDOM}};
  image_761 = _RAND_573[3:0];
  _RAND_574 = {1{`RANDOM}};
  image_762 = _RAND_574[3:0];
  _RAND_575 = {1{`RANDOM}};
  image_763 = _RAND_575[3:0];
  _RAND_576 = {1{`RANDOM}};
  image_765 = _RAND_576[3:0];
  _RAND_577 = {1{`RANDOM}};
  image_766 = _RAND_577[3:0];
  _RAND_578 = {1{`RANDOM}};
  image_767 = _RAND_578[3:0];
  _RAND_579 = {1{`RANDOM}};
  image_768 = _RAND_579[3:0];
  _RAND_580 = {1{`RANDOM}};
  image_769 = _RAND_580[3:0];
  _RAND_581 = {1{`RANDOM}};
  image_770 = _RAND_581[3:0];
  _RAND_582 = {1{`RANDOM}};
  image_771 = _RAND_582[3:0];
  _RAND_583 = {1{`RANDOM}};
  image_772 = _RAND_583[3:0];
  _RAND_584 = {1{`RANDOM}};
  image_773 = _RAND_584[3:0];
  _RAND_585 = {1{`RANDOM}};
  image_774 = _RAND_585[3:0];
  _RAND_586 = {1{`RANDOM}};
  image_775 = _RAND_586[3:0];
  _RAND_587 = {1{`RANDOM}};
  image_776 = _RAND_587[3:0];
  _RAND_588 = {1{`RANDOM}};
  image_777 = _RAND_588[3:0];
  _RAND_589 = {1{`RANDOM}};
  image_778 = _RAND_589[3:0];
  _RAND_590 = {1{`RANDOM}};
  image_779 = _RAND_590[3:0];
  _RAND_591 = {1{`RANDOM}};
  image_780 = _RAND_591[3:0];
  _RAND_592 = {1{`RANDOM}};
  image_781 = _RAND_592[3:0];
  _RAND_593 = {1{`RANDOM}};
  image_782 = _RAND_593[3:0];
  _RAND_594 = {1{`RANDOM}};
  image_783 = _RAND_594[3:0];
  _RAND_595 = {1{`RANDOM}};
  image_784 = _RAND_595[3:0];
  _RAND_596 = {1{`RANDOM}};
  image_785 = _RAND_596[3:0];
  _RAND_597 = {1{`RANDOM}};
  image_786 = _RAND_597[3:0];
  _RAND_598 = {1{`RANDOM}};
  image_787 = _RAND_598[3:0];
  _RAND_599 = {1{`RANDOM}};
  image_788 = _RAND_599[3:0];
  _RAND_600 = {1{`RANDOM}};
  image_789 = _RAND_600[3:0];
  _RAND_601 = {1{`RANDOM}};
  image_790 = _RAND_601[3:0];
  _RAND_602 = {1{`RANDOM}};
  image_791 = _RAND_602[3:0];
  _RAND_603 = {1{`RANDOM}};
  image_792 = _RAND_603[3:0];
  _RAND_604 = {1{`RANDOM}};
  image_793 = _RAND_604[3:0];
  _RAND_605 = {1{`RANDOM}};
  image_794 = _RAND_605[3:0];
  _RAND_606 = {1{`RANDOM}};
  image_795 = _RAND_606[3:0];
  _RAND_607 = {1{`RANDOM}};
  image_796 = _RAND_607[3:0];
  _RAND_608 = {1{`RANDOM}};
  image_797 = _RAND_608[3:0];
  _RAND_609 = {1{`RANDOM}};
  image_800 = _RAND_609[3:0];
  _RAND_610 = {1{`RANDOM}};
  image_801 = _RAND_610[3:0];
  _RAND_611 = {1{`RANDOM}};
  image_802 = _RAND_611[3:0];
  _RAND_612 = {1{`RANDOM}};
  image_803 = _RAND_612[3:0];
  _RAND_613 = {1{`RANDOM}};
  image_804 = _RAND_613[3:0];
  _RAND_614 = {1{`RANDOM}};
  image_805 = _RAND_614[3:0];
  _RAND_615 = {1{`RANDOM}};
  image_806 = _RAND_615[3:0];
  _RAND_616 = {1{`RANDOM}};
  image_808 = _RAND_616[3:0];
  _RAND_617 = {1{`RANDOM}};
  image_809 = _RAND_617[3:0];
  _RAND_618 = {1{`RANDOM}};
  image_810 = _RAND_618[3:0];
  _RAND_619 = {1{`RANDOM}};
  image_811 = _RAND_619[3:0];
  _RAND_620 = {1{`RANDOM}};
  image_812 = _RAND_620[3:0];
  _RAND_621 = {1{`RANDOM}};
  image_813 = _RAND_621[3:0];
  _RAND_622 = {1{`RANDOM}};
  image_814 = _RAND_622[3:0];
  _RAND_623 = {1{`RANDOM}};
  image_815 = _RAND_623[3:0];
  _RAND_624 = {1{`RANDOM}};
  image_816 = _RAND_624[3:0];
  _RAND_625 = {1{`RANDOM}};
  image_817 = _RAND_625[3:0];
  _RAND_626 = {1{`RANDOM}};
  image_818 = _RAND_626[3:0];
  _RAND_627 = {1{`RANDOM}};
  image_819 = _RAND_627[3:0];
  _RAND_628 = {1{`RANDOM}};
  image_820 = _RAND_628[3:0];
  _RAND_629 = {1{`RANDOM}};
  image_822 = _RAND_629[3:0];
  _RAND_630 = {1{`RANDOM}};
  image_823 = _RAND_630[3:0];
  _RAND_631 = {1{`RANDOM}};
  image_824 = _RAND_631[3:0];
  _RAND_632 = {1{`RANDOM}};
  image_825 = _RAND_632[3:0];
  _RAND_633 = {1{`RANDOM}};
  image_826 = _RAND_633[3:0];
  _RAND_634 = {1{`RANDOM}};
  image_828 = _RAND_634[3:0];
  _RAND_635 = {1{`RANDOM}};
  image_829 = _RAND_635[3:0];
  _RAND_636 = {1{`RANDOM}};
  image_830 = _RAND_636[3:0];
  _RAND_637 = {1{`RANDOM}};
  image_831 = _RAND_637[3:0];
  _RAND_638 = {1{`RANDOM}};
  image_833 = _RAND_638[3:0];
  _RAND_639 = {1{`RANDOM}};
  image_834 = _RAND_639[3:0];
  _RAND_640 = {1{`RANDOM}};
  image_835 = _RAND_640[3:0];
  _RAND_641 = {1{`RANDOM}};
  image_836 = _RAND_641[3:0];
  _RAND_642 = {1{`RANDOM}};
  image_837 = _RAND_642[3:0];
  _RAND_643 = {1{`RANDOM}};
  image_838 = _RAND_643[3:0];
  _RAND_644 = {1{`RANDOM}};
  image_839 = _RAND_644[3:0];
  _RAND_645 = {1{`RANDOM}};
  image_840 = _RAND_645[3:0];
  _RAND_646 = {1{`RANDOM}};
  image_841 = _RAND_646[3:0];
  _RAND_647 = {1{`RANDOM}};
  image_842 = _RAND_647[3:0];
  _RAND_648 = {1{`RANDOM}};
  image_843 = _RAND_648[3:0];
  _RAND_649 = {1{`RANDOM}};
  image_844 = _RAND_649[3:0];
  _RAND_650 = {1{`RANDOM}};
  image_845 = _RAND_650[3:0];
  _RAND_651 = {1{`RANDOM}};
  image_846 = _RAND_651[3:0];
  _RAND_652 = {1{`RANDOM}};
  image_847 = _RAND_652[3:0];
  _RAND_653 = {1{`RANDOM}};
  image_848 = _RAND_653[3:0];
  _RAND_654 = {1{`RANDOM}};
  image_849 = _RAND_654[3:0];
  _RAND_655 = {1{`RANDOM}};
  image_850 = _RAND_655[3:0];
  _RAND_656 = {1{`RANDOM}};
  image_851 = _RAND_656[3:0];
  _RAND_657 = {1{`RANDOM}};
  image_852 = _RAND_657[3:0];
  _RAND_658 = {1{`RANDOM}};
  image_853 = _RAND_658[3:0];
  _RAND_659 = {1{`RANDOM}};
  image_854 = _RAND_659[3:0];
  _RAND_660 = {1{`RANDOM}};
  image_855 = _RAND_660[3:0];
  _RAND_661 = {1{`RANDOM}};
  image_856 = _RAND_661[3:0];
  _RAND_662 = {1{`RANDOM}};
  image_857 = _RAND_662[3:0];
  _RAND_663 = {1{`RANDOM}};
  image_858 = _RAND_663[3:0];
  _RAND_664 = {1{`RANDOM}};
  image_859 = _RAND_664[3:0];
  _RAND_665 = {1{`RANDOM}};
  image_860 = _RAND_665[3:0];
  _RAND_666 = {1{`RANDOM}};
  image_861 = _RAND_666[3:0];
  _RAND_667 = {1{`RANDOM}};
  image_862 = _RAND_667[3:0];
  _RAND_668 = {1{`RANDOM}};
  image_865 = _RAND_668[3:0];
  _RAND_669 = {1{`RANDOM}};
  image_866 = _RAND_669[3:0];
  _RAND_670 = {1{`RANDOM}};
  image_867 = _RAND_670[3:0];
  _RAND_671 = {1{`RANDOM}};
  image_868 = _RAND_671[3:0];
  _RAND_672 = {1{`RANDOM}};
  image_869 = _RAND_672[3:0];
  _RAND_673 = {1{`RANDOM}};
  image_872 = _RAND_673[3:0];
  _RAND_674 = {1{`RANDOM}};
  image_873 = _RAND_674[3:0];
  _RAND_675 = {1{`RANDOM}};
  image_874 = _RAND_675[3:0];
  _RAND_676 = {1{`RANDOM}};
  image_875 = _RAND_676[3:0];
  _RAND_677 = {1{`RANDOM}};
  image_876 = _RAND_677[3:0];
  _RAND_678 = {1{`RANDOM}};
  image_877 = _RAND_678[3:0];
  _RAND_679 = {1{`RANDOM}};
  image_878 = _RAND_679[3:0];
  _RAND_680 = {1{`RANDOM}};
  image_879 = _RAND_680[3:0];
  _RAND_681 = {1{`RANDOM}};
  image_880 = _RAND_681[3:0];
  _RAND_682 = {1{`RANDOM}};
  image_881 = _RAND_682[3:0];
  _RAND_683 = {1{`RANDOM}};
  image_882 = _RAND_683[3:0];
  _RAND_684 = {1{`RANDOM}};
  image_883 = _RAND_684[3:0];
  _RAND_685 = {1{`RANDOM}};
  image_884 = _RAND_685[3:0];
  _RAND_686 = {1{`RANDOM}};
  image_885 = _RAND_686[3:0];
  _RAND_687 = {1{`RANDOM}};
  image_891 = _RAND_687[3:0];
  _RAND_688 = {1{`RANDOM}};
  image_892 = _RAND_688[3:0];
  _RAND_689 = {1{`RANDOM}};
  image_893 = _RAND_689[3:0];
  _RAND_690 = {1{`RANDOM}};
  image_894 = _RAND_690[3:0];
  _RAND_691 = {1{`RANDOM}};
  image_895 = _RAND_691[3:0];
  _RAND_692 = {1{`RANDOM}};
  image_897 = _RAND_692[3:0];
  _RAND_693 = {1{`RANDOM}};
  image_898 = _RAND_693[3:0];
  _RAND_694 = {1{`RANDOM}};
  image_899 = _RAND_694[3:0];
  _RAND_695 = {1{`RANDOM}};
  image_900 = _RAND_695[3:0];
  _RAND_696 = {1{`RANDOM}};
  image_901 = _RAND_696[3:0];
  _RAND_697 = {1{`RANDOM}};
  image_902 = _RAND_697[3:0];
  _RAND_698 = {1{`RANDOM}};
  image_903 = _RAND_698[3:0];
  _RAND_699 = {1{`RANDOM}};
  image_904 = _RAND_699[3:0];
  _RAND_700 = {1{`RANDOM}};
  image_905 = _RAND_700[3:0];
  _RAND_701 = {1{`RANDOM}};
  image_906 = _RAND_701[3:0];
  _RAND_702 = {1{`RANDOM}};
  image_907 = _RAND_702[3:0];
  _RAND_703 = {1{`RANDOM}};
  image_908 = _RAND_703[3:0];
  _RAND_704 = {1{`RANDOM}};
  image_909 = _RAND_704[3:0];
  _RAND_705 = {1{`RANDOM}};
  image_910 = _RAND_705[3:0];
  _RAND_706 = {1{`RANDOM}};
  image_911 = _RAND_706[3:0];
  _RAND_707 = {1{`RANDOM}};
  image_912 = _RAND_707[3:0];
  _RAND_708 = {1{`RANDOM}};
  image_913 = _RAND_708[3:0];
  _RAND_709 = {1{`RANDOM}};
  image_914 = _RAND_709[3:0];
  _RAND_710 = {1{`RANDOM}};
  image_915 = _RAND_710[3:0];
  _RAND_711 = {1{`RANDOM}};
  image_916 = _RAND_711[3:0];
  _RAND_712 = {1{`RANDOM}};
  image_917 = _RAND_712[3:0];
  _RAND_713 = {1{`RANDOM}};
  image_918 = _RAND_713[3:0];
  _RAND_714 = {1{`RANDOM}};
  image_919 = _RAND_714[3:0];
  _RAND_715 = {1{`RANDOM}};
  image_920 = _RAND_715[3:0];
  _RAND_716 = {1{`RANDOM}};
  image_921 = _RAND_716[3:0];
  _RAND_717 = {1{`RANDOM}};
  image_922 = _RAND_717[3:0];
  _RAND_718 = {1{`RANDOM}};
  image_923 = _RAND_718[3:0];
  _RAND_719 = {1{`RANDOM}};
  image_924 = _RAND_719[3:0];
  _RAND_720 = {1{`RANDOM}};
  image_925 = _RAND_720[3:0];
  _RAND_721 = {1{`RANDOM}};
  image_926 = _RAND_721[3:0];
  _RAND_722 = {1{`RANDOM}};
  image_927 = _RAND_722[3:0];
  _RAND_723 = {1{`RANDOM}};
  image_929 = _RAND_723[3:0];
  _RAND_724 = {1{`RANDOM}};
  image_930 = _RAND_724[3:0];
  _RAND_725 = {1{`RANDOM}};
  image_935 = _RAND_725[3:0];
  _RAND_726 = {1{`RANDOM}};
  image_936 = _RAND_726[3:0];
  _RAND_727 = {1{`RANDOM}};
  image_937 = _RAND_727[3:0];
  _RAND_728 = {1{`RANDOM}};
  image_938 = _RAND_728[3:0];
  _RAND_729 = {1{`RANDOM}};
  image_939 = _RAND_729[3:0];
  _RAND_730 = {1{`RANDOM}};
  image_940 = _RAND_730[3:0];
  _RAND_731 = {1{`RANDOM}};
  image_941 = _RAND_731[3:0];
  _RAND_732 = {1{`RANDOM}};
  image_942 = _RAND_732[3:0];
  _RAND_733 = {1{`RANDOM}};
  image_943 = _RAND_733[3:0];
  _RAND_734 = {1{`RANDOM}};
  image_944 = _RAND_734[3:0];
  _RAND_735 = {1{`RANDOM}};
  image_945 = _RAND_735[3:0];
  _RAND_736 = {1{`RANDOM}};
  image_946 = _RAND_736[3:0];
  _RAND_737 = {1{`RANDOM}};
  image_947 = _RAND_737[3:0];
  _RAND_738 = {1{`RANDOM}};
  image_948 = _RAND_738[3:0];
  _RAND_739 = {1{`RANDOM}};
  image_949 = _RAND_739[3:0];
  _RAND_740 = {1{`RANDOM}};
  image_950 = _RAND_740[3:0];
  _RAND_741 = {1{`RANDOM}};
  image_951 = _RAND_741[3:0];
  _RAND_742 = {1{`RANDOM}};
  image_952 = _RAND_742[3:0];
  _RAND_743 = {1{`RANDOM}};
  image_953 = _RAND_743[3:0];
  _RAND_744 = {1{`RANDOM}};
  image_954 = _RAND_744[3:0];
  _RAND_745 = {1{`RANDOM}};
  image_955 = _RAND_745[3:0];
  _RAND_746 = {1{`RANDOM}};
  image_956 = _RAND_746[3:0];
  _RAND_747 = {1{`RANDOM}};
  image_957 = _RAND_747[3:0];
  _RAND_748 = {1{`RANDOM}};
  image_958 = _RAND_748[3:0];
  _RAND_749 = {1{`RANDOM}};
  image_959 = _RAND_749[3:0];
  _RAND_750 = {1{`RANDOM}};
  image_961 = _RAND_750[3:0];
  _RAND_751 = {1{`RANDOM}};
  image_962 = _RAND_751[3:0];
  _RAND_752 = {1{`RANDOM}};
  image_963 = _RAND_752[3:0];
  _RAND_753 = {1{`RANDOM}};
  image_964 = _RAND_753[3:0];
  _RAND_754 = {1{`RANDOM}};
  image_965 = _RAND_754[3:0];
  _RAND_755 = {1{`RANDOM}};
  image_966 = _RAND_755[3:0];
  _RAND_756 = {1{`RANDOM}};
  image_967 = _RAND_756[3:0];
  _RAND_757 = {1{`RANDOM}};
  image_968 = _RAND_757[3:0];
  _RAND_758 = {1{`RANDOM}};
  image_969 = _RAND_758[3:0];
  _RAND_759 = {1{`RANDOM}};
  image_970 = _RAND_759[3:0];
  _RAND_760 = {1{`RANDOM}};
  image_971 = _RAND_760[3:0];
  _RAND_761 = {1{`RANDOM}};
  image_972 = _RAND_761[3:0];
  _RAND_762 = {1{`RANDOM}};
  image_973 = _RAND_762[3:0];
  _RAND_763 = {1{`RANDOM}};
  image_974 = _RAND_763[3:0];
  _RAND_764 = {1{`RANDOM}};
  image_975 = _RAND_764[3:0];
  _RAND_765 = {1{`RANDOM}};
  image_976 = _RAND_765[3:0];
  _RAND_766 = {1{`RANDOM}};
  image_977 = _RAND_766[3:0];
  _RAND_767 = {1{`RANDOM}};
  image_978 = _RAND_767[3:0];
  _RAND_768 = {1{`RANDOM}};
  image_979 = _RAND_768[3:0];
  _RAND_769 = {1{`RANDOM}};
  image_980 = _RAND_769[3:0];
  _RAND_770 = {1{`RANDOM}};
  image_981 = _RAND_770[3:0];
  _RAND_771 = {1{`RANDOM}};
  image_982 = _RAND_771[3:0];
  _RAND_772 = {1{`RANDOM}};
  image_983 = _RAND_772[3:0];
  _RAND_773 = {1{`RANDOM}};
  image_984 = _RAND_773[3:0];
  _RAND_774 = {1{`RANDOM}};
  image_985 = _RAND_774[3:0];
  _RAND_775 = {1{`RANDOM}};
  image_986 = _RAND_775[3:0];
  _RAND_776 = {1{`RANDOM}};
  image_987 = _RAND_776[3:0];
  _RAND_777 = {1{`RANDOM}};
  image_988 = _RAND_777[3:0];
  _RAND_778 = {1{`RANDOM}};
  image_989 = _RAND_778[3:0];
  _RAND_779 = {1{`RANDOM}};
  image_990 = _RAND_779[3:0];
  _RAND_780 = {1{`RANDOM}};
  image_991 = _RAND_780[3:0];
  _RAND_781 = {1{`RANDOM}};
  image_992 = _RAND_781[3:0];
  _RAND_782 = {1{`RANDOM}};
  image_997 = _RAND_782[3:0];
  _RAND_783 = {1{`RANDOM}};
  image_998 = _RAND_783[3:0];
  _RAND_784 = {1{`RANDOM}};
  image_999 = _RAND_784[3:0];
  _RAND_785 = {1{`RANDOM}};
  image_1000 = _RAND_785[3:0];
  _RAND_786 = {1{`RANDOM}};
  image_1001 = _RAND_786[3:0];
  _RAND_787 = {1{`RANDOM}};
  image_1002 = _RAND_787[3:0];
  _RAND_788 = {1{`RANDOM}};
  image_1003 = _RAND_788[3:0];
  _RAND_789 = {1{`RANDOM}};
  image_1004 = _RAND_789[3:0];
  _RAND_790 = {1{`RANDOM}};
  image_1005 = _RAND_790[3:0];
  _RAND_791 = {1{`RANDOM}};
  image_1006 = _RAND_791[3:0];
  _RAND_792 = {1{`RANDOM}};
  image_1007 = _RAND_792[3:0];
  _RAND_793 = {1{`RANDOM}};
  image_1008 = _RAND_793[3:0];
  _RAND_794 = {1{`RANDOM}};
  image_1009 = _RAND_794[3:0];
  _RAND_795 = {1{`RANDOM}};
  image_1010 = _RAND_795[3:0];
  _RAND_796 = {1{`RANDOM}};
  image_1011 = _RAND_796[3:0];
  _RAND_797 = {1{`RANDOM}};
  image_1012 = _RAND_797[3:0];
  _RAND_798 = {1{`RANDOM}};
  image_1013 = _RAND_798[3:0];
  _RAND_799 = {1{`RANDOM}};
  image_1014 = _RAND_799[3:0];
  _RAND_800 = {1{`RANDOM}};
  image_1015 = _RAND_800[3:0];
  _RAND_801 = {1{`RANDOM}};
  image_1016 = _RAND_801[3:0];
  _RAND_802 = {1{`RANDOM}};
  image_1017 = _RAND_802[3:0];
  _RAND_803 = {1{`RANDOM}};
  image_1018 = _RAND_803[3:0];
  _RAND_804 = {1{`RANDOM}};
  image_1019 = _RAND_804[3:0];
  _RAND_805 = {1{`RANDOM}};
  image_1020 = _RAND_805[3:0];
  _RAND_806 = {1{`RANDOM}};
  image_1024 = _RAND_806[3:0];
  _RAND_807 = {1{`RANDOM}};
  image_1025 = _RAND_807[3:0];
  _RAND_808 = {1{`RANDOM}};
  image_1026 = _RAND_808[3:0];
  _RAND_809 = {1{`RANDOM}};
  image_1027 = _RAND_809[3:0];
  _RAND_810 = {1{`RANDOM}};
  image_1028 = _RAND_810[3:0];
  _RAND_811 = {1{`RANDOM}};
  image_1029 = _RAND_811[3:0];
  _RAND_812 = {1{`RANDOM}};
  image_1030 = _RAND_812[3:0];
  _RAND_813 = {1{`RANDOM}};
  image_1031 = _RAND_813[3:0];
  _RAND_814 = {1{`RANDOM}};
  image_1032 = _RAND_814[3:0];
  _RAND_815 = {1{`RANDOM}};
  image_1033 = _RAND_815[3:0];
  _RAND_816 = {1{`RANDOM}};
  image_1034 = _RAND_816[3:0];
  _RAND_817 = {1{`RANDOM}};
  image_1035 = _RAND_817[3:0];
  _RAND_818 = {1{`RANDOM}};
  image_1036 = _RAND_818[3:0];
  _RAND_819 = {1{`RANDOM}};
  image_1037 = _RAND_819[3:0];
  _RAND_820 = {1{`RANDOM}};
  image_1038 = _RAND_820[3:0];
  _RAND_821 = {1{`RANDOM}};
  image_1039 = _RAND_821[3:0];
  _RAND_822 = {1{`RANDOM}};
  image_1040 = _RAND_822[3:0];
  _RAND_823 = {1{`RANDOM}};
  image_1041 = _RAND_823[3:0];
  _RAND_824 = {1{`RANDOM}};
  image_1042 = _RAND_824[3:0];
  _RAND_825 = {1{`RANDOM}};
  image_1043 = _RAND_825[3:0];
  _RAND_826 = {1{`RANDOM}};
  image_1044 = _RAND_826[3:0];
  _RAND_827 = {1{`RANDOM}};
  image_1045 = _RAND_827[3:0];
  _RAND_828 = {1{`RANDOM}};
  image_1046 = _RAND_828[3:0];
  _RAND_829 = {1{`RANDOM}};
  image_1047 = _RAND_829[3:0];
  _RAND_830 = {1{`RANDOM}};
  image_1048 = _RAND_830[3:0];
  _RAND_831 = {1{`RANDOM}};
  image_1049 = _RAND_831[3:0];
  _RAND_832 = {1{`RANDOM}};
  image_1050 = _RAND_832[3:0];
  _RAND_833 = {1{`RANDOM}};
  image_1051 = _RAND_833[3:0];
  _RAND_834 = {1{`RANDOM}};
  image_1052 = _RAND_834[3:0];
  _RAND_835 = {1{`RANDOM}};
  image_1053 = _RAND_835[3:0];
  _RAND_836 = {1{`RANDOM}};
  image_1054 = _RAND_836[3:0];
  _RAND_837 = {1{`RANDOM}};
  image_1055 = _RAND_837[3:0];
  _RAND_838 = {1{`RANDOM}};
  image_1056 = _RAND_838[3:0];
  _RAND_839 = {1{`RANDOM}};
  image_1057 = _RAND_839[3:0];
  _RAND_840 = {1{`RANDOM}};
  image_1058 = _RAND_840[3:0];
  _RAND_841 = {1{`RANDOM}};
  image_1059 = _RAND_841[3:0];
  _RAND_842 = {1{`RANDOM}};
  image_1060 = _RAND_842[3:0];
  _RAND_843 = {1{`RANDOM}};
  image_1061 = _RAND_843[3:0];
  _RAND_844 = {1{`RANDOM}};
  image_1062 = _RAND_844[3:0];
  _RAND_845 = {1{`RANDOM}};
  image_1063 = _RAND_845[3:0];
  _RAND_846 = {1{`RANDOM}};
  image_1064 = _RAND_846[3:0];
  _RAND_847 = {1{`RANDOM}};
  image_1065 = _RAND_847[3:0];
  _RAND_848 = {1{`RANDOM}};
  image_1066 = _RAND_848[3:0];
  _RAND_849 = {1{`RANDOM}};
  image_1067 = _RAND_849[3:0];
  _RAND_850 = {1{`RANDOM}};
  image_1068 = _RAND_850[3:0];
  _RAND_851 = {1{`RANDOM}};
  image_1069 = _RAND_851[3:0];
  _RAND_852 = {1{`RANDOM}};
  image_1070 = _RAND_852[3:0];
  _RAND_853 = {1{`RANDOM}};
  image_1071 = _RAND_853[3:0];
  _RAND_854 = {1{`RANDOM}};
  image_1072 = _RAND_854[3:0];
  _RAND_855 = {1{`RANDOM}};
  image_1073 = _RAND_855[3:0];
  _RAND_856 = {1{`RANDOM}};
  image_1074 = _RAND_856[3:0];
  _RAND_857 = {1{`RANDOM}};
  image_1075 = _RAND_857[3:0];
  _RAND_858 = {1{`RANDOM}};
  image_1076 = _RAND_858[3:0];
  _RAND_859 = {1{`RANDOM}};
  image_1077 = _RAND_859[3:0];
  _RAND_860 = {1{`RANDOM}};
  image_1078 = _RAND_860[3:0];
  _RAND_861 = {1{`RANDOM}};
  image_1079 = _RAND_861[3:0];
  _RAND_862 = {1{`RANDOM}};
  image_1080 = _RAND_862[3:0];
  _RAND_863 = {1{`RANDOM}};
  image_1081 = _RAND_863[3:0];
  _RAND_864 = {1{`RANDOM}};
  image_1082 = _RAND_864[3:0];
  _RAND_865 = {1{`RANDOM}};
  image_1083 = _RAND_865[3:0];
  _RAND_866 = {1{`RANDOM}};
  image_1084 = _RAND_866[3:0];
  _RAND_867 = {1{`RANDOM}};
  image_1085 = _RAND_867[3:0];
  _RAND_868 = {1{`RANDOM}};
  image_1088 = _RAND_868[3:0];
  _RAND_869 = {1{`RANDOM}};
  image_1089 = _RAND_869[3:0];
  _RAND_870 = {1{`RANDOM}};
  image_1090 = _RAND_870[3:0];
  _RAND_871 = {1{`RANDOM}};
  image_1091 = _RAND_871[3:0];
  _RAND_872 = {1{`RANDOM}};
  image_1092 = _RAND_872[3:0];
  _RAND_873 = {1{`RANDOM}};
  image_1093 = _RAND_873[3:0];
  _RAND_874 = {1{`RANDOM}};
  image_1094 = _RAND_874[3:0];
  _RAND_875 = {1{`RANDOM}};
  image_1095 = _RAND_875[3:0];
  _RAND_876 = {1{`RANDOM}};
  image_1096 = _RAND_876[3:0];
  _RAND_877 = {1{`RANDOM}};
  image_1097 = _RAND_877[3:0];
  _RAND_878 = {1{`RANDOM}};
  image_1098 = _RAND_878[3:0];
  _RAND_879 = {1{`RANDOM}};
  image_1099 = _RAND_879[3:0];
  _RAND_880 = {1{`RANDOM}};
  image_1100 = _RAND_880[3:0];
  _RAND_881 = {1{`RANDOM}};
  image_1101 = _RAND_881[3:0];
  _RAND_882 = {1{`RANDOM}};
  image_1102 = _RAND_882[3:0];
  _RAND_883 = {1{`RANDOM}};
  image_1103 = _RAND_883[3:0];
  _RAND_884 = {1{`RANDOM}};
  image_1104 = _RAND_884[3:0];
  _RAND_885 = {1{`RANDOM}};
  image_1105 = _RAND_885[3:0];
  _RAND_886 = {1{`RANDOM}};
  image_1106 = _RAND_886[3:0];
  _RAND_887 = {1{`RANDOM}};
  image_1107 = _RAND_887[3:0];
  _RAND_888 = {1{`RANDOM}};
  image_1108 = _RAND_888[3:0];
  _RAND_889 = {1{`RANDOM}};
  image_1109 = _RAND_889[3:0];
  _RAND_890 = {1{`RANDOM}};
  image_1110 = _RAND_890[3:0];
  _RAND_891 = {1{`RANDOM}};
  image_1111 = _RAND_891[3:0];
  _RAND_892 = {1{`RANDOM}};
  image_1112 = _RAND_892[3:0];
  _RAND_893 = {1{`RANDOM}};
  image_1113 = _RAND_893[3:0];
  _RAND_894 = {1{`RANDOM}};
  image_1114 = _RAND_894[3:0];
  _RAND_895 = {1{`RANDOM}};
  image_1115 = _RAND_895[3:0];
  _RAND_896 = {1{`RANDOM}};
  image_1116 = _RAND_896[3:0];
  _RAND_897 = {1{`RANDOM}};
  image_1117 = _RAND_897[3:0];
  _RAND_898 = {1{`RANDOM}};
  image_1118 = _RAND_898[3:0];
  _RAND_899 = {1{`RANDOM}};
  image_1119 = _RAND_899[3:0];
  _RAND_900 = {1{`RANDOM}};
  image_1120 = _RAND_900[3:0];
  _RAND_901 = {1{`RANDOM}};
  image_1121 = _RAND_901[3:0];
  _RAND_902 = {1{`RANDOM}};
  image_1122 = _RAND_902[3:0];
  _RAND_903 = {1{`RANDOM}};
  image_1123 = _RAND_903[3:0];
  _RAND_904 = {1{`RANDOM}};
  image_1124 = _RAND_904[3:0];
  _RAND_905 = {1{`RANDOM}};
  image_1125 = _RAND_905[3:0];
  _RAND_906 = {1{`RANDOM}};
  image_1126 = _RAND_906[3:0];
  _RAND_907 = {1{`RANDOM}};
  image_1127 = _RAND_907[3:0];
  _RAND_908 = {1{`RANDOM}};
  image_1128 = _RAND_908[3:0];
  _RAND_909 = {1{`RANDOM}};
  image_1129 = _RAND_909[3:0];
  _RAND_910 = {1{`RANDOM}};
  image_1130 = _RAND_910[3:0];
  _RAND_911 = {1{`RANDOM}};
  image_1131 = _RAND_911[3:0];
  _RAND_912 = {1{`RANDOM}};
  image_1132 = _RAND_912[3:0];
  _RAND_913 = {1{`RANDOM}};
  image_1133 = _RAND_913[3:0];
  _RAND_914 = {1{`RANDOM}};
  image_1134 = _RAND_914[3:0];
  _RAND_915 = {1{`RANDOM}};
  image_1135 = _RAND_915[3:0];
  _RAND_916 = {1{`RANDOM}};
  image_1136 = _RAND_916[3:0];
  _RAND_917 = {1{`RANDOM}};
  image_1137 = _RAND_917[3:0];
  _RAND_918 = {1{`RANDOM}};
  image_1138 = _RAND_918[3:0];
  _RAND_919 = {1{`RANDOM}};
  image_1139 = _RAND_919[3:0];
  _RAND_920 = {1{`RANDOM}};
  image_1140 = _RAND_920[3:0];
  _RAND_921 = {1{`RANDOM}};
  image_1141 = _RAND_921[3:0];
  _RAND_922 = {1{`RANDOM}};
  image_1142 = _RAND_922[3:0];
  _RAND_923 = {1{`RANDOM}};
  image_1143 = _RAND_923[3:0];
  _RAND_924 = {1{`RANDOM}};
  image_1144 = _RAND_924[3:0];
  _RAND_925 = {1{`RANDOM}};
  image_1145 = _RAND_925[3:0];
  _RAND_926 = {1{`RANDOM}};
  image_1146 = _RAND_926[3:0];
  _RAND_927 = {1{`RANDOM}};
  image_1147 = _RAND_927[3:0];
  _RAND_928 = {1{`RANDOM}};
  image_1148 = _RAND_928[3:0];
  _RAND_929 = {1{`RANDOM}};
  image_1152 = _RAND_929[3:0];
  _RAND_930 = {1{`RANDOM}};
  image_1153 = _RAND_930[3:0];
  _RAND_931 = {1{`RANDOM}};
  image_1154 = _RAND_931[3:0];
  _RAND_932 = {1{`RANDOM}};
  image_1155 = _RAND_932[3:0];
  _RAND_933 = {1{`RANDOM}};
  image_1156 = _RAND_933[3:0];
  _RAND_934 = {1{`RANDOM}};
  image_1157 = _RAND_934[3:0];
  _RAND_935 = {1{`RANDOM}};
  image_1158 = _RAND_935[3:0];
  _RAND_936 = {1{`RANDOM}};
  image_1159 = _RAND_936[3:0];
  _RAND_937 = {1{`RANDOM}};
  image_1160 = _RAND_937[3:0];
  _RAND_938 = {1{`RANDOM}};
  image_1161 = _RAND_938[3:0];
  _RAND_939 = {1{`RANDOM}};
  image_1162 = _RAND_939[3:0];
  _RAND_940 = {1{`RANDOM}};
  image_1163 = _RAND_940[3:0];
  _RAND_941 = {1{`RANDOM}};
  image_1164 = _RAND_941[3:0];
  _RAND_942 = {1{`RANDOM}};
  image_1165 = _RAND_942[3:0];
  _RAND_943 = {1{`RANDOM}};
  image_1166 = _RAND_943[3:0];
  _RAND_944 = {1{`RANDOM}};
  image_1167 = _RAND_944[3:0];
  _RAND_945 = {1{`RANDOM}};
  image_1168 = _RAND_945[3:0];
  _RAND_946 = {1{`RANDOM}};
  image_1169 = _RAND_946[3:0];
  _RAND_947 = {1{`RANDOM}};
  image_1170 = _RAND_947[3:0];
  _RAND_948 = {1{`RANDOM}};
  image_1171 = _RAND_948[3:0];
  _RAND_949 = {1{`RANDOM}};
  image_1172 = _RAND_949[3:0];
  _RAND_950 = {1{`RANDOM}};
  image_1173 = _RAND_950[3:0];
  _RAND_951 = {1{`RANDOM}};
  image_1174 = _RAND_951[3:0];
  _RAND_952 = {1{`RANDOM}};
  image_1175 = _RAND_952[3:0];
  _RAND_953 = {1{`RANDOM}};
  image_1176 = _RAND_953[3:0];
  _RAND_954 = {1{`RANDOM}};
  image_1177 = _RAND_954[3:0];
  _RAND_955 = {1{`RANDOM}};
  image_1178 = _RAND_955[3:0];
  _RAND_956 = {1{`RANDOM}};
  image_1179 = _RAND_956[3:0];
  _RAND_957 = {1{`RANDOM}};
  image_1180 = _RAND_957[3:0];
  _RAND_958 = {1{`RANDOM}};
  image_1181 = _RAND_958[3:0];
  _RAND_959 = {1{`RANDOM}};
  image_1182 = _RAND_959[3:0];
  _RAND_960 = {1{`RANDOM}};
  image_1183 = _RAND_960[3:0];
  _RAND_961 = {1{`RANDOM}};
  image_1184 = _RAND_961[3:0];
  _RAND_962 = {1{`RANDOM}};
  image_1185 = _RAND_962[3:0];
  _RAND_963 = {1{`RANDOM}};
  image_1186 = _RAND_963[3:0];
  _RAND_964 = {1{`RANDOM}};
  image_1187 = _RAND_964[3:0];
  _RAND_965 = {1{`RANDOM}};
  image_1188 = _RAND_965[3:0];
  _RAND_966 = {1{`RANDOM}};
  image_1189 = _RAND_966[3:0];
  _RAND_967 = {1{`RANDOM}};
  image_1190 = _RAND_967[3:0];
  _RAND_968 = {1{`RANDOM}};
  image_1191 = _RAND_968[3:0];
  _RAND_969 = {1{`RANDOM}};
  image_1192 = _RAND_969[3:0];
  _RAND_970 = {1{`RANDOM}};
  image_1193 = _RAND_970[3:0];
  _RAND_971 = {1{`RANDOM}};
  image_1194 = _RAND_971[3:0];
  _RAND_972 = {1{`RANDOM}};
  image_1195 = _RAND_972[3:0];
  _RAND_973 = {1{`RANDOM}};
  image_1196 = _RAND_973[3:0];
  _RAND_974 = {1{`RANDOM}};
  image_1197 = _RAND_974[3:0];
  _RAND_975 = {1{`RANDOM}};
  image_1198 = _RAND_975[3:0];
  _RAND_976 = {1{`RANDOM}};
  image_1199 = _RAND_976[3:0];
  _RAND_977 = {1{`RANDOM}};
  image_1200 = _RAND_977[3:0];
  _RAND_978 = {1{`RANDOM}};
  image_1201 = _RAND_978[3:0];
  _RAND_979 = {1{`RANDOM}};
  image_1202 = _RAND_979[3:0];
  _RAND_980 = {1{`RANDOM}};
  image_1203 = _RAND_980[3:0];
  _RAND_981 = {1{`RANDOM}};
  image_1204 = _RAND_981[3:0];
  _RAND_982 = {1{`RANDOM}};
  image_1205 = _RAND_982[3:0];
  _RAND_983 = {1{`RANDOM}};
  image_1206 = _RAND_983[3:0];
  _RAND_984 = {1{`RANDOM}};
  image_1207 = _RAND_984[3:0];
  _RAND_985 = {1{`RANDOM}};
  image_1208 = _RAND_985[3:0];
  _RAND_986 = {1{`RANDOM}};
  image_1216 = _RAND_986[3:0];
  _RAND_987 = {1{`RANDOM}};
  image_1217 = _RAND_987[3:0];
  _RAND_988 = {1{`RANDOM}};
  image_1218 = _RAND_988[3:0];
  _RAND_989 = {1{`RANDOM}};
  image_1219 = _RAND_989[3:0];
  _RAND_990 = {1{`RANDOM}};
  image_1220 = _RAND_990[3:0];
  _RAND_991 = {1{`RANDOM}};
  image_1221 = _RAND_991[3:0];
  _RAND_992 = {1{`RANDOM}};
  image_1222 = _RAND_992[3:0];
  _RAND_993 = {1{`RANDOM}};
  image_1223 = _RAND_993[3:0];
  _RAND_994 = {1{`RANDOM}};
  image_1224 = _RAND_994[3:0];
  _RAND_995 = {1{`RANDOM}};
  image_1225 = _RAND_995[3:0];
  _RAND_996 = {1{`RANDOM}};
  image_1226 = _RAND_996[3:0];
  _RAND_997 = {1{`RANDOM}};
  image_1227 = _RAND_997[3:0];
  _RAND_998 = {1{`RANDOM}};
  image_1228 = _RAND_998[3:0];
  _RAND_999 = {1{`RANDOM}};
  image_1229 = _RAND_999[3:0];
  _RAND_1000 = {1{`RANDOM}};
  image_1230 = _RAND_1000[3:0];
  _RAND_1001 = {1{`RANDOM}};
  image_1231 = _RAND_1001[3:0];
  _RAND_1002 = {1{`RANDOM}};
  image_1232 = _RAND_1002[3:0];
  _RAND_1003 = {1{`RANDOM}};
  image_1233 = _RAND_1003[3:0];
  _RAND_1004 = {1{`RANDOM}};
  image_1234 = _RAND_1004[3:0];
  _RAND_1005 = {1{`RANDOM}};
  image_1235 = _RAND_1005[3:0];
  _RAND_1006 = {1{`RANDOM}};
  image_1236 = _RAND_1006[3:0];
  _RAND_1007 = {1{`RANDOM}};
  image_1237 = _RAND_1007[3:0];
  _RAND_1008 = {1{`RANDOM}};
  image_1238 = _RAND_1008[3:0];
  _RAND_1009 = {1{`RANDOM}};
  image_1239 = _RAND_1009[3:0];
  _RAND_1010 = {1{`RANDOM}};
  image_1240 = _RAND_1010[3:0];
  _RAND_1011 = {1{`RANDOM}};
  image_1241 = _RAND_1011[3:0];
  _RAND_1012 = {1{`RANDOM}};
  image_1242 = _RAND_1012[3:0];
  _RAND_1013 = {1{`RANDOM}};
  image_1243 = _RAND_1013[3:0];
  _RAND_1014 = {1{`RANDOM}};
  image_1244 = _RAND_1014[3:0];
  _RAND_1015 = {1{`RANDOM}};
  image_1245 = _RAND_1015[3:0];
  _RAND_1016 = {1{`RANDOM}};
  image_1246 = _RAND_1016[3:0];
  _RAND_1017 = {1{`RANDOM}};
  image_1247 = _RAND_1017[3:0];
  _RAND_1018 = {1{`RANDOM}};
  image_1248 = _RAND_1018[3:0];
  _RAND_1019 = {1{`RANDOM}};
  image_1249 = _RAND_1019[3:0];
  _RAND_1020 = {1{`RANDOM}};
  image_1250 = _RAND_1020[3:0];
  _RAND_1021 = {1{`RANDOM}};
  image_1251 = _RAND_1021[3:0];
  _RAND_1022 = {1{`RANDOM}};
  image_1252 = _RAND_1022[3:0];
  _RAND_1023 = {1{`RANDOM}};
  image_1253 = _RAND_1023[3:0];
  _RAND_1024 = {1{`RANDOM}};
  image_1254 = _RAND_1024[3:0];
  _RAND_1025 = {1{`RANDOM}};
  image_1255 = _RAND_1025[3:0];
  _RAND_1026 = {1{`RANDOM}};
  image_1256 = _RAND_1026[3:0];
  _RAND_1027 = {1{`RANDOM}};
  image_1257 = _RAND_1027[3:0];
  _RAND_1028 = {1{`RANDOM}};
  image_1258 = _RAND_1028[3:0];
  _RAND_1029 = {1{`RANDOM}};
  image_1259 = _RAND_1029[3:0];
  _RAND_1030 = {1{`RANDOM}};
  image_1260 = _RAND_1030[3:0];
  _RAND_1031 = {1{`RANDOM}};
  image_1261 = _RAND_1031[3:0];
  _RAND_1032 = {1{`RANDOM}};
  image_1262 = _RAND_1032[3:0];
  _RAND_1033 = {1{`RANDOM}};
  image_1263 = _RAND_1033[3:0];
  _RAND_1034 = {1{`RANDOM}};
  image_1264 = _RAND_1034[3:0];
  _RAND_1035 = {1{`RANDOM}};
  image_1265 = _RAND_1035[3:0];
  _RAND_1036 = {1{`RANDOM}};
  image_1266 = _RAND_1036[3:0];
  _RAND_1037 = {1{`RANDOM}};
  image_1267 = _RAND_1037[3:0];
  _RAND_1038 = {1{`RANDOM}};
  image_1268 = _RAND_1038[3:0];
  _RAND_1039 = {1{`RANDOM}};
  image_1269 = _RAND_1039[3:0];
  _RAND_1040 = {1{`RANDOM}};
  image_1270 = _RAND_1040[3:0];
  _RAND_1041 = {1{`RANDOM}};
  image_1271 = _RAND_1041[3:0];
  _RAND_1042 = {1{`RANDOM}};
  image_1272 = _RAND_1042[3:0];
  _RAND_1043 = {1{`RANDOM}};
  image_1273 = _RAND_1043[3:0];
  _RAND_1044 = {1{`RANDOM}};
  image_1274 = _RAND_1044[3:0];
  _RAND_1045 = {1{`RANDOM}};
  image_1275 = _RAND_1045[3:0];
  _RAND_1046 = {1{`RANDOM}};
  image_1280 = _RAND_1046[3:0];
  _RAND_1047 = {1{`RANDOM}};
  image_1281 = _RAND_1047[3:0];
  _RAND_1048 = {1{`RANDOM}};
  image_1282 = _RAND_1048[3:0];
  _RAND_1049 = {1{`RANDOM}};
  image_1283 = _RAND_1049[3:0];
  _RAND_1050 = {1{`RANDOM}};
  image_1284 = _RAND_1050[3:0];
  _RAND_1051 = {1{`RANDOM}};
  image_1285 = _RAND_1051[3:0];
  _RAND_1052 = {1{`RANDOM}};
  image_1286 = _RAND_1052[3:0];
  _RAND_1053 = {1{`RANDOM}};
  image_1287 = _RAND_1053[3:0];
  _RAND_1054 = {1{`RANDOM}};
  image_1288 = _RAND_1054[3:0];
  _RAND_1055 = {1{`RANDOM}};
  image_1289 = _RAND_1055[3:0];
  _RAND_1056 = {1{`RANDOM}};
  image_1290 = _RAND_1056[3:0];
  _RAND_1057 = {1{`RANDOM}};
  image_1291 = _RAND_1057[3:0];
  _RAND_1058 = {1{`RANDOM}};
  image_1292 = _RAND_1058[3:0];
  _RAND_1059 = {1{`RANDOM}};
  image_1293 = _RAND_1059[3:0];
  _RAND_1060 = {1{`RANDOM}};
  image_1294 = _RAND_1060[3:0];
  _RAND_1061 = {1{`RANDOM}};
  image_1295 = _RAND_1061[3:0];
  _RAND_1062 = {1{`RANDOM}};
  image_1296 = _RAND_1062[3:0];
  _RAND_1063 = {1{`RANDOM}};
  image_1297 = _RAND_1063[3:0];
  _RAND_1064 = {1{`RANDOM}};
  image_1298 = _RAND_1064[3:0];
  _RAND_1065 = {1{`RANDOM}};
  image_1299 = _RAND_1065[3:0];
  _RAND_1066 = {1{`RANDOM}};
  image_1300 = _RAND_1066[3:0];
  _RAND_1067 = {1{`RANDOM}};
  image_1301 = _RAND_1067[3:0];
  _RAND_1068 = {1{`RANDOM}};
  image_1302 = _RAND_1068[3:0];
  _RAND_1069 = {1{`RANDOM}};
  image_1303 = _RAND_1069[3:0];
  _RAND_1070 = {1{`RANDOM}};
  image_1304 = _RAND_1070[3:0];
  _RAND_1071 = {1{`RANDOM}};
  image_1305 = _RAND_1071[3:0];
  _RAND_1072 = {1{`RANDOM}};
  image_1306 = _RAND_1072[3:0];
  _RAND_1073 = {1{`RANDOM}};
  image_1307 = _RAND_1073[3:0];
  _RAND_1074 = {1{`RANDOM}};
  image_1308 = _RAND_1074[3:0];
  _RAND_1075 = {1{`RANDOM}};
  image_1309 = _RAND_1075[3:0];
  _RAND_1076 = {1{`RANDOM}};
  image_1310 = _RAND_1076[3:0];
  _RAND_1077 = {1{`RANDOM}};
  image_1311 = _RAND_1077[3:0];
  _RAND_1078 = {1{`RANDOM}};
  image_1312 = _RAND_1078[3:0];
  _RAND_1079 = {1{`RANDOM}};
  image_1313 = _RAND_1079[3:0];
  _RAND_1080 = {1{`RANDOM}};
  image_1314 = _RAND_1080[3:0];
  _RAND_1081 = {1{`RANDOM}};
  image_1315 = _RAND_1081[3:0];
  _RAND_1082 = {1{`RANDOM}};
  image_1316 = _RAND_1082[3:0];
  _RAND_1083 = {1{`RANDOM}};
  image_1317 = _RAND_1083[3:0];
  _RAND_1084 = {1{`RANDOM}};
  image_1318 = _RAND_1084[3:0];
  _RAND_1085 = {1{`RANDOM}};
  image_1319 = _RAND_1085[3:0];
  _RAND_1086 = {1{`RANDOM}};
  image_1320 = _RAND_1086[3:0];
  _RAND_1087 = {1{`RANDOM}};
  image_1321 = _RAND_1087[3:0];
  _RAND_1088 = {1{`RANDOM}};
  image_1322 = _RAND_1088[3:0];
  _RAND_1089 = {1{`RANDOM}};
  image_1323 = _RAND_1089[3:0];
  _RAND_1090 = {1{`RANDOM}};
  image_1324 = _RAND_1090[3:0];
  _RAND_1091 = {1{`RANDOM}};
  image_1325 = _RAND_1091[3:0];
  _RAND_1092 = {1{`RANDOM}};
  image_1326 = _RAND_1092[3:0];
  _RAND_1093 = {1{`RANDOM}};
  image_1327 = _RAND_1093[3:0];
  _RAND_1094 = {1{`RANDOM}};
  image_1328 = _RAND_1094[3:0];
  _RAND_1095 = {1{`RANDOM}};
  image_1329 = _RAND_1095[3:0];
  _RAND_1096 = {1{`RANDOM}};
  image_1330 = _RAND_1096[3:0];
  _RAND_1097 = {1{`RANDOM}};
  image_1331 = _RAND_1097[3:0];
  _RAND_1098 = {1{`RANDOM}};
  image_1332 = _RAND_1098[3:0];
  _RAND_1099 = {1{`RANDOM}};
  image_1333 = _RAND_1099[3:0];
  _RAND_1100 = {1{`RANDOM}};
  image_1334 = _RAND_1100[3:0];
  _RAND_1101 = {1{`RANDOM}};
  image_1335 = _RAND_1101[3:0];
  _RAND_1102 = {1{`RANDOM}};
  image_1336 = _RAND_1102[3:0];
  _RAND_1103 = {1{`RANDOM}};
  image_1337 = _RAND_1103[3:0];
  _RAND_1104 = {1{`RANDOM}};
  image_1338 = _RAND_1104[3:0];
  _RAND_1105 = {1{`RANDOM}};
  image_1339 = _RAND_1105[3:0];
  _RAND_1106 = {1{`RANDOM}};
  image_1340 = _RAND_1106[3:0];
  _RAND_1107 = {1{`RANDOM}};
  image_1341 = _RAND_1107[3:0];
  _RAND_1108 = {1{`RANDOM}};
  image_1344 = _RAND_1108[3:0];
  _RAND_1109 = {1{`RANDOM}};
  image_1345 = _RAND_1109[3:0];
  _RAND_1110 = {1{`RANDOM}};
  image_1346 = _RAND_1110[3:0];
  _RAND_1111 = {1{`RANDOM}};
  image_1347 = _RAND_1111[3:0];
  _RAND_1112 = {1{`RANDOM}};
  image_1348 = _RAND_1112[3:0];
  _RAND_1113 = {1{`RANDOM}};
  image_1349 = _RAND_1113[3:0];
  _RAND_1114 = {1{`RANDOM}};
  image_1350 = _RAND_1114[3:0];
  _RAND_1115 = {1{`RANDOM}};
  image_1351 = _RAND_1115[3:0];
  _RAND_1116 = {1{`RANDOM}};
  image_1352 = _RAND_1116[3:0];
  _RAND_1117 = {1{`RANDOM}};
  image_1353 = _RAND_1117[3:0];
  _RAND_1118 = {1{`RANDOM}};
  image_1354 = _RAND_1118[3:0];
  _RAND_1119 = {1{`RANDOM}};
  image_1355 = _RAND_1119[3:0];
  _RAND_1120 = {1{`RANDOM}};
  image_1356 = _RAND_1120[3:0];
  _RAND_1121 = {1{`RANDOM}};
  image_1357 = _RAND_1121[3:0];
  _RAND_1122 = {1{`RANDOM}};
  image_1358 = _RAND_1122[3:0];
  _RAND_1123 = {1{`RANDOM}};
  image_1359 = _RAND_1123[3:0];
  _RAND_1124 = {1{`RANDOM}};
  image_1360 = _RAND_1124[3:0];
  _RAND_1125 = {1{`RANDOM}};
  image_1361 = _RAND_1125[3:0];
  _RAND_1126 = {1{`RANDOM}};
  image_1362 = _RAND_1126[3:0];
  _RAND_1127 = {1{`RANDOM}};
  image_1363 = _RAND_1127[3:0];
  _RAND_1128 = {1{`RANDOM}};
  image_1364 = _RAND_1128[3:0];
  _RAND_1129 = {1{`RANDOM}};
  image_1365 = _RAND_1129[3:0];
  _RAND_1130 = {1{`RANDOM}};
  image_1366 = _RAND_1130[3:0];
  _RAND_1131 = {1{`RANDOM}};
  image_1367 = _RAND_1131[3:0];
  _RAND_1132 = {1{`RANDOM}};
  image_1368 = _RAND_1132[3:0];
  _RAND_1133 = {1{`RANDOM}};
  image_1369 = _RAND_1133[3:0];
  _RAND_1134 = {1{`RANDOM}};
  image_1370 = _RAND_1134[3:0];
  _RAND_1135 = {1{`RANDOM}};
  image_1371 = _RAND_1135[3:0];
  _RAND_1136 = {1{`RANDOM}};
  image_1372 = _RAND_1136[3:0];
  _RAND_1137 = {1{`RANDOM}};
  image_1373 = _RAND_1137[3:0];
  _RAND_1138 = {1{`RANDOM}};
  image_1374 = _RAND_1138[3:0];
  _RAND_1139 = {1{`RANDOM}};
  image_1375 = _RAND_1139[3:0];
  _RAND_1140 = {1{`RANDOM}};
  image_1376 = _RAND_1140[3:0];
  _RAND_1141 = {1{`RANDOM}};
  image_1377 = _RAND_1141[3:0];
  _RAND_1142 = {1{`RANDOM}};
  image_1378 = _RAND_1142[3:0];
  _RAND_1143 = {1{`RANDOM}};
  image_1379 = _RAND_1143[3:0];
  _RAND_1144 = {1{`RANDOM}};
  image_1380 = _RAND_1144[3:0];
  _RAND_1145 = {1{`RANDOM}};
  image_1381 = _RAND_1145[3:0];
  _RAND_1146 = {1{`RANDOM}};
  image_1382 = _RAND_1146[3:0];
  _RAND_1147 = {1{`RANDOM}};
  image_1383 = _RAND_1147[3:0];
  _RAND_1148 = {1{`RANDOM}};
  image_1384 = _RAND_1148[3:0];
  _RAND_1149 = {1{`RANDOM}};
  image_1385 = _RAND_1149[3:0];
  _RAND_1150 = {1{`RANDOM}};
  image_1386 = _RAND_1150[3:0];
  _RAND_1151 = {1{`RANDOM}};
  image_1387 = _RAND_1151[3:0];
  _RAND_1152 = {1{`RANDOM}};
  image_1388 = _RAND_1152[3:0];
  _RAND_1153 = {1{`RANDOM}};
  image_1389 = _RAND_1153[3:0];
  _RAND_1154 = {1{`RANDOM}};
  image_1390 = _RAND_1154[3:0];
  _RAND_1155 = {1{`RANDOM}};
  image_1391 = _RAND_1155[3:0];
  _RAND_1156 = {1{`RANDOM}};
  image_1392 = _RAND_1156[3:0];
  _RAND_1157 = {1{`RANDOM}};
  image_1393 = _RAND_1157[3:0];
  _RAND_1158 = {1{`RANDOM}};
  image_1394 = _RAND_1158[3:0];
  _RAND_1159 = {1{`RANDOM}};
  image_1395 = _RAND_1159[3:0];
  _RAND_1160 = {1{`RANDOM}};
  image_1396 = _RAND_1160[3:0];
  _RAND_1161 = {1{`RANDOM}};
  image_1397 = _RAND_1161[3:0];
  _RAND_1162 = {1{`RANDOM}};
  image_1398 = _RAND_1162[3:0];
  _RAND_1163 = {1{`RANDOM}};
  image_1399 = _RAND_1163[3:0];
  _RAND_1164 = {1{`RANDOM}};
  image_1400 = _RAND_1164[3:0];
  _RAND_1165 = {1{`RANDOM}};
  image_1401 = _RAND_1165[3:0];
  _RAND_1166 = {1{`RANDOM}};
  image_1402 = _RAND_1166[3:0];
  _RAND_1167 = {1{`RANDOM}};
  image_1403 = _RAND_1167[3:0];
  _RAND_1168 = {1{`RANDOM}};
  image_1404 = _RAND_1168[3:0];
  _RAND_1169 = {1{`RANDOM}};
  image_1405 = _RAND_1169[3:0];
  _RAND_1170 = {1{`RANDOM}};
  image_1408 = _RAND_1170[3:0];
  _RAND_1171 = {1{`RANDOM}};
  image_1409 = _RAND_1171[3:0];
  _RAND_1172 = {1{`RANDOM}};
  image_1410 = _RAND_1172[3:0];
  _RAND_1173 = {1{`RANDOM}};
  image_1411 = _RAND_1173[3:0];
  _RAND_1174 = {1{`RANDOM}};
  image_1412 = _RAND_1174[3:0];
  _RAND_1175 = {1{`RANDOM}};
  image_1413 = _RAND_1175[3:0];
  _RAND_1176 = {1{`RANDOM}};
  image_1414 = _RAND_1176[3:0];
  _RAND_1177 = {1{`RANDOM}};
  image_1415 = _RAND_1177[3:0];
  _RAND_1178 = {1{`RANDOM}};
  image_1416 = _RAND_1178[3:0];
  _RAND_1179 = {1{`RANDOM}};
  image_1417 = _RAND_1179[3:0];
  _RAND_1180 = {1{`RANDOM}};
  image_1418 = _RAND_1180[3:0];
  _RAND_1181 = {1{`RANDOM}};
  image_1419 = _RAND_1181[3:0];
  _RAND_1182 = {1{`RANDOM}};
  image_1420 = _RAND_1182[3:0];
  _RAND_1183 = {1{`RANDOM}};
  image_1421 = _RAND_1183[3:0];
  _RAND_1184 = {1{`RANDOM}};
  image_1422 = _RAND_1184[3:0];
  _RAND_1185 = {1{`RANDOM}};
  image_1423 = _RAND_1185[3:0];
  _RAND_1186 = {1{`RANDOM}};
  image_1424 = _RAND_1186[3:0];
  _RAND_1187 = {1{`RANDOM}};
  image_1425 = _RAND_1187[3:0];
  _RAND_1188 = {1{`RANDOM}};
  image_1426 = _RAND_1188[3:0];
  _RAND_1189 = {1{`RANDOM}};
  image_1427 = _RAND_1189[3:0];
  _RAND_1190 = {1{`RANDOM}};
  image_1428 = _RAND_1190[3:0];
  _RAND_1191 = {1{`RANDOM}};
  image_1429 = _RAND_1191[3:0];
  _RAND_1192 = {1{`RANDOM}};
  image_1430 = _RAND_1192[3:0];
  _RAND_1193 = {1{`RANDOM}};
  image_1431 = _RAND_1193[3:0];
  _RAND_1194 = {1{`RANDOM}};
  image_1432 = _RAND_1194[3:0];
  _RAND_1195 = {1{`RANDOM}};
  image_1433 = _RAND_1195[3:0];
  _RAND_1196 = {1{`RANDOM}};
  image_1434 = _RAND_1196[3:0];
  _RAND_1197 = {1{`RANDOM}};
  image_1435 = _RAND_1197[3:0];
  _RAND_1198 = {1{`RANDOM}};
  image_1436 = _RAND_1198[3:0];
  _RAND_1199 = {1{`RANDOM}};
  image_1437 = _RAND_1199[3:0];
  _RAND_1200 = {1{`RANDOM}};
  image_1438 = _RAND_1200[3:0];
  _RAND_1201 = {1{`RANDOM}};
  image_1439 = _RAND_1201[3:0];
  _RAND_1202 = {1{`RANDOM}};
  image_1440 = _RAND_1202[3:0];
  _RAND_1203 = {1{`RANDOM}};
  image_1441 = _RAND_1203[3:0];
  _RAND_1204 = {1{`RANDOM}};
  image_1442 = _RAND_1204[3:0];
  _RAND_1205 = {1{`RANDOM}};
  image_1443 = _RAND_1205[3:0];
  _RAND_1206 = {1{`RANDOM}};
  image_1444 = _RAND_1206[3:0];
  _RAND_1207 = {1{`RANDOM}};
  image_1445 = _RAND_1207[3:0];
  _RAND_1208 = {1{`RANDOM}};
  image_1446 = _RAND_1208[3:0];
  _RAND_1209 = {1{`RANDOM}};
  image_1447 = _RAND_1209[3:0];
  _RAND_1210 = {1{`RANDOM}};
  image_1448 = _RAND_1210[3:0];
  _RAND_1211 = {1{`RANDOM}};
  image_1449 = _RAND_1211[3:0];
  _RAND_1212 = {1{`RANDOM}};
  image_1450 = _RAND_1212[3:0];
  _RAND_1213 = {1{`RANDOM}};
  image_1451 = _RAND_1213[3:0];
  _RAND_1214 = {1{`RANDOM}};
  image_1452 = _RAND_1214[3:0];
  _RAND_1215 = {1{`RANDOM}};
  image_1453 = _RAND_1215[3:0];
  _RAND_1216 = {1{`RANDOM}};
  image_1454 = _RAND_1216[3:0];
  _RAND_1217 = {1{`RANDOM}};
  image_1455 = _RAND_1217[3:0];
  _RAND_1218 = {1{`RANDOM}};
  image_1456 = _RAND_1218[3:0];
  _RAND_1219 = {1{`RANDOM}};
  image_1457 = _RAND_1219[3:0];
  _RAND_1220 = {1{`RANDOM}};
  image_1458 = _RAND_1220[3:0];
  _RAND_1221 = {1{`RANDOM}};
  image_1459 = _RAND_1221[3:0];
  _RAND_1222 = {1{`RANDOM}};
  image_1460 = _RAND_1222[3:0];
  _RAND_1223 = {1{`RANDOM}};
  image_1461 = _RAND_1223[3:0];
  _RAND_1224 = {1{`RANDOM}};
  image_1462 = _RAND_1224[3:0];
  _RAND_1225 = {1{`RANDOM}};
  image_1463 = _RAND_1225[3:0];
  _RAND_1226 = {1{`RANDOM}};
  image_1464 = _RAND_1226[3:0];
  _RAND_1227 = {1{`RANDOM}};
  image_1465 = _RAND_1227[3:0];
  _RAND_1228 = {1{`RANDOM}};
  image_1466 = _RAND_1228[3:0];
  _RAND_1229 = {1{`RANDOM}};
  image_1467 = _RAND_1229[3:0];
  _RAND_1230 = {1{`RANDOM}};
  image_1468 = _RAND_1230[3:0];
  _RAND_1231 = {1{`RANDOM}};
  image_1469 = _RAND_1231[3:0];
  _RAND_1232 = {1{`RANDOM}};
  image_1472 = _RAND_1232[3:0];
  _RAND_1233 = {1{`RANDOM}};
  image_1473 = _RAND_1233[3:0];
  _RAND_1234 = {1{`RANDOM}};
  image_1474 = _RAND_1234[3:0];
  _RAND_1235 = {1{`RANDOM}};
  image_1475 = _RAND_1235[3:0];
  _RAND_1236 = {1{`RANDOM}};
  image_1476 = _RAND_1236[3:0];
  _RAND_1237 = {1{`RANDOM}};
  image_1477 = _RAND_1237[3:0];
  _RAND_1238 = {1{`RANDOM}};
  image_1478 = _RAND_1238[3:0];
  _RAND_1239 = {1{`RANDOM}};
  image_1479 = _RAND_1239[3:0];
  _RAND_1240 = {1{`RANDOM}};
  image_1480 = _RAND_1240[3:0];
  _RAND_1241 = {1{`RANDOM}};
  image_1481 = _RAND_1241[3:0];
  _RAND_1242 = {1{`RANDOM}};
  image_1482 = _RAND_1242[3:0];
  _RAND_1243 = {1{`RANDOM}};
  image_1483 = _RAND_1243[3:0];
  _RAND_1244 = {1{`RANDOM}};
  image_1484 = _RAND_1244[3:0];
  _RAND_1245 = {1{`RANDOM}};
  image_1485 = _RAND_1245[3:0];
  _RAND_1246 = {1{`RANDOM}};
  image_1486 = _RAND_1246[3:0];
  _RAND_1247 = {1{`RANDOM}};
  image_1487 = _RAND_1247[3:0];
  _RAND_1248 = {1{`RANDOM}};
  image_1488 = _RAND_1248[3:0];
  _RAND_1249 = {1{`RANDOM}};
  image_1489 = _RAND_1249[3:0];
  _RAND_1250 = {1{`RANDOM}};
  image_1490 = _RAND_1250[3:0];
  _RAND_1251 = {1{`RANDOM}};
  image_1491 = _RAND_1251[3:0];
  _RAND_1252 = {1{`RANDOM}};
  image_1492 = _RAND_1252[3:0];
  _RAND_1253 = {1{`RANDOM}};
  image_1493 = _RAND_1253[3:0];
  _RAND_1254 = {1{`RANDOM}};
  image_1494 = _RAND_1254[3:0];
  _RAND_1255 = {1{`RANDOM}};
  image_1495 = _RAND_1255[3:0];
  _RAND_1256 = {1{`RANDOM}};
  image_1496 = _RAND_1256[3:0];
  _RAND_1257 = {1{`RANDOM}};
  image_1497 = _RAND_1257[3:0];
  _RAND_1258 = {1{`RANDOM}};
  image_1498 = _RAND_1258[3:0];
  _RAND_1259 = {1{`RANDOM}};
  image_1499 = _RAND_1259[3:0];
  _RAND_1260 = {1{`RANDOM}};
  image_1500 = _RAND_1260[3:0];
  _RAND_1261 = {1{`RANDOM}};
  image_1501 = _RAND_1261[3:0];
  _RAND_1262 = {1{`RANDOM}};
  image_1502 = _RAND_1262[3:0];
  _RAND_1263 = {1{`RANDOM}};
  image_1503 = _RAND_1263[3:0];
  _RAND_1264 = {1{`RANDOM}};
  image_1504 = _RAND_1264[3:0];
  _RAND_1265 = {1{`RANDOM}};
  image_1505 = _RAND_1265[3:0];
  _RAND_1266 = {1{`RANDOM}};
  image_1506 = _RAND_1266[3:0];
  _RAND_1267 = {1{`RANDOM}};
  image_1507 = _RAND_1267[3:0];
  _RAND_1268 = {1{`RANDOM}};
  image_1508 = _RAND_1268[3:0];
  _RAND_1269 = {1{`RANDOM}};
  image_1509 = _RAND_1269[3:0];
  _RAND_1270 = {1{`RANDOM}};
  image_1510 = _RAND_1270[3:0];
  _RAND_1271 = {1{`RANDOM}};
  image_1511 = _RAND_1271[3:0];
  _RAND_1272 = {1{`RANDOM}};
  image_1512 = _RAND_1272[3:0];
  _RAND_1273 = {1{`RANDOM}};
  image_1513 = _RAND_1273[3:0];
  _RAND_1274 = {1{`RANDOM}};
  image_1514 = _RAND_1274[3:0];
  _RAND_1275 = {1{`RANDOM}};
  image_1515 = _RAND_1275[3:0];
  _RAND_1276 = {1{`RANDOM}};
  image_1516 = _RAND_1276[3:0];
  _RAND_1277 = {1{`RANDOM}};
  image_1517 = _RAND_1277[3:0];
  _RAND_1278 = {1{`RANDOM}};
  image_1518 = _RAND_1278[3:0];
  _RAND_1279 = {1{`RANDOM}};
  image_1519 = _RAND_1279[3:0];
  _RAND_1280 = {1{`RANDOM}};
  image_1520 = _RAND_1280[3:0];
  _RAND_1281 = {1{`RANDOM}};
  image_1521 = _RAND_1281[3:0];
  _RAND_1282 = {1{`RANDOM}};
  image_1522 = _RAND_1282[3:0];
  _RAND_1283 = {1{`RANDOM}};
  image_1523 = _RAND_1283[3:0];
  _RAND_1284 = {1{`RANDOM}};
  image_1524 = _RAND_1284[3:0];
  _RAND_1285 = {1{`RANDOM}};
  image_1525 = _RAND_1285[3:0];
  _RAND_1286 = {1{`RANDOM}};
  image_1526 = _RAND_1286[3:0];
  _RAND_1287 = {1{`RANDOM}};
  image_1527 = _RAND_1287[3:0];
  _RAND_1288 = {1{`RANDOM}};
  image_1528 = _RAND_1288[3:0];
  _RAND_1289 = {1{`RANDOM}};
  image_1529 = _RAND_1289[3:0];
  _RAND_1290 = {1{`RANDOM}};
  image_1530 = _RAND_1290[3:0];
  _RAND_1291 = {1{`RANDOM}};
  image_1531 = _RAND_1291[3:0];
  _RAND_1292 = {1{`RANDOM}};
  image_1532 = _RAND_1292[3:0];
  _RAND_1293 = {1{`RANDOM}};
  image_1533 = _RAND_1293[3:0];
  _RAND_1294 = {1{`RANDOM}};
  image_1536 = _RAND_1294[3:0];
  _RAND_1295 = {1{`RANDOM}};
  image_1537 = _RAND_1295[3:0];
  _RAND_1296 = {1{`RANDOM}};
  image_1538 = _RAND_1296[3:0];
  _RAND_1297 = {1{`RANDOM}};
  image_1539 = _RAND_1297[3:0];
  _RAND_1298 = {1{`RANDOM}};
  image_1540 = _RAND_1298[3:0];
  _RAND_1299 = {1{`RANDOM}};
  image_1541 = _RAND_1299[3:0];
  _RAND_1300 = {1{`RANDOM}};
  image_1542 = _RAND_1300[3:0];
  _RAND_1301 = {1{`RANDOM}};
  image_1543 = _RAND_1301[3:0];
  _RAND_1302 = {1{`RANDOM}};
  image_1544 = _RAND_1302[3:0];
  _RAND_1303 = {1{`RANDOM}};
  image_1545 = _RAND_1303[3:0];
  _RAND_1304 = {1{`RANDOM}};
  image_1546 = _RAND_1304[3:0];
  _RAND_1305 = {1{`RANDOM}};
  image_1547 = _RAND_1305[3:0];
  _RAND_1306 = {1{`RANDOM}};
  image_1548 = _RAND_1306[3:0];
  _RAND_1307 = {1{`RANDOM}};
  image_1549 = _RAND_1307[3:0];
  _RAND_1308 = {1{`RANDOM}};
  image_1550 = _RAND_1308[3:0];
  _RAND_1309 = {1{`RANDOM}};
  image_1551 = _RAND_1309[3:0];
  _RAND_1310 = {1{`RANDOM}};
  image_1552 = _RAND_1310[3:0];
  _RAND_1311 = {1{`RANDOM}};
  image_1553 = _RAND_1311[3:0];
  _RAND_1312 = {1{`RANDOM}};
  image_1554 = _RAND_1312[3:0];
  _RAND_1313 = {1{`RANDOM}};
  image_1555 = _RAND_1313[3:0];
  _RAND_1314 = {1{`RANDOM}};
  image_1556 = _RAND_1314[3:0];
  _RAND_1315 = {1{`RANDOM}};
  image_1557 = _RAND_1315[3:0];
  _RAND_1316 = {1{`RANDOM}};
  image_1558 = _RAND_1316[3:0];
  _RAND_1317 = {1{`RANDOM}};
  image_1559 = _RAND_1317[3:0];
  _RAND_1318 = {1{`RANDOM}};
  image_1560 = _RAND_1318[3:0];
  _RAND_1319 = {1{`RANDOM}};
  image_1561 = _RAND_1319[3:0];
  _RAND_1320 = {1{`RANDOM}};
  image_1562 = _RAND_1320[3:0];
  _RAND_1321 = {1{`RANDOM}};
  image_1563 = _RAND_1321[3:0];
  _RAND_1322 = {1{`RANDOM}};
  image_1564 = _RAND_1322[3:0];
  _RAND_1323 = {1{`RANDOM}};
  image_1565 = _RAND_1323[3:0];
  _RAND_1324 = {1{`RANDOM}};
  image_1566 = _RAND_1324[3:0];
  _RAND_1325 = {1{`RANDOM}};
  image_1567 = _RAND_1325[3:0];
  _RAND_1326 = {1{`RANDOM}};
  image_1568 = _RAND_1326[3:0];
  _RAND_1327 = {1{`RANDOM}};
  image_1569 = _RAND_1327[3:0];
  _RAND_1328 = {1{`RANDOM}};
  image_1570 = _RAND_1328[3:0];
  _RAND_1329 = {1{`RANDOM}};
  image_1571 = _RAND_1329[3:0];
  _RAND_1330 = {1{`RANDOM}};
  image_1572 = _RAND_1330[3:0];
  _RAND_1331 = {1{`RANDOM}};
  image_1573 = _RAND_1331[3:0];
  _RAND_1332 = {1{`RANDOM}};
  image_1574 = _RAND_1332[3:0];
  _RAND_1333 = {1{`RANDOM}};
  image_1575 = _RAND_1333[3:0];
  _RAND_1334 = {1{`RANDOM}};
  image_1576 = _RAND_1334[3:0];
  _RAND_1335 = {1{`RANDOM}};
  image_1577 = _RAND_1335[3:0];
  _RAND_1336 = {1{`RANDOM}};
  image_1578 = _RAND_1336[3:0];
  _RAND_1337 = {1{`RANDOM}};
  image_1579 = _RAND_1337[3:0];
  _RAND_1338 = {1{`RANDOM}};
  image_1580 = _RAND_1338[3:0];
  _RAND_1339 = {1{`RANDOM}};
  image_1581 = _RAND_1339[3:0];
  _RAND_1340 = {1{`RANDOM}};
  image_1582 = _RAND_1340[3:0];
  _RAND_1341 = {1{`RANDOM}};
  image_1583 = _RAND_1341[3:0];
  _RAND_1342 = {1{`RANDOM}};
  image_1584 = _RAND_1342[3:0];
  _RAND_1343 = {1{`RANDOM}};
  image_1585 = _RAND_1343[3:0];
  _RAND_1344 = {1{`RANDOM}};
  image_1586 = _RAND_1344[3:0];
  _RAND_1345 = {1{`RANDOM}};
  image_1587 = _RAND_1345[3:0];
  _RAND_1346 = {1{`RANDOM}};
  image_1588 = _RAND_1346[3:0];
  _RAND_1347 = {1{`RANDOM}};
  image_1589 = _RAND_1347[3:0];
  _RAND_1348 = {1{`RANDOM}};
  image_1590 = _RAND_1348[3:0];
  _RAND_1349 = {1{`RANDOM}};
  image_1591 = _RAND_1349[3:0];
  _RAND_1350 = {1{`RANDOM}};
  image_1592 = _RAND_1350[3:0];
  _RAND_1351 = {1{`RANDOM}};
  image_1593 = _RAND_1351[3:0];
  _RAND_1352 = {1{`RANDOM}};
  image_1594 = _RAND_1352[3:0];
  _RAND_1353 = {1{`RANDOM}};
  image_1595 = _RAND_1353[3:0];
  _RAND_1354 = {1{`RANDOM}};
  image_1596 = _RAND_1354[3:0];
  _RAND_1355 = {1{`RANDOM}};
  image_1597 = _RAND_1355[3:0];
  _RAND_1356 = {1{`RANDOM}};
  image_1600 = _RAND_1356[3:0];
  _RAND_1357 = {1{`RANDOM}};
  image_1601 = _RAND_1357[3:0];
  _RAND_1358 = {1{`RANDOM}};
  image_1602 = _RAND_1358[3:0];
  _RAND_1359 = {1{`RANDOM}};
  image_1603 = _RAND_1359[3:0];
  _RAND_1360 = {1{`RANDOM}};
  image_1604 = _RAND_1360[3:0];
  _RAND_1361 = {1{`RANDOM}};
  image_1605 = _RAND_1361[3:0];
  _RAND_1362 = {1{`RANDOM}};
  image_1606 = _RAND_1362[3:0];
  _RAND_1363 = {1{`RANDOM}};
  image_1607 = _RAND_1363[3:0];
  _RAND_1364 = {1{`RANDOM}};
  image_1608 = _RAND_1364[3:0];
  _RAND_1365 = {1{`RANDOM}};
  image_1609 = _RAND_1365[3:0];
  _RAND_1366 = {1{`RANDOM}};
  image_1610 = _RAND_1366[3:0];
  _RAND_1367 = {1{`RANDOM}};
  image_1611 = _RAND_1367[3:0];
  _RAND_1368 = {1{`RANDOM}};
  image_1612 = _RAND_1368[3:0];
  _RAND_1369 = {1{`RANDOM}};
  image_1613 = _RAND_1369[3:0];
  _RAND_1370 = {1{`RANDOM}};
  image_1614 = _RAND_1370[3:0];
  _RAND_1371 = {1{`RANDOM}};
  image_1615 = _RAND_1371[3:0];
  _RAND_1372 = {1{`RANDOM}};
  image_1616 = _RAND_1372[3:0];
  _RAND_1373 = {1{`RANDOM}};
  image_1617 = _RAND_1373[3:0];
  _RAND_1374 = {1{`RANDOM}};
  image_1618 = _RAND_1374[3:0];
  _RAND_1375 = {1{`RANDOM}};
  image_1619 = _RAND_1375[3:0];
  _RAND_1376 = {1{`RANDOM}};
  image_1620 = _RAND_1376[3:0];
  _RAND_1377 = {1{`RANDOM}};
  image_1621 = _RAND_1377[3:0];
  _RAND_1378 = {1{`RANDOM}};
  image_1622 = _RAND_1378[3:0];
  _RAND_1379 = {1{`RANDOM}};
  image_1623 = _RAND_1379[3:0];
  _RAND_1380 = {1{`RANDOM}};
  image_1624 = _RAND_1380[3:0];
  _RAND_1381 = {1{`RANDOM}};
  image_1625 = _RAND_1381[3:0];
  _RAND_1382 = {1{`RANDOM}};
  image_1626 = _RAND_1382[3:0];
  _RAND_1383 = {1{`RANDOM}};
  image_1627 = _RAND_1383[3:0];
  _RAND_1384 = {1{`RANDOM}};
  image_1628 = _RAND_1384[3:0];
  _RAND_1385 = {1{`RANDOM}};
  image_1629 = _RAND_1385[3:0];
  _RAND_1386 = {1{`RANDOM}};
  image_1630 = _RAND_1386[3:0];
  _RAND_1387 = {1{`RANDOM}};
  image_1631 = _RAND_1387[3:0];
  _RAND_1388 = {1{`RANDOM}};
  image_1632 = _RAND_1388[3:0];
  _RAND_1389 = {1{`RANDOM}};
  image_1633 = _RAND_1389[3:0];
  _RAND_1390 = {1{`RANDOM}};
  image_1634 = _RAND_1390[3:0];
  _RAND_1391 = {1{`RANDOM}};
  image_1635 = _RAND_1391[3:0];
  _RAND_1392 = {1{`RANDOM}};
  image_1636 = _RAND_1392[3:0];
  _RAND_1393 = {1{`RANDOM}};
  image_1637 = _RAND_1393[3:0];
  _RAND_1394 = {1{`RANDOM}};
  image_1638 = _RAND_1394[3:0];
  _RAND_1395 = {1{`RANDOM}};
  image_1639 = _RAND_1395[3:0];
  _RAND_1396 = {1{`RANDOM}};
  image_1640 = _RAND_1396[3:0];
  _RAND_1397 = {1{`RANDOM}};
  image_1641 = _RAND_1397[3:0];
  _RAND_1398 = {1{`RANDOM}};
  image_1642 = _RAND_1398[3:0];
  _RAND_1399 = {1{`RANDOM}};
  image_1643 = _RAND_1399[3:0];
  _RAND_1400 = {1{`RANDOM}};
  image_1644 = _RAND_1400[3:0];
  _RAND_1401 = {1{`RANDOM}};
  image_1645 = _RAND_1401[3:0];
  _RAND_1402 = {1{`RANDOM}};
  image_1646 = _RAND_1402[3:0];
  _RAND_1403 = {1{`RANDOM}};
  image_1647 = _RAND_1403[3:0];
  _RAND_1404 = {1{`RANDOM}};
  image_1648 = _RAND_1404[3:0];
  _RAND_1405 = {1{`RANDOM}};
  image_1649 = _RAND_1405[3:0];
  _RAND_1406 = {1{`RANDOM}};
  image_1650 = _RAND_1406[3:0];
  _RAND_1407 = {1{`RANDOM}};
  image_1651 = _RAND_1407[3:0];
  _RAND_1408 = {1{`RANDOM}};
  image_1652 = _RAND_1408[3:0];
  _RAND_1409 = {1{`RANDOM}};
  image_1653 = _RAND_1409[3:0];
  _RAND_1410 = {1{`RANDOM}};
  image_1654 = _RAND_1410[3:0];
  _RAND_1411 = {1{`RANDOM}};
  image_1655 = _RAND_1411[3:0];
  _RAND_1412 = {1{`RANDOM}};
  image_1656 = _RAND_1412[3:0];
  _RAND_1413 = {1{`RANDOM}};
  image_1657 = _RAND_1413[3:0];
  _RAND_1414 = {1{`RANDOM}};
  image_1658 = _RAND_1414[3:0];
  _RAND_1415 = {1{`RANDOM}};
  image_1659 = _RAND_1415[3:0];
  _RAND_1416 = {1{`RANDOM}};
  image_1660 = _RAND_1416[3:0];
  _RAND_1417 = {1{`RANDOM}};
  image_1664 = _RAND_1417[3:0];
  _RAND_1418 = {1{`RANDOM}};
  image_1665 = _RAND_1418[3:0];
  _RAND_1419 = {1{`RANDOM}};
  image_1666 = _RAND_1419[3:0];
  _RAND_1420 = {1{`RANDOM}};
  image_1667 = _RAND_1420[3:0];
  _RAND_1421 = {1{`RANDOM}};
  image_1668 = _RAND_1421[3:0];
  _RAND_1422 = {1{`RANDOM}};
  image_1669 = _RAND_1422[3:0];
  _RAND_1423 = {1{`RANDOM}};
  image_1670 = _RAND_1423[3:0];
  _RAND_1424 = {1{`RANDOM}};
  image_1671 = _RAND_1424[3:0];
  _RAND_1425 = {1{`RANDOM}};
  image_1672 = _RAND_1425[3:0];
  _RAND_1426 = {1{`RANDOM}};
  image_1673 = _RAND_1426[3:0];
  _RAND_1427 = {1{`RANDOM}};
  image_1674 = _RAND_1427[3:0];
  _RAND_1428 = {1{`RANDOM}};
  image_1675 = _RAND_1428[3:0];
  _RAND_1429 = {1{`RANDOM}};
  image_1676 = _RAND_1429[3:0];
  _RAND_1430 = {1{`RANDOM}};
  image_1677 = _RAND_1430[3:0];
  _RAND_1431 = {1{`RANDOM}};
  image_1678 = _RAND_1431[3:0];
  _RAND_1432 = {1{`RANDOM}};
  image_1679 = _RAND_1432[3:0];
  _RAND_1433 = {1{`RANDOM}};
  image_1680 = _RAND_1433[3:0];
  _RAND_1434 = {1{`RANDOM}};
  image_1681 = _RAND_1434[3:0];
  _RAND_1435 = {1{`RANDOM}};
  image_1682 = _RAND_1435[3:0];
  _RAND_1436 = {1{`RANDOM}};
  image_1683 = _RAND_1436[3:0];
  _RAND_1437 = {1{`RANDOM}};
  image_1684 = _RAND_1437[3:0];
  _RAND_1438 = {1{`RANDOM}};
  image_1685 = _RAND_1438[3:0];
  _RAND_1439 = {1{`RANDOM}};
  image_1686 = _RAND_1439[3:0];
  _RAND_1440 = {1{`RANDOM}};
  image_1687 = _RAND_1440[3:0];
  _RAND_1441 = {1{`RANDOM}};
  image_1688 = _RAND_1441[3:0];
  _RAND_1442 = {1{`RANDOM}};
  image_1689 = _RAND_1442[3:0];
  _RAND_1443 = {1{`RANDOM}};
  image_1690 = _RAND_1443[3:0];
  _RAND_1444 = {1{`RANDOM}};
  image_1691 = _RAND_1444[3:0];
  _RAND_1445 = {1{`RANDOM}};
  image_1692 = _RAND_1445[3:0];
  _RAND_1446 = {1{`RANDOM}};
  image_1693 = _RAND_1446[3:0];
  _RAND_1447 = {1{`RANDOM}};
  image_1694 = _RAND_1447[3:0];
  _RAND_1448 = {1{`RANDOM}};
  image_1695 = _RAND_1448[3:0];
  _RAND_1449 = {1{`RANDOM}};
  image_1696 = _RAND_1449[3:0];
  _RAND_1450 = {1{`RANDOM}};
  image_1697 = _RAND_1450[3:0];
  _RAND_1451 = {1{`RANDOM}};
  image_1698 = _RAND_1451[3:0];
  _RAND_1452 = {1{`RANDOM}};
  image_1699 = _RAND_1452[3:0];
  _RAND_1453 = {1{`RANDOM}};
  image_1700 = _RAND_1453[3:0];
  _RAND_1454 = {1{`RANDOM}};
  image_1701 = _RAND_1454[3:0];
  _RAND_1455 = {1{`RANDOM}};
  image_1702 = _RAND_1455[3:0];
  _RAND_1456 = {1{`RANDOM}};
  image_1703 = _RAND_1456[3:0];
  _RAND_1457 = {1{`RANDOM}};
  image_1704 = _RAND_1457[3:0];
  _RAND_1458 = {1{`RANDOM}};
  image_1705 = _RAND_1458[3:0];
  _RAND_1459 = {1{`RANDOM}};
  image_1706 = _RAND_1459[3:0];
  _RAND_1460 = {1{`RANDOM}};
  image_1707 = _RAND_1460[3:0];
  _RAND_1461 = {1{`RANDOM}};
  image_1708 = _RAND_1461[3:0];
  _RAND_1462 = {1{`RANDOM}};
  image_1709 = _RAND_1462[3:0];
  _RAND_1463 = {1{`RANDOM}};
  image_1710 = _RAND_1463[3:0];
  _RAND_1464 = {1{`RANDOM}};
  image_1711 = _RAND_1464[3:0];
  _RAND_1465 = {1{`RANDOM}};
  image_1712 = _RAND_1465[3:0];
  _RAND_1466 = {1{`RANDOM}};
  image_1713 = _RAND_1466[3:0];
  _RAND_1467 = {1{`RANDOM}};
  image_1714 = _RAND_1467[3:0];
  _RAND_1468 = {1{`RANDOM}};
  image_1715 = _RAND_1468[3:0];
  _RAND_1469 = {1{`RANDOM}};
  image_1716 = _RAND_1469[3:0];
  _RAND_1470 = {1{`RANDOM}};
  image_1717 = _RAND_1470[3:0];
  _RAND_1471 = {1{`RANDOM}};
  image_1718 = _RAND_1471[3:0];
  _RAND_1472 = {1{`RANDOM}};
  image_1719 = _RAND_1472[3:0];
  _RAND_1473 = {1{`RANDOM}};
  image_1720 = _RAND_1473[3:0];
  _RAND_1474 = {1{`RANDOM}};
  image_1721 = _RAND_1474[3:0];
  _RAND_1475 = {1{`RANDOM}};
  image_1722 = _RAND_1475[3:0];
  _RAND_1476 = {1{`RANDOM}};
  image_1723 = _RAND_1476[3:0];
  _RAND_1477 = {1{`RANDOM}};
  image_1728 = _RAND_1477[3:0];
  _RAND_1478 = {1{`RANDOM}};
  image_1729 = _RAND_1478[3:0];
  _RAND_1479 = {1{`RANDOM}};
  image_1730 = _RAND_1479[3:0];
  _RAND_1480 = {1{`RANDOM}};
  image_1731 = _RAND_1480[3:0];
  _RAND_1481 = {1{`RANDOM}};
  image_1732 = _RAND_1481[3:0];
  _RAND_1482 = {1{`RANDOM}};
  image_1733 = _RAND_1482[3:0];
  _RAND_1483 = {1{`RANDOM}};
  image_1734 = _RAND_1483[3:0];
  _RAND_1484 = {1{`RANDOM}};
  image_1735 = _RAND_1484[3:0];
  _RAND_1485 = {1{`RANDOM}};
  image_1736 = _RAND_1485[3:0];
  _RAND_1486 = {1{`RANDOM}};
  image_1737 = _RAND_1486[3:0];
  _RAND_1487 = {1{`RANDOM}};
  image_1738 = _RAND_1487[3:0];
  _RAND_1488 = {1{`RANDOM}};
  image_1739 = _RAND_1488[3:0];
  _RAND_1489 = {1{`RANDOM}};
  image_1740 = _RAND_1489[3:0];
  _RAND_1490 = {1{`RANDOM}};
  image_1741 = _RAND_1490[3:0];
  _RAND_1491 = {1{`RANDOM}};
  image_1742 = _RAND_1491[3:0];
  _RAND_1492 = {1{`RANDOM}};
  image_1743 = _RAND_1492[3:0];
  _RAND_1493 = {1{`RANDOM}};
  image_1744 = _RAND_1493[3:0];
  _RAND_1494 = {1{`RANDOM}};
  image_1745 = _RAND_1494[3:0];
  _RAND_1495 = {1{`RANDOM}};
  image_1746 = _RAND_1495[3:0];
  _RAND_1496 = {1{`RANDOM}};
  image_1747 = _RAND_1496[3:0];
  _RAND_1497 = {1{`RANDOM}};
  image_1748 = _RAND_1497[3:0];
  _RAND_1498 = {1{`RANDOM}};
  image_1749 = _RAND_1498[3:0];
  _RAND_1499 = {1{`RANDOM}};
  image_1750 = _RAND_1499[3:0];
  _RAND_1500 = {1{`RANDOM}};
  image_1751 = _RAND_1500[3:0];
  _RAND_1501 = {1{`RANDOM}};
  image_1752 = _RAND_1501[3:0];
  _RAND_1502 = {1{`RANDOM}};
  image_1753 = _RAND_1502[3:0];
  _RAND_1503 = {1{`RANDOM}};
  image_1754 = _RAND_1503[3:0];
  _RAND_1504 = {1{`RANDOM}};
  image_1755 = _RAND_1504[3:0];
  _RAND_1505 = {1{`RANDOM}};
  image_1756 = _RAND_1505[3:0];
  _RAND_1506 = {1{`RANDOM}};
  image_1757 = _RAND_1506[3:0];
  _RAND_1507 = {1{`RANDOM}};
  image_1758 = _RAND_1507[3:0];
  _RAND_1508 = {1{`RANDOM}};
  image_1759 = _RAND_1508[3:0];
  _RAND_1509 = {1{`RANDOM}};
  image_1760 = _RAND_1509[3:0];
  _RAND_1510 = {1{`RANDOM}};
  image_1761 = _RAND_1510[3:0];
  _RAND_1511 = {1{`RANDOM}};
  image_1762 = _RAND_1511[3:0];
  _RAND_1512 = {1{`RANDOM}};
  image_1763 = _RAND_1512[3:0];
  _RAND_1513 = {1{`RANDOM}};
  image_1764 = _RAND_1513[3:0];
  _RAND_1514 = {1{`RANDOM}};
  image_1765 = _RAND_1514[3:0];
  _RAND_1515 = {1{`RANDOM}};
  image_1766 = _RAND_1515[3:0];
  _RAND_1516 = {1{`RANDOM}};
  image_1767 = _RAND_1516[3:0];
  _RAND_1517 = {1{`RANDOM}};
  image_1768 = _RAND_1517[3:0];
  _RAND_1518 = {1{`RANDOM}};
  image_1769 = _RAND_1518[3:0];
  _RAND_1519 = {1{`RANDOM}};
  image_1770 = _RAND_1519[3:0];
  _RAND_1520 = {1{`RANDOM}};
  image_1771 = _RAND_1520[3:0];
  _RAND_1521 = {1{`RANDOM}};
  image_1772 = _RAND_1521[3:0];
  _RAND_1522 = {1{`RANDOM}};
  image_1773 = _RAND_1522[3:0];
  _RAND_1523 = {1{`RANDOM}};
  image_1774 = _RAND_1523[3:0];
  _RAND_1524 = {1{`RANDOM}};
  image_1775 = _RAND_1524[3:0];
  _RAND_1525 = {1{`RANDOM}};
  image_1776 = _RAND_1525[3:0];
  _RAND_1526 = {1{`RANDOM}};
  image_1777 = _RAND_1526[3:0];
  _RAND_1527 = {1{`RANDOM}};
  image_1778 = _RAND_1527[3:0];
  _RAND_1528 = {1{`RANDOM}};
  image_1779 = _RAND_1528[3:0];
  _RAND_1529 = {1{`RANDOM}};
  image_1780 = _RAND_1529[3:0];
  _RAND_1530 = {1{`RANDOM}};
  image_1781 = _RAND_1530[3:0];
  _RAND_1531 = {1{`RANDOM}};
  image_1782 = _RAND_1531[3:0];
  _RAND_1532 = {1{`RANDOM}};
  image_1783 = _RAND_1532[3:0];
  _RAND_1533 = {1{`RANDOM}};
  image_1784 = _RAND_1533[3:0];
  _RAND_1534 = {1{`RANDOM}};
  image_1785 = _RAND_1534[3:0];
  _RAND_1535 = {1{`RANDOM}};
  image_1786 = _RAND_1535[3:0];
  _RAND_1536 = {1{`RANDOM}};
  image_1793 = _RAND_1536[3:0];
  _RAND_1537 = {1{`RANDOM}};
  image_1794 = _RAND_1537[3:0];
  _RAND_1538 = {1{`RANDOM}};
  image_1795 = _RAND_1538[3:0];
  _RAND_1539 = {1{`RANDOM}};
  image_1796 = _RAND_1539[3:0];
  _RAND_1540 = {1{`RANDOM}};
  image_1797 = _RAND_1540[3:0];
  _RAND_1541 = {1{`RANDOM}};
  image_1798 = _RAND_1541[3:0];
  _RAND_1542 = {1{`RANDOM}};
  image_1799 = _RAND_1542[3:0];
  _RAND_1543 = {1{`RANDOM}};
  image_1800 = _RAND_1543[3:0];
  _RAND_1544 = {1{`RANDOM}};
  image_1801 = _RAND_1544[3:0];
  _RAND_1545 = {1{`RANDOM}};
  image_1802 = _RAND_1545[3:0];
  _RAND_1546 = {1{`RANDOM}};
  image_1803 = _RAND_1546[3:0];
  _RAND_1547 = {1{`RANDOM}};
  image_1804 = _RAND_1547[3:0];
  _RAND_1548 = {1{`RANDOM}};
  image_1805 = _RAND_1548[3:0];
  _RAND_1549 = {1{`RANDOM}};
  image_1806 = _RAND_1549[3:0];
  _RAND_1550 = {1{`RANDOM}};
  image_1807 = _RAND_1550[3:0];
  _RAND_1551 = {1{`RANDOM}};
  image_1808 = _RAND_1551[3:0];
  _RAND_1552 = {1{`RANDOM}};
  image_1809 = _RAND_1552[3:0];
  _RAND_1553 = {1{`RANDOM}};
  image_1810 = _RAND_1553[3:0];
  _RAND_1554 = {1{`RANDOM}};
  image_1811 = _RAND_1554[3:0];
  _RAND_1555 = {1{`RANDOM}};
  image_1812 = _RAND_1555[3:0];
  _RAND_1556 = {1{`RANDOM}};
  image_1813 = _RAND_1556[3:0];
  _RAND_1557 = {1{`RANDOM}};
  image_1814 = _RAND_1557[3:0];
  _RAND_1558 = {1{`RANDOM}};
  image_1815 = _RAND_1558[3:0];
  _RAND_1559 = {1{`RANDOM}};
  image_1816 = _RAND_1559[3:0];
  _RAND_1560 = {1{`RANDOM}};
  image_1817 = _RAND_1560[3:0];
  _RAND_1561 = {1{`RANDOM}};
  image_1818 = _RAND_1561[3:0];
  _RAND_1562 = {1{`RANDOM}};
  image_1819 = _RAND_1562[3:0];
  _RAND_1563 = {1{`RANDOM}};
  image_1820 = _RAND_1563[3:0];
  _RAND_1564 = {1{`RANDOM}};
  image_1821 = _RAND_1564[3:0];
  _RAND_1565 = {1{`RANDOM}};
  image_1822 = _RAND_1565[3:0];
  _RAND_1566 = {1{`RANDOM}};
  image_1823 = _RAND_1566[3:0];
  _RAND_1567 = {1{`RANDOM}};
  image_1824 = _RAND_1567[3:0];
  _RAND_1568 = {1{`RANDOM}};
  image_1825 = _RAND_1568[3:0];
  _RAND_1569 = {1{`RANDOM}};
  image_1826 = _RAND_1569[3:0];
  _RAND_1570 = {1{`RANDOM}};
  image_1827 = _RAND_1570[3:0];
  _RAND_1571 = {1{`RANDOM}};
  image_1828 = _RAND_1571[3:0];
  _RAND_1572 = {1{`RANDOM}};
  image_1829 = _RAND_1572[3:0];
  _RAND_1573 = {1{`RANDOM}};
  image_1830 = _RAND_1573[3:0];
  _RAND_1574 = {1{`RANDOM}};
  image_1831 = _RAND_1574[3:0];
  _RAND_1575 = {1{`RANDOM}};
  image_1832 = _RAND_1575[3:0];
  _RAND_1576 = {1{`RANDOM}};
  image_1833 = _RAND_1576[3:0];
  _RAND_1577 = {1{`RANDOM}};
  image_1834 = _RAND_1577[3:0];
  _RAND_1578 = {1{`RANDOM}};
  image_1835 = _RAND_1578[3:0];
  _RAND_1579 = {1{`RANDOM}};
  image_1836 = _RAND_1579[3:0];
  _RAND_1580 = {1{`RANDOM}};
  image_1837 = _RAND_1580[3:0];
  _RAND_1581 = {1{`RANDOM}};
  image_1838 = _RAND_1581[3:0];
  _RAND_1582 = {1{`RANDOM}};
  image_1839 = _RAND_1582[3:0];
  _RAND_1583 = {1{`RANDOM}};
  image_1840 = _RAND_1583[3:0];
  _RAND_1584 = {1{`RANDOM}};
  image_1841 = _RAND_1584[3:0];
  _RAND_1585 = {1{`RANDOM}};
  image_1842 = _RAND_1585[3:0];
  _RAND_1586 = {1{`RANDOM}};
  image_1843 = _RAND_1586[3:0];
  _RAND_1587 = {1{`RANDOM}};
  image_1844 = _RAND_1587[3:0];
  _RAND_1588 = {1{`RANDOM}};
  image_1845 = _RAND_1588[3:0];
  _RAND_1589 = {1{`RANDOM}};
  image_1846 = _RAND_1589[3:0];
  _RAND_1590 = {1{`RANDOM}};
  image_1847 = _RAND_1590[3:0];
  _RAND_1591 = {1{`RANDOM}};
  image_1848 = _RAND_1591[3:0];
  _RAND_1592 = {1{`RANDOM}};
  image_1849 = _RAND_1592[3:0];
  _RAND_1593 = {1{`RANDOM}};
  image_1857 = _RAND_1593[3:0];
  _RAND_1594 = {1{`RANDOM}};
  image_1858 = _RAND_1594[3:0];
  _RAND_1595 = {1{`RANDOM}};
  image_1859 = _RAND_1595[3:0];
  _RAND_1596 = {1{`RANDOM}};
  image_1860 = _RAND_1596[3:0];
  _RAND_1597 = {1{`RANDOM}};
  image_1861 = _RAND_1597[3:0];
  _RAND_1598 = {1{`RANDOM}};
  image_1862 = _RAND_1598[3:0];
  _RAND_1599 = {1{`RANDOM}};
  image_1863 = _RAND_1599[3:0];
  _RAND_1600 = {1{`RANDOM}};
  image_1864 = _RAND_1600[3:0];
  _RAND_1601 = {1{`RANDOM}};
  image_1865 = _RAND_1601[3:0];
  _RAND_1602 = {1{`RANDOM}};
  image_1866 = _RAND_1602[3:0];
  _RAND_1603 = {1{`RANDOM}};
  image_1867 = _RAND_1603[3:0];
  _RAND_1604 = {1{`RANDOM}};
  image_1868 = _RAND_1604[3:0];
  _RAND_1605 = {1{`RANDOM}};
  image_1869 = _RAND_1605[3:0];
  _RAND_1606 = {1{`RANDOM}};
  image_1870 = _RAND_1606[3:0];
  _RAND_1607 = {1{`RANDOM}};
  image_1871 = _RAND_1607[3:0];
  _RAND_1608 = {1{`RANDOM}};
  image_1872 = _RAND_1608[3:0];
  _RAND_1609 = {1{`RANDOM}};
  image_1873 = _RAND_1609[3:0];
  _RAND_1610 = {1{`RANDOM}};
  image_1874 = _RAND_1610[3:0];
  _RAND_1611 = {1{`RANDOM}};
  image_1875 = _RAND_1611[3:0];
  _RAND_1612 = {1{`RANDOM}};
  image_1876 = _RAND_1612[3:0];
  _RAND_1613 = {1{`RANDOM}};
  image_1877 = _RAND_1613[3:0];
  _RAND_1614 = {1{`RANDOM}};
  image_1878 = _RAND_1614[3:0];
  _RAND_1615 = {1{`RANDOM}};
  image_1879 = _RAND_1615[3:0];
  _RAND_1616 = {1{`RANDOM}};
  image_1880 = _RAND_1616[3:0];
  _RAND_1617 = {1{`RANDOM}};
  image_1881 = _RAND_1617[3:0];
  _RAND_1618 = {1{`RANDOM}};
  image_1882 = _RAND_1618[3:0];
  _RAND_1619 = {1{`RANDOM}};
  image_1883 = _RAND_1619[3:0];
  _RAND_1620 = {1{`RANDOM}};
  image_1884 = _RAND_1620[3:0];
  _RAND_1621 = {1{`RANDOM}};
  image_1885 = _RAND_1621[3:0];
  _RAND_1622 = {1{`RANDOM}};
  image_1886 = _RAND_1622[3:0];
  _RAND_1623 = {1{`RANDOM}};
  image_1887 = _RAND_1623[3:0];
  _RAND_1624 = {1{`RANDOM}};
  image_1888 = _RAND_1624[3:0];
  _RAND_1625 = {1{`RANDOM}};
  image_1889 = _RAND_1625[3:0];
  _RAND_1626 = {1{`RANDOM}};
  image_1890 = _RAND_1626[3:0];
  _RAND_1627 = {1{`RANDOM}};
  image_1891 = _RAND_1627[3:0];
  _RAND_1628 = {1{`RANDOM}};
  image_1892 = _RAND_1628[3:0];
  _RAND_1629 = {1{`RANDOM}};
  image_1893 = _RAND_1629[3:0];
  _RAND_1630 = {1{`RANDOM}};
  image_1894 = _RAND_1630[3:0];
  _RAND_1631 = {1{`RANDOM}};
  image_1895 = _RAND_1631[3:0];
  _RAND_1632 = {1{`RANDOM}};
  image_1896 = _RAND_1632[3:0];
  _RAND_1633 = {1{`RANDOM}};
  image_1897 = _RAND_1633[3:0];
  _RAND_1634 = {1{`RANDOM}};
  image_1898 = _RAND_1634[3:0];
  _RAND_1635 = {1{`RANDOM}};
  image_1899 = _RAND_1635[3:0];
  _RAND_1636 = {1{`RANDOM}};
  image_1900 = _RAND_1636[3:0];
  _RAND_1637 = {1{`RANDOM}};
  image_1901 = _RAND_1637[3:0];
  _RAND_1638 = {1{`RANDOM}};
  image_1902 = _RAND_1638[3:0];
  _RAND_1639 = {1{`RANDOM}};
  image_1903 = _RAND_1639[3:0];
  _RAND_1640 = {1{`RANDOM}};
  image_1904 = _RAND_1640[3:0];
  _RAND_1641 = {1{`RANDOM}};
  image_1905 = _RAND_1641[3:0];
  _RAND_1642 = {1{`RANDOM}};
  image_1906 = _RAND_1642[3:0];
  _RAND_1643 = {1{`RANDOM}};
  image_1907 = _RAND_1643[3:0];
  _RAND_1644 = {1{`RANDOM}};
  image_1908 = _RAND_1644[3:0];
  _RAND_1645 = {1{`RANDOM}};
  image_1909 = _RAND_1645[3:0];
  _RAND_1646 = {1{`RANDOM}};
  image_1910 = _RAND_1646[3:0];
  _RAND_1647 = {1{`RANDOM}};
  image_1911 = _RAND_1647[3:0];
  _RAND_1648 = {1{`RANDOM}};
  image_1912 = _RAND_1648[3:0];
  _RAND_1649 = {1{`RANDOM}};
  image_1913 = _RAND_1649[3:0];
  _RAND_1650 = {1{`RANDOM}};
  image_1921 = _RAND_1650[3:0];
  _RAND_1651 = {1{`RANDOM}};
  image_1922 = _RAND_1651[3:0];
  _RAND_1652 = {1{`RANDOM}};
  image_1923 = _RAND_1652[3:0];
  _RAND_1653 = {1{`RANDOM}};
  image_1924 = _RAND_1653[3:0];
  _RAND_1654 = {1{`RANDOM}};
  image_1925 = _RAND_1654[3:0];
  _RAND_1655 = {1{`RANDOM}};
  image_1926 = _RAND_1655[3:0];
  _RAND_1656 = {1{`RANDOM}};
  image_1927 = _RAND_1656[3:0];
  _RAND_1657 = {1{`RANDOM}};
  image_1928 = _RAND_1657[3:0];
  _RAND_1658 = {1{`RANDOM}};
  image_1929 = _RAND_1658[3:0];
  _RAND_1659 = {1{`RANDOM}};
  image_1930 = _RAND_1659[3:0];
  _RAND_1660 = {1{`RANDOM}};
  image_1931 = _RAND_1660[3:0];
  _RAND_1661 = {1{`RANDOM}};
  image_1932 = _RAND_1661[3:0];
  _RAND_1662 = {1{`RANDOM}};
  image_1933 = _RAND_1662[3:0];
  _RAND_1663 = {1{`RANDOM}};
  image_1934 = _RAND_1663[3:0];
  _RAND_1664 = {1{`RANDOM}};
  image_1935 = _RAND_1664[3:0];
  _RAND_1665 = {1{`RANDOM}};
  image_1936 = _RAND_1665[3:0];
  _RAND_1666 = {1{`RANDOM}};
  image_1937 = _RAND_1666[3:0];
  _RAND_1667 = {1{`RANDOM}};
  image_1938 = _RAND_1667[3:0];
  _RAND_1668 = {1{`RANDOM}};
  image_1939 = _RAND_1668[3:0];
  _RAND_1669 = {1{`RANDOM}};
  image_1940 = _RAND_1669[3:0];
  _RAND_1670 = {1{`RANDOM}};
  image_1941 = _RAND_1670[3:0];
  _RAND_1671 = {1{`RANDOM}};
  image_1942 = _RAND_1671[3:0];
  _RAND_1672 = {1{`RANDOM}};
  image_1943 = _RAND_1672[3:0];
  _RAND_1673 = {1{`RANDOM}};
  image_1944 = _RAND_1673[3:0];
  _RAND_1674 = {1{`RANDOM}};
  image_1945 = _RAND_1674[3:0];
  _RAND_1675 = {1{`RANDOM}};
  image_1946 = _RAND_1675[3:0];
  _RAND_1676 = {1{`RANDOM}};
  image_1947 = _RAND_1676[3:0];
  _RAND_1677 = {1{`RANDOM}};
  image_1948 = _RAND_1677[3:0];
  _RAND_1678 = {1{`RANDOM}};
  image_1949 = _RAND_1678[3:0];
  _RAND_1679 = {1{`RANDOM}};
  image_1950 = _RAND_1679[3:0];
  _RAND_1680 = {1{`RANDOM}};
  image_1951 = _RAND_1680[3:0];
  _RAND_1681 = {1{`RANDOM}};
  image_1952 = _RAND_1681[3:0];
  _RAND_1682 = {1{`RANDOM}};
  image_1953 = _RAND_1682[3:0];
  _RAND_1683 = {1{`RANDOM}};
  image_1954 = _RAND_1683[3:0];
  _RAND_1684 = {1{`RANDOM}};
  image_1955 = _RAND_1684[3:0];
  _RAND_1685 = {1{`RANDOM}};
  image_1956 = _RAND_1685[3:0];
  _RAND_1686 = {1{`RANDOM}};
  image_1957 = _RAND_1686[3:0];
  _RAND_1687 = {1{`RANDOM}};
  image_1958 = _RAND_1687[3:0];
  _RAND_1688 = {1{`RANDOM}};
  image_1959 = _RAND_1688[3:0];
  _RAND_1689 = {1{`RANDOM}};
  image_1960 = _RAND_1689[3:0];
  _RAND_1690 = {1{`RANDOM}};
  image_1961 = _RAND_1690[3:0];
  _RAND_1691 = {1{`RANDOM}};
  image_1962 = _RAND_1691[3:0];
  _RAND_1692 = {1{`RANDOM}};
  image_1963 = _RAND_1692[3:0];
  _RAND_1693 = {1{`RANDOM}};
  image_1964 = _RAND_1693[3:0];
  _RAND_1694 = {1{`RANDOM}};
  image_1965 = _RAND_1694[3:0];
  _RAND_1695 = {1{`RANDOM}};
  image_1966 = _RAND_1695[3:0];
  _RAND_1696 = {1{`RANDOM}};
  image_1967 = _RAND_1696[3:0];
  _RAND_1697 = {1{`RANDOM}};
  image_1968 = _RAND_1697[3:0];
  _RAND_1698 = {1{`RANDOM}};
  image_1969 = _RAND_1698[3:0];
  _RAND_1699 = {1{`RANDOM}};
  image_1970 = _RAND_1699[3:0];
  _RAND_1700 = {1{`RANDOM}};
  image_1971 = _RAND_1700[3:0];
  _RAND_1701 = {1{`RANDOM}};
  image_1972 = _RAND_1701[3:0];
  _RAND_1702 = {1{`RANDOM}};
  image_1973 = _RAND_1702[3:0];
  _RAND_1703 = {1{`RANDOM}};
  image_1974 = _RAND_1703[3:0];
  _RAND_1704 = {1{`RANDOM}};
  image_1975 = _RAND_1704[3:0];
  _RAND_1705 = {1{`RANDOM}};
  image_1976 = _RAND_1705[3:0];
  _RAND_1706 = {1{`RANDOM}};
  image_1977 = _RAND_1706[3:0];
  _RAND_1707 = {1{`RANDOM}};
  image_1985 = _RAND_1707[3:0];
  _RAND_1708 = {1{`RANDOM}};
  image_1986 = _RAND_1708[3:0];
  _RAND_1709 = {1{`RANDOM}};
  image_1987 = _RAND_1709[3:0];
  _RAND_1710 = {1{`RANDOM}};
  image_1988 = _RAND_1710[3:0];
  _RAND_1711 = {1{`RANDOM}};
  image_1989 = _RAND_1711[3:0];
  _RAND_1712 = {1{`RANDOM}};
  image_1990 = _RAND_1712[3:0];
  _RAND_1713 = {1{`RANDOM}};
  image_1991 = _RAND_1713[3:0];
  _RAND_1714 = {1{`RANDOM}};
  image_1992 = _RAND_1714[3:0];
  _RAND_1715 = {1{`RANDOM}};
  image_1993 = _RAND_1715[3:0];
  _RAND_1716 = {1{`RANDOM}};
  image_1994 = _RAND_1716[3:0];
  _RAND_1717 = {1{`RANDOM}};
  image_1995 = _RAND_1717[3:0];
  _RAND_1718 = {1{`RANDOM}};
  image_1996 = _RAND_1718[3:0];
  _RAND_1719 = {1{`RANDOM}};
  image_1997 = _RAND_1719[3:0];
  _RAND_1720 = {1{`RANDOM}};
  image_1998 = _RAND_1720[3:0];
  _RAND_1721 = {1{`RANDOM}};
  image_1999 = _RAND_1721[3:0];
  _RAND_1722 = {1{`RANDOM}};
  image_2000 = _RAND_1722[3:0];
  _RAND_1723 = {1{`RANDOM}};
  image_2001 = _RAND_1723[3:0];
  _RAND_1724 = {1{`RANDOM}};
  image_2002 = _RAND_1724[3:0];
  _RAND_1725 = {1{`RANDOM}};
  image_2003 = _RAND_1725[3:0];
  _RAND_1726 = {1{`RANDOM}};
  image_2004 = _RAND_1726[3:0];
  _RAND_1727 = {1{`RANDOM}};
  image_2005 = _RAND_1727[3:0];
  _RAND_1728 = {1{`RANDOM}};
  image_2006 = _RAND_1728[3:0];
  _RAND_1729 = {1{`RANDOM}};
  image_2007 = _RAND_1729[3:0];
  _RAND_1730 = {1{`RANDOM}};
  image_2008 = _RAND_1730[3:0];
  _RAND_1731 = {1{`RANDOM}};
  image_2009 = _RAND_1731[3:0];
  _RAND_1732 = {1{`RANDOM}};
  image_2010 = _RAND_1732[3:0];
  _RAND_1733 = {1{`RANDOM}};
  image_2011 = _RAND_1733[3:0];
  _RAND_1734 = {1{`RANDOM}};
  image_2012 = _RAND_1734[3:0];
  _RAND_1735 = {1{`RANDOM}};
  image_2013 = _RAND_1735[3:0];
  _RAND_1736 = {1{`RANDOM}};
  image_2014 = _RAND_1736[3:0];
  _RAND_1737 = {1{`RANDOM}};
  image_2015 = _RAND_1737[3:0];
  _RAND_1738 = {1{`RANDOM}};
  image_2016 = _RAND_1738[3:0];
  _RAND_1739 = {1{`RANDOM}};
  image_2017 = _RAND_1739[3:0];
  _RAND_1740 = {1{`RANDOM}};
  image_2018 = _RAND_1740[3:0];
  _RAND_1741 = {1{`RANDOM}};
  image_2019 = _RAND_1741[3:0];
  _RAND_1742 = {1{`RANDOM}};
  image_2020 = _RAND_1742[3:0];
  _RAND_1743 = {1{`RANDOM}};
  image_2021 = _RAND_1743[3:0];
  _RAND_1744 = {1{`RANDOM}};
  image_2022 = _RAND_1744[3:0];
  _RAND_1745 = {1{`RANDOM}};
  image_2023 = _RAND_1745[3:0];
  _RAND_1746 = {1{`RANDOM}};
  image_2024 = _RAND_1746[3:0];
  _RAND_1747 = {1{`RANDOM}};
  image_2025 = _RAND_1747[3:0];
  _RAND_1748 = {1{`RANDOM}};
  image_2026 = _RAND_1748[3:0];
  _RAND_1749 = {1{`RANDOM}};
  image_2027 = _RAND_1749[3:0];
  _RAND_1750 = {1{`RANDOM}};
  image_2028 = _RAND_1750[3:0];
  _RAND_1751 = {1{`RANDOM}};
  image_2029 = _RAND_1751[3:0];
  _RAND_1752 = {1{`RANDOM}};
  image_2030 = _RAND_1752[3:0];
  _RAND_1753 = {1{`RANDOM}};
  image_2031 = _RAND_1753[3:0];
  _RAND_1754 = {1{`RANDOM}};
  image_2032 = _RAND_1754[3:0];
  _RAND_1755 = {1{`RANDOM}};
  image_2033 = _RAND_1755[3:0];
  _RAND_1756 = {1{`RANDOM}};
  image_2034 = _RAND_1756[3:0];
  _RAND_1757 = {1{`RANDOM}};
  image_2035 = _RAND_1757[3:0];
  _RAND_1758 = {1{`RANDOM}};
  image_2036 = _RAND_1758[3:0];
  _RAND_1759 = {1{`RANDOM}};
  image_2037 = _RAND_1759[3:0];
  _RAND_1760 = {1{`RANDOM}};
  image_2038 = _RAND_1760[3:0];
  _RAND_1761 = {1{`RANDOM}};
  image_2039 = _RAND_1761[3:0];
  _RAND_1762 = {1{`RANDOM}};
  image_2040 = _RAND_1762[3:0];
  _RAND_1763 = {1{`RANDOM}};
  image_2041 = _RAND_1763[3:0];
  _RAND_1764 = {1{`RANDOM}};
  image_2049 = _RAND_1764[3:0];
  _RAND_1765 = {1{`RANDOM}};
  image_2050 = _RAND_1765[3:0];
  _RAND_1766 = {1{`RANDOM}};
  image_2051 = _RAND_1766[3:0];
  _RAND_1767 = {1{`RANDOM}};
  image_2052 = _RAND_1767[3:0];
  _RAND_1768 = {1{`RANDOM}};
  image_2053 = _RAND_1768[3:0];
  _RAND_1769 = {1{`RANDOM}};
  image_2054 = _RAND_1769[3:0];
  _RAND_1770 = {1{`RANDOM}};
  image_2055 = _RAND_1770[3:0];
  _RAND_1771 = {1{`RANDOM}};
  image_2056 = _RAND_1771[3:0];
  _RAND_1772 = {1{`RANDOM}};
  image_2057 = _RAND_1772[3:0];
  _RAND_1773 = {1{`RANDOM}};
  image_2058 = _RAND_1773[3:0];
  _RAND_1774 = {1{`RANDOM}};
  image_2059 = _RAND_1774[3:0];
  _RAND_1775 = {1{`RANDOM}};
  image_2060 = _RAND_1775[3:0];
  _RAND_1776 = {1{`RANDOM}};
  image_2061 = _RAND_1776[3:0];
  _RAND_1777 = {1{`RANDOM}};
  image_2062 = _RAND_1777[3:0];
  _RAND_1778 = {1{`RANDOM}};
  image_2063 = _RAND_1778[3:0];
  _RAND_1779 = {1{`RANDOM}};
  image_2064 = _RAND_1779[3:0];
  _RAND_1780 = {1{`RANDOM}};
  image_2065 = _RAND_1780[3:0];
  _RAND_1781 = {1{`RANDOM}};
  image_2066 = _RAND_1781[3:0];
  _RAND_1782 = {1{`RANDOM}};
  image_2067 = _RAND_1782[3:0];
  _RAND_1783 = {1{`RANDOM}};
  image_2068 = _RAND_1783[3:0];
  _RAND_1784 = {1{`RANDOM}};
  image_2069 = _RAND_1784[3:0];
  _RAND_1785 = {1{`RANDOM}};
  image_2070 = _RAND_1785[3:0];
  _RAND_1786 = {1{`RANDOM}};
  image_2071 = _RAND_1786[3:0];
  _RAND_1787 = {1{`RANDOM}};
  image_2072 = _RAND_1787[3:0];
  _RAND_1788 = {1{`RANDOM}};
  image_2073 = _RAND_1788[3:0];
  _RAND_1789 = {1{`RANDOM}};
  image_2074 = _RAND_1789[3:0];
  _RAND_1790 = {1{`RANDOM}};
  image_2075 = _RAND_1790[3:0];
  _RAND_1791 = {1{`RANDOM}};
  image_2076 = _RAND_1791[3:0];
  _RAND_1792 = {1{`RANDOM}};
  image_2077 = _RAND_1792[3:0];
  _RAND_1793 = {1{`RANDOM}};
  image_2078 = _RAND_1793[3:0];
  _RAND_1794 = {1{`RANDOM}};
  image_2079 = _RAND_1794[3:0];
  _RAND_1795 = {1{`RANDOM}};
  image_2080 = _RAND_1795[3:0];
  _RAND_1796 = {1{`RANDOM}};
  image_2081 = _RAND_1796[3:0];
  _RAND_1797 = {1{`RANDOM}};
  image_2082 = _RAND_1797[3:0];
  _RAND_1798 = {1{`RANDOM}};
  image_2083 = _RAND_1798[3:0];
  _RAND_1799 = {1{`RANDOM}};
  image_2084 = _RAND_1799[3:0];
  _RAND_1800 = {1{`RANDOM}};
  image_2085 = _RAND_1800[3:0];
  _RAND_1801 = {1{`RANDOM}};
  image_2086 = _RAND_1801[3:0];
  _RAND_1802 = {1{`RANDOM}};
  image_2087 = _RAND_1802[3:0];
  _RAND_1803 = {1{`RANDOM}};
  image_2088 = _RAND_1803[3:0];
  _RAND_1804 = {1{`RANDOM}};
  image_2089 = _RAND_1804[3:0];
  _RAND_1805 = {1{`RANDOM}};
  image_2090 = _RAND_1805[3:0];
  _RAND_1806 = {1{`RANDOM}};
  image_2091 = _RAND_1806[3:0];
  _RAND_1807 = {1{`RANDOM}};
  image_2092 = _RAND_1807[3:0];
  _RAND_1808 = {1{`RANDOM}};
  image_2093 = _RAND_1808[3:0];
  _RAND_1809 = {1{`RANDOM}};
  image_2094 = _RAND_1809[3:0];
  _RAND_1810 = {1{`RANDOM}};
  image_2095 = _RAND_1810[3:0];
  _RAND_1811 = {1{`RANDOM}};
  image_2096 = _RAND_1811[3:0];
  _RAND_1812 = {1{`RANDOM}};
  image_2097 = _RAND_1812[3:0];
  _RAND_1813 = {1{`RANDOM}};
  image_2098 = _RAND_1813[3:0];
  _RAND_1814 = {1{`RANDOM}};
  image_2099 = _RAND_1814[3:0];
  _RAND_1815 = {1{`RANDOM}};
  image_2100 = _RAND_1815[3:0];
  _RAND_1816 = {1{`RANDOM}};
  image_2101 = _RAND_1816[3:0];
  _RAND_1817 = {1{`RANDOM}};
  image_2102 = _RAND_1817[3:0];
  _RAND_1818 = {1{`RANDOM}};
  image_2103 = _RAND_1818[3:0];
  _RAND_1819 = {1{`RANDOM}};
  image_2104 = _RAND_1819[3:0];
  _RAND_1820 = {1{`RANDOM}};
  image_2105 = _RAND_1820[3:0];
  _RAND_1821 = {1{`RANDOM}};
  image_2106 = _RAND_1821[3:0];
  _RAND_1822 = {1{`RANDOM}};
  image_2114 = _RAND_1822[3:0];
  _RAND_1823 = {1{`RANDOM}};
  image_2115 = _RAND_1823[3:0];
  _RAND_1824 = {1{`RANDOM}};
  image_2116 = _RAND_1824[3:0];
  _RAND_1825 = {1{`RANDOM}};
  image_2117 = _RAND_1825[3:0];
  _RAND_1826 = {1{`RANDOM}};
  image_2118 = _RAND_1826[3:0];
  _RAND_1827 = {1{`RANDOM}};
  image_2119 = _RAND_1827[3:0];
  _RAND_1828 = {1{`RANDOM}};
  image_2120 = _RAND_1828[3:0];
  _RAND_1829 = {1{`RANDOM}};
  image_2121 = _RAND_1829[3:0];
  _RAND_1830 = {1{`RANDOM}};
  image_2122 = _RAND_1830[3:0];
  _RAND_1831 = {1{`RANDOM}};
  image_2123 = _RAND_1831[3:0];
  _RAND_1832 = {1{`RANDOM}};
  image_2124 = _RAND_1832[3:0];
  _RAND_1833 = {1{`RANDOM}};
  image_2125 = _RAND_1833[3:0];
  _RAND_1834 = {1{`RANDOM}};
  image_2126 = _RAND_1834[3:0];
  _RAND_1835 = {1{`RANDOM}};
  image_2127 = _RAND_1835[3:0];
  _RAND_1836 = {1{`RANDOM}};
  image_2128 = _RAND_1836[3:0];
  _RAND_1837 = {1{`RANDOM}};
  image_2129 = _RAND_1837[3:0];
  _RAND_1838 = {1{`RANDOM}};
  image_2130 = _RAND_1838[3:0];
  _RAND_1839 = {1{`RANDOM}};
  image_2131 = _RAND_1839[3:0];
  _RAND_1840 = {1{`RANDOM}};
  image_2132 = _RAND_1840[3:0];
  _RAND_1841 = {1{`RANDOM}};
  image_2133 = _RAND_1841[3:0];
  _RAND_1842 = {1{`RANDOM}};
  image_2134 = _RAND_1842[3:0];
  _RAND_1843 = {1{`RANDOM}};
  image_2135 = _RAND_1843[3:0];
  _RAND_1844 = {1{`RANDOM}};
  image_2136 = _RAND_1844[3:0];
  _RAND_1845 = {1{`RANDOM}};
  image_2137 = _RAND_1845[3:0];
  _RAND_1846 = {1{`RANDOM}};
  image_2138 = _RAND_1846[3:0];
  _RAND_1847 = {1{`RANDOM}};
  image_2139 = _RAND_1847[3:0];
  _RAND_1848 = {1{`RANDOM}};
  image_2140 = _RAND_1848[3:0];
  _RAND_1849 = {1{`RANDOM}};
  image_2141 = _RAND_1849[3:0];
  _RAND_1850 = {1{`RANDOM}};
  image_2142 = _RAND_1850[3:0];
  _RAND_1851 = {1{`RANDOM}};
  image_2143 = _RAND_1851[3:0];
  _RAND_1852 = {1{`RANDOM}};
  image_2144 = _RAND_1852[3:0];
  _RAND_1853 = {1{`RANDOM}};
  image_2145 = _RAND_1853[3:0];
  _RAND_1854 = {1{`RANDOM}};
  image_2146 = _RAND_1854[3:0];
  _RAND_1855 = {1{`RANDOM}};
  image_2147 = _RAND_1855[3:0];
  _RAND_1856 = {1{`RANDOM}};
  image_2148 = _RAND_1856[3:0];
  _RAND_1857 = {1{`RANDOM}};
  image_2149 = _RAND_1857[3:0];
  _RAND_1858 = {1{`RANDOM}};
  image_2150 = _RAND_1858[3:0];
  _RAND_1859 = {1{`RANDOM}};
  image_2151 = _RAND_1859[3:0];
  _RAND_1860 = {1{`RANDOM}};
  image_2152 = _RAND_1860[3:0];
  _RAND_1861 = {1{`RANDOM}};
  image_2153 = _RAND_1861[3:0];
  _RAND_1862 = {1{`RANDOM}};
  image_2154 = _RAND_1862[3:0];
  _RAND_1863 = {1{`RANDOM}};
  image_2155 = _RAND_1863[3:0];
  _RAND_1864 = {1{`RANDOM}};
  image_2156 = _RAND_1864[3:0];
  _RAND_1865 = {1{`RANDOM}};
  image_2157 = _RAND_1865[3:0];
  _RAND_1866 = {1{`RANDOM}};
  image_2158 = _RAND_1866[3:0];
  _RAND_1867 = {1{`RANDOM}};
  image_2159 = _RAND_1867[3:0];
  _RAND_1868 = {1{`RANDOM}};
  image_2160 = _RAND_1868[3:0];
  _RAND_1869 = {1{`RANDOM}};
  image_2161 = _RAND_1869[3:0];
  _RAND_1870 = {1{`RANDOM}};
  image_2162 = _RAND_1870[3:0];
  _RAND_1871 = {1{`RANDOM}};
  image_2163 = _RAND_1871[3:0];
  _RAND_1872 = {1{`RANDOM}};
  image_2164 = _RAND_1872[3:0];
  _RAND_1873 = {1{`RANDOM}};
  image_2165 = _RAND_1873[3:0];
  _RAND_1874 = {1{`RANDOM}};
  image_2166 = _RAND_1874[3:0];
  _RAND_1875 = {1{`RANDOM}};
  image_2167 = _RAND_1875[3:0];
  _RAND_1876 = {1{`RANDOM}};
  image_2168 = _RAND_1876[3:0];
  _RAND_1877 = {1{`RANDOM}};
  image_2169 = _RAND_1877[3:0];
  _RAND_1878 = {1{`RANDOM}};
  image_2170 = _RAND_1878[3:0];
  _RAND_1879 = {1{`RANDOM}};
  image_2177 = _RAND_1879[3:0];
  _RAND_1880 = {1{`RANDOM}};
  image_2178 = _RAND_1880[3:0];
  _RAND_1881 = {1{`RANDOM}};
  image_2179 = _RAND_1881[3:0];
  _RAND_1882 = {1{`RANDOM}};
  image_2180 = _RAND_1882[3:0];
  _RAND_1883 = {1{`RANDOM}};
  image_2181 = _RAND_1883[3:0];
  _RAND_1884 = {1{`RANDOM}};
  image_2182 = _RAND_1884[3:0];
  _RAND_1885 = {1{`RANDOM}};
  image_2183 = _RAND_1885[3:0];
  _RAND_1886 = {1{`RANDOM}};
  image_2184 = _RAND_1886[3:0];
  _RAND_1887 = {1{`RANDOM}};
  image_2185 = _RAND_1887[3:0];
  _RAND_1888 = {1{`RANDOM}};
  image_2186 = _RAND_1888[3:0];
  _RAND_1889 = {1{`RANDOM}};
  image_2187 = _RAND_1889[3:0];
  _RAND_1890 = {1{`RANDOM}};
  image_2188 = _RAND_1890[3:0];
  _RAND_1891 = {1{`RANDOM}};
  image_2189 = _RAND_1891[3:0];
  _RAND_1892 = {1{`RANDOM}};
  image_2190 = _RAND_1892[3:0];
  _RAND_1893 = {1{`RANDOM}};
  image_2191 = _RAND_1893[3:0];
  _RAND_1894 = {1{`RANDOM}};
  image_2192 = _RAND_1894[3:0];
  _RAND_1895 = {1{`RANDOM}};
  image_2193 = _RAND_1895[3:0];
  _RAND_1896 = {1{`RANDOM}};
  image_2194 = _RAND_1896[3:0];
  _RAND_1897 = {1{`RANDOM}};
  image_2195 = _RAND_1897[3:0];
  _RAND_1898 = {1{`RANDOM}};
  image_2196 = _RAND_1898[3:0];
  _RAND_1899 = {1{`RANDOM}};
  image_2197 = _RAND_1899[3:0];
  _RAND_1900 = {1{`RANDOM}};
  image_2198 = _RAND_1900[3:0];
  _RAND_1901 = {1{`RANDOM}};
  image_2199 = _RAND_1901[3:0];
  _RAND_1902 = {1{`RANDOM}};
  image_2200 = _RAND_1902[3:0];
  _RAND_1903 = {1{`RANDOM}};
  image_2201 = _RAND_1903[3:0];
  _RAND_1904 = {1{`RANDOM}};
  image_2202 = _RAND_1904[3:0];
  _RAND_1905 = {1{`RANDOM}};
  image_2203 = _RAND_1905[3:0];
  _RAND_1906 = {1{`RANDOM}};
  image_2204 = _RAND_1906[3:0];
  _RAND_1907 = {1{`RANDOM}};
  image_2205 = _RAND_1907[3:0];
  _RAND_1908 = {1{`RANDOM}};
  image_2206 = _RAND_1908[3:0];
  _RAND_1909 = {1{`RANDOM}};
  image_2207 = _RAND_1909[3:0];
  _RAND_1910 = {1{`RANDOM}};
  image_2208 = _RAND_1910[3:0];
  _RAND_1911 = {1{`RANDOM}};
  image_2209 = _RAND_1911[3:0];
  _RAND_1912 = {1{`RANDOM}};
  image_2210 = _RAND_1912[3:0];
  _RAND_1913 = {1{`RANDOM}};
  image_2211 = _RAND_1913[3:0];
  _RAND_1914 = {1{`RANDOM}};
  image_2212 = _RAND_1914[3:0];
  _RAND_1915 = {1{`RANDOM}};
  image_2213 = _RAND_1915[3:0];
  _RAND_1916 = {1{`RANDOM}};
  image_2214 = _RAND_1916[3:0];
  _RAND_1917 = {1{`RANDOM}};
  image_2215 = _RAND_1917[3:0];
  _RAND_1918 = {1{`RANDOM}};
  image_2216 = _RAND_1918[3:0];
  _RAND_1919 = {1{`RANDOM}};
  image_2217 = _RAND_1919[3:0];
  _RAND_1920 = {1{`RANDOM}};
  image_2218 = _RAND_1920[3:0];
  _RAND_1921 = {1{`RANDOM}};
  image_2219 = _RAND_1921[3:0];
  _RAND_1922 = {1{`RANDOM}};
  image_2220 = _RAND_1922[3:0];
  _RAND_1923 = {1{`RANDOM}};
  image_2221 = _RAND_1923[3:0];
  _RAND_1924 = {1{`RANDOM}};
  image_2222 = _RAND_1924[3:0];
  _RAND_1925 = {1{`RANDOM}};
  image_2223 = _RAND_1925[3:0];
  _RAND_1926 = {1{`RANDOM}};
  image_2224 = _RAND_1926[3:0];
  _RAND_1927 = {1{`RANDOM}};
  image_2225 = _RAND_1927[3:0];
  _RAND_1928 = {1{`RANDOM}};
  image_2226 = _RAND_1928[3:0];
  _RAND_1929 = {1{`RANDOM}};
  image_2227 = _RAND_1929[3:0];
  _RAND_1930 = {1{`RANDOM}};
  image_2228 = _RAND_1930[3:0];
  _RAND_1931 = {1{`RANDOM}};
  image_2229 = _RAND_1931[3:0];
  _RAND_1932 = {1{`RANDOM}};
  image_2230 = _RAND_1932[3:0];
  _RAND_1933 = {1{`RANDOM}};
  image_2231 = _RAND_1933[3:0];
  _RAND_1934 = {1{`RANDOM}};
  image_2232 = _RAND_1934[3:0];
  _RAND_1935 = {1{`RANDOM}};
  image_2233 = _RAND_1935[3:0];
  _RAND_1936 = {1{`RANDOM}};
  image_2234 = _RAND_1936[3:0];
  _RAND_1937 = {1{`RANDOM}};
  image_2243 = _RAND_1937[3:0];
  _RAND_1938 = {1{`RANDOM}};
  image_2244 = _RAND_1938[3:0];
  _RAND_1939 = {1{`RANDOM}};
  image_2245 = _RAND_1939[3:0];
  _RAND_1940 = {1{`RANDOM}};
  image_2246 = _RAND_1940[3:0];
  _RAND_1941 = {1{`RANDOM}};
  image_2247 = _RAND_1941[3:0];
  _RAND_1942 = {1{`RANDOM}};
  image_2248 = _RAND_1942[3:0];
  _RAND_1943 = {1{`RANDOM}};
  image_2249 = _RAND_1943[3:0];
  _RAND_1944 = {1{`RANDOM}};
  image_2250 = _RAND_1944[3:0];
  _RAND_1945 = {1{`RANDOM}};
  image_2251 = _RAND_1945[3:0];
  _RAND_1946 = {1{`RANDOM}};
  image_2252 = _RAND_1946[3:0];
  _RAND_1947 = {1{`RANDOM}};
  image_2253 = _RAND_1947[3:0];
  _RAND_1948 = {1{`RANDOM}};
  image_2254 = _RAND_1948[3:0];
  _RAND_1949 = {1{`RANDOM}};
  image_2255 = _RAND_1949[3:0];
  _RAND_1950 = {1{`RANDOM}};
  image_2256 = _RAND_1950[3:0];
  _RAND_1951 = {1{`RANDOM}};
  image_2257 = _RAND_1951[3:0];
  _RAND_1952 = {1{`RANDOM}};
  image_2258 = _RAND_1952[3:0];
  _RAND_1953 = {1{`RANDOM}};
  image_2259 = _RAND_1953[3:0];
  _RAND_1954 = {1{`RANDOM}};
  image_2260 = _RAND_1954[3:0];
  _RAND_1955 = {1{`RANDOM}};
  image_2261 = _RAND_1955[3:0];
  _RAND_1956 = {1{`RANDOM}};
  image_2262 = _RAND_1956[3:0];
  _RAND_1957 = {1{`RANDOM}};
  image_2263 = _RAND_1957[3:0];
  _RAND_1958 = {1{`RANDOM}};
  image_2264 = _RAND_1958[3:0];
  _RAND_1959 = {1{`RANDOM}};
  image_2265 = _RAND_1959[3:0];
  _RAND_1960 = {1{`RANDOM}};
  image_2266 = _RAND_1960[3:0];
  _RAND_1961 = {1{`RANDOM}};
  image_2267 = _RAND_1961[3:0];
  _RAND_1962 = {1{`RANDOM}};
  image_2268 = _RAND_1962[3:0];
  _RAND_1963 = {1{`RANDOM}};
  image_2269 = _RAND_1963[3:0];
  _RAND_1964 = {1{`RANDOM}};
  image_2270 = _RAND_1964[3:0];
  _RAND_1965 = {1{`RANDOM}};
  image_2271 = _RAND_1965[3:0];
  _RAND_1966 = {1{`RANDOM}};
  image_2272 = _RAND_1966[3:0];
  _RAND_1967 = {1{`RANDOM}};
  image_2273 = _RAND_1967[3:0];
  _RAND_1968 = {1{`RANDOM}};
  image_2274 = _RAND_1968[3:0];
  _RAND_1969 = {1{`RANDOM}};
  image_2275 = _RAND_1969[3:0];
  _RAND_1970 = {1{`RANDOM}};
  image_2276 = _RAND_1970[3:0];
  _RAND_1971 = {1{`RANDOM}};
  image_2277 = _RAND_1971[3:0];
  _RAND_1972 = {1{`RANDOM}};
  image_2278 = _RAND_1972[3:0];
  _RAND_1973 = {1{`RANDOM}};
  image_2279 = _RAND_1973[3:0];
  _RAND_1974 = {1{`RANDOM}};
  image_2280 = _RAND_1974[3:0];
  _RAND_1975 = {1{`RANDOM}};
  image_2281 = _RAND_1975[3:0];
  _RAND_1976 = {1{`RANDOM}};
  image_2282 = _RAND_1976[3:0];
  _RAND_1977 = {1{`RANDOM}};
  image_2283 = _RAND_1977[3:0];
  _RAND_1978 = {1{`RANDOM}};
  image_2284 = _RAND_1978[3:0];
  _RAND_1979 = {1{`RANDOM}};
  image_2285 = _RAND_1979[3:0];
  _RAND_1980 = {1{`RANDOM}};
  image_2286 = _RAND_1980[3:0];
  _RAND_1981 = {1{`RANDOM}};
  image_2287 = _RAND_1981[3:0];
  _RAND_1982 = {1{`RANDOM}};
  image_2288 = _RAND_1982[3:0];
  _RAND_1983 = {1{`RANDOM}};
  image_2289 = _RAND_1983[3:0];
  _RAND_1984 = {1{`RANDOM}};
  image_2290 = _RAND_1984[3:0];
  _RAND_1985 = {1{`RANDOM}};
  image_2291 = _RAND_1985[3:0];
  _RAND_1986 = {1{`RANDOM}};
  image_2292 = _RAND_1986[3:0];
  _RAND_1987 = {1{`RANDOM}};
  image_2293 = _RAND_1987[3:0];
  _RAND_1988 = {1{`RANDOM}};
  image_2294 = _RAND_1988[3:0];
  _RAND_1989 = {1{`RANDOM}};
  image_2295 = _RAND_1989[3:0];
  _RAND_1990 = {1{`RANDOM}};
  image_2296 = _RAND_1990[3:0];
  _RAND_1991 = {1{`RANDOM}};
  image_2297 = _RAND_1991[3:0];
  _RAND_1992 = {1{`RANDOM}};
  image_2298 = _RAND_1992[3:0];
  _RAND_1993 = {1{`RANDOM}};
  image_2307 = _RAND_1993[3:0];
  _RAND_1994 = {1{`RANDOM}};
  image_2308 = _RAND_1994[3:0];
  _RAND_1995 = {1{`RANDOM}};
  image_2309 = _RAND_1995[3:0];
  _RAND_1996 = {1{`RANDOM}};
  image_2310 = _RAND_1996[3:0];
  _RAND_1997 = {1{`RANDOM}};
  image_2311 = _RAND_1997[3:0];
  _RAND_1998 = {1{`RANDOM}};
  image_2312 = _RAND_1998[3:0];
  _RAND_1999 = {1{`RANDOM}};
  image_2313 = _RAND_1999[3:0];
  _RAND_2000 = {1{`RANDOM}};
  image_2314 = _RAND_2000[3:0];
  _RAND_2001 = {1{`RANDOM}};
  image_2315 = _RAND_2001[3:0];
  _RAND_2002 = {1{`RANDOM}};
  image_2316 = _RAND_2002[3:0];
  _RAND_2003 = {1{`RANDOM}};
  image_2317 = _RAND_2003[3:0];
  _RAND_2004 = {1{`RANDOM}};
  image_2318 = _RAND_2004[3:0];
  _RAND_2005 = {1{`RANDOM}};
  image_2319 = _RAND_2005[3:0];
  _RAND_2006 = {1{`RANDOM}};
  image_2320 = _RAND_2006[3:0];
  _RAND_2007 = {1{`RANDOM}};
  image_2321 = _RAND_2007[3:0];
  _RAND_2008 = {1{`RANDOM}};
  image_2322 = _RAND_2008[3:0];
  _RAND_2009 = {1{`RANDOM}};
  image_2323 = _RAND_2009[3:0];
  _RAND_2010 = {1{`RANDOM}};
  image_2324 = _RAND_2010[3:0];
  _RAND_2011 = {1{`RANDOM}};
  image_2325 = _RAND_2011[3:0];
  _RAND_2012 = {1{`RANDOM}};
  image_2326 = _RAND_2012[3:0];
  _RAND_2013 = {1{`RANDOM}};
  image_2327 = _RAND_2013[3:0];
  _RAND_2014 = {1{`RANDOM}};
  image_2328 = _RAND_2014[3:0];
  _RAND_2015 = {1{`RANDOM}};
  image_2329 = _RAND_2015[3:0];
  _RAND_2016 = {1{`RANDOM}};
  image_2330 = _RAND_2016[3:0];
  _RAND_2017 = {1{`RANDOM}};
  image_2331 = _RAND_2017[3:0];
  _RAND_2018 = {1{`RANDOM}};
  image_2332 = _RAND_2018[3:0];
  _RAND_2019 = {1{`RANDOM}};
  image_2333 = _RAND_2019[3:0];
  _RAND_2020 = {1{`RANDOM}};
  image_2334 = _RAND_2020[3:0];
  _RAND_2021 = {1{`RANDOM}};
  image_2335 = _RAND_2021[3:0];
  _RAND_2022 = {1{`RANDOM}};
  image_2336 = _RAND_2022[3:0];
  _RAND_2023 = {1{`RANDOM}};
  image_2337 = _RAND_2023[3:0];
  _RAND_2024 = {1{`RANDOM}};
  image_2338 = _RAND_2024[3:0];
  _RAND_2025 = {1{`RANDOM}};
  image_2339 = _RAND_2025[3:0];
  _RAND_2026 = {1{`RANDOM}};
  image_2340 = _RAND_2026[3:0];
  _RAND_2027 = {1{`RANDOM}};
  image_2341 = _RAND_2027[3:0];
  _RAND_2028 = {1{`RANDOM}};
  image_2342 = _RAND_2028[3:0];
  _RAND_2029 = {1{`RANDOM}};
  image_2343 = _RAND_2029[3:0];
  _RAND_2030 = {1{`RANDOM}};
  image_2344 = _RAND_2030[3:0];
  _RAND_2031 = {1{`RANDOM}};
  image_2345 = _RAND_2031[3:0];
  _RAND_2032 = {1{`RANDOM}};
  image_2346 = _RAND_2032[3:0];
  _RAND_2033 = {1{`RANDOM}};
  image_2347 = _RAND_2033[3:0];
  _RAND_2034 = {1{`RANDOM}};
  image_2348 = _RAND_2034[3:0];
  _RAND_2035 = {1{`RANDOM}};
  image_2349 = _RAND_2035[3:0];
  _RAND_2036 = {1{`RANDOM}};
  image_2350 = _RAND_2036[3:0];
  _RAND_2037 = {1{`RANDOM}};
  image_2351 = _RAND_2037[3:0];
  _RAND_2038 = {1{`RANDOM}};
  image_2352 = _RAND_2038[3:0];
  _RAND_2039 = {1{`RANDOM}};
  image_2353 = _RAND_2039[3:0];
  _RAND_2040 = {1{`RANDOM}};
  image_2354 = _RAND_2040[3:0];
  _RAND_2041 = {1{`RANDOM}};
  image_2355 = _RAND_2041[3:0];
  _RAND_2042 = {1{`RANDOM}};
  image_2356 = _RAND_2042[3:0];
  _RAND_2043 = {1{`RANDOM}};
  image_2357 = _RAND_2043[3:0];
  _RAND_2044 = {1{`RANDOM}};
  image_2358 = _RAND_2044[3:0];
  _RAND_2045 = {1{`RANDOM}};
  image_2359 = _RAND_2045[3:0];
  _RAND_2046 = {1{`RANDOM}};
  image_2360 = _RAND_2046[3:0];
  _RAND_2047 = {1{`RANDOM}};
  image_2361 = _RAND_2047[3:0];
  _RAND_2048 = {1{`RANDOM}};
  image_2362 = _RAND_2048[3:0];
  _RAND_2049 = {1{`RANDOM}};
  image_2372 = _RAND_2049[3:0];
  _RAND_2050 = {1{`RANDOM}};
  image_2373 = _RAND_2050[3:0];
  _RAND_2051 = {1{`RANDOM}};
  image_2374 = _RAND_2051[3:0];
  _RAND_2052 = {1{`RANDOM}};
  image_2375 = _RAND_2052[3:0];
  _RAND_2053 = {1{`RANDOM}};
  image_2376 = _RAND_2053[3:0];
  _RAND_2054 = {1{`RANDOM}};
  image_2377 = _RAND_2054[3:0];
  _RAND_2055 = {1{`RANDOM}};
  image_2378 = _RAND_2055[3:0];
  _RAND_2056 = {1{`RANDOM}};
  image_2379 = _RAND_2056[3:0];
  _RAND_2057 = {1{`RANDOM}};
  image_2380 = _RAND_2057[3:0];
  _RAND_2058 = {1{`RANDOM}};
  image_2381 = _RAND_2058[3:0];
  _RAND_2059 = {1{`RANDOM}};
  image_2382 = _RAND_2059[3:0];
  _RAND_2060 = {1{`RANDOM}};
  image_2383 = _RAND_2060[3:0];
  _RAND_2061 = {1{`RANDOM}};
  image_2384 = _RAND_2061[3:0];
  _RAND_2062 = {1{`RANDOM}};
  image_2385 = _RAND_2062[3:0];
  _RAND_2063 = {1{`RANDOM}};
  image_2386 = _RAND_2063[3:0];
  _RAND_2064 = {1{`RANDOM}};
  image_2387 = _RAND_2064[3:0];
  _RAND_2065 = {1{`RANDOM}};
  image_2388 = _RAND_2065[3:0];
  _RAND_2066 = {1{`RANDOM}};
  image_2389 = _RAND_2066[3:0];
  _RAND_2067 = {1{`RANDOM}};
  image_2390 = _RAND_2067[3:0];
  _RAND_2068 = {1{`RANDOM}};
  image_2391 = _RAND_2068[3:0];
  _RAND_2069 = {1{`RANDOM}};
  image_2392 = _RAND_2069[3:0];
  _RAND_2070 = {1{`RANDOM}};
  image_2393 = _RAND_2070[3:0];
  _RAND_2071 = {1{`RANDOM}};
  image_2394 = _RAND_2071[3:0];
  _RAND_2072 = {1{`RANDOM}};
  image_2395 = _RAND_2072[3:0];
  _RAND_2073 = {1{`RANDOM}};
  image_2396 = _RAND_2073[3:0];
  _RAND_2074 = {1{`RANDOM}};
  image_2397 = _RAND_2074[3:0];
  _RAND_2075 = {1{`RANDOM}};
  image_2398 = _RAND_2075[3:0];
  _RAND_2076 = {1{`RANDOM}};
  image_2399 = _RAND_2076[3:0];
  _RAND_2077 = {1{`RANDOM}};
  image_2400 = _RAND_2077[3:0];
  _RAND_2078 = {1{`RANDOM}};
  image_2401 = _RAND_2078[3:0];
  _RAND_2079 = {1{`RANDOM}};
  image_2402 = _RAND_2079[3:0];
  _RAND_2080 = {1{`RANDOM}};
  image_2403 = _RAND_2080[3:0];
  _RAND_2081 = {1{`RANDOM}};
  image_2404 = _RAND_2081[3:0];
  _RAND_2082 = {1{`RANDOM}};
  image_2405 = _RAND_2082[3:0];
  _RAND_2083 = {1{`RANDOM}};
  image_2406 = _RAND_2083[3:0];
  _RAND_2084 = {1{`RANDOM}};
  image_2407 = _RAND_2084[3:0];
  _RAND_2085 = {1{`RANDOM}};
  image_2408 = _RAND_2085[3:0];
  _RAND_2086 = {1{`RANDOM}};
  image_2409 = _RAND_2086[3:0];
  _RAND_2087 = {1{`RANDOM}};
  image_2410 = _RAND_2087[3:0];
  _RAND_2088 = {1{`RANDOM}};
  image_2411 = _RAND_2088[3:0];
  _RAND_2089 = {1{`RANDOM}};
  image_2412 = _RAND_2089[3:0];
  _RAND_2090 = {1{`RANDOM}};
  image_2413 = _RAND_2090[3:0];
  _RAND_2091 = {1{`RANDOM}};
  image_2414 = _RAND_2091[3:0];
  _RAND_2092 = {1{`RANDOM}};
  image_2415 = _RAND_2092[3:0];
  _RAND_2093 = {1{`RANDOM}};
  image_2416 = _RAND_2093[3:0];
  _RAND_2094 = {1{`RANDOM}};
  image_2417 = _RAND_2094[3:0];
  _RAND_2095 = {1{`RANDOM}};
  image_2418 = _RAND_2095[3:0];
  _RAND_2096 = {1{`RANDOM}};
  image_2419 = _RAND_2096[3:0];
  _RAND_2097 = {1{`RANDOM}};
  image_2420 = _RAND_2097[3:0];
  _RAND_2098 = {1{`RANDOM}};
  image_2421 = _RAND_2098[3:0];
  _RAND_2099 = {1{`RANDOM}};
  image_2422 = _RAND_2099[3:0];
  _RAND_2100 = {1{`RANDOM}};
  image_2423 = _RAND_2100[3:0];
  _RAND_2101 = {1{`RANDOM}};
  image_2424 = _RAND_2101[3:0];
  _RAND_2102 = {1{`RANDOM}};
  image_2425 = _RAND_2102[3:0];
  _RAND_2103 = {1{`RANDOM}};
  image_2426 = _RAND_2103[3:0];
  _RAND_2104 = {1{`RANDOM}};
  image_2437 = _RAND_2104[3:0];
  _RAND_2105 = {1{`RANDOM}};
  image_2438 = _RAND_2105[3:0];
  _RAND_2106 = {1{`RANDOM}};
  image_2439 = _RAND_2106[3:0];
  _RAND_2107 = {1{`RANDOM}};
  image_2440 = _RAND_2107[3:0];
  _RAND_2108 = {1{`RANDOM}};
  image_2441 = _RAND_2108[3:0];
  _RAND_2109 = {1{`RANDOM}};
  image_2442 = _RAND_2109[3:0];
  _RAND_2110 = {1{`RANDOM}};
  image_2443 = _RAND_2110[3:0];
  _RAND_2111 = {1{`RANDOM}};
  image_2444 = _RAND_2111[3:0];
  _RAND_2112 = {1{`RANDOM}};
  image_2445 = _RAND_2112[3:0];
  _RAND_2113 = {1{`RANDOM}};
  image_2446 = _RAND_2113[3:0];
  _RAND_2114 = {1{`RANDOM}};
  image_2447 = _RAND_2114[3:0];
  _RAND_2115 = {1{`RANDOM}};
  image_2448 = _RAND_2115[3:0];
  _RAND_2116 = {1{`RANDOM}};
  image_2449 = _RAND_2116[3:0];
  _RAND_2117 = {1{`RANDOM}};
  image_2450 = _RAND_2117[3:0];
  _RAND_2118 = {1{`RANDOM}};
  image_2451 = _RAND_2118[3:0];
  _RAND_2119 = {1{`RANDOM}};
  image_2452 = _RAND_2119[3:0];
  _RAND_2120 = {1{`RANDOM}};
  image_2453 = _RAND_2120[3:0];
  _RAND_2121 = {1{`RANDOM}};
  image_2454 = _RAND_2121[3:0];
  _RAND_2122 = {1{`RANDOM}};
  image_2455 = _RAND_2122[3:0];
  _RAND_2123 = {1{`RANDOM}};
  image_2456 = _RAND_2123[3:0];
  _RAND_2124 = {1{`RANDOM}};
  image_2457 = _RAND_2124[3:0];
  _RAND_2125 = {1{`RANDOM}};
  image_2458 = _RAND_2125[3:0];
  _RAND_2126 = {1{`RANDOM}};
  image_2459 = _RAND_2126[3:0];
  _RAND_2127 = {1{`RANDOM}};
  image_2460 = _RAND_2127[3:0];
  _RAND_2128 = {1{`RANDOM}};
  image_2461 = _RAND_2128[3:0];
  _RAND_2129 = {1{`RANDOM}};
  image_2462 = _RAND_2129[3:0];
  _RAND_2130 = {1{`RANDOM}};
  image_2463 = _RAND_2130[3:0];
  _RAND_2131 = {1{`RANDOM}};
  image_2464 = _RAND_2131[3:0];
  _RAND_2132 = {1{`RANDOM}};
  image_2465 = _RAND_2132[3:0];
  _RAND_2133 = {1{`RANDOM}};
  image_2466 = _RAND_2133[3:0];
  _RAND_2134 = {1{`RANDOM}};
  image_2467 = _RAND_2134[3:0];
  _RAND_2135 = {1{`RANDOM}};
  image_2468 = _RAND_2135[3:0];
  _RAND_2136 = {1{`RANDOM}};
  image_2469 = _RAND_2136[3:0];
  _RAND_2137 = {1{`RANDOM}};
  image_2470 = _RAND_2137[3:0];
  _RAND_2138 = {1{`RANDOM}};
  image_2471 = _RAND_2138[3:0];
  _RAND_2139 = {1{`RANDOM}};
  image_2472 = _RAND_2139[3:0];
  _RAND_2140 = {1{`RANDOM}};
  image_2473 = _RAND_2140[3:0];
  _RAND_2141 = {1{`RANDOM}};
  image_2474 = _RAND_2141[3:0];
  _RAND_2142 = {1{`RANDOM}};
  image_2475 = _RAND_2142[3:0];
  _RAND_2143 = {1{`RANDOM}};
  image_2476 = _RAND_2143[3:0];
  _RAND_2144 = {1{`RANDOM}};
  image_2477 = _RAND_2144[3:0];
  _RAND_2145 = {1{`RANDOM}};
  image_2478 = _RAND_2145[3:0];
  _RAND_2146 = {1{`RANDOM}};
  image_2479 = _RAND_2146[3:0];
  _RAND_2147 = {1{`RANDOM}};
  image_2480 = _RAND_2147[3:0];
  _RAND_2148 = {1{`RANDOM}};
  image_2481 = _RAND_2148[3:0];
  _RAND_2149 = {1{`RANDOM}};
  image_2482 = _RAND_2149[3:0];
  _RAND_2150 = {1{`RANDOM}};
  image_2483 = _RAND_2150[3:0];
  _RAND_2151 = {1{`RANDOM}};
  image_2484 = _RAND_2151[3:0];
  _RAND_2152 = {1{`RANDOM}};
  image_2485 = _RAND_2152[3:0];
  _RAND_2153 = {1{`RANDOM}};
  image_2486 = _RAND_2153[3:0];
  _RAND_2154 = {1{`RANDOM}};
  image_2487 = _RAND_2154[3:0];
  _RAND_2155 = {1{`RANDOM}};
  image_2488 = _RAND_2155[3:0];
  _RAND_2156 = {1{`RANDOM}};
  image_2489 = _RAND_2156[3:0];
  _RAND_2157 = {1{`RANDOM}};
  image_2490 = _RAND_2157[3:0];
  _RAND_2158 = {1{`RANDOM}};
  image_2502 = _RAND_2158[3:0];
  _RAND_2159 = {1{`RANDOM}};
  image_2503 = _RAND_2159[3:0];
  _RAND_2160 = {1{`RANDOM}};
  image_2504 = _RAND_2160[3:0];
  _RAND_2161 = {1{`RANDOM}};
  image_2505 = _RAND_2161[3:0];
  _RAND_2162 = {1{`RANDOM}};
  image_2506 = _RAND_2162[3:0];
  _RAND_2163 = {1{`RANDOM}};
  image_2507 = _RAND_2163[3:0];
  _RAND_2164 = {1{`RANDOM}};
  image_2508 = _RAND_2164[3:0];
  _RAND_2165 = {1{`RANDOM}};
  image_2509 = _RAND_2165[3:0];
  _RAND_2166 = {1{`RANDOM}};
  image_2510 = _RAND_2166[3:0];
  _RAND_2167 = {1{`RANDOM}};
  image_2511 = _RAND_2167[3:0];
  _RAND_2168 = {1{`RANDOM}};
  image_2512 = _RAND_2168[3:0];
  _RAND_2169 = {1{`RANDOM}};
  image_2513 = _RAND_2169[3:0];
  _RAND_2170 = {1{`RANDOM}};
  image_2514 = _RAND_2170[3:0];
  _RAND_2171 = {1{`RANDOM}};
  image_2515 = _RAND_2171[3:0];
  _RAND_2172 = {1{`RANDOM}};
  image_2516 = _RAND_2172[3:0];
  _RAND_2173 = {1{`RANDOM}};
  image_2517 = _RAND_2173[3:0];
  _RAND_2174 = {1{`RANDOM}};
  image_2518 = _RAND_2174[3:0];
  _RAND_2175 = {1{`RANDOM}};
  image_2519 = _RAND_2175[3:0];
  _RAND_2176 = {1{`RANDOM}};
  image_2520 = _RAND_2176[3:0];
  _RAND_2177 = {1{`RANDOM}};
  image_2521 = _RAND_2177[3:0];
  _RAND_2178 = {1{`RANDOM}};
  image_2522 = _RAND_2178[3:0];
  _RAND_2179 = {1{`RANDOM}};
  image_2523 = _RAND_2179[3:0];
  _RAND_2180 = {1{`RANDOM}};
  image_2524 = _RAND_2180[3:0];
  _RAND_2181 = {1{`RANDOM}};
  image_2525 = _RAND_2181[3:0];
  _RAND_2182 = {1{`RANDOM}};
  image_2526 = _RAND_2182[3:0];
  _RAND_2183 = {1{`RANDOM}};
  image_2527 = _RAND_2183[3:0];
  _RAND_2184 = {1{`RANDOM}};
  image_2528 = _RAND_2184[3:0];
  _RAND_2185 = {1{`RANDOM}};
  image_2529 = _RAND_2185[3:0];
  _RAND_2186 = {1{`RANDOM}};
  image_2530 = _RAND_2186[3:0];
  _RAND_2187 = {1{`RANDOM}};
  image_2531 = _RAND_2187[3:0];
  _RAND_2188 = {1{`RANDOM}};
  image_2532 = _RAND_2188[3:0];
  _RAND_2189 = {1{`RANDOM}};
  image_2533 = _RAND_2189[3:0];
  _RAND_2190 = {1{`RANDOM}};
  image_2534 = _RAND_2190[3:0];
  _RAND_2191 = {1{`RANDOM}};
  image_2535 = _RAND_2191[3:0];
  _RAND_2192 = {1{`RANDOM}};
  image_2536 = _RAND_2192[3:0];
  _RAND_2193 = {1{`RANDOM}};
  image_2537 = _RAND_2193[3:0];
  _RAND_2194 = {1{`RANDOM}};
  image_2538 = _RAND_2194[3:0];
  _RAND_2195 = {1{`RANDOM}};
  image_2539 = _RAND_2195[3:0];
  _RAND_2196 = {1{`RANDOM}};
  image_2540 = _RAND_2196[3:0];
  _RAND_2197 = {1{`RANDOM}};
  image_2541 = _RAND_2197[3:0];
  _RAND_2198 = {1{`RANDOM}};
  image_2542 = _RAND_2198[3:0];
  _RAND_2199 = {1{`RANDOM}};
  image_2543 = _RAND_2199[3:0];
  _RAND_2200 = {1{`RANDOM}};
  image_2544 = _RAND_2200[3:0];
  _RAND_2201 = {1{`RANDOM}};
  image_2545 = _RAND_2201[3:0];
  _RAND_2202 = {1{`RANDOM}};
  image_2546 = _RAND_2202[3:0];
  _RAND_2203 = {1{`RANDOM}};
  image_2547 = _RAND_2203[3:0];
  _RAND_2204 = {1{`RANDOM}};
  image_2548 = _RAND_2204[3:0];
  _RAND_2205 = {1{`RANDOM}};
  image_2549 = _RAND_2205[3:0];
  _RAND_2206 = {1{`RANDOM}};
  image_2550 = _RAND_2206[3:0];
  _RAND_2207 = {1{`RANDOM}};
  image_2551 = _RAND_2207[3:0];
  _RAND_2208 = {1{`RANDOM}};
  image_2552 = _RAND_2208[3:0];
  _RAND_2209 = {1{`RANDOM}};
  image_2553 = _RAND_2209[3:0];
  _RAND_2210 = {1{`RANDOM}};
  image_2554 = _RAND_2210[3:0];
  _RAND_2211 = {1{`RANDOM}};
  image_2567 = _RAND_2211[3:0];
  _RAND_2212 = {1{`RANDOM}};
  image_2568 = _RAND_2212[3:0];
  _RAND_2213 = {1{`RANDOM}};
  image_2569 = _RAND_2213[3:0];
  _RAND_2214 = {1{`RANDOM}};
  image_2570 = _RAND_2214[3:0];
  _RAND_2215 = {1{`RANDOM}};
  image_2571 = _RAND_2215[3:0];
  _RAND_2216 = {1{`RANDOM}};
  image_2572 = _RAND_2216[3:0];
  _RAND_2217 = {1{`RANDOM}};
  image_2573 = _RAND_2217[3:0];
  _RAND_2218 = {1{`RANDOM}};
  image_2574 = _RAND_2218[3:0];
  _RAND_2219 = {1{`RANDOM}};
  image_2575 = _RAND_2219[3:0];
  _RAND_2220 = {1{`RANDOM}};
  image_2576 = _RAND_2220[3:0];
  _RAND_2221 = {1{`RANDOM}};
  image_2577 = _RAND_2221[3:0];
  _RAND_2222 = {1{`RANDOM}};
  image_2578 = _RAND_2222[3:0];
  _RAND_2223 = {1{`RANDOM}};
  image_2579 = _RAND_2223[3:0];
  _RAND_2224 = {1{`RANDOM}};
  image_2580 = _RAND_2224[3:0];
  _RAND_2225 = {1{`RANDOM}};
  image_2581 = _RAND_2225[3:0];
  _RAND_2226 = {1{`RANDOM}};
  image_2582 = _RAND_2226[3:0];
  _RAND_2227 = {1{`RANDOM}};
  image_2583 = _RAND_2227[3:0];
  _RAND_2228 = {1{`RANDOM}};
  image_2584 = _RAND_2228[3:0];
  _RAND_2229 = {1{`RANDOM}};
  image_2585 = _RAND_2229[3:0];
  _RAND_2230 = {1{`RANDOM}};
  image_2586 = _RAND_2230[3:0];
  _RAND_2231 = {1{`RANDOM}};
  image_2587 = _RAND_2231[3:0];
  _RAND_2232 = {1{`RANDOM}};
  image_2588 = _RAND_2232[3:0];
  _RAND_2233 = {1{`RANDOM}};
  image_2589 = _RAND_2233[3:0];
  _RAND_2234 = {1{`RANDOM}};
  image_2590 = _RAND_2234[3:0];
  _RAND_2235 = {1{`RANDOM}};
  image_2591 = _RAND_2235[3:0];
  _RAND_2236 = {1{`RANDOM}};
  image_2592 = _RAND_2236[3:0];
  _RAND_2237 = {1{`RANDOM}};
  image_2593 = _RAND_2237[3:0];
  _RAND_2238 = {1{`RANDOM}};
  image_2594 = _RAND_2238[3:0];
  _RAND_2239 = {1{`RANDOM}};
  image_2595 = _RAND_2239[3:0];
  _RAND_2240 = {1{`RANDOM}};
  image_2596 = _RAND_2240[3:0];
  _RAND_2241 = {1{`RANDOM}};
  image_2597 = _RAND_2241[3:0];
  _RAND_2242 = {1{`RANDOM}};
  image_2598 = _RAND_2242[3:0];
  _RAND_2243 = {1{`RANDOM}};
  image_2599 = _RAND_2243[3:0];
  _RAND_2244 = {1{`RANDOM}};
  image_2600 = _RAND_2244[3:0];
  _RAND_2245 = {1{`RANDOM}};
  image_2601 = _RAND_2245[3:0];
  _RAND_2246 = {1{`RANDOM}};
  image_2602 = _RAND_2246[3:0];
  _RAND_2247 = {1{`RANDOM}};
  image_2603 = _RAND_2247[3:0];
  _RAND_2248 = {1{`RANDOM}};
  image_2604 = _RAND_2248[3:0];
  _RAND_2249 = {1{`RANDOM}};
  image_2605 = _RAND_2249[3:0];
  _RAND_2250 = {1{`RANDOM}};
  image_2606 = _RAND_2250[3:0];
  _RAND_2251 = {1{`RANDOM}};
  image_2607 = _RAND_2251[3:0];
  _RAND_2252 = {1{`RANDOM}};
  image_2608 = _RAND_2252[3:0];
  _RAND_2253 = {1{`RANDOM}};
  image_2609 = _RAND_2253[3:0];
  _RAND_2254 = {1{`RANDOM}};
  image_2610 = _RAND_2254[3:0];
  _RAND_2255 = {1{`RANDOM}};
  image_2611 = _RAND_2255[3:0];
  _RAND_2256 = {1{`RANDOM}};
  image_2612 = _RAND_2256[3:0];
  _RAND_2257 = {1{`RANDOM}};
  image_2613 = _RAND_2257[3:0];
  _RAND_2258 = {1{`RANDOM}};
  image_2614 = _RAND_2258[3:0];
  _RAND_2259 = {1{`RANDOM}};
  image_2615 = _RAND_2259[3:0];
  _RAND_2260 = {1{`RANDOM}};
  image_2616 = _RAND_2260[3:0];
  _RAND_2261 = {1{`RANDOM}};
  image_2617 = _RAND_2261[3:0];
  _RAND_2262 = {1{`RANDOM}};
  image_2618 = _RAND_2262[3:0];
  _RAND_2263 = {1{`RANDOM}};
  image_2632 = _RAND_2263[3:0];
  _RAND_2264 = {1{`RANDOM}};
  image_2633 = _RAND_2264[3:0];
  _RAND_2265 = {1{`RANDOM}};
  image_2634 = _RAND_2265[3:0];
  _RAND_2266 = {1{`RANDOM}};
  image_2635 = _RAND_2266[3:0];
  _RAND_2267 = {1{`RANDOM}};
  image_2636 = _RAND_2267[3:0];
  _RAND_2268 = {1{`RANDOM}};
  image_2637 = _RAND_2268[3:0];
  _RAND_2269 = {1{`RANDOM}};
  image_2638 = _RAND_2269[3:0];
  _RAND_2270 = {1{`RANDOM}};
  image_2639 = _RAND_2270[3:0];
  _RAND_2271 = {1{`RANDOM}};
  image_2640 = _RAND_2271[3:0];
  _RAND_2272 = {1{`RANDOM}};
  image_2641 = _RAND_2272[3:0];
  _RAND_2273 = {1{`RANDOM}};
  image_2642 = _RAND_2273[3:0];
  _RAND_2274 = {1{`RANDOM}};
  image_2643 = _RAND_2274[3:0];
  _RAND_2275 = {1{`RANDOM}};
  image_2644 = _RAND_2275[3:0];
  _RAND_2276 = {1{`RANDOM}};
  image_2645 = _RAND_2276[3:0];
  _RAND_2277 = {1{`RANDOM}};
  image_2646 = _RAND_2277[3:0];
  _RAND_2278 = {1{`RANDOM}};
  image_2647 = _RAND_2278[3:0];
  _RAND_2279 = {1{`RANDOM}};
  image_2648 = _RAND_2279[3:0];
  _RAND_2280 = {1{`RANDOM}};
  image_2649 = _RAND_2280[3:0];
  _RAND_2281 = {1{`RANDOM}};
  image_2650 = _RAND_2281[3:0];
  _RAND_2282 = {1{`RANDOM}};
  image_2651 = _RAND_2282[3:0];
  _RAND_2283 = {1{`RANDOM}};
  image_2652 = _RAND_2283[3:0];
  _RAND_2284 = {1{`RANDOM}};
  image_2653 = _RAND_2284[3:0];
  _RAND_2285 = {1{`RANDOM}};
  image_2654 = _RAND_2285[3:0];
  _RAND_2286 = {1{`RANDOM}};
  image_2655 = _RAND_2286[3:0];
  _RAND_2287 = {1{`RANDOM}};
  image_2656 = _RAND_2287[3:0];
  _RAND_2288 = {1{`RANDOM}};
  image_2657 = _RAND_2288[3:0];
  _RAND_2289 = {1{`RANDOM}};
  image_2658 = _RAND_2289[3:0];
  _RAND_2290 = {1{`RANDOM}};
  image_2659 = _RAND_2290[3:0];
  _RAND_2291 = {1{`RANDOM}};
  image_2660 = _RAND_2291[3:0];
  _RAND_2292 = {1{`RANDOM}};
  image_2661 = _RAND_2292[3:0];
  _RAND_2293 = {1{`RANDOM}};
  image_2662 = _RAND_2293[3:0];
  _RAND_2294 = {1{`RANDOM}};
  image_2663 = _RAND_2294[3:0];
  _RAND_2295 = {1{`RANDOM}};
  image_2664 = _RAND_2295[3:0];
  _RAND_2296 = {1{`RANDOM}};
  image_2665 = _RAND_2296[3:0];
  _RAND_2297 = {1{`RANDOM}};
  image_2666 = _RAND_2297[3:0];
  _RAND_2298 = {1{`RANDOM}};
  image_2667 = _RAND_2298[3:0];
  _RAND_2299 = {1{`RANDOM}};
  image_2668 = _RAND_2299[3:0];
  _RAND_2300 = {1{`RANDOM}};
  image_2669 = _RAND_2300[3:0];
  _RAND_2301 = {1{`RANDOM}};
  image_2670 = _RAND_2301[3:0];
  _RAND_2302 = {1{`RANDOM}};
  image_2671 = _RAND_2302[3:0];
  _RAND_2303 = {1{`RANDOM}};
  image_2672 = _RAND_2303[3:0];
  _RAND_2304 = {1{`RANDOM}};
  image_2673 = _RAND_2304[3:0];
  _RAND_2305 = {1{`RANDOM}};
  image_2674 = _RAND_2305[3:0];
  _RAND_2306 = {1{`RANDOM}};
  image_2675 = _RAND_2306[3:0];
  _RAND_2307 = {1{`RANDOM}};
  image_2676 = _RAND_2307[3:0];
  _RAND_2308 = {1{`RANDOM}};
  image_2677 = _RAND_2308[3:0];
  _RAND_2309 = {1{`RANDOM}};
  image_2678 = _RAND_2309[3:0];
  _RAND_2310 = {1{`RANDOM}};
  image_2679 = _RAND_2310[3:0];
  _RAND_2311 = {1{`RANDOM}};
  image_2680 = _RAND_2311[3:0];
  _RAND_2312 = {1{`RANDOM}};
  image_2681 = _RAND_2312[3:0];
  _RAND_2313 = {1{`RANDOM}};
  image_2682 = _RAND_2313[3:0];
  _RAND_2314 = {1{`RANDOM}};
  image_2697 = _RAND_2314[3:0];
  _RAND_2315 = {1{`RANDOM}};
  image_2698 = _RAND_2315[3:0];
  _RAND_2316 = {1{`RANDOM}};
  image_2699 = _RAND_2316[3:0];
  _RAND_2317 = {1{`RANDOM}};
  image_2700 = _RAND_2317[3:0];
  _RAND_2318 = {1{`RANDOM}};
  image_2701 = _RAND_2318[3:0];
  _RAND_2319 = {1{`RANDOM}};
  image_2702 = _RAND_2319[3:0];
  _RAND_2320 = {1{`RANDOM}};
  image_2703 = _RAND_2320[3:0];
  _RAND_2321 = {1{`RANDOM}};
  image_2704 = _RAND_2321[3:0];
  _RAND_2322 = {1{`RANDOM}};
  image_2705 = _RAND_2322[3:0];
  _RAND_2323 = {1{`RANDOM}};
  image_2706 = _RAND_2323[3:0];
  _RAND_2324 = {1{`RANDOM}};
  image_2707 = _RAND_2324[3:0];
  _RAND_2325 = {1{`RANDOM}};
  image_2708 = _RAND_2325[3:0];
  _RAND_2326 = {1{`RANDOM}};
  image_2709 = _RAND_2326[3:0];
  _RAND_2327 = {1{`RANDOM}};
  image_2710 = _RAND_2327[3:0];
  _RAND_2328 = {1{`RANDOM}};
  image_2711 = _RAND_2328[3:0];
  _RAND_2329 = {1{`RANDOM}};
  image_2712 = _RAND_2329[3:0];
  _RAND_2330 = {1{`RANDOM}};
  image_2713 = _RAND_2330[3:0];
  _RAND_2331 = {1{`RANDOM}};
  image_2714 = _RAND_2331[3:0];
  _RAND_2332 = {1{`RANDOM}};
  image_2715 = _RAND_2332[3:0];
  _RAND_2333 = {1{`RANDOM}};
  image_2716 = _RAND_2333[3:0];
  _RAND_2334 = {1{`RANDOM}};
  image_2717 = _RAND_2334[3:0];
  _RAND_2335 = {1{`RANDOM}};
  image_2718 = _RAND_2335[3:0];
  _RAND_2336 = {1{`RANDOM}};
  image_2719 = _RAND_2336[3:0];
  _RAND_2337 = {1{`RANDOM}};
  image_2720 = _RAND_2337[3:0];
  _RAND_2338 = {1{`RANDOM}};
  image_2721 = _RAND_2338[3:0];
  _RAND_2339 = {1{`RANDOM}};
  image_2722 = _RAND_2339[3:0];
  _RAND_2340 = {1{`RANDOM}};
  image_2723 = _RAND_2340[3:0];
  _RAND_2341 = {1{`RANDOM}};
  image_2724 = _RAND_2341[3:0];
  _RAND_2342 = {1{`RANDOM}};
  image_2725 = _RAND_2342[3:0];
  _RAND_2343 = {1{`RANDOM}};
  image_2726 = _RAND_2343[3:0];
  _RAND_2344 = {1{`RANDOM}};
  image_2727 = _RAND_2344[3:0];
  _RAND_2345 = {1{`RANDOM}};
  image_2728 = _RAND_2345[3:0];
  _RAND_2346 = {1{`RANDOM}};
  image_2729 = _RAND_2346[3:0];
  _RAND_2347 = {1{`RANDOM}};
  image_2730 = _RAND_2347[3:0];
  _RAND_2348 = {1{`RANDOM}};
  image_2731 = _RAND_2348[3:0];
  _RAND_2349 = {1{`RANDOM}};
  image_2732 = _RAND_2349[3:0];
  _RAND_2350 = {1{`RANDOM}};
  image_2733 = _RAND_2350[3:0];
  _RAND_2351 = {1{`RANDOM}};
  image_2734 = _RAND_2351[3:0];
  _RAND_2352 = {1{`RANDOM}};
  image_2735 = _RAND_2352[3:0];
  _RAND_2353 = {1{`RANDOM}};
  image_2736 = _RAND_2353[3:0];
  _RAND_2354 = {1{`RANDOM}};
  image_2737 = _RAND_2354[3:0];
  _RAND_2355 = {1{`RANDOM}};
  image_2738 = _RAND_2355[3:0];
  _RAND_2356 = {1{`RANDOM}};
  image_2739 = _RAND_2356[3:0];
  _RAND_2357 = {1{`RANDOM}};
  image_2740 = _RAND_2357[3:0];
  _RAND_2358 = {1{`RANDOM}};
  image_2741 = _RAND_2358[3:0];
  _RAND_2359 = {1{`RANDOM}};
  image_2742 = _RAND_2359[3:0];
  _RAND_2360 = {1{`RANDOM}};
  image_2743 = _RAND_2360[3:0];
  _RAND_2361 = {1{`RANDOM}};
  image_2744 = _RAND_2361[3:0];
  _RAND_2362 = {1{`RANDOM}};
  image_2745 = _RAND_2362[3:0];
  _RAND_2363 = {1{`RANDOM}};
  image_2763 = _RAND_2363[3:0];
  _RAND_2364 = {1{`RANDOM}};
  image_2764 = _RAND_2364[3:0];
  _RAND_2365 = {1{`RANDOM}};
  image_2765 = _RAND_2365[3:0];
  _RAND_2366 = {1{`RANDOM}};
  image_2766 = _RAND_2366[3:0];
  _RAND_2367 = {1{`RANDOM}};
  image_2767 = _RAND_2367[3:0];
  _RAND_2368 = {1{`RANDOM}};
  image_2768 = _RAND_2368[3:0];
  _RAND_2369 = {1{`RANDOM}};
  image_2769 = _RAND_2369[3:0];
  _RAND_2370 = {1{`RANDOM}};
  image_2770 = _RAND_2370[3:0];
  _RAND_2371 = {1{`RANDOM}};
  image_2771 = _RAND_2371[3:0];
  _RAND_2372 = {1{`RANDOM}};
  image_2772 = _RAND_2372[3:0];
  _RAND_2373 = {1{`RANDOM}};
  image_2773 = _RAND_2373[3:0];
  _RAND_2374 = {1{`RANDOM}};
  image_2774 = _RAND_2374[3:0];
  _RAND_2375 = {1{`RANDOM}};
  image_2775 = _RAND_2375[3:0];
  _RAND_2376 = {1{`RANDOM}};
  image_2776 = _RAND_2376[3:0];
  _RAND_2377 = {1{`RANDOM}};
  image_2777 = _RAND_2377[3:0];
  _RAND_2378 = {1{`RANDOM}};
  image_2778 = _RAND_2378[3:0];
  _RAND_2379 = {1{`RANDOM}};
  image_2779 = _RAND_2379[3:0];
  _RAND_2380 = {1{`RANDOM}};
  image_2780 = _RAND_2380[3:0];
  _RAND_2381 = {1{`RANDOM}};
  image_2781 = _RAND_2381[3:0];
  _RAND_2382 = {1{`RANDOM}};
  image_2782 = _RAND_2382[3:0];
  _RAND_2383 = {1{`RANDOM}};
  image_2783 = _RAND_2383[3:0];
  _RAND_2384 = {1{`RANDOM}};
  image_2784 = _RAND_2384[3:0];
  _RAND_2385 = {1{`RANDOM}};
  image_2785 = _RAND_2385[3:0];
  _RAND_2386 = {1{`RANDOM}};
  image_2786 = _RAND_2386[3:0];
  _RAND_2387 = {1{`RANDOM}};
  image_2787 = _RAND_2387[3:0];
  _RAND_2388 = {1{`RANDOM}};
  image_2788 = _RAND_2388[3:0];
  _RAND_2389 = {1{`RANDOM}};
  image_2789 = _RAND_2389[3:0];
  _RAND_2390 = {1{`RANDOM}};
  image_2790 = _RAND_2390[3:0];
  _RAND_2391 = {1{`RANDOM}};
  image_2791 = _RAND_2391[3:0];
  _RAND_2392 = {1{`RANDOM}};
  image_2792 = _RAND_2392[3:0];
  _RAND_2393 = {1{`RANDOM}};
  image_2793 = _RAND_2393[3:0];
  _RAND_2394 = {1{`RANDOM}};
  image_2794 = _RAND_2394[3:0];
  _RAND_2395 = {1{`RANDOM}};
  image_2795 = _RAND_2395[3:0];
  _RAND_2396 = {1{`RANDOM}};
  image_2796 = _RAND_2396[3:0];
  _RAND_2397 = {1{`RANDOM}};
  image_2797 = _RAND_2397[3:0];
  _RAND_2398 = {1{`RANDOM}};
  image_2798 = _RAND_2398[3:0];
  _RAND_2399 = {1{`RANDOM}};
  image_2799 = _RAND_2399[3:0];
  _RAND_2400 = {1{`RANDOM}};
  image_2800 = _RAND_2400[3:0];
  _RAND_2401 = {1{`RANDOM}};
  image_2801 = _RAND_2401[3:0];
  _RAND_2402 = {1{`RANDOM}};
  image_2802 = _RAND_2402[3:0];
  _RAND_2403 = {1{`RANDOM}};
  image_2803 = _RAND_2403[3:0];
  _RAND_2404 = {1{`RANDOM}};
  image_2804 = _RAND_2404[3:0];
  _RAND_2405 = {1{`RANDOM}};
  image_2805 = _RAND_2405[3:0];
  _RAND_2406 = {1{`RANDOM}};
  image_2806 = _RAND_2406[3:0];
  _RAND_2407 = {1{`RANDOM}};
  image_2807 = _RAND_2407[3:0];
  _RAND_2408 = {1{`RANDOM}};
  image_2808 = _RAND_2408[3:0];
  _RAND_2409 = {1{`RANDOM}};
  image_2828 = _RAND_2409[3:0];
  _RAND_2410 = {1{`RANDOM}};
  image_2829 = _RAND_2410[3:0];
  _RAND_2411 = {1{`RANDOM}};
  image_2830 = _RAND_2411[3:0];
  _RAND_2412 = {1{`RANDOM}};
  image_2831 = _RAND_2412[3:0];
  _RAND_2413 = {1{`RANDOM}};
  image_2832 = _RAND_2413[3:0];
  _RAND_2414 = {1{`RANDOM}};
  image_2833 = _RAND_2414[3:0];
  _RAND_2415 = {1{`RANDOM}};
  image_2834 = _RAND_2415[3:0];
  _RAND_2416 = {1{`RANDOM}};
  image_2835 = _RAND_2416[3:0];
  _RAND_2417 = {1{`RANDOM}};
  image_2836 = _RAND_2417[3:0];
  _RAND_2418 = {1{`RANDOM}};
  image_2837 = _RAND_2418[3:0];
  _RAND_2419 = {1{`RANDOM}};
  image_2838 = _RAND_2419[3:0];
  _RAND_2420 = {1{`RANDOM}};
  image_2839 = _RAND_2420[3:0];
  _RAND_2421 = {1{`RANDOM}};
  image_2840 = _RAND_2421[3:0];
  _RAND_2422 = {1{`RANDOM}};
  image_2841 = _RAND_2422[3:0];
  _RAND_2423 = {1{`RANDOM}};
  image_2842 = _RAND_2423[3:0];
  _RAND_2424 = {1{`RANDOM}};
  image_2843 = _RAND_2424[3:0];
  _RAND_2425 = {1{`RANDOM}};
  image_2844 = _RAND_2425[3:0];
  _RAND_2426 = {1{`RANDOM}};
  image_2845 = _RAND_2426[3:0];
  _RAND_2427 = {1{`RANDOM}};
  image_2846 = _RAND_2427[3:0];
  _RAND_2428 = {1{`RANDOM}};
  image_2847 = _RAND_2428[3:0];
  _RAND_2429 = {1{`RANDOM}};
  image_2848 = _RAND_2429[3:0];
  _RAND_2430 = {1{`RANDOM}};
  image_2849 = _RAND_2430[3:0];
  _RAND_2431 = {1{`RANDOM}};
  image_2850 = _RAND_2431[3:0];
  _RAND_2432 = {1{`RANDOM}};
  image_2851 = _RAND_2432[3:0];
  _RAND_2433 = {1{`RANDOM}};
  image_2852 = _RAND_2433[3:0];
  _RAND_2434 = {1{`RANDOM}};
  image_2853 = _RAND_2434[3:0];
  _RAND_2435 = {1{`RANDOM}};
  image_2854 = _RAND_2435[3:0];
  _RAND_2436 = {1{`RANDOM}};
  image_2855 = _RAND_2436[3:0];
  _RAND_2437 = {1{`RANDOM}};
  image_2856 = _RAND_2437[3:0];
  _RAND_2438 = {1{`RANDOM}};
  image_2857 = _RAND_2438[3:0];
  _RAND_2439 = {1{`RANDOM}};
  image_2858 = _RAND_2439[3:0];
  _RAND_2440 = {1{`RANDOM}};
  image_2859 = _RAND_2440[3:0];
  _RAND_2441 = {1{`RANDOM}};
  image_2860 = _RAND_2441[3:0];
  _RAND_2442 = {1{`RANDOM}};
  image_2861 = _RAND_2442[3:0];
  _RAND_2443 = {1{`RANDOM}};
  image_2862 = _RAND_2443[3:0];
  _RAND_2444 = {1{`RANDOM}};
  image_2863 = _RAND_2444[3:0];
  _RAND_2445 = {1{`RANDOM}};
  image_2864 = _RAND_2445[3:0];
  _RAND_2446 = {1{`RANDOM}};
  image_2865 = _RAND_2446[3:0];
  _RAND_2447 = {1{`RANDOM}};
  image_2866 = _RAND_2447[3:0];
  _RAND_2448 = {1{`RANDOM}};
  image_2867 = _RAND_2448[3:0];
  _RAND_2449 = {1{`RANDOM}};
  image_2868 = _RAND_2449[3:0];
  _RAND_2450 = {1{`RANDOM}};
  image_2869 = _RAND_2450[3:0];
  _RAND_2451 = {1{`RANDOM}};
  image_2870 = _RAND_2451[3:0];
  _RAND_2452 = {1{`RANDOM}};
  image_2871 = _RAND_2452[3:0];
  _RAND_2453 = {1{`RANDOM}};
  image_2895 = _RAND_2453[3:0];
  _RAND_2454 = {1{`RANDOM}};
  image_2896 = _RAND_2454[3:0];
  _RAND_2455 = {1{`RANDOM}};
  image_2897 = _RAND_2455[3:0];
  _RAND_2456 = {1{`RANDOM}};
  image_2898 = _RAND_2456[3:0];
  _RAND_2457 = {1{`RANDOM}};
  image_2899 = _RAND_2457[3:0];
  _RAND_2458 = {1{`RANDOM}};
  image_2900 = _RAND_2458[3:0];
  _RAND_2459 = {1{`RANDOM}};
  image_2901 = _RAND_2459[3:0];
  _RAND_2460 = {1{`RANDOM}};
  image_2902 = _RAND_2460[3:0];
  _RAND_2461 = {1{`RANDOM}};
  image_2903 = _RAND_2461[3:0];
  _RAND_2462 = {1{`RANDOM}};
  image_2904 = _RAND_2462[3:0];
  _RAND_2463 = {1{`RANDOM}};
  image_2905 = _RAND_2463[3:0];
  _RAND_2464 = {1{`RANDOM}};
  image_2906 = _RAND_2464[3:0];
  _RAND_2465 = {1{`RANDOM}};
  image_2907 = _RAND_2465[3:0];
  _RAND_2466 = {1{`RANDOM}};
  image_2908 = _RAND_2466[3:0];
  _RAND_2467 = {1{`RANDOM}};
  image_2909 = _RAND_2467[3:0];
  _RAND_2468 = {1{`RANDOM}};
  image_2910 = _RAND_2468[3:0];
  _RAND_2469 = {1{`RANDOM}};
  image_2911 = _RAND_2469[3:0];
  _RAND_2470 = {1{`RANDOM}};
  image_2912 = _RAND_2470[3:0];
  _RAND_2471 = {1{`RANDOM}};
  image_2913 = _RAND_2471[3:0];
  _RAND_2472 = {1{`RANDOM}};
  image_2914 = _RAND_2472[3:0];
  _RAND_2473 = {1{`RANDOM}};
  image_2915 = _RAND_2473[3:0];
  _RAND_2474 = {1{`RANDOM}};
  image_2916 = _RAND_2474[3:0];
  _RAND_2475 = {1{`RANDOM}};
  image_2917 = _RAND_2475[3:0];
  _RAND_2476 = {1{`RANDOM}};
  image_2918 = _RAND_2476[3:0];
  _RAND_2477 = {1{`RANDOM}};
  image_2919 = _RAND_2477[3:0];
  _RAND_2478 = {1{`RANDOM}};
  image_2920 = _RAND_2478[3:0];
  _RAND_2479 = {1{`RANDOM}};
  image_2921 = _RAND_2479[3:0];
  _RAND_2480 = {1{`RANDOM}};
  image_2922 = _RAND_2480[3:0];
  _RAND_2481 = {1{`RANDOM}};
  image_2923 = _RAND_2481[3:0];
  _RAND_2482 = {1{`RANDOM}};
  image_2924 = _RAND_2482[3:0];
  _RAND_2483 = {1{`RANDOM}};
  image_2925 = _RAND_2483[3:0];
  _RAND_2484 = {1{`RANDOM}};
  image_2926 = _RAND_2484[3:0];
  _RAND_2485 = {1{`RANDOM}};
  image_2927 = _RAND_2485[3:0];
  _RAND_2486 = {1{`RANDOM}};
  image_2928 = _RAND_2486[3:0];
  _RAND_2487 = {1{`RANDOM}};
  image_2929 = _RAND_2487[3:0];
  _RAND_2488 = {1{`RANDOM}};
  image_2930 = _RAND_2488[3:0];
  _RAND_2489 = {1{`RANDOM}};
  image_2931 = _RAND_2489[3:0];
  _RAND_2490 = {1{`RANDOM}};
  image_2932 = _RAND_2490[3:0];
  _RAND_2491 = {1{`RANDOM}};
  image_2933 = _RAND_2491[3:0];
  _RAND_2492 = {1{`RANDOM}};
  image_2934 = _RAND_2492[3:0];
  _RAND_2493 = {1{`RANDOM}};
  image_2965 = _RAND_2493[3:0];
  _RAND_2494 = {1{`RANDOM}};
  image_2966 = _RAND_2494[3:0];
  _RAND_2495 = {1{`RANDOM}};
  image_2967 = _RAND_2495[3:0];
  _RAND_2496 = {1{`RANDOM}};
  image_2968 = _RAND_2496[3:0];
  _RAND_2497 = {1{`RANDOM}};
  image_2969 = _RAND_2497[3:0];
  _RAND_2498 = {1{`RANDOM}};
  image_2970 = _RAND_2498[3:0];
  _RAND_2499 = {1{`RANDOM}};
  image_2971 = _RAND_2499[3:0];
  _RAND_2500 = {1{`RANDOM}};
  image_2972 = _RAND_2500[3:0];
  _RAND_2501 = {1{`RANDOM}};
  image_2973 = _RAND_2501[3:0];
  _RAND_2502 = {1{`RANDOM}};
  image_2974 = _RAND_2502[3:0];
  _RAND_2503 = {1{`RANDOM}};
  image_2975 = _RAND_2503[3:0];
  _RAND_2504 = {1{`RANDOM}};
  image_2976 = _RAND_2504[3:0];
  _RAND_2505 = {1{`RANDOM}};
  image_2977 = _RAND_2505[3:0];
  _RAND_2506 = {1{`RANDOM}};
  image_2978 = _RAND_2506[3:0];
  _RAND_2507 = {1{`RANDOM}};
  image_2979 = _RAND_2507[3:0];
  _RAND_2508 = {1{`RANDOM}};
  image_2980 = _RAND_2508[3:0];
  _RAND_2509 = {1{`RANDOM}};
  image_2981 = _RAND_2509[3:0];
  _RAND_2510 = {1{`RANDOM}};
  image_2982 = _RAND_2510[3:0];
  _RAND_2511 = {1{`RANDOM}};
  image_2983 = _RAND_2511[3:0];
  _RAND_2512 = {1{`RANDOM}};
  image_2984 = _RAND_2512[3:0];
  _RAND_2513 = {1{`RANDOM}};
  image_2985 = _RAND_2513[3:0];
  _RAND_2514 = {1{`RANDOM}};
  image_2986 = _RAND_2514[3:0];
  _RAND_2515 = {1{`RANDOM}};
  image_2987 = _RAND_2515[3:0];
  _RAND_2516 = {1{`RANDOM}};
  image_2988 = _RAND_2516[3:0];
  _RAND_2517 = {1{`RANDOM}};
  image_2989 = _RAND_2517[3:0];
  _RAND_2518 = {1{`RANDOM}};
  image_2990 = _RAND_2518[3:0];
  _RAND_2519 = {1{`RANDOM}};
  image_2991 = _RAND_2519[3:0];
  _RAND_2520 = {1{`RANDOM}};
  image_2992 = _RAND_2520[3:0];
  _RAND_2521 = {1{`RANDOM}};
  image_2993 = _RAND_2521[3:0];
  _RAND_2522 = {1{`RANDOM}};
  image_2994 = _RAND_2522[3:0];
  _RAND_2523 = {1{`RANDOM}};
  image_2995 = _RAND_2523[3:0];
  _RAND_2524 = {1{`RANDOM}};
  image_2996 = _RAND_2524[3:0];
  _RAND_2525 = {1{`RANDOM}};
  image_3035 = _RAND_2525[3:0];
  _RAND_2526 = {1{`RANDOM}};
  image_3036 = _RAND_2526[3:0];
  _RAND_2527 = {1{`RANDOM}};
  image_3037 = _RAND_2527[3:0];
  _RAND_2528 = {1{`RANDOM}};
  image_3038 = _RAND_2528[3:0];
  _RAND_2529 = {1{`RANDOM}};
  image_3039 = _RAND_2529[3:0];
  _RAND_2530 = {1{`RANDOM}};
  image_3040 = _RAND_2530[3:0];
  _RAND_2531 = {1{`RANDOM}};
  image_3041 = _RAND_2531[3:0];
  _RAND_2532 = {1{`RANDOM}};
  image_3042 = _RAND_2532[3:0];
  _RAND_2533 = {1{`RANDOM}};
  image_3043 = _RAND_2533[3:0];
  _RAND_2534 = {1{`RANDOM}};
  image_3044 = _RAND_2534[3:0];
  _RAND_2535 = {1{`RANDOM}};
  image_3045 = _RAND_2535[3:0];
  _RAND_2536 = {1{`RANDOM}};
  image_3046 = _RAND_2536[3:0];
  _RAND_2537 = {1{`RANDOM}};
  image_3047 = _RAND_2537[3:0];
  _RAND_2538 = {1{`RANDOM}};
  image_3048 = _RAND_2538[3:0];
  _RAND_2539 = {1{`RANDOM}};
  image_3049 = _RAND_2539[3:0];
  _RAND_2540 = {1{`RANDOM}};
  image_3050 = _RAND_2540[3:0];
  _RAND_2541 = {1{`RANDOM}};
  image_3051 = _RAND_2541[3:0];
  _RAND_2542 = {1{`RANDOM}};
  image_3052 = _RAND_2542[3:0];
  _RAND_2543 = {1{`RANDOM}};
  image_3053 = _RAND_2543[3:0];
  _RAND_2544 = {1{`RANDOM}};
  image_3054 = _RAND_2544[3:0];
  _RAND_2545 = {1{`RANDOM}};
  image_3055 = _RAND_2545[3:0];
  _RAND_2546 = {1{`RANDOM}};
  image_3056 = _RAND_2546[3:0];
  _RAND_2547 = {1{`RANDOM}};
  kernelCounter = _RAND_2547[3:0];
  _RAND_2548 = {1{`RANDOM}};
  imageCounterX = _RAND_2548[1:0];
  _RAND_2549 = {1{`RANDOM}};
  imageCounterY = _RAND_2549[1:0];
  _RAND_2550 = {1{`RANDOM}};
  pixelIndex = _RAND_2550[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      image_12 <= 4'h0;
    end else begin
      image_12 <= 4'h1;
    end
    if (reset) begin
      image_14 <= 4'h0;
    end else begin
      image_14 <= 4'h2;
    end
    if (reset) begin
      image_15 <= 4'h0;
    end else begin
      image_15 <= 4'h4;
    end
    if (reset) begin
      image_16 <= 4'h0;
    end else begin
      image_16 <= 4'h4;
    end
    if (reset) begin
      image_17 <= 4'h0;
    end else begin
      image_17 <= 4'h5;
    end
    if (reset) begin
      image_18 <= 4'h0;
    end else begin
      image_18 <= 4'h5;
    end
    if (reset) begin
      image_19 <= 4'h0;
    end else begin
      image_19 <= 4'h5;
    end
    if (reset) begin
      image_20 <= 4'h0;
    end else begin
      image_20 <= 4'h5;
    end
    if (reset) begin
      image_21 <= 4'h0;
    end else begin
      image_21 <= 4'h5;
    end
    if (reset) begin
      image_22 <= 4'h0;
    end else begin
      image_22 <= 4'h5;
    end
    if (reset) begin
      image_23 <= 4'h0;
    end else begin
      image_23 <= 4'h3;
    end
    if (reset) begin
      image_35 <= 4'h0;
    end else begin
      image_35 <= 4'h1;
    end
    if (reset) begin
      image_36 <= 4'h0;
    end else begin
      image_36 <= 4'h3;
    end
    if (reset) begin
      image_37 <= 4'h0;
    end else begin
      image_37 <= 4'h4;
    end
    if (reset) begin
      image_38 <= 4'h0;
    end else begin
      image_38 <= 4'h4;
    end
    if (reset) begin
      image_39 <= 4'h0;
    end else begin
      image_39 <= 4'h4;
    end
    if (reset) begin
      image_40 <= 4'h0;
    end else begin
      image_40 <= 4'h4;
    end
    if (reset) begin
      image_41 <= 4'h0;
    end else begin
      image_41 <= 4'h4;
    end
    if (reset) begin
      image_42 <= 4'h0;
    end else begin
      image_42 <= 4'h2;
    end
    if (reset) begin
      image_75 <= 4'h0;
    end else begin
      image_75 <= 4'h3;
    end
    if (reset) begin
      image_76 <= 4'h0;
    end else begin
      image_76 <= 4'h5;
    end
    if (reset) begin
      image_77 <= 4'h0;
    end else begin
      image_77 <= 4'h6;
    end
    if (reset) begin
      image_78 <= 4'h0;
    end else begin
      image_78 <= 4'h6;
    end
    if (reset) begin
      image_79 <= 4'h0;
    end else begin
      image_79 <= 4'h6;
    end
    if (reset) begin
      image_80 <= 4'h0;
    end else begin
      image_80 <= 4'h6;
    end
    if (reset) begin
      image_81 <= 4'h0;
    end else begin
      image_81 <= 4'h6;
    end
    if (reset) begin
      image_82 <= 4'h0;
    end else begin
      image_82 <= 4'h6;
    end
    if (reset) begin
      image_83 <= 4'h0;
    end else begin
      image_83 <= 4'h6;
    end
    if (reset) begin
      image_84 <= 4'h0;
    end else begin
      image_84 <= 4'h6;
    end
    if (reset) begin
      image_85 <= 4'h0;
    end else begin
      image_85 <= 4'h6;
    end
    if (reset) begin
      image_86 <= 4'h0;
    end else begin
      image_86 <= 4'h6;
    end
    if (reset) begin
      image_87 <= 4'h0;
    end else begin
      image_87 <= 4'h6;
    end
    if (reset) begin
      image_88 <= 4'h0;
    end else begin
      image_88 <= 4'h6;
    end
    if (reset) begin
      image_89 <= 4'h0;
    end else begin
      image_89 <= 4'h5;
    end
    if (reset) begin
      image_90 <= 4'h0;
    end else begin
      image_90 <= 4'h3;
    end
    if (reset) begin
      image_93 <= 4'h0;
    end else begin
      image_93 <= 4'h1;
    end
    if (reset) begin
      image_95 <= 4'h0;
    end else begin
      image_95 <= 4'h3;
    end
    if (reset) begin
      image_96 <= 4'h0;
    end else begin
      image_96 <= 4'h4;
    end
    if (reset) begin
      image_97 <= 4'h0;
    end else begin
      image_97 <= 4'h5;
    end
    if (reset) begin
      image_98 <= 4'h0;
    end else begin
      image_98 <= 4'h6;
    end
    if (reset) begin
      image_99 <= 4'h0;
    end else begin
      image_99 <= 4'h6;
    end
    if (reset) begin
      image_100 <= 4'h0;
    end else begin
      image_100 <= 4'h6;
    end
    if (reset) begin
      image_101 <= 4'h0;
    end else begin
      image_101 <= 4'h6;
    end
    if (reset) begin
      image_102 <= 4'h0;
    end else begin
      image_102 <= 4'h6;
    end
    if (reset) begin
      image_103 <= 4'h0;
    end else begin
      image_103 <= 4'h6;
    end
    if (reset) begin
      image_104 <= 4'h0;
    end else begin
      image_104 <= 4'h6;
    end
    if (reset) begin
      image_105 <= 4'h0;
    end else begin
      image_105 <= 4'h6;
    end
    if (reset) begin
      image_106 <= 4'h0;
    end else begin
      image_106 <= 4'h6;
    end
    if (reset) begin
      image_107 <= 4'h0;
    end else begin
      image_107 <= 4'h4;
    end
    if (reset) begin
      image_108 <= 4'h0;
    end else begin
      image_108 <= 4'h3;
    end
    if (reset) begin
      image_136 <= 4'h0;
    end else begin
      image_136 <= 4'h1;
    end
    if (reset) begin
      image_137 <= 4'h0;
    end else begin
      image_137 <= 4'h2;
    end
    if (reset) begin
      image_138 <= 4'h0;
    end else begin
      image_138 <= 4'h5;
    end
    if (reset) begin
      image_139 <= 4'h0;
    end else begin
      image_139 <= 4'h6;
    end
    if (reset) begin
      image_140 <= 4'h0;
    end else begin
      image_140 <= 4'h6;
    end
    if (reset) begin
      image_141 <= 4'h0;
    end else begin
      image_141 <= 4'h6;
    end
    if (reset) begin
      image_142 <= 4'h0;
    end else begin
      image_142 <= 4'h6;
    end
    if (reset) begin
      image_143 <= 4'h0;
    end else begin
      image_143 <= 4'h6;
    end
    if (reset) begin
      image_144 <= 4'h0;
    end else begin
      image_144 <= 4'h6;
    end
    if (reset) begin
      image_145 <= 4'h0;
    end else begin
      image_145 <= 4'h6;
    end
    if (reset) begin
      image_146 <= 4'h0;
    end else begin
      image_146 <= 4'h6;
    end
    if (reset) begin
      image_147 <= 4'h0;
    end else begin
      image_147 <= 4'h6;
    end
    if (reset) begin
      image_148 <= 4'h0;
    end else begin
      image_148 <= 4'h6;
    end
    if (reset) begin
      image_149 <= 4'h0;
    end else begin
      image_149 <= 4'h6;
    end
    if (reset) begin
      image_150 <= 4'h0;
    end else begin
      image_150 <= 4'h5;
    end
    if (reset) begin
      image_151 <= 4'h0;
    end else begin
      image_151 <= 4'h5;
    end
    if (reset) begin
      image_152 <= 4'h0;
    end else begin
      image_152 <= 4'h5;
    end
    if (reset) begin
      image_153 <= 4'h0;
    end else begin
      image_153 <= 4'h4;
    end
    if (reset) begin
      image_154 <= 4'h0;
    end else begin
      image_154 <= 4'h4;
    end
    if (reset) begin
      image_155 <= 4'h0;
    end else begin
      image_155 <= 4'h3;
    end
    if (reset) begin
      image_157 <= 4'h0;
    end else begin
      image_157 <= 4'h1;
    end
    if (reset) begin
      image_158 <= 4'h0;
    end else begin
      image_158 <= 4'h4;
    end
    if (reset) begin
      image_159 <= 4'h0;
    end else begin
      image_159 <= 4'h6;
    end
    if (reset) begin
      image_160 <= 4'h0;
    end else begin
      image_160 <= 4'h6;
    end
    if (reset) begin
      image_161 <= 4'h0;
    end else begin
      image_161 <= 4'h6;
    end
    if (reset) begin
      image_162 <= 4'h0;
    end else begin
      image_162 <= 4'h6;
    end
    if (reset) begin
      image_163 <= 4'h0;
    end else begin
      image_163 <= 4'h6;
    end
    if (reset) begin
      image_164 <= 4'h0;
    end else begin
      image_164 <= 4'h6;
    end
    if (reset) begin
      image_165 <= 4'h0;
    end else begin
      image_165 <= 4'h6;
    end
    if (reset) begin
      image_166 <= 4'h0;
    end else begin
      image_166 <= 4'h6;
    end
    if (reset) begin
      image_167 <= 4'h0;
    end else begin
      image_167 <= 4'h6;
    end
    if (reset) begin
      image_168 <= 4'h0;
    end else begin
      image_168 <= 4'h6;
    end
    if (reset) begin
      image_169 <= 4'h0;
    end else begin
      image_169 <= 4'h6;
    end
    if (reset) begin
      image_170 <= 4'h0;
    end else begin
      image_170 <= 4'h5;
    end
    if (reset) begin
      image_171 <= 4'h0;
    end else begin
      image_171 <= 4'h4;
    end
    if (reset) begin
      image_172 <= 4'h0;
    end else begin
      image_172 <= 4'h4;
    end
    if (reset) begin
      image_173 <= 4'h0;
    end else begin
      image_173 <= 4'h5;
    end
    if (reset) begin
      image_174 <= 4'h0;
    end else begin
      image_174 <= 4'h5;
    end
    if (reset) begin
      image_175 <= 4'h0;
    end else begin
      image_175 <= 4'h5;
    end
    if (reset) begin
      image_176 <= 4'h0;
    end else begin
      image_176 <= 4'h5;
    end
    if (reset) begin
      image_177 <= 4'h0;
    end else begin
      image_177 <= 4'h5;
    end
    if (reset) begin
      image_178 <= 4'h0;
    end else begin
      image_178 <= 4'h3;
    end
    if (reset) begin
      image_179 <= 4'h0;
    end else begin
      image_179 <= 4'h1;
    end
    if (reset) begin
      image_199 <= 4'h0;
    end else begin
      image_199 <= 4'h1;
    end
    if (reset) begin
      image_200 <= 4'h0;
    end else begin
      image_200 <= 4'h4;
    end
    if (reset) begin
      image_201 <= 4'h0;
    end else begin
      image_201 <= 4'h6;
    end
    if (reset) begin
      image_202 <= 4'h0;
    end else begin
      image_202 <= 4'h6;
    end
    if (reset) begin
      image_203 <= 4'h0;
    end else begin
      image_203 <= 4'h6;
    end
    if (reset) begin
      image_204 <= 4'h0;
    end else begin
      image_204 <= 4'h6;
    end
    if (reset) begin
      image_205 <= 4'h0;
    end else begin
      image_205 <= 4'h6;
    end
    if (reset) begin
      image_206 <= 4'h0;
    end else begin
      image_206 <= 4'h6;
    end
    if (reset) begin
      image_207 <= 4'h0;
    end else begin
      image_207 <= 4'h6;
    end
    if (reset) begin
      image_208 <= 4'h0;
    end else begin
      image_208 <= 4'h5;
    end
    if (reset) begin
      image_209 <= 4'h0;
    end else begin
      image_209 <= 4'h4;
    end
    if (reset) begin
      image_210 <= 4'h0;
    end else begin
      image_210 <= 4'h4;
    end
    if (reset) begin
      image_211 <= 4'h0;
    end else begin
      image_211 <= 4'h4;
    end
    if (reset) begin
      image_212 <= 4'h0;
    end else begin
      image_212 <= 4'h5;
    end
    if (reset) begin
      image_213 <= 4'h0;
    end else begin
      image_213 <= 4'h5;
    end
    if (reset) begin
      image_214 <= 4'h0;
    end else begin
      image_214 <= 4'h6;
    end
    if (reset) begin
      image_215 <= 4'h0;
    end else begin
      image_215 <= 4'h6;
    end
    if (reset) begin
      image_216 <= 4'h0;
    end else begin
      image_216 <= 4'h6;
    end
    if (reset) begin
      image_217 <= 4'h0;
    end else begin
      image_217 <= 4'h6;
    end
    if (reset) begin
      image_218 <= 4'h0;
    end else begin
      image_218 <= 4'h6;
    end
    if (reset) begin
      image_219 <= 4'h0;
    end else begin
      image_219 <= 4'h6;
    end
    if (reset) begin
      image_220 <= 4'h0;
    end else begin
      image_220 <= 4'h6;
    end
    if (reset) begin
      image_221 <= 4'h0;
    end else begin
      image_221 <= 4'h6;
    end
    if (reset) begin
      image_222 <= 4'h0;
    end else begin
      image_222 <= 4'h6;
    end
    if (reset) begin
      image_223 <= 4'h0;
    end else begin
      image_223 <= 4'h5;
    end
    if (reset) begin
      image_224 <= 4'h0;
    end else begin
      image_224 <= 4'h4;
    end
    if (reset) begin
      image_225 <= 4'h0;
    end else begin
      image_225 <= 4'h5;
    end
    if (reset) begin
      image_226 <= 4'h0;
    end else begin
      image_226 <= 4'h6;
    end
    if (reset) begin
      image_227 <= 4'h0;
    end else begin
      image_227 <= 4'h6;
    end
    if (reset) begin
      image_228 <= 4'h0;
    end else begin
      image_228 <= 4'h6;
    end
    if (reset) begin
      image_229 <= 4'h0;
    end else begin
      image_229 <= 4'h6;
    end
    if (reset) begin
      image_230 <= 4'h0;
    end else begin
      image_230 <= 4'h6;
    end
    if (reset) begin
      image_231 <= 4'h0;
    end else begin
      image_231 <= 4'h6;
    end
    if (reset) begin
      image_232 <= 4'h0;
    end else begin
      image_232 <= 4'h5;
    end
    if (reset) begin
      image_233 <= 4'h0;
    end else begin
      image_233 <= 4'h5;
    end
    if (reset) begin
      image_234 <= 4'h0;
    end else begin
      image_234 <= 4'h6;
    end
    if (reset) begin
      image_235 <= 4'h0;
    end else begin
      image_235 <= 4'h6;
    end
    if (reset) begin
      image_236 <= 4'h0;
    end else begin
      image_236 <= 4'h6;
    end
    if (reset) begin
      image_237 <= 4'h0;
    end else begin
      image_237 <= 4'h6;
    end
    if (reset) begin
      image_238 <= 4'h0;
    end else begin
      image_238 <= 4'h5;
    end
    if (reset) begin
      image_239 <= 4'h0;
    end else begin
      image_239 <= 4'h4;
    end
    if (reset) begin
      image_240 <= 4'h0;
    end else begin
      image_240 <= 4'h4;
    end
    if (reset) begin
      image_241 <= 4'h0;
    end else begin
      image_241 <= 4'h4;
    end
    if (reset) begin
      image_242 <= 4'h0;
    end else begin
      image_242 <= 4'h5;
    end
    if (reset) begin
      image_243 <= 4'h0;
    end else begin
      image_243 <= 4'h5;
    end
    if (reset) begin
      image_244 <= 4'h0;
    end else begin
      image_244 <= 4'h5;
    end
    if (reset) begin
      image_245 <= 4'h0;
    end else begin
      image_245 <= 4'h4;
    end
    if (reset) begin
      image_246 <= 4'h0;
    end else begin
      image_246 <= 4'h3;
    end
    if (reset) begin
      image_262 <= 4'h0;
    end else begin
      image_262 <= 4'h2;
    end
    if (reset) begin
      image_263 <= 4'h0;
    end else begin
      image_263 <= 4'h5;
    end
    if (reset) begin
      image_264 <= 4'h0;
    end else begin
      image_264 <= 4'h6;
    end
    if (reset) begin
      image_265 <= 4'h0;
    end else begin
      image_265 <= 4'h6;
    end
    if (reset) begin
      image_266 <= 4'h0;
    end else begin
      image_266 <= 4'h6;
    end
    if (reset) begin
      image_267 <= 4'h0;
    end else begin
      image_267 <= 4'h6;
    end
    if (reset) begin
      image_268 <= 4'h0;
    end else begin
      image_268 <= 4'h6;
    end
    if (reset) begin
      image_269 <= 4'h0;
    end else begin
      image_269 <= 4'h5;
    end
    if (reset) begin
      image_270 <= 4'h0;
    end else begin
      image_270 <= 4'h4;
    end
    if (reset) begin
      image_271 <= 4'h0;
    end else begin
      image_271 <= 4'h5;
    end
    if (reset) begin
      image_272 <= 4'h0;
    end else begin
      image_272 <= 4'h6;
    end
    if (reset) begin
      image_273 <= 4'h0;
    end else begin
      image_273 <= 4'h6;
    end
    if (reset) begin
      image_274 <= 4'h0;
    end else begin
      image_274 <= 4'h6;
    end
    if (reset) begin
      image_275 <= 4'h0;
    end else begin
      image_275 <= 4'h6;
    end
    if (reset) begin
      image_276 <= 4'h0;
    end else begin
      image_276 <= 4'h6;
    end
    if (reset) begin
      image_277 <= 4'h0;
    end else begin
      image_277 <= 4'h6;
    end
    if (reset) begin
      image_278 <= 4'h0;
    end else begin
      image_278 <= 4'h6;
    end
    if (reset) begin
      image_279 <= 4'h0;
    end else begin
      image_279 <= 4'h6;
    end
    if (reset) begin
      image_280 <= 4'h0;
    end else begin
      image_280 <= 4'h5;
    end
    if (reset) begin
      image_281 <= 4'h0;
    end else begin
      image_281 <= 4'h4;
    end
    if (reset) begin
      image_282 <= 4'h0;
    end else begin
      image_282 <= 4'h5;
    end
    if (reset) begin
      image_283 <= 4'h0;
    end else begin
      image_283 <= 4'h4;
    end
    if (reset) begin
      image_284 <= 4'h0;
    end else begin
      image_284 <= 4'h4;
    end
    if (reset) begin
      image_285 <= 4'h0;
    end else begin
      image_285 <= 4'h4;
    end
    if (reset) begin
      image_286 <= 4'h0;
    end else begin
      image_286 <= 4'h4;
    end
    if (reset) begin
      image_287 <= 4'h0;
    end else begin
      image_287 <= 4'h4;
    end
    if (reset) begin
      image_288 <= 4'h0;
    end else begin
      image_288 <= 4'h4;
    end
    if (reset) begin
      image_289 <= 4'h0;
    end else begin
      image_289 <= 4'h2;
    end
    if (reset) begin
      image_290 <= 4'h0;
    end else begin
      image_290 <= 4'h3;
    end
    if (reset) begin
      image_291 <= 4'h0;
    end else begin
      image_291 <= 4'h4;
    end
    if (reset) begin
      image_292 <= 4'h0;
    end else begin
      image_292 <= 4'h5;
    end
    if (reset) begin
      image_293 <= 4'h0;
    end else begin
      image_293 <= 4'h6;
    end
    if (reset) begin
      image_294 <= 4'h0;
    end else begin
      image_294 <= 4'h6;
    end
    if (reset) begin
      image_295 <= 4'h0;
    end else begin
      image_295 <= 4'h6;
    end
    if (reset) begin
      image_296 <= 4'h0;
    end else begin
      image_296 <= 4'h6;
    end
    if (reset) begin
      image_297 <= 4'h0;
    end else begin
      image_297 <= 4'h6;
    end
    if (reset) begin
      image_298 <= 4'h0;
    end else begin
      image_298 <= 4'h6;
    end
    if (reset) begin
      image_299 <= 4'h0;
    end else begin
      image_299 <= 4'h5;
    end
    if (reset) begin
      image_300 <= 4'h0;
    end else begin
      image_300 <= 4'h4;
    end
    if (reset) begin
      image_301 <= 4'h0;
    end else begin
      image_301 <= 4'h5;
    end
    if (reset) begin
      image_302 <= 4'h0;
    end else begin
      image_302 <= 4'h6;
    end
    if (reset) begin
      image_303 <= 4'h0;
    end else begin
      image_303 <= 4'h6;
    end
    if (reset) begin
      image_304 <= 4'h0;
    end else begin
      image_304 <= 4'h6;
    end
    if (reset) begin
      image_305 <= 4'h0;
    end else begin
      image_305 <= 4'h6;
    end
    if (reset) begin
      image_306 <= 4'h0;
    end else begin
      image_306 <= 4'h6;
    end
    if (reset) begin
      image_307 <= 4'h0;
    end else begin
      image_307 <= 4'h6;
    end
    if (reset) begin
      image_308 <= 4'h0;
    end else begin
      image_308 <= 4'h6;
    end
    if (reset) begin
      image_309 <= 4'h0;
    end else begin
      image_309 <= 4'h6;
    end
    if (reset) begin
      image_310 <= 4'h0;
    end else begin
      image_310 <= 4'h6;
    end
    if (reset) begin
      image_311 <= 4'h0;
    end else begin
      image_311 <= 4'h6;
    end
    if (reset) begin
      image_312 <= 4'h0;
    end else begin
      image_312 <= 4'h5;
    end
    if (reset) begin
      image_313 <= 4'h0;
    end else begin
      image_313 <= 4'h3;
    end
    if (reset) begin
      image_314 <= 4'h0;
    end else begin
      image_314 <= 4'h1;
    end
    if (reset) begin
      image_315 <= 4'h0;
    end else begin
      image_315 <= 4'h1;
    end
    if (reset) begin
      image_325 <= 4'h0;
    end else begin
      image_325 <= 4'h2;
    end
    if (reset) begin
      image_326 <= 4'h0;
    end else begin
      image_326 <= 4'h5;
    end
    if (reset) begin
      image_327 <= 4'h0;
    end else begin
      image_327 <= 4'h6;
    end
    if (reset) begin
      image_328 <= 4'h0;
    end else begin
      image_328 <= 4'h6;
    end
    if (reset) begin
      image_329 <= 4'h0;
    end else begin
      image_329 <= 4'h6;
    end
    if (reset) begin
      image_330 <= 4'h0;
    end else begin
      image_330 <= 4'h6;
    end
    if (reset) begin
      image_331 <= 4'h0;
    end else begin
      image_331 <= 4'h5;
    end
    if (reset) begin
      image_332 <= 4'h0;
    end else begin
      image_332 <= 4'h4;
    end
    if (reset) begin
      image_333 <= 4'h0;
    end else begin
      image_333 <= 4'h6;
    end
    if (reset) begin
      image_334 <= 4'h0;
    end else begin
      image_334 <= 4'h6;
    end
    if (reset) begin
      image_335 <= 4'h0;
    end else begin
      image_335 <= 4'h6;
    end
    if (reset) begin
      image_336 <= 4'h0;
    end else begin
      image_336 <= 4'h6;
    end
    if (reset) begin
      image_337 <= 4'h0;
    end else begin
      image_337 <= 4'h6;
    end
    if (reset) begin
      image_338 <= 4'h0;
    end else begin
      image_338 <= 4'h6;
    end
    if (reset) begin
      image_339 <= 4'h0;
    end else begin
      image_339 <= 4'h6;
    end
    if (reset) begin
      image_340 <= 4'h0;
    end else begin
      image_340 <= 4'h5;
    end
    if (reset) begin
      image_341 <= 4'h0;
    end else begin
      image_341 <= 4'h4;
    end
    if (reset) begin
      image_342 <= 4'h0;
    end else begin
      image_342 <= 4'h4;
    end
    if (reset) begin
      image_343 <= 4'h0;
    end else begin
      image_343 <= 4'h5;
    end
    if (reset) begin
      image_344 <= 4'h0;
    end else begin
      image_344 <= 4'h6;
    end
    if (reset) begin
      image_345 <= 4'h0;
    end else begin
      image_345 <= 4'h6;
    end
    if (reset) begin
      image_346 <= 4'h0;
    end else begin
      image_346 <= 4'h5;
    end
    if (reset) begin
      image_347 <= 4'h0;
    end else begin
      image_347 <= 4'h5;
    end
    if (reset) begin
      image_348 <= 4'h0;
    end else begin
      image_348 <= 4'h5;
    end
    if (reset) begin
      image_349 <= 4'h0;
    end else begin
      image_349 <= 4'h5;
    end
    if (reset) begin
      image_350 <= 4'h0;
    end else begin
      image_350 <= 4'h5;
    end
    if (reset) begin
      image_351 <= 4'h0;
    end else begin
      image_351 <= 4'h5;
    end
    if (reset) begin
      image_352 <= 4'h0;
    end else begin
      image_352 <= 4'h5;
    end
    if (reset) begin
      image_353 <= 4'h0;
    end else begin
      image_353 <= 4'h6;
    end
    if (reset) begin
      image_354 <= 4'h0;
    end else begin
      image_354 <= 4'h6;
    end
    if (reset) begin
      image_355 <= 4'h0;
    end else begin
      image_355 <= 4'h6;
    end
    if (reset) begin
      image_356 <= 4'h0;
    end else begin
      image_356 <= 4'h5;
    end
    if (reset) begin
      image_357 <= 4'h0;
    end else begin
      image_357 <= 4'h4;
    end
    if (reset) begin
      image_358 <= 4'h0;
    end else begin
      image_358 <= 4'h4;
    end
    if (reset) begin
      image_359 <= 4'h0;
    end else begin
      image_359 <= 4'h6;
    end
    if (reset) begin
      image_360 <= 4'h0;
    end else begin
      image_360 <= 4'h6;
    end
    if (reset) begin
      image_361 <= 4'h0;
    end else begin
      image_361 <= 4'h4;
    end
    if (reset) begin
      image_362 <= 4'h0;
    end else begin
      image_362 <= 4'h4;
    end
    if (reset) begin
      image_363 <= 4'h0;
    end else begin
      image_363 <= 4'h6;
    end
    if (reset) begin
      image_364 <= 4'h0;
    end else begin
      image_364 <= 4'h6;
    end
    if (reset) begin
      image_365 <= 4'h0;
    end else begin
      image_365 <= 4'h5;
    end
    if (reset) begin
      image_366 <= 4'h0;
    end else begin
      image_366 <= 4'h5;
    end
    if (reset) begin
      image_367 <= 4'h0;
    end else begin
      image_367 <= 4'h8;
    end
    if (reset) begin
      image_368 <= 4'h0;
    end else begin
      image_368 <= 4'ha;
    end
    if (reset) begin
      image_369 <= 4'h0;
    end else begin
      image_369 <= 4'hb;
    end
    if (reset) begin
      image_370 <= 4'h0;
    end else begin
      image_370 <= 4'hb;
    end
    if (reset) begin
      image_371 <= 4'h0;
    end else begin
      image_371 <= 4'hb;
    end
    if (reset) begin
      image_372 <= 4'h0;
    end else begin
      image_372 <= 4'hb;
    end
    if (reset) begin
      image_373 <= 4'h0;
    end else begin
      image_373 <= 4'ha;
    end
    if (reset) begin
      image_374 <= 4'h0;
    end else begin
      image_374 <= 4'h9;
    end
    if (reset) begin
      image_375 <= 4'h0;
    end else begin
      image_375 <= 4'h8;
    end
    if (reset) begin
      image_376 <= 4'h0;
    end else begin
      image_376 <= 4'h5;
    end
    if (reset) begin
      image_377 <= 4'h0;
    end else begin
      image_377 <= 4'h5;
    end
    if (reset) begin
      image_378 <= 4'h0;
    end else begin
      image_378 <= 4'h5;
    end
    if (reset) begin
      image_379 <= 4'h0;
    end else begin
      image_379 <= 4'h3;
    end
    if (reset) begin
      image_388 <= 4'h0;
    end else begin
      image_388 <= 4'h3;
    end
    if (reset) begin
      image_389 <= 4'h0;
    end else begin
      image_389 <= 4'h5;
    end
    if (reset) begin
      image_390 <= 4'h0;
    end else begin
      image_390 <= 4'h5;
    end
    if (reset) begin
      image_391 <= 4'h0;
    end else begin
      image_391 <= 4'h6;
    end
    if (reset) begin
      image_392 <= 4'h0;
    end else begin
      image_392 <= 4'h6;
    end
    if (reset) begin
      image_393 <= 4'h0;
    end else begin
      image_393 <= 4'h6;
    end
    if (reset) begin
      image_394 <= 4'h0;
    end else begin
      image_394 <= 4'h5;
    end
    if (reset) begin
      image_395 <= 4'h0;
    end else begin
      image_395 <= 4'h5;
    end
    if (reset) begin
      image_396 <= 4'h0;
    end else begin
      image_396 <= 4'h6;
    end
    if (reset) begin
      image_397 <= 4'h0;
    end else begin
      image_397 <= 4'h6;
    end
    if (reset) begin
      image_398 <= 4'h0;
    end else begin
      image_398 <= 4'h6;
    end
    if (reset) begin
      image_399 <= 4'h0;
    end else begin
      image_399 <= 4'h6;
    end
    if (reset) begin
      image_400 <= 4'h0;
    end else begin
      image_400 <= 4'h6;
    end
    if (reset) begin
      image_401 <= 4'h0;
    end else begin
      image_401 <= 4'h6;
    end
    if (reset) begin
      image_402 <= 4'h0;
    end else begin
      image_402 <= 4'h5;
    end
    if (reset) begin
      image_403 <= 4'h0;
    end else begin
      image_403 <= 4'h4;
    end
    if (reset) begin
      image_404 <= 4'h0;
    end else begin
      image_404 <= 4'h5;
    end
    if (reset) begin
      image_405 <= 4'h0;
    end else begin
      image_405 <= 4'h6;
    end
    if (reset) begin
      image_406 <= 4'h0;
    end else begin
      image_406 <= 4'h5;
    end
    if (reset) begin
      image_407 <= 4'h0;
    end else begin
      image_407 <= 4'h6;
    end
    if (reset) begin
      image_408 <= 4'h0;
    end else begin
      image_408 <= 4'h9;
    end
    if (reset) begin
      image_409 <= 4'h0;
    end else begin
      image_409 <= 4'hb;
    end
    if (reset) begin
      image_410 <= 4'h0;
    end else begin
      image_410 <= 4'hc;
    end
    if (reset) begin
      image_411 <= 4'h0;
    end else begin
      image_411 <= 4'hd;
    end
    if (reset) begin
      image_412 <= 4'h0;
    end else begin
      image_412 <= 4'he;
    end
    if (reset) begin
      image_413 <= 4'h0;
    end else begin
      image_413 <= 4'he;
    end
    if (reset) begin
      image_414 <= 4'h0;
    end else begin
      image_414 <= 4'hd;
    end
    if (reset) begin
      image_415 <= 4'h0;
    end else begin
      image_415 <= 4'hd;
    end
    if (reset) begin
      image_416 <= 4'h0;
    end else begin
      image_416 <= 4'hc;
    end
    if (reset) begin
      image_417 <= 4'h0;
    end else begin
      image_417 <= 4'hb;
    end
    if (reset) begin
      image_418 <= 4'h0;
    end else begin
      image_418 <= 4'h8;
    end
    if (reset) begin
      image_419 <= 4'h0;
    end else begin
      image_419 <= 4'h5;
    end
    if (reset) begin
      image_420 <= 4'h0;
    end else begin
      image_420 <= 4'h5;
    end
    if (reset) begin
      image_421 <= 4'h0;
    end else begin
      image_421 <= 4'h6;
    end
    if (reset) begin
      image_422 <= 4'h0;
    end else begin
      image_422 <= 4'h5;
    end
    if (reset) begin
      image_423 <= 4'h0;
    end else begin
      image_423 <= 4'h3;
    end
    if (reset) begin
      image_424 <= 4'h0;
    end else begin
      image_424 <= 4'h5;
    end
    if (reset) begin
      image_425 <= 4'h0;
    end else begin
      image_425 <= 4'h6;
    end
    if (reset) begin
      image_426 <= 4'h0;
    end else begin
      image_426 <= 4'h6;
    end
    if (reset) begin
      image_427 <= 4'h0;
    end else begin
      image_427 <= 4'h5;
    end
    if (reset) begin
      image_428 <= 4'h0;
    end else begin
      image_428 <= 4'h9;
    end
    if (reset) begin
      image_429 <= 4'h0;
    end else begin
      image_429 <= 4'hd;
    end
    if (reset) begin
      image_430 <= 4'h0;
    end else begin
      image_430 <= 4'he;
    end
    if (reset) begin
      image_431 <= 4'h0;
    end else begin
      image_431 <= 4'he;
    end
    if (reset) begin
      image_432 <= 4'h0;
    end else begin
      image_432 <= 4'he;
    end
    if (reset) begin
      image_433 <= 4'h0;
    end else begin
      image_433 <= 4'he;
    end
    if (reset) begin
      image_434 <= 4'h0;
    end else begin
      image_434 <= 4'he;
    end
    if (reset) begin
      image_435 <= 4'h0;
    end else begin
      image_435 <= 4'he;
    end
    if (reset) begin
      image_436 <= 4'h0;
    end else begin
      image_436 <= 4'he;
    end
    if (reset) begin
      image_437 <= 4'h0;
    end else begin
      image_437 <= 4'he;
    end
    if (reset) begin
      image_438 <= 4'h0;
    end else begin
      image_438 <= 4'he;
    end
    if (reset) begin
      image_439 <= 4'h0;
    end else begin
      image_439 <= 4'he;
    end
    if (reset) begin
      image_440 <= 4'h0;
    end else begin
      image_440 <= 4'he;
    end
    if (reset) begin
      image_441 <= 4'h0;
    end else begin
      image_441 <= 4'hc;
    end
    if (reset) begin
      image_442 <= 4'h0;
    end else begin
      image_442 <= 4'h9;
    end
    if (reset) begin
      image_443 <= 4'h0;
    end else begin
      image_443 <= 4'h4;
    end
    if (reset) begin
      image_444 <= 4'h0;
    end else begin
      image_444 <= 4'h3;
    end
    if (reset) begin
      image_451 <= 4'h0;
    end else begin
      image_451 <= 4'h2;
    end
    if (reset) begin
      image_452 <= 4'h0;
    end else begin
      image_452 <= 4'h5;
    end
    if (reset) begin
      image_453 <= 4'h0;
    end else begin
      image_453 <= 4'h5;
    end
    if (reset) begin
      image_454 <= 4'h0;
    end else begin
      image_454 <= 4'h6;
    end
    if (reset) begin
      image_455 <= 4'h0;
    end else begin
      image_455 <= 4'h6;
    end
    if (reset) begin
      image_456 <= 4'h0;
    end else begin
      image_456 <= 4'h6;
    end
    if (reset) begin
      image_457 <= 4'h0;
    end else begin
      image_457 <= 4'h6;
    end
    if (reset) begin
      image_458 <= 4'h0;
    end else begin
      image_458 <= 4'h6;
    end
    if (reset) begin
      image_459 <= 4'h0;
    end else begin
      image_459 <= 4'h6;
    end
    if (reset) begin
      image_460 <= 4'h0;
    end else begin
      image_460 <= 4'h6;
    end
    if (reset) begin
      image_461 <= 4'h0;
    end else begin
      image_461 <= 4'h6;
    end
    if (reset) begin
      image_462 <= 4'h0;
    end else begin
      image_462 <= 4'h6;
    end
    if (reset) begin
      image_463 <= 4'h0;
    end else begin
      image_463 <= 4'h6;
    end
    if (reset) begin
      image_464 <= 4'h0;
    end else begin
      image_464 <= 4'h5;
    end
    if (reset) begin
      image_465 <= 4'h0;
    end else begin
      image_465 <= 4'h4;
    end
    if (reset) begin
      image_466 <= 4'h0;
    end else begin
      image_466 <= 4'h5;
    end
    if (reset) begin
      image_467 <= 4'h0;
    end else begin
      image_467 <= 4'h6;
    end
    if (reset) begin
      image_468 <= 4'h0;
    end else begin
      image_468 <= 4'h5;
    end
    if (reset) begin
      image_469 <= 4'h0;
    end else begin
      image_469 <= 4'h9;
    end
    if (reset) begin
      image_470 <= 4'h0;
    end else begin
      image_470 <= 4'hd;
    end
    if (reset) begin
      image_471 <= 4'h0;
    end else begin
      image_471 <= 4'he;
    end
    if (reset) begin
      image_472 <= 4'h0;
    end else begin
      image_472 <= 4'he;
    end
    if (reset) begin
      image_473 <= 4'h0;
    end else begin
      image_473 <= 4'he;
    end
    if (reset) begin
      image_474 <= 4'h0;
    end else begin
      image_474 <= 4'he;
    end
    if (reset) begin
      image_475 <= 4'h0;
    end else begin
      image_475 <= 4'he;
    end
    if (reset) begin
      image_476 <= 4'h0;
    end else begin
      image_476 <= 4'he;
    end
    if (reset) begin
      image_477 <= 4'h0;
    end else begin
      image_477 <= 4'he;
    end
    if (reset) begin
      image_478 <= 4'h0;
    end else begin
      image_478 <= 4'hf;
    end
    if (reset) begin
      image_479 <= 4'h0;
    end else begin
      image_479 <= 4'hf;
    end
    if (reset) begin
      image_480 <= 4'h0;
    end else begin
      image_480 <= 4'he;
    end
    if (reset) begin
      image_481 <= 4'h0;
    end else begin
      image_481 <= 4'he;
    end
    if (reset) begin
      image_482 <= 4'h0;
    end else begin
      image_482 <= 4'he;
    end
    if (reset) begin
      image_483 <= 4'h0;
    end else begin
      image_483 <= 4'he;
    end
    if (reset) begin
      image_484 <= 4'h0;
    end else begin
      image_484 <= 4'hc;
    end
    if (reset) begin
      image_485 <= 4'h0;
    end else begin
      image_485 <= 4'h8;
    end
    if (reset) begin
      image_486 <= 4'h0;
    end else begin
      image_486 <= 4'h3;
    end
    if (reset) begin
      image_487 <= 4'h0;
    end else begin
      image_487 <= 4'h5;
    end
    if (reset) begin
      image_488 <= 4'h0;
    end else begin
      image_488 <= 4'h6;
    end
    if (reset) begin
      image_489 <= 4'h0;
    end else begin
      image_489 <= 4'h6;
    end
    if (reset) begin
      image_490 <= 4'h0;
    end else begin
      image_490 <= 4'h6;
    end
    if (reset) begin
      image_491 <= 4'h0;
    end else begin
      image_491 <= 4'hd;
    end
    if (reset) begin
      image_492 <= 4'h0;
    end else begin
      image_492 <= 4'he;
    end
    if (reset) begin
      image_493 <= 4'h0;
    end else begin
      image_493 <= 4'he;
    end
    if (reset) begin
      image_494 <= 4'h0;
    end else begin
      image_494 <= 4'he;
    end
    if (reset) begin
      image_495 <= 4'h0;
    end else begin
      image_495 <= 4'hf;
    end
    if (reset) begin
      image_496 <= 4'h0;
    end else begin
      image_496 <= 4'he;
    end
    if (reset) begin
      image_497 <= 4'h0;
    end else begin
      image_497 <= 4'hf;
    end
    if (reset) begin
      image_498 <= 4'h0;
    end else begin
      image_498 <= 4'hf;
    end
    if (reset) begin
      image_499 <= 4'h0;
    end else begin
      image_499 <= 4'he;
    end
    if (reset) begin
      image_500 <= 4'h0;
    end else begin
      image_500 <= 4'he;
    end
    if (reset) begin
      image_501 <= 4'h0;
    end else begin
      image_501 <= 4'he;
    end
    if (reset) begin
      image_502 <= 4'h0;
    end else begin
      image_502 <= 4'he;
    end
    if (reset) begin
      image_503 <= 4'h0;
    end else begin
      image_503 <= 4'hc;
    end
    if (reset) begin
      image_504 <= 4'h0;
    end else begin
      image_504 <= 4'ha;
    end
    if (reset) begin
      image_505 <= 4'h0;
    end else begin
      image_505 <= 4'hb;
    end
    if (reset) begin
      image_506 <= 4'h0;
    end else begin
      image_506 <= 4'hd;
    end
    if (reset) begin
      image_507 <= 4'h0;
    end else begin
      image_507 <= 4'he;
    end
    if (reset) begin
      image_508 <= 4'h0;
    end else begin
      image_508 <= 4'h9;
    end
    if (reset) begin
      image_509 <= 4'h0;
    end else begin
      image_509 <= 4'h2;
    end
    if (reset) begin
      image_515 <= 4'h0;
    end else begin
      image_515 <= 4'h4;
    end
    if (reset) begin
      image_516 <= 4'h0;
    end else begin
      image_516 <= 4'h5;
    end
    if (reset) begin
      image_517 <= 4'h0;
    end else begin
      image_517 <= 4'h5;
    end
    if (reset) begin
      image_518 <= 4'h0;
    end else begin
      image_518 <= 4'h6;
    end
    if (reset) begin
      image_519 <= 4'h0;
    end else begin
      image_519 <= 4'h6;
    end
    if (reset) begin
      image_520 <= 4'h0;
    end else begin
      image_520 <= 4'h6;
    end
    if (reset) begin
      image_521 <= 4'h0;
    end else begin
      image_521 <= 4'h6;
    end
    if (reset) begin
      image_522 <= 4'h0;
    end else begin
      image_522 <= 4'h6;
    end
    if (reset) begin
      image_523 <= 4'h0;
    end else begin
      image_523 <= 4'h6;
    end
    if (reset) begin
      image_524 <= 4'h0;
    end else begin
      image_524 <= 4'h6;
    end
    if (reset) begin
      image_525 <= 4'h0;
    end else begin
      image_525 <= 4'h6;
    end
    if (reset) begin
      image_526 <= 4'h0;
    end else begin
      image_526 <= 4'h6;
    end
    if (reset) begin
      image_527 <= 4'h0;
    end else begin
      image_527 <= 4'h4;
    end
    if (reset) begin
      image_528 <= 4'h0;
    end else begin
      image_528 <= 4'h5;
    end
    if (reset) begin
      image_529 <= 4'h0;
    end else begin
      image_529 <= 4'h6;
    end
    if (reset) begin
      image_530 <= 4'h0;
    end else begin
      image_530 <= 4'h6;
    end
    if (reset) begin
      image_531 <= 4'h0;
    end else begin
      image_531 <= 4'h6;
    end
    if (reset) begin
      image_532 <= 4'h0;
    end else begin
      image_532 <= 4'hd;
    end
    if (reset) begin
      image_533 <= 4'h0;
    end else begin
      image_533 <= 4'he;
    end
    if (reset) begin
      image_534 <= 4'h0;
    end else begin
      image_534 <= 4'he;
    end
    if (reset) begin
      image_535 <= 4'h0;
    end else begin
      image_535 <= 4'he;
    end
    if (reset) begin
      image_536 <= 4'h0;
    end else begin
      image_536 <= 4'hf;
    end
    if (reset) begin
      image_537 <= 4'h0;
    end else begin
      image_537 <= 4'he;
    end
    if (reset) begin
      image_538 <= 4'h0;
    end else begin
      image_538 <= 4'hf;
    end
    if (reset) begin
      image_539 <= 4'h0;
    end else begin
      image_539 <= 4'hf;
    end
    if (reset) begin
      image_540 <= 4'h0;
    end else begin
      image_540 <= 4'he;
    end
    if (reset) begin
      image_541 <= 4'h0;
    end else begin
      image_541 <= 4'hf;
    end
    if (reset) begin
      image_542 <= 4'h0;
    end else begin
      image_542 <= 4'hf;
    end
    if (reset) begin
      image_543 <= 4'h0;
    end else begin
      image_543 <= 4'he;
    end
    if (reset) begin
      image_544 <= 4'h0;
    end else begin
      image_544 <= 4'hd;
    end
    if (reset) begin
      image_545 <= 4'h0;
    end else begin
      image_545 <= 4'ha;
    end
    if (reset) begin
      image_546 <= 4'h0;
    end else begin
      image_546 <= 4'h7;
    end
    if (reset) begin
      image_547 <= 4'h0;
    end else begin
      image_547 <= 4'h7;
    end
    if (reset) begin
      image_548 <= 4'h0;
    end else begin
      image_548 <= 4'h9;
    end
    if (reset) begin
      image_549 <= 4'h0;
    end else begin
      image_549 <= 4'hc;
    end
    if (reset) begin
      image_550 <= 4'h0;
    end else begin
      image_550 <= 4'hd;
    end
    if (reset) begin
      image_551 <= 4'h0;
    end else begin
      image_551 <= 4'h8;
    end
    if (reset) begin
      image_552 <= 4'h0;
    end else begin
      image_552 <= 4'h5;
    end
    if (reset) begin
      image_553 <= 4'h0;
    end else begin
      image_553 <= 4'h6;
    end
    if (reset) begin
      image_554 <= 4'h0;
    end else begin
      image_554 <= 4'he;
    end
    if (reset) begin
      image_555 <= 4'h0;
    end else begin
      image_555 <= 4'he;
    end
    if (reset) begin
      image_556 <= 4'h0;
    end else begin
      image_556 <= 4'he;
    end
    if (reset) begin
      image_557 <= 4'h0;
    end else begin
      image_557 <= 4'he;
    end
    if (reset) begin
      image_558 <= 4'h0;
    end else begin
      image_558 <= 4'hf;
    end
    if (reset) begin
      image_559 <= 4'h0;
    end else begin
      image_559 <= 4'hf;
    end
    if (reset) begin
      image_560 <= 4'h0;
    end else begin
      image_560 <= 4'hf;
    end
    if (reset) begin
      image_561 <= 4'h0;
    end else begin
      image_561 <= 4'hf;
    end
    if (reset) begin
      image_562 <= 4'h0;
    end else begin
      image_562 <= 4'hf;
    end
    if (reset) begin
      image_563 <= 4'h0;
    end else begin
      image_563 <= 4'hf;
    end
    if (reset) begin
      image_564 <= 4'h0;
    end else begin
      image_564 <= 4'he;
    end
    if (reset) begin
      image_565 <= 4'h0;
    end else begin
      image_565 <= 4'hb;
    end
    if (reset) begin
      image_566 <= 4'h0;
    end else begin
      image_566 <= 4'h3;
    end
    if (reset) begin
      image_571 <= 4'h0;
    end else begin
      image_571 <= 4'h7;
    end
    if (reset) begin
      image_572 <= 4'h0;
    end else begin
      image_572 <= 4'he;
    end
    if (reset) begin
      image_573 <= 4'h0;
    end else begin
      image_573 <= 4'hc;
    end
    if (reset) begin
      image_574 <= 4'h0;
    end else begin
      image_574 <= 4'h6;
    end
    if (reset) begin
      image_578 <= 4'h0;
    end else begin
      image_578 <= 4'h3;
    end
    if (reset) begin
      image_579 <= 4'h0;
    end else begin
      image_579 <= 4'h5;
    end
    if (reset) begin
      image_580 <= 4'h0;
    end else begin
      image_580 <= 4'h5;
    end
    if (reset) begin
      image_581 <= 4'h0;
    end else begin
      image_581 <= 4'h5;
    end
    if (reset) begin
      image_582 <= 4'h0;
    end else begin
      image_582 <= 4'h6;
    end
    if (reset) begin
      image_583 <= 4'h0;
    end else begin
      image_583 <= 4'h6;
    end
    if (reset) begin
      image_584 <= 4'h0;
    end else begin
      image_584 <= 4'h6;
    end
    if (reset) begin
      image_585 <= 4'h0;
    end else begin
      image_585 <= 4'h6;
    end
    if (reset) begin
      image_586 <= 4'h0;
    end else begin
      image_586 <= 4'h6;
    end
    if (reset) begin
      image_587 <= 4'h0;
    end else begin
      image_587 <= 4'h6;
    end
    if (reset) begin
      image_588 <= 4'h0;
    end else begin
      image_588 <= 4'h6;
    end
    if (reset) begin
      image_589 <= 4'h0;
    end else begin
      image_589 <= 4'h6;
    end
    if (reset) begin
      image_590 <= 4'h0;
    end else begin
      image_590 <= 4'h6;
    end
    if (reset) begin
      image_591 <= 4'h0;
    end else begin
      image_591 <= 4'h6;
    end
    if (reset) begin
      image_592 <= 4'h0;
    end else begin
      image_592 <= 4'h6;
    end
    if (reset) begin
      image_593 <= 4'h0;
    end else begin
      image_593 <= 4'h5;
    end
    if (reset) begin
      image_594 <= 4'h0;
    end else begin
      image_594 <= 4'h8;
    end
    if (reset) begin
      image_595 <= 4'h0;
    end else begin
      image_595 <= 4'he;
    end
    if (reset) begin
      image_596 <= 4'h0;
    end else begin
      image_596 <= 4'he;
    end
    if (reset) begin
      image_597 <= 4'h0;
    end else begin
      image_597 <= 4'he;
    end
    if (reset) begin
      image_598 <= 4'h0;
    end else begin
      image_598 <= 4'he;
    end
    if (reset) begin
      image_599 <= 4'h0;
    end else begin
      image_599 <= 4'he;
    end
    if (reset) begin
      image_600 <= 4'h0;
    end else begin
      image_600 <= 4'hf;
    end
    if (reset) begin
      image_601 <= 4'h0;
    end else begin
      image_601 <= 4'hf;
    end
    if (reset) begin
      image_602 <= 4'h0;
    end else begin
      image_602 <= 4'hf;
    end
    if (reset) begin
      image_603 <= 4'h0;
    end else begin
      image_603 <= 4'hf;
    end
    if (reset) begin
      image_604 <= 4'h0;
    end else begin
      image_604 <= 4'hf;
    end
    if (reset) begin
      image_605 <= 4'h0;
    end else begin
      image_605 <= 4'hf;
    end
    if (reset) begin
      image_606 <= 4'h0;
    end else begin
      image_606 <= 4'he;
    end
    if (reset) begin
      image_607 <= 4'h0;
    end else begin
      image_607 <= 4'h9;
    end
    if (reset) begin
      image_614 <= 4'h0;
    end else begin
      image_614 <= 4'h5;
    end
    if (reset) begin
      image_615 <= 4'h0;
    end else begin
      image_615 <= 4'hd;
    end
    if (reset) begin
      image_616 <= 4'h0;
    end else begin
      image_616 <= 4'ha;
    end
    if (reset) begin
      image_617 <= 4'h0;
    end else begin
      image_617 <= 4'h9;
    end
    if (reset) begin
      image_618 <= 4'h0;
    end else begin
      image_618 <= 4'he;
    end
    if (reset) begin
      image_619 <= 4'h0;
    end else begin
      image_619 <= 4'he;
    end
    if (reset) begin
      image_620 <= 4'h0;
    end else begin
      image_620 <= 4'he;
    end
    if (reset) begin
      image_621 <= 4'h0;
    end else begin
      image_621 <= 4'he;
    end
    if (reset) begin
      image_622 <= 4'h0;
    end else begin
      image_622 <= 4'hf;
    end
    if (reset) begin
      image_623 <= 4'h0;
    end else begin
      image_623 <= 4'hf;
    end
    if (reset) begin
      image_624 <= 4'h0;
    end else begin
      image_624 <= 4'hf;
    end
    if (reset) begin
      image_625 <= 4'h0;
    end else begin
      image_625 <= 4'hf;
    end
    if (reset) begin
      image_626 <= 4'h0;
    end else begin
      image_626 <= 4'hf;
    end
    if (reset) begin
      image_627 <= 4'h0;
    end else begin
      image_627 <= 4'hf;
    end
    if (reset) begin
      image_628 <= 4'h0;
    end else begin
      image_628 <= 4'hb;
    end
    if (reset) begin
      image_636 <= 4'h0;
    end else begin
      image_636 <= 4'h6;
    end
    if (reset) begin
      image_637 <= 4'h0;
    end else begin
      image_637 <= 4'he;
    end
    if (reset) begin
      image_638 <= 4'h0;
    end else begin
      image_638 <= 4'hb;
    end
    if (reset) begin
      image_639 <= 4'h0;
    end else begin
      image_639 <= 4'h3;
    end
    if (reset) begin
      image_642 <= 4'h0;
    end else begin
      image_642 <= 4'h4;
    end
    if (reset) begin
      image_643 <= 4'h0;
    end else begin
      image_643 <= 4'h5;
    end
    if (reset) begin
      image_644 <= 4'h0;
    end else begin
      image_644 <= 4'h5;
    end
    if (reset) begin
      image_645 <= 4'h0;
    end else begin
      image_645 <= 4'h5;
    end
    if (reset) begin
      image_646 <= 4'h0;
    end else begin
      image_646 <= 4'h6;
    end
    if (reset) begin
      image_647 <= 4'h0;
    end else begin
      image_647 <= 4'h6;
    end
    if (reset) begin
      image_648 <= 4'h0;
    end else begin
      image_648 <= 4'h6;
    end
    if (reset) begin
      image_649 <= 4'h0;
    end else begin
      image_649 <= 4'h6;
    end
    if (reset) begin
      image_650 <= 4'h0;
    end else begin
      image_650 <= 4'h6;
    end
    if (reset) begin
      image_651 <= 4'h0;
    end else begin
      image_651 <= 4'h6;
    end
    if (reset) begin
      image_652 <= 4'h0;
    end else begin
      image_652 <= 4'h6;
    end
    if (reset) begin
      image_653 <= 4'h0;
    end else begin
      image_653 <= 4'h6;
    end
    if (reset) begin
      image_654 <= 4'h0;
    end else begin
      image_654 <= 4'h5;
    end
    if (reset) begin
      image_655 <= 4'h0;
    end else begin
      image_655 <= 4'h4;
    end
    if (reset) begin
      image_656 <= 4'h0;
    end else begin
      image_656 <= 4'h7;
    end
    if (reset) begin
      image_657 <= 4'h0;
    end else begin
      image_657 <= 4'hb;
    end
    if (reset) begin
      image_658 <= 4'h0;
    end else begin
      image_658 <= 4'he;
    end
    if (reset) begin
      image_659 <= 4'h0;
    end else begin
      image_659 <= 4'he;
    end
    if (reset) begin
      image_660 <= 4'h0;
    end else begin
      image_660 <= 4'hf;
    end
    if (reset) begin
      image_661 <= 4'h0;
    end else begin
      image_661 <= 4'hf;
    end
    if (reset) begin
      image_662 <= 4'h0;
    end else begin
      image_662 <= 4'hf;
    end
    if (reset) begin
      image_663 <= 4'h0;
    end else begin
      image_663 <= 4'hf;
    end
    if (reset) begin
      image_664 <= 4'h0;
    end else begin
      image_664 <= 4'hf;
    end
    if (reset) begin
      image_665 <= 4'h0;
    end else begin
      image_665 <= 4'hf;
    end
    if (reset) begin
      image_666 <= 4'h0;
    end else begin
      image_666 <= 4'hf;
    end
    if (reset) begin
      image_667 <= 4'h0;
    end else begin
      image_667 <= 4'hf;
    end
    if (reset) begin
      image_668 <= 4'h0;
    end else begin
      image_668 <= 4'hf;
    end
    if (reset) begin
      image_669 <= 4'h0;
    end else begin
      image_669 <= 4'he;
    end
    if (reset) begin
      image_670 <= 4'h0;
    end else begin
      image_670 <= 4'h9;
    end
    if (reset) begin
      image_679 <= 4'h0;
    end else begin
      image_679 <= 4'h5;
    end
    if (reset) begin
      image_680 <= 4'h0;
    end else begin
      image_680 <= 4'he;
    end
    if (reset) begin
      image_681 <= 4'h0;
    end else begin
      image_681 <= 4'h9;
    end
    if (reset) begin
      image_682 <= 4'h0;
    end else begin
      image_682 <= 4'hc;
    end
    if (reset) begin
      image_683 <= 4'h0;
    end else begin
      image_683 <= 4'he;
    end
    if (reset) begin
      image_684 <= 4'h0;
    end else begin
      image_684 <= 4'hf;
    end
    if (reset) begin
      image_685 <= 4'h0;
    end else begin
      image_685 <= 4'hf;
    end
    if (reset) begin
      image_686 <= 4'h0;
    end else begin
      image_686 <= 4'hf;
    end
    if (reset) begin
      image_687 <= 4'h0;
    end else begin
      image_687 <= 4'hf;
    end
    if (reset) begin
      image_688 <= 4'h0;
    end else begin
      image_688 <= 4'hf;
    end
    if (reset) begin
      image_689 <= 4'h0;
    end else begin
      image_689 <= 4'hf;
    end
    if (reset) begin
      image_690 <= 4'h0;
    end else begin
      image_690 <= 4'hf;
    end
    if (reset) begin
      image_691 <= 4'h0;
    end else begin
      image_691 <= 4'he;
    end
    if (reset) begin
      image_692 <= 4'h0;
    end else begin
      image_692 <= 4'h6;
    end
    if (reset) begin
      image_693 <= 4'h0;
    end else begin
      image_693 <= 4'h5;
    end
    if (reset) begin
      image_694 <= 4'h0;
    end else begin
      image_694 <= 4'hd;
    end
    if (reset) begin
      image_695 <= 4'h0;
    end else begin
      image_695 <= 4'h5;
    end
    if (reset) begin
      image_696 <= 4'h0;
    end else begin
      image_696 <= 4'h7;
    end
    if (reset) begin
      image_697 <= 4'h0;
    end else begin
      image_697 <= 4'hc;
    end
    if (reset) begin
      image_698 <= 4'h0;
    end else begin
      image_698 <= 4'h9;
    end
    if (reset) begin
      image_701 <= 4'h0;
    end else begin
      image_701 <= 4'hd;
    end
    if (reset) begin
      image_702 <= 4'h0;
    end else begin
      image_702 <= 4'hd;
    end
    if (reset) begin
      image_703 <= 4'h0;
    end else begin
      image_703 <= 4'h8;
    end
    if (reset) begin
      image_705 <= 4'h0;
    end else begin
      image_705 <= 4'h2;
    end
    if (reset) begin
      image_706 <= 4'h0;
    end else begin
      image_706 <= 4'h5;
    end
    if (reset) begin
      image_707 <= 4'h0;
    end else begin
      image_707 <= 4'h5;
    end
    if (reset) begin
      image_708 <= 4'h0;
    end else begin
      image_708 <= 4'h5;
    end
    if (reset) begin
      image_709 <= 4'h0;
    end else begin
      image_709 <= 4'h6;
    end
    if (reset) begin
      image_710 <= 4'h0;
    end else begin
      image_710 <= 4'h6;
    end
    if (reset) begin
      image_711 <= 4'h0;
    end else begin
      image_711 <= 4'h6;
    end
    if (reset) begin
      image_712 <= 4'h0;
    end else begin
      image_712 <= 4'h6;
    end
    if (reset) begin
      image_713 <= 4'h0;
    end else begin
      image_713 <= 4'h6;
    end
    if (reset) begin
      image_714 <= 4'h0;
    end else begin
      image_714 <= 4'h6;
    end
    if (reset) begin
      image_715 <= 4'h0;
    end else begin
      image_715 <= 4'h6;
    end
    if (reset) begin
      image_716 <= 4'h0;
    end else begin
      image_716 <= 4'h6;
    end
    if (reset) begin
      image_717 <= 4'h0;
    end else begin
      image_717 <= 4'h7;
    end
    if (reset) begin
      image_718 <= 4'h0;
    end else begin
      image_718 <= 4'hd;
    end
    if (reset) begin
      image_719 <= 4'h0;
    end else begin
      image_719 <= 4'he;
    end
    if (reset) begin
      image_720 <= 4'h0;
    end else begin
      image_720 <= 4'he;
    end
    if (reset) begin
      image_721 <= 4'h0;
    end else begin
      image_721 <= 4'he;
    end
    if (reset) begin
      image_722 <= 4'h0;
    end else begin
      image_722 <= 4'hf;
    end
    if (reset) begin
      image_723 <= 4'h0;
    end else begin
      image_723 <= 4'hf;
    end
    if (reset) begin
      image_724 <= 4'h0;
    end else begin
      image_724 <= 4'hf;
    end
    if (reset) begin
      image_725 <= 4'h0;
    end else begin
      image_725 <= 4'hf;
    end
    if (reset) begin
      image_726 <= 4'h0;
    end else begin
      image_726 <= 4'hf;
    end
    if (reset) begin
      image_727 <= 4'h0;
    end else begin
      image_727 <= 4'hf;
    end
    if (reset) begin
      image_728 <= 4'h0;
    end else begin
      image_728 <= 4'hf;
    end
    if (reset) begin
      image_729 <= 4'h0;
    end else begin
      image_729 <= 4'hf;
    end
    if (reset) begin
      image_730 <= 4'h0;
    end else begin
      image_730 <= 4'hf;
    end
    if (reset) begin
      image_731 <= 4'h0;
    end else begin
      image_731 <= 4'hf;
    end
    if (reset) begin
      image_732 <= 4'h0;
    end else begin
      image_732 <= 4'hf;
    end
    if (reset) begin
      image_733 <= 4'h0;
    end else begin
      image_733 <= 4'hd;
    end
    if (reset) begin
      image_734 <= 4'h0;
    end else begin
      image_734 <= 4'h1;
    end
    if (reset) begin
      image_736 <= 4'h0;
    end else begin
      image_736 <= 4'hc;
    end
    if (reset) begin
      image_737 <= 4'h0;
    end else begin
      image_737 <= 4'hc;
    end
    if (reset) begin
      image_739 <= 4'h0;
    end else begin
      image_739 <= 4'ha;
    end
    if (reset) begin
      image_740 <= 4'h0;
    end else begin
      image_740 <= 4'hd;
    end
    if (reset) begin
      image_741 <= 4'h0;
    end else begin
      image_741 <= 4'h9;
    end
    if (reset) begin
      image_744 <= 4'h0;
    end else begin
      image_744 <= 4'hb;
    end
    if (reset) begin
      image_745 <= 4'h0;
    end else begin
      image_745 <= 4'he;
    end
    if (reset) begin
      image_746 <= 4'h0;
    end else begin
      image_746 <= 4'h7;
    end
    if (reset) begin
      image_747 <= 4'h0;
    end else begin
      image_747 <= 4'he;
    end
    if (reset) begin
      image_748 <= 4'h0;
    end else begin
      image_748 <= 4'hf;
    end
    if (reset) begin
      image_749 <= 4'h0;
    end else begin
      image_749 <= 4'hf;
    end
    if (reset) begin
      image_750 <= 4'h0;
    end else begin
      image_750 <= 4'hf;
    end
    if (reset) begin
      image_751 <= 4'h0;
    end else begin
      image_751 <= 4'hf;
    end
    if (reset) begin
      image_752 <= 4'h0;
    end else begin
      image_752 <= 4'hf;
    end
    if (reset) begin
      image_753 <= 4'h0;
    end else begin
      image_753 <= 4'hf;
    end
    if (reset) begin
      image_754 <= 4'h0;
    end else begin
      image_754 <= 4'hf;
    end
    if (reset) begin
      image_755 <= 4'h0;
    end else begin
      image_755 <= 4'he;
    end
    if (reset) begin
      image_756 <= 4'h0;
    end else begin
      image_756 <= 4'h5;
    end
    if (reset) begin
      image_758 <= 4'h0;
    end else begin
      image_758 <= 4'h4;
    end
    if (reset) begin
      image_760 <= 4'h0;
    end else begin
      image_760 <= 4'hc;
    end
    if (reset) begin
      image_761 <= 4'h0;
    end else begin
      image_761 <= 4'he;
    end
    if (reset) begin
      image_762 <= 4'h0;
    end else begin
      image_762 <= 4'hd;
    end
    if (reset) begin
      image_763 <= 4'h0;
    end else begin
      image_763 <= 4'h1;
    end
    if (reset) begin
      image_765 <= 4'h0;
    end else begin
      image_765 <= 4'hc;
    end
    if (reset) begin
      image_766 <= 4'h0;
    end else begin
      image_766 <= 4'he;
    end
    if (reset) begin
      image_767 <= 4'h0;
    end else begin
      image_767 <= 4'h9;
    end
    if (reset) begin
      image_768 <= 4'h0;
    end else begin
      image_768 <= 4'h1;
    end
    if (reset) begin
      image_769 <= 4'h0;
    end else begin
      image_769 <= 4'h3;
    end
    if (reset) begin
      image_770 <= 4'h0;
    end else begin
      image_770 <= 4'h5;
    end
    if (reset) begin
      image_771 <= 4'h0;
    end else begin
      image_771 <= 4'h5;
    end
    if (reset) begin
      image_772 <= 4'h0;
    end else begin
      image_772 <= 4'h5;
    end
    if (reset) begin
      image_773 <= 4'h0;
    end else begin
      image_773 <= 4'h6;
    end
    if (reset) begin
      image_774 <= 4'h0;
    end else begin
      image_774 <= 4'h6;
    end
    if (reset) begin
      image_775 <= 4'h0;
    end else begin
      image_775 <= 4'h6;
    end
    if (reset) begin
      image_776 <= 4'h0;
    end else begin
      image_776 <= 4'h6;
    end
    if (reset) begin
      image_777 <= 4'h0;
    end else begin
      image_777 <= 4'h6;
    end
    if (reset) begin
      image_778 <= 4'h0;
    end else begin
      image_778 <= 4'h6;
    end
    if (reset) begin
      image_779 <= 4'h0;
    end else begin
      image_779 <= 4'h6;
    end
    if (reset) begin
      image_780 <= 4'h0;
    end else begin
      image_780 <= 4'h4;
    end
    if (reset) begin
      image_781 <= 4'h0;
    end else begin
      image_781 <= 4'hb;
    end
    if (reset) begin
      image_782 <= 4'h0;
    end else begin
      image_782 <= 4'he;
    end
    if (reset) begin
      image_783 <= 4'h0;
    end else begin
      image_783 <= 4'he;
    end
    if (reset) begin
      image_784 <= 4'h0;
    end else begin
      image_784 <= 4'he;
    end
    if (reset) begin
      image_785 <= 4'h0;
    end else begin
      image_785 <= 4'he;
    end
    if (reset) begin
      image_786 <= 4'h0;
    end else begin
      image_786 <= 4'hf;
    end
    if (reset) begin
      image_787 <= 4'h0;
    end else begin
      image_787 <= 4'hf;
    end
    if (reset) begin
      image_788 <= 4'h0;
    end else begin
      image_788 <= 4'hf;
    end
    if (reset) begin
      image_789 <= 4'h0;
    end else begin
      image_789 <= 4'hf;
    end
    if (reset) begin
      image_790 <= 4'h0;
    end else begin
      image_790 <= 4'hf;
    end
    if (reset) begin
      image_791 <= 4'h0;
    end else begin
      image_791 <= 4'hf;
    end
    if (reset) begin
      image_792 <= 4'h0;
    end else begin
      image_792 <= 4'hf;
    end
    if (reset) begin
      image_793 <= 4'h0;
    end else begin
      image_793 <= 4'hf;
    end
    if (reset) begin
      image_794 <= 4'h0;
    end else begin
      image_794 <= 4'hf;
    end
    if (reset) begin
      image_795 <= 4'h0;
    end else begin
      image_795 <= 4'hf;
    end
    if (reset) begin
      image_796 <= 4'h0;
    end else begin
      image_796 <= 4'hf;
    end
    if (reset) begin
      image_797 <= 4'h0;
    end else begin
      image_797 <= 4'hd;
    end
    if (reset) begin
      image_800 <= 4'h0;
    end else begin
      image_800 <= 4'h6;
    end
    if (reset) begin
      image_801 <= 4'h0;
    end else begin
      image_801 <= 4'h6;
    end
    if (reset) begin
      image_802 <= 4'h0;
    end else begin
      image_802 <= 4'h4;
    end
    if (reset) begin
      image_803 <= 4'h0;
    end else begin
      image_803 <= 4'he;
    end
    if (reset) begin
      image_804 <= 4'h0;
    end else begin
      image_804 <= 4'he;
    end
    if (reset) begin
      image_805 <= 4'h0;
    end else begin
      image_805 <= 4'he;
    end
    if (reset) begin
      image_806 <= 4'h0;
    end else begin
      image_806 <= 4'h2;
    end
    if (reset) begin
      image_808 <= 4'h0;
    end else begin
      image_808 <= 4'hb;
    end
    if (reset) begin
      image_809 <= 4'h0;
    end else begin
      image_809 <= 4'he;
    end
    if (reset) begin
      image_810 <= 4'h0;
    end else begin
      image_810 <= 4'h7;
    end
    if (reset) begin
      image_811 <= 4'h0;
    end else begin
      image_811 <= 4'he;
    end
    if (reset) begin
      image_812 <= 4'h0;
    end else begin
      image_812 <= 4'hf;
    end
    if (reset) begin
      image_813 <= 4'h0;
    end else begin
      image_813 <= 4'hf;
    end
    if (reset) begin
      image_814 <= 4'h0;
    end else begin
      image_814 <= 4'hf;
    end
    if (reset) begin
      image_815 <= 4'h0;
    end else begin
      image_815 <= 4'hf;
    end
    if (reset) begin
      image_816 <= 4'h0;
    end else begin
      image_816 <= 4'hf;
    end
    if (reset) begin
      image_817 <= 4'h0;
    end else begin
      image_817 <= 4'hf;
    end
    if (reset) begin
      image_818 <= 4'h0;
    end else begin
      image_818 <= 4'hf;
    end
    if (reset) begin
      image_819 <= 4'h0;
    end else begin
      image_819 <= 4'he;
    end
    if (reset) begin
      image_820 <= 4'h0;
    end else begin
      image_820 <= 4'ha;
    end
    if (reset) begin
      image_822 <= 4'h0;
    end else begin
      image_822 <= 4'h5;
    end
    if (reset) begin
      image_823 <= 4'h0;
    end else begin
      image_823 <= 4'h7;
    end
    if (reset) begin
      image_824 <= 4'h0;
    end else begin
      image_824 <= 4'h3;
    end
    if (reset) begin
      image_825 <= 4'h0;
    end else begin
      image_825 <= 4'h8;
    end
    if (reset) begin
      image_826 <= 4'h0;
    end else begin
      image_826 <= 4'h5;
    end
    if (reset) begin
      image_828 <= 4'h0;
    end else begin
      image_828 <= 4'h5;
    end
    if (reset) begin
      image_829 <= 4'h0;
    end else begin
      image_829 <= 4'he;
    end
    if (reset) begin
      image_830 <= 4'h0;
    end else begin
      image_830 <= 4'hd;
    end
    if (reset) begin
      image_831 <= 4'h0;
    end else begin
      image_831 <= 4'h8;
    end
    if (reset) begin
      image_833 <= 4'h0;
    end else begin
      image_833 <= 4'h4;
    end
    if (reset) begin
      image_834 <= 4'h0;
    end else begin
      image_834 <= 4'h5;
    end
    if (reset) begin
      image_835 <= 4'h0;
    end else begin
      image_835 <= 4'h5;
    end
    if (reset) begin
      image_836 <= 4'h0;
    end else begin
      image_836 <= 4'h5;
    end
    if (reset) begin
      image_837 <= 4'h0;
    end else begin
      image_837 <= 4'h6;
    end
    if (reset) begin
      image_838 <= 4'h0;
    end else begin
      image_838 <= 4'h6;
    end
    if (reset) begin
      image_839 <= 4'h0;
    end else begin
      image_839 <= 4'h6;
    end
    if (reset) begin
      image_840 <= 4'h0;
    end else begin
      image_840 <= 4'h6;
    end
    if (reset) begin
      image_841 <= 4'h0;
    end else begin
      image_841 <= 4'h6;
    end
    if (reset) begin
      image_842 <= 4'h0;
    end else begin
      image_842 <= 4'h6;
    end
    if (reset) begin
      image_843 <= 4'h0;
    end else begin
      image_843 <= 4'h6;
    end
    if (reset) begin
      image_844 <= 4'h0;
    end else begin
      image_844 <= 4'h6;
    end
    if (reset) begin
      image_845 <= 4'h0;
    end else begin
      image_845 <= 4'h5;
    end
    if (reset) begin
      image_846 <= 4'h0;
    end else begin
      image_846 <= 4'h6;
    end
    if (reset) begin
      image_847 <= 4'h0;
    end else begin
      image_847 <= 4'h8;
    end
    if (reset) begin
      image_848 <= 4'h0;
    end else begin
      image_848 <= 4'hb;
    end
    if (reset) begin
      image_849 <= 4'h0;
    end else begin
      image_849 <= 4'he;
    end
    if (reset) begin
      image_850 <= 4'h0;
    end else begin
      image_850 <= 4'he;
    end
    if (reset) begin
      image_851 <= 4'h0;
    end else begin
      image_851 <= 4'he;
    end
    if (reset) begin
      image_852 <= 4'h0;
    end else begin
      image_852 <= 4'hf;
    end
    if (reset) begin
      image_853 <= 4'h0;
    end else begin
      image_853 <= 4'hf;
    end
    if (reset) begin
      image_854 <= 4'h0;
    end else begin
      image_854 <= 4'hf;
    end
    if (reset) begin
      image_855 <= 4'h0;
    end else begin
      image_855 <= 4'hf;
    end
    if (reset) begin
      image_856 <= 4'h0;
    end else begin
      image_856 <= 4'hf;
    end
    if (reset) begin
      image_857 <= 4'h0;
    end else begin
      image_857 <= 4'hf;
    end
    if (reset) begin
      image_858 <= 4'h0;
    end else begin
      image_858 <= 4'hf;
    end
    if (reset) begin
      image_859 <= 4'h0;
    end else begin
      image_859 <= 4'hf;
    end
    if (reset) begin
      image_860 <= 4'h0;
    end else begin
      image_860 <= 4'hf;
    end
    if (reset) begin
      image_861 <= 4'h0;
    end else begin
      image_861 <= 4'he;
    end
    if (reset) begin
      image_862 <= 4'h0;
    end else begin
      image_862 <= 4'h3;
    end
    if (reset) begin
      image_865 <= 4'h0;
    end else begin
      image_865 <= 4'h6;
    end
    if (reset) begin
      image_866 <= 4'h0;
    end else begin
      image_866 <= 4'h1;
    end
    if (reset) begin
      image_867 <= 4'h0;
    end else begin
      image_867 <= 4'h9;
    end
    if (reset) begin
      image_868 <= 4'h0;
    end else begin
      image_868 <= 4'hb;
    end
    if (reset) begin
      image_869 <= 4'h0;
    end else begin
      image_869 <= 4'h8;
    end
    if (reset) begin
      image_872 <= 4'h0;
    end else begin
      image_872 <= 4'hc;
    end
    if (reset) begin
      image_873 <= 4'h0;
    end else begin
      image_873 <= 4'he;
    end
    if (reset) begin
      image_874 <= 4'h0;
    end else begin
      image_874 <= 4'h5;
    end
    if (reset) begin
      image_875 <= 4'h0;
    end else begin
      image_875 <= 4'hd;
    end
    if (reset) begin
      image_876 <= 4'h0;
    end else begin
      image_876 <= 4'he;
    end
    if (reset) begin
      image_877 <= 4'h0;
    end else begin
      image_877 <= 4'he;
    end
    if (reset) begin
      image_878 <= 4'h0;
    end else begin
      image_878 <= 4'hf;
    end
    if (reset) begin
      image_879 <= 4'h0;
    end else begin
      image_879 <= 4'hf;
    end
    if (reset) begin
      image_880 <= 4'h0;
    end else begin
      image_880 <= 4'hf;
    end
    if (reset) begin
      image_881 <= 4'h0;
    end else begin
      image_881 <= 4'hf;
    end
    if (reset) begin
      image_882 <= 4'h0;
    end else begin
      image_882 <= 4'hf;
    end
    if (reset) begin
      image_883 <= 4'h0;
    end else begin
      image_883 <= 4'hf;
    end
    if (reset) begin
      image_884 <= 4'h0;
    end else begin
      image_884 <= 4'he;
    end
    if (reset) begin
      image_885 <= 4'h0;
    end else begin
      image_885 <= 4'h9;
    end
    if (reset) begin
      image_891 <= 4'h0;
    end else begin
      image_891 <= 4'h5;
    end
    if (reset) begin
      image_892 <= 4'h0;
    end else begin
      image_892 <= 4'hd;
    end
    if (reset) begin
      image_893 <= 4'h0;
    end else begin
      image_893 <= 4'he;
    end
    if (reset) begin
      image_894 <= 4'h0;
    end else begin
      image_894 <= 4'hb;
    end
    if (reset) begin
      image_895 <= 4'h0;
    end else begin
      image_895 <= 4'h3;
    end
    if (reset) begin
      image_897 <= 4'h0;
    end else begin
      image_897 <= 4'h4;
    end
    if (reset) begin
      image_898 <= 4'h0;
    end else begin
      image_898 <= 4'h5;
    end
    if (reset) begin
      image_899 <= 4'h0;
    end else begin
      image_899 <= 4'h5;
    end
    if (reset) begin
      image_900 <= 4'h0;
    end else begin
      image_900 <= 4'h5;
    end
    if (reset) begin
      image_901 <= 4'h0;
    end else begin
      image_901 <= 4'h6;
    end
    if (reset) begin
      image_902 <= 4'h0;
    end else begin
      image_902 <= 4'h6;
    end
    if (reset) begin
      image_903 <= 4'h0;
    end else begin
      image_903 <= 4'h6;
    end
    if (reset) begin
      image_904 <= 4'h0;
    end else begin
      image_904 <= 4'h6;
    end
    if (reset) begin
      image_905 <= 4'h0;
    end else begin
      image_905 <= 4'h6;
    end
    if (reset) begin
      image_906 <= 4'h0;
    end else begin
      image_906 <= 4'h6;
    end
    if (reset) begin
      image_907 <= 4'h0;
    end else begin
      image_907 <= 4'h6;
    end
    if (reset) begin
      image_908 <= 4'h0;
    end else begin
      image_908 <= 4'h6;
    end
    if (reset) begin
      image_909 <= 4'h0;
    end else begin
      image_909 <= 4'h6;
    end
    if (reset) begin
      image_910 <= 4'h0;
    end else begin
      image_910 <= 4'h6;
    end
    if (reset) begin
      image_911 <= 4'h0;
    end else begin
      image_911 <= 4'h6;
    end
    if (reset) begin
      image_912 <= 4'h0;
    end else begin
      image_912 <= 4'h5;
    end
    if (reset) begin
      image_913 <= 4'h0;
    end else begin
      image_913 <= 4'h6;
    end
    if (reset) begin
      image_914 <= 4'h0;
    end else begin
      image_914 <= 4'hc;
    end
    if (reset) begin
      image_915 <= 4'h0;
    end else begin
      image_915 <= 4'he;
    end
    if (reset) begin
      image_916 <= 4'h0;
    end else begin
      image_916 <= 4'hf;
    end
    if (reset) begin
      image_917 <= 4'h0;
    end else begin
      image_917 <= 4'hf;
    end
    if (reset) begin
      image_918 <= 4'h0;
    end else begin
      image_918 <= 4'hf;
    end
    if (reset) begin
      image_919 <= 4'h0;
    end else begin
      image_919 <= 4'hf;
    end
    if (reset) begin
      image_920 <= 4'h0;
    end else begin
      image_920 <= 4'hf;
    end
    if (reset) begin
      image_921 <= 4'h0;
    end else begin
      image_921 <= 4'hf;
    end
    if (reset) begin
      image_922 <= 4'h0;
    end else begin
      image_922 <= 4'hf;
    end
    if (reset) begin
      image_923 <= 4'h0;
    end else begin
      image_923 <= 4'hf;
    end
    if (reset) begin
      image_924 <= 4'h0;
    end else begin
      image_924 <= 4'hf;
    end
    if (reset) begin
      image_925 <= 4'h0;
    end else begin
      image_925 <= 4'he;
    end
    if (reset) begin
      image_926 <= 4'h0;
    end else begin
      image_926 <= 4'hb;
    end
    if (reset) begin
      image_927 <= 4'h0;
    end else begin
      image_927 <= 4'h1;
    end
    if (reset) begin
      image_929 <= 4'h0;
    end else begin
      image_929 <= 4'h9;
    end
    if (reset) begin
      image_930 <= 4'h0;
    end else begin
      image_930 <= 4'h3;
    end
    if (reset) begin
      image_935 <= 4'h0;
    end else begin
      image_935 <= 4'h8;
    end
    if (reset) begin
      image_936 <= 4'h0;
    end else begin
      image_936 <= 4'he;
    end
    if (reset) begin
      image_937 <= 4'h0;
    end else begin
      image_937 <= 4'hc;
    end
    if (reset) begin
      image_938 <= 4'h0;
    end else begin
      image_938 <= 4'h4;
    end
    if (reset) begin
      image_939 <= 4'h0;
    end else begin
      image_939 <= 4'h5;
    end
    if (reset) begin
      image_940 <= 4'h0;
    end else begin
      image_940 <= 4'h9;
    end
    if (reset) begin
      image_941 <= 4'h0;
    end else begin
      image_941 <= 4'he;
    end
    if (reset) begin
      image_942 <= 4'h0;
    end else begin
      image_942 <= 4'he;
    end
    if (reset) begin
      image_943 <= 4'h0;
    end else begin
      image_943 <= 4'he;
    end
    if (reset) begin
      image_944 <= 4'h0;
    end else begin
      image_944 <= 4'hf;
    end
    if (reset) begin
      image_945 <= 4'h0;
    end else begin
      image_945 <= 4'hf;
    end
    if (reset) begin
      image_946 <= 4'h0;
    end else begin
      image_946 <= 4'hf;
    end
    if (reset) begin
      image_947 <= 4'h0;
    end else begin
      image_947 <= 4'hf;
    end
    if (reset) begin
      image_948 <= 4'h0;
    end else begin
      image_948 <= 4'hf;
    end
    if (reset) begin
      image_949 <= 4'h0;
    end else begin
      image_949 <= 4'he;
    end
    if (reset) begin
      image_950 <= 4'h0;
    end else begin
      image_950 <= 4'hc;
    end
    if (reset) begin
      image_951 <= 4'h0;
    end else begin
      image_951 <= 4'ha;
    end
    if (reset) begin
      image_952 <= 4'h0;
    end else begin
      image_952 <= 4'h8;
    end
    if (reset) begin
      image_953 <= 4'h0;
    end else begin
      image_953 <= 4'h9;
    end
    if (reset) begin
      image_954 <= 4'h0;
    end else begin
      image_954 <= 4'hb;
    end
    if (reset) begin
      image_955 <= 4'h0;
    end else begin
      image_955 <= 4'he;
    end
    if (reset) begin
      image_956 <= 4'h0;
    end else begin
      image_956 <= 4'he;
    end
    if (reset) begin
      image_957 <= 4'h0;
    end else begin
      image_957 <= 4'hb;
    end
    if (reset) begin
      image_958 <= 4'h0;
    end else begin
      image_958 <= 4'h4;
    end
    if (reset) begin
      image_959 <= 4'h0;
    end else begin
      image_959 <= 4'h2;
    end
    if (reset) begin
      image_961 <= 4'h0;
    end else begin
      image_961 <= 4'h5;
    end
    if (reset) begin
      image_962 <= 4'h0;
    end else begin
      image_962 <= 4'h5;
    end
    if (reset) begin
      image_963 <= 4'h0;
    end else begin
      image_963 <= 4'h5;
    end
    if (reset) begin
      image_964 <= 4'h0;
    end else begin
      image_964 <= 4'h5;
    end
    if (reset) begin
      image_965 <= 4'h0;
    end else begin
      image_965 <= 4'h6;
    end
    if (reset) begin
      image_966 <= 4'h0;
    end else begin
      image_966 <= 4'h6;
    end
    if (reset) begin
      image_967 <= 4'h0;
    end else begin
      image_967 <= 4'h6;
    end
    if (reset) begin
      image_968 <= 4'h0;
    end else begin
      image_968 <= 4'h6;
    end
    if (reset) begin
      image_969 <= 4'h0;
    end else begin
      image_969 <= 4'h6;
    end
    if (reset) begin
      image_970 <= 4'h0;
    end else begin
      image_970 <= 4'h6;
    end
    if (reset) begin
      image_971 <= 4'h0;
    end else begin
      image_971 <= 4'h6;
    end
    if (reset) begin
      image_972 <= 4'h0;
    end else begin
      image_972 <= 4'h6;
    end
    if (reset) begin
      image_973 <= 4'h0;
    end else begin
      image_973 <= 4'h6;
    end
    if (reset) begin
      image_974 <= 4'h0;
    end else begin
      image_974 <= 4'h6;
    end
    if (reset) begin
      image_975 <= 4'h0;
    end else begin
      image_975 <= 4'h6;
    end
    if (reset) begin
      image_976 <= 4'h0;
    end else begin
      image_976 <= 4'h6;
    end
    if (reset) begin
      image_977 <= 4'h0;
    end else begin
      image_977 <= 4'h6;
    end
    if (reset) begin
      image_978 <= 4'h0;
    end else begin
      image_978 <= 4'h5;
    end
    if (reset) begin
      image_979 <= 4'h0;
    end else begin
      image_979 <= 4'h9;
    end
    if (reset) begin
      image_980 <= 4'h0;
    end else begin
      image_980 <= 4'he;
    end
    if (reset) begin
      image_981 <= 4'h0;
    end else begin
      image_981 <= 4'hf;
    end
    if (reset) begin
      image_982 <= 4'h0;
    end else begin
      image_982 <= 4'hf;
    end
    if (reset) begin
      image_983 <= 4'h0;
    end else begin
      image_983 <= 4'hf;
    end
    if (reset) begin
      image_984 <= 4'h0;
    end else begin
      image_984 <= 4'hf;
    end
    if (reset) begin
      image_985 <= 4'h0;
    end else begin
      image_985 <= 4'hf;
    end
    if (reset) begin
      image_986 <= 4'h0;
    end else begin
      image_986 <= 4'hf;
    end
    if (reset) begin
      image_987 <= 4'h0;
    end else begin
      image_987 <= 4'hf;
    end
    if (reset) begin
      image_988 <= 4'h0;
    end else begin
      image_988 <= 4'hf;
    end
    if (reset) begin
      image_989 <= 4'h0;
    end else begin
      image_989 <= 4'hf;
    end
    if (reset) begin
      image_990 <= 4'h0;
    end else begin
      image_990 <= 4'he;
    end
    if (reset) begin
      image_991 <= 4'h0;
    end else begin
      image_991 <= 4'hc;
    end
    if (reset) begin
      image_992 <= 4'h0;
    end else begin
      image_992 <= 4'h5;
    end
    if (reset) begin
      image_997 <= 4'h0;
    end else begin
      image_997 <= 4'h3;
    end
    if (reset) begin
      image_998 <= 4'h0;
    end else begin
      image_998 <= 4'ha;
    end
    if (reset) begin
      image_999 <= 4'h0;
    end else begin
      image_999 <= 4'he;
    end
    if (reset) begin
      image_1000 <= 4'h0;
    end else begin
      image_1000 <= 4'hd;
    end
    if (reset) begin
      image_1001 <= 4'h0;
    end else begin
      image_1001 <= 4'h5;
    end
    if (reset) begin
      image_1002 <= 4'h0;
    end else begin
      image_1002 <= 4'h6;
    end
    if (reset) begin
      image_1003 <= 4'h0;
    end else begin
      image_1003 <= 4'h6;
    end
    if (reset) begin
      image_1004 <= 4'h0;
    end else begin
      image_1004 <= 4'h6;
    end
    if (reset) begin
      image_1005 <= 4'h0;
    end else begin
      image_1005 <= 4'h5;
    end
    if (reset) begin
      image_1006 <= 4'h0;
    end else begin
      image_1006 <= 4'h9;
    end
    if (reset) begin
      image_1007 <= 4'h0;
    end else begin
      image_1007 <= 4'hc;
    end
    if (reset) begin
      image_1008 <= 4'h0;
    end else begin
      image_1008 <= 4'he;
    end
    if (reset) begin
      image_1009 <= 4'h0;
    end else begin
      image_1009 <= 4'he;
    end
    if (reset) begin
      image_1010 <= 4'h0;
    end else begin
      image_1010 <= 4'he;
    end
    if (reset) begin
      image_1011 <= 4'h0;
    end else begin
      image_1011 <= 4'he;
    end
    if (reset) begin
      image_1012 <= 4'h0;
    end else begin
      image_1012 <= 4'he;
    end
    if (reset) begin
      image_1013 <= 4'h0;
    end else begin
      image_1013 <= 4'he;
    end
    if (reset) begin
      image_1014 <= 4'h0;
    end else begin
      image_1014 <= 4'he;
    end
    if (reset) begin
      image_1015 <= 4'h0;
    end else begin
      image_1015 <= 4'he;
    end
    if (reset) begin
      image_1016 <= 4'h0;
    end else begin
      image_1016 <= 4'he;
    end
    if (reset) begin
      image_1017 <= 4'h0;
    end else begin
      image_1017 <= 4'he;
    end
    if (reset) begin
      image_1018 <= 4'h0;
    end else begin
      image_1018 <= 4'he;
    end
    if (reset) begin
      image_1019 <= 4'h0;
    end else begin
      image_1019 <= 4'hb;
    end
    if (reset) begin
      image_1020 <= 4'h0;
    end else begin
      image_1020 <= 4'h6;
    end
    if (reset) begin
      image_1024 <= 4'h0;
    end else begin
      image_1024 <= 4'h1;
    end
    if (reset) begin
      image_1025 <= 4'h0;
    end else begin
      image_1025 <= 4'h5;
    end
    if (reset) begin
      image_1026 <= 4'h0;
    end else begin
      image_1026 <= 4'h5;
    end
    if (reset) begin
      image_1027 <= 4'h0;
    end else begin
      image_1027 <= 4'h5;
    end
    if (reset) begin
      image_1028 <= 4'h0;
    end else begin
      image_1028 <= 4'h5;
    end
    if (reset) begin
      image_1029 <= 4'h0;
    end else begin
      image_1029 <= 4'h6;
    end
    if (reset) begin
      image_1030 <= 4'h0;
    end else begin
      image_1030 <= 4'h6;
    end
    if (reset) begin
      image_1031 <= 4'h0;
    end else begin
      image_1031 <= 4'h6;
    end
    if (reset) begin
      image_1032 <= 4'h0;
    end else begin
      image_1032 <= 4'h6;
    end
    if (reset) begin
      image_1033 <= 4'h0;
    end else begin
      image_1033 <= 4'h6;
    end
    if (reset) begin
      image_1034 <= 4'h0;
    end else begin
      image_1034 <= 4'h6;
    end
    if (reset) begin
      image_1035 <= 4'h0;
    end else begin
      image_1035 <= 4'h6;
    end
    if (reset) begin
      image_1036 <= 4'h0;
    end else begin
      image_1036 <= 4'h6;
    end
    if (reset) begin
      image_1037 <= 4'h0;
    end else begin
      image_1037 <= 4'h6;
    end
    if (reset) begin
      image_1038 <= 4'h0;
    end else begin
      image_1038 <= 4'h6;
    end
    if (reset) begin
      image_1039 <= 4'h0;
    end else begin
      image_1039 <= 4'h6;
    end
    if (reset) begin
      image_1040 <= 4'h0;
    end else begin
      image_1040 <= 4'h5;
    end
    if (reset) begin
      image_1041 <= 4'h0;
    end else begin
      image_1041 <= 4'h6;
    end
    if (reset) begin
      image_1042 <= 4'h0;
    end else begin
      image_1042 <= 4'h6;
    end
    if (reset) begin
      image_1043 <= 4'h0;
    end else begin
      image_1043 <= 4'h6;
    end
    if (reset) begin
      image_1044 <= 4'h0;
    end else begin
      image_1044 <= 4'h5;
    end
    if (reset) begin
      image_1045 <= 4'h0;
    end else begin
      image_1045 <= 4'hb;
    end
    if (reset) begin
      image_1046 <= 4'h0;
    end else begin
      image_1046 <= 4'he;
    end
    if (reset) begin
      image_1047 <= 4'h0;
    end else begin
      image_1047 <= 4'he;
    end
    if (reset) begin
      image_1048 <= 4'h0;
    end else begin
      image_1048 <= 4'hf;
    end
    if (reset) begin
      image_1049 <= 4'h0;
    end else begin
      image_1049 <= 4'hf;
    end
    if (reset) begin
      image_1050 <= 4'h0;
    end else begin
      image_1050 <= 4'hf;
    end
    if (reset) begin
      image_1051 <= 4'h0;
    end else begin
      image_1051 <= 4'hf;
    end
    if (reset) begin
      image_1052 <= 4'h0;
    end else begin
      image_1052 <= 4'hf;
    end
    if (reset) begin
      image_1053 <= 4'h0;
    end else begin
      image_1053 <= 4'hf;
    end
    if (reset) begin
      image_1054 <= 4'h0;
    end else begin
      image_1054 <= 4'hf;
    end
    if (reset) begin
      image_1055 <= 4'h0;
    end else begin
      image_1055 <= 4'hf;
    end
    if (reset) begin
      image_1056 <= 4'h0;
    end else begin
      image_1056 <= 4'he;
    end
    if (reset) begin
      image_1057 <= 4'h0;
    end else begin
      image_1057 <= 4'hd;
    end
    if (reset) begin
      image_1058 <= 4'h0;
    end else begin
      image_1058 <= 4'hb;
    end
    if (reset) begin
      image_1059 <= 4'h0;
    end else begin
      image_1059 <= 4'hb;
    end
    if (reset) begin
      image_1060 <= 4'h0;
    end else begin
      image_1060 <= 4'hc;
    end
    if (reset) begin
      image_1061 <= 4'h0;
    end else begin
      image_1061 <= 4'he;
    end
    if (reset) begin
      image_1062 <= 4'h0;
    end else begin
      image_1062 <= 4'he;
    end
    if (reset) begin
      image_1063 <= 4'h0;
    end else begin
      image_1063 <= 4'hb;
    end
    if (reset) begin
      image_1064 <= 4'h0;
    end else begin
      image_1064 <= 4'h4;
    end
    if (reset) begin
      image_1065 <= 4'h0;
    end else begin
      image_1065 <= 4'h6;
    end
    if (reset) begin
      image_1066 <= 4'h0;
    end else begin
      image_1066 <= 4'h6;
    end
    if (reset) begin
      image_1067 <= 4'h0;
    end else begin
      image_1067 <= 4'h6;
    end
    if (reset) begin
      image_1068 <= 4'h0;
    end else begin
      image_1068 <= 4'h6;
    end
    if (reset) begin
      image_1069 <= 4'h0;
    end else begin
      image_1069 <= 4'h6;
    end
    if (reset) begin
      image_1070 <= 4'h0;
    end else begin
      image_1070 <= 4'h6;
    end
    if (reset) begin
      image_1071 <= 4'h0;
    end else begin
      image_1071 <= 4'h5;
    end
    if (reset) begin
      image_1072 <= 4'h0;
    end else begin
      image_1072 <= 4'h5;
    end
    if (reset) begin
      image_1073 <= 4'h0;
    end else begin
      image_1073 <= 4'h6;
    end
    if (reset) begin
      image_1074 <= 4'h0;
    end else begin
      image_1074 <= 4'h8;
    end
    if (reset) begin
      image_1075 <= 4'h0;
    end else begin
      image_1075 <= 4'ha;
    end
    if (reset) begin
      image_1076 <= 4'h0;
    end else begin
      image_1076 <= 4'hb;
    end
    if (reset) begin
      image_1077 <= 4'h0;
    end else begin
      image_1077 <= 4'hb;
    end
    if (reset) begin
      image_1078 <= 4'h0;
    end else begin
      image_1078 <= 4'hb;
    end
    if (reset) begin
      image_1079 <= 4'h0;
    end else begin
      image_1079 <= 4'ha;
    end
    if (reset) begin
      image_1080 <= 4'h0;
    end else begin
      image_1080 <= 4'h9;
    end
    if (reset) begin
      image_1081 <= 4'h0;
    end else begin
      image_1081 <= 4'h7;
    end
    if (reset) begin
      image_1082 <= 4'h0;
    end else begin
      image_1082 <= 4'h5;
    end
    if (reset) begin
      image_1083 <= 4'h0;
    end else begin
      image_1083 <= 4'h5;
    end
    if (reset) begin
      image_1084 <= 4'h0;
    end else begin
      image_1084 <= 4'h6;
    end
    if (reset) begin
      image_1085 <= 4'h0;
    end else begin
      image_1085 <= 4'h1;
    end
    if (reset) begin
      image_1088 <= 4'h0;
    end else begin
      image_1088 <= 4'h2;
    end
    if (reset) begin
      image_1089 <= 4'h0;
    end else begin
      image_1089 <= 4'h5;
    end
    if (reset) begin
      image_1090 <= 4'h0;
    end else begin
      image_1090 <= 4'h5;
    end
    if (reset) begin
      image_1091 <= 4'h0;
    end else begin
      image_1091 <= 4'h5;
    end
    if (reset) begin
      image_1092 <= 4'h0;
    end else begin
      image_1092 <= 4'h5;
    end
    if (reset) begin
      image_1093 <= 4'h0;
    end else begin
      image_1093 <= 4'h6;
    end
    if (reset) begin
      image_1094 <= 4'h0;
    end else begin
      image_1094 <= 4'h6;
    end
    if (reset) begin
      image_1095 <= 4'h0;
    end else begin
      image_1095 <= 4'h6;
    end
    if (reset) begin
      image_1096 <= 4'h0;
    end else begin
      image_1096 <= 4'h6;
    end
    if (reset) begin
      image_1097 <= 4'h0;
    end else begin
      image_1097 <= 4'h6;
    end
    if (reset) begin
      image_1098 <= 4'h0;
    end else begin
      image_1098 <= 4'h6;
    end
    if (reset) begin
      image_1099 <= 4'h0;
    end else begin
      image_1099 <= 4'h6;
    end
    if (reset) begin
      image_1100 <= 4'h0;
    end else begin
      image_1100 <= 4'h6;
    end
    if (reset) begin
      image_1101 <= 4'h0;
    end else begin
      image_1101 <= 4'h6;
    end
    if (reset) begin
      image_1102 <= 4'h0;
    end else begin
      image_1102 <= 4'h6;
    end
    if (reset) begin
      image_1103 <= 4'h0;
    end else begin
      image_1103 <= 4'h6;
    end
    if (reset) begin
      image_1104 <= 4'h0;
    end else begin
      image_1104 <= 4'h6;
    end
    if (reset) begin
      image_1105 <= 4'h0;
    end else begin
      image_1105 <= 4'h4;
    end
    if (reset) begin
      image_1106 <= 4'h0;
    end else begin
      image_1106 <= 4'h5;
    end
    if (reset) begin
      image_1107 <= 4'h0;
    end else begin
      image_1107 <= 4'h6;
    end
    if (reset) begin
      image_1108 <= 4'h0;
    end else begin
      image_1108 <= 4'h6;
    end
    if (reset) begin
      image_1109 <= 4'h0;
    end else begin
      image_1109 <= 4'h5;
    end
    if (reset) begin
      image_1110 <= 4'h0;
    end else begin
      image_1110 <= 4'h6;
    end
    if (reset) begin
      image_1111 <= 4'h0;
    end else begin
      image_1111 <= 4'ha;
    end
    if (reset) begin
      image_1112 <= 4'h0;
    end else begin
      image_1112 <= 4'hd;
    end
    if (reset) begin
      image_1113 <= 4'h0;
    end else begin
      image_1113 <= 4'he;
    end
    if (reset) begin
      image_1114 <= 4'h0;
    end else begin
      image_1114 <= 4'he;
    end
    if (reset) begin
      image_1115 <= 4'h0;
    end else begin
      image_1115 <= 4'he;
    end
    if (reset) begin
      image_1116 <= 4'h0;
    end else begin
      image_1116 <= 4'hf;
    end
    if (reset) begin
      image_1117 <= 4'h0;
    end else begin
      image_1117 <= 4'he;
    end
    if (reset) begin
      image_1118 <= 4'h0;
    end else begin
      image_1118 <= 4'he;
    end
    if (reset) begin
      image_1119 <= 4'h0;
    end else begin
      image_1119 <= 4'hf;
    end
    if (reset) begin
      image_1120 <= 4'h0;
    end else begin
      image_1120 <= 4'he;
    end
    if (reset) begin
      image_1121 <= 4'h0;
    end else begin
      image_1121 <= 4'he;
    end
    if (reset) begin
      image_1122 <= 4'h0;
    end else begin
      image_1122 <= 4'he;
    end
    if (reset) begin
      image_1123 <= 4'h0;
    end else begin
      image_1123 <= 4'he;
    end
    if (reset) begin
      image_1124 <= 4'h0;
    end else begin
      image_1124 <= 4'hd;
    end
    if (reset) begin
      image_1125 <= 4'h0;
    end else begin
      image_1125 <= 4'hb;
    end
    if (reset) begin
      image_1126 <= 4'h0;
    end else begin
      image_1126 <= 4'h6;
    end
    if (reset) begin
      image_1127 <= 4'h0;
    end else begin
      image_1127 <= 4'h4;
    end
    if (reset) begin
      image_1128 <= 4'h0;
    end else begin
      image_1128 <= 4'h5;
    end
    if (reset) begin
      image_1129 <= 4'h0;
    end else begin
      image_1129 <= 4'h6;
    end
    if (reset) begin
      image_1130 <= 4'h0;
    end else begin
      image_1130 <= 4'h6;
    end
    if (reset) begin
      image_1131 <= 4'h0;
    end else begin
      image_1131 <= 4'h6;
    end
    if (reset) begin
      image_1132 <= 4'h0;
    end else begin
      image_1132 <= 4'h6;
    end
    if (reset) begin
      image_1133 <= 4'h0;
    end else begin
      image_1133 <= 4'h6;
    end
    if (reset) begin
      image_1134 <= 4'h0;
    end else begin
      image_1134 <= 4'h6;
    end
    if (reset) begin
      image_1135 <= 4'h0;
    end else begin
      image_1135 <= 4'h5;
    end
    if (reset) begin
      image_1136 <= 4'h0;
    end else begin
      image_1136 <= 4'h5;
    end
    if (reset) begin
      image_1137 <= 4'h0;
    end else begin
      image_1137 <= 4'h6;
    end
    if (reset) begin
      image_1138 <= 4'h0;
    end else begin
      image_1138 <= 4'h6;
    end
    if (reset) begin
      image_1139 <= 4'h0;
    end else begin
      image_1139 <= 4'h6;
    end
    if (reset) begin
      image_1140 <= 4'h0;
    end else begin
      image_1140 <= 4'h6;
    end
    if (reset) begin
      image_1141 <= 4'h0;
    end else begin
      image_1141 <= 4'h6;
    end
    if (reset) begin
      image_1142 <= 4'h0;
    end else begin
      image_1142 <= 4'h6;
    end
    if (reset) begin
      image_1143 <= 4'h0;
    end else begin
      image_1143 <= 4'h6;
    end
    if (reset) begin
      image_1144 <= 4'h0;
    end else begin
      image_1144 <= 4'h7;
    end
    if (reset) begin
      image_1145 <= 4'h0;
    end else begin
      image_1145 <= 4'h6;
    end
    if (reset) begin
      image_1146 <= 4'h0;
    end else begin
      image_1146 <= 4'h5;
    end
    if (reset) begin
      image_1147 <= 4'h0;
    end else begin
      image_1147 <= 4'h4;
    end
    if (reset) begin
      image_1148 <= 4'h0;
    end else begin
      image_1148 <= 4'h2;
    end
    if (reset) begin
      image_1152 <= 4'h0;
    end else begin
      image_1152 <= 4'h3;
    end
    if (reset) begin
      image_1153 <= 4'h0;
    end else begin
      image_1153 <= 4'h5;
    end
    if (reset) begin
      image_1154 <= 4'h0;
    end else begin
      image_1154 <= 4'h5;
    end
    if (reset) begin
      image_1155 <= 4'h0;
    end else begin
      image_1155 <= 4'h5;
    end
    if (reset) begin
      image_1156 <= 4'h0;
    end else begin
      image_1156 <= 4'h5;
    end
    if (reset) begin
      image_1157 <= 4'h0;
    end else begin
      image_1157 <= 4'h6;
    end
    if (reset) begin
      image_1158 <= 4'h0;
    end else begin
      image_1158 <= 4'h6;
    end
    if (reset) begin
      image_1159 <= 4'h0;
    end else begin
      image_1159 <= 4'h6;
    end
    if (reset) begin
      image_1160 <= 4'h0;
    end else begin
      image_1160 <= 4'h6;
    end
    if (reset) begin
      image_1161 <= 4'h0;
    end else begin
      image_1161 <= 4'h6;
    end
    if (reset) begin
      image_1162 <= 4'h0;
    end else begin
      image_1162 <= 4'h6;
    end
    if (reset) begin
      image_1163 <= 4'h0;
    end else begin
      image_1163 <= 4'h6;
    end
    if (reset) begin
      image_1164 <= 4'h0;
    end else begin
      image_1164 <= 4'h6;
    end
    if (reset) begin
      image_1165 <= 4'h0;
    end else begin
      image_1165 <= 4'h6;
    end
    if (reset) begin
      image_1166 <= 4'h0;
    end else begin
      image_1166 <= 4'h6;
    end
    if (reset) begin
      image_1167 <= 4'h0;
    end else begin
      image_1167 <= 4'h6;
    end
    if (reset) begin
      image_1168 <= 4'h0;
    end else begin
      image_1168 <= 4'h6;
    end
    if (reset) begin
      image_1169 <= 4'h0;
    end else begin
      image_1169 <= 4'h6;
    end
    if (reset) begin
      image_1170 <= 4'h0;
    end else begin
      image_1170 <= 4'h6;
    end
    if (reset) begin
      image_1171 <= 4'h0;
    end else begin
      image_1171 <= 4'h4;
    end
    if (reset) begin
      image_1172 <= 4'h0;
    end else begin
      image_1172 <= 4'h5;
    end
    if (reset) begin
      image_1173 <= 4'h0;
    end else begin
      image_1173 <= 4'h6;
    end
    if (reset) begin
      image_1174 <= 4'h0;
    end else begin
      image_1174 <= 4'h6;
    end
    if (reset) begin
      image_1175 <= 4'h0;
    end else begin
      image_1175 <= 4'h6;
    end
    if (reset) begin
      image_1176 <= 4'h0;
    end else begin
      image_1176 <= 4'h5;
    end
    if (reset) begin
      image_1177 <= 4'h0;
    end else begin
      image_1177 <= 4'h5;
    end
    if (reset) begin
      image_1178 <= 4'h0;
    end else begin
      image_1178 <= 4'h8;
    end
    if (reset) begin
      image_1179 <= 4'h0;
    end else begin
      image_1179 <= 4'ha;
    end
    if (reset) begin
      image_1180 <= 4'h0;
    end else begin
      image_1180 <= 4'hb;
    end
    if (reset) begin
      image_1181 <= 4'h0;
    end else begin
      image_1181 <= 4'hb;
    end
    if (reset) begin
      image_1182 <= 4'h0;
    end else begin
      image_1182 <= 4'hc;
    end
    if (reset) begin
      image_1183 <= 4'h0;
    end else begin
      image_1183 <= 4'hc;
    end
    if (reset) begin
      image_1184 <= 4'h0;
    end else begin
      image_1184 <= 4'hb;
    end
    if (reset) begin
      image_1185 <= 4'h0;
    end else begin
      image_1185 <= 4'ha;
    end
    if (reset) begin
      image_1186 <= 4'h0;
    end else begin
      image_1186 <= 4'h8;
    end
    if (reset) begin
      image_1187 <= 4'h0;
    end else begin
      image_1187 <= 4'h6;
    end
    if (reset) begin
      image_1188 <= 4'h0;
    end else begin
      image_1188 <= 4'h4;
    end
    if (reset) begin
      image_1189 <= 4'h0;
    end else begin
      image_1189 <= 4'h5;
    end
    if (reset) begin
      image_1190 <= 4'h0;
    end else begin
      image_1190 <= 4'h6;
    end
    if (reset) begin
      image_1191 <= 4'h0;
    end else begin
      image_1191 <= 4'h3;
    end
    if (reset) begin
      image_1192 <= 4'h0;
    end else begin
      image_1192 <= 4'h6;
    end
    if (reset) begin
      image_1193 <= 4'h0;
    end else begin
      image_1193 <= 4'h6;
    end
    if (reset) begin
      image_1194 <= 4'h0;
    end else begin
      image_1194 <= 4'h6;
    end
    if (reset) begin
      image_1195 <= 4'h0;
    end else begin
      image_1195 <= 4'h6;
    end
    if (reset) begin
      image_1196 <= 4'h0;
    end else begin
      image_1196 <= 4'h6;
    end
    if (reset) begin
      image_1197 <= 4'h0;
    end else begin
      image_1197 <= 4'h6;
    end
    if (reset) begin
      image_1198 <= 4'h0;
    end else begin
      image_1198 <= 4'h6;
    end
    if (reset) begin
      image_1199 <= 4'h0;
    end else begin
      image_1199 <= 4'h6;
    end
    if (reset) begin
      image_1200 <= 4'h0;
    end else begin
      image_1200 <= 4'h6;
    end
    if (reset) begin
      image_1201 <= 4'h0;
    end else begin
      image_1201 <= 4'h5;
    end
    if (reset) begin
      image_1202 <= 4'h0;
    end else begin
      image_1202 <= 4'h4;
    end
    if (reset) begin
      image_1203 <= 4'h0;
    end else begin
      image_1203 <= 4'h4;
    end
    if (reset) begin
      image_1204 <= 4'h0;
    end else begin
      image_1204 <= 4'h4;
    end
    if (reset) begin
      image_1205 <= 4'h0;
    end else begin
      image_1205 <= 4'h4;
    end
    if (reset) begin
      image_1206 <= 4'h0;
    end else begin
      image_1206 <= 4'h4;
    end
    if (reset) begin
      image_1207 <= 4'h0;
    end else begin
      image_1207 <= 4'h4;
    end
    if (reset) begin
      image_1208 <= 4'h0;
    end else begin
      image_1208 <= 4'h3;
    end
    if (reset) begin
      image_1216 <= 4'h0;
    end else begin
      image_1216 <= 4'h3;
    end
    if (reset) begin
      image_1217 <= 4'h0;
    end else begin
      image_1217 <= 4'h5;
    end
    if (reset) begin
      image_1218 <= 4'h0;
    end else begin
      image_1218 <= 4'h5;
    end
    if (reset) begin
      image_1219 <= 4'h0;
    end else begin
      image_1219 <= 4'h5;
    end
    if (reset) begin
      image_1220 <= 4'h0;
    end else begin
      image_1220 <= 4'h5;
    end
    if (reset) begin
      image_1221 <= 4'h0;
    end else begin
      image_1221 <= 4'h6;
    end
    if (reset) begin
      image_1222 <= 4'h0;
    end else begin
      image_1222 <= 4'h6;
    end
    if (reset) begin
      image_1223 <= 4'h0;
    end else begin
      image_1223 <= 4'h6;
    end
    if (reset) begin
      image_1224 <= 4'h0;
    end else begin
      image_1224 <= 4'h6;
    end
    if (reset) begin
      image_1225 <= 4'h0;
    end else begin
      image_1225 <= 4'h6;
    end
    if (reset) begin
      image_1226 <= 4'h0;
    end else begin
      image_1226 <= 4'h6;
    end
    if (reset) begin
      image_1227 <= 4'h0;
    end else begin
      image_1227 <= 4'h6;
    end
    if (reset) begin
      image_1228 <= 4'h0;
    end else begin
      image_1228 <= 4'h6;
    end
    if (reset) begin
      image_1229 <= 4'h0;
    end else begin
      image_1229 <= 4'h6;
    end
    if (reset) begin
      image_1230 <= 4'h0;
    end else begin
      image_1230 <= 4'h6;
    end
    if (reset) begin
      image_1231 <= 4'h0;
    end else begin
      image_1231 <= 4'h6;
    end
    if (reset) begin
      image_1232 <= 4'h0;
    end else begin
      image_1232 <= 4'h6;
    end
    if (reset) begin
      image_1233 <= 4'h0;
    end else begin
      image_1233 <= 4'h6;
    end
    if (reset) begin
      image_1234 <= 4'h0;
    end else begin
      image_1234 <= 4'h6;
    end
    if (reset) begin
      image_1235 <= 4'h0;
    end else begin
      image_1235 <= 4'h6;
    end
    if (reset) begin
      image_1236 <= 4'h0;
    end else begin
      image_1236 <= 4'h6;
    end
    if (reset) begin
      image_1237 <= 4'h0;
    end else begin
      image_1237 <= 4'h5;
    end
    if (reset) begin
      image_1238 <= 4'h0;
    end else begin
      image_1238 <= 4'h4;
    end
    if (reset) begin
      image_1239 <= 4'h0;
    end else begin
      image_1239 <= 4'h4;
    end
    if (reset) begin
      image_1240 <= 4'h0;
    end else begin
      image_1240 <= 4'h5;
    end
    if (reset) begin
      image_1241 <= 4'h0;
    end else begin
      image_1241 <= 4'h6;
    end
    if (reset) begin
      image_1242 <= 4'h0;
    end else begin
      image_1242 <= 4'h6;
    end
    if (reset) begin
      image_1243 <= 4'h0;
    end else begin
      image_1243 <= 4'h6;
    end
    if (reset) begin
      image_1244 <= 4'h0;
    end else begin
      image_1244 <= 4'h6;
    end
    if (reset) begin
      image_1245 <= 4'h0;
    end else begin
      image_1245 <= 4'h6;
    end
    if (reset) begin
      image_1246 <= 4'h0;
    end else begin
      image_1246 <= 4'h5;
    end
    if (reset) begin
      image_1247 <= 4'h0;
    end else begin
      image_1247 <= 4'h5;
    end
    if (reset) begin
      image_1248 <= 4'h0;
    end else begin
      image_1248 <= 4'h6;
    end
    if (reset) begin
      image_1249 <= 4'h0;
    end else begin
      image_1249 <= 4'h6;
    end
    if (reset) begin
      image_1250 <= 4'h0;
    end else begin
      image_1250 <= 4'h6;
    end
    if (reset) begin
      image_1251 <= 4'h0;
    end else begin
      image_1251 <= 4'h6;
    end
    if (reset) begin
      image_1252 <= 4'h0;
    end else begin
      image_1252 <= 4'h6;
    end
    if (reset) begin
      image_1253 <= 4'h0;
    end else begin
      image_1253 <= 4'h5;
    end
    if (reset) begin
      image_1254 <= 4'h0;
    end else begin
      image_1254 <= 4'h3;
    end
    if (reset) begin
      image_1255 <= 4'h0;
    end else begin
      image_1255 <= 4'h5;
    end
    if (reset) begin
      image_1256 <= 4'h0;
    end else begin
      image_1256 <= 4'h6;
    end
    if (reset) begin
      image_1257 <= 4'h0;
    end else begin
      image_1257 <= 4'h6;
    end
    if (reset) begin
      image_1258 <= 4'h0;
    end else begin
      image_1258 <= 4'h6;
    end
    if (reset) begin
      image_1259 <= 4'h0;
    end else begin
      image_1259 <= 4'h6;
    end
    if (reset) begin
      image_1260 <= 4'h0;
    end else begin
      image_1260 <= 4'h6;
    end
    if (reset) begin
      image_1261 <= 4'h0;
    end else begin
      image_1261 <= 4'h6;
    end
    if (reset) begin
      image_1262 <= 4'h0;
    end else begin
      image_1262 <= 4'h6;
    end
    if (reset) begin
      image_1263 <= 4'h0;
    end else begin
      image_1263 <= 4'h6;
    end
    if (reset) begin
      image_1264 <= 4'h0;
    end else begin
      image_1264 <= 4'h6;
    end
    if (reset) begin
      image_1265 <= 4'h0;
    end else begin
      image_1265 <= 4'h6;
    end
    if (reset) begin
      image_1266 <= 4'h0;
    end else begin
      image_1266 <= 4'h6;
    end
    if (reset) begin
      image_1267 <= 4'h0;
    end else begin
      image_1267 <= 4'h6;
    end
    if (reset) begin
      image_1268 <= 4'h0;
    end else begin
      image_1268 <= 4'h6;
    end
    if (reset) begin
      image_1269 <= 4'h0;
    end else begin
      image_1269 <= 4'h6;
    end
    if (reset) begin
      image_1270 <= 4'h0;
    end else begin
      image_1270 <= 4'h6;
    end
    if (reset) begin
      image_1271 <= 4'h0;
    end else begin
      image_1271 <= 4'h6;
    end
    if (reset) begin
      image_1272 <= 4'h0;
    end else begin
      image_1272 <= 4'h6;
    end
    if (reset) begin
      image_1273 <= 4'h0;
    end else begin
      image_1273 <= 4'h5;
    end
    if (reset) begin
      image_1274 <= 4'h0;
    end else begin
      image_1274 <= 4'h3;
    end
    if (reset) begin
      image_1275 <= 4'h0;
    end else begin
      image_1275 <= 4'h1;
    end
    if (reset) begin
      image_1280 <= 4'h0;
    end else begin
      image_1280 <= 4'h3;
    end
    if (reset) begin
      image_1281 <= 4'h0;
    end else begin
      image_1281 <= 4'h5;
    end
    if (reset) begin
      image_1282 <= 4'h0;
    end else begin
      image_1282 <= 4'h5;
    end
    if (reset) begin
      image_1283 <= 4'h0;
    end else begin
      image_1283 <= 4'h5;
    end
    if (reset) begin
      image_1284 <= 4'h0;
    end else begin
      image_1284 <= 4'h5;
    end
    if (reset) begin
      image_1285 <= 4'h0;
    end else begin
      image_1285 <= 4'h6;
    end
    if (reset) begin
      image_1286 <= 4'h0;
    end else begin
      image_1286 <= 4'h6;
    end
    if (reset) begin
      image_1287 <= 4'h0;
    end else begin
      image_1287 <= 4'h6;
    end
    if (reset) begin
      image_1288 <= 4'h0;
    end else begin
      image_1288 <= 4'h6;
    end
    if (reset) begin
      image_1289 <= 4'h0;
    end else begin
      image_1289 <= 4'h6;
    end
    if (reset) begin
      image_1290 <= 4'h0;
    end else begin
      image_1290 <= 4'h6;
    end
    if (reset) begin
      image_1291 <= 4'h0;
    end else begin
      image_1291 <= 4'h6;
    end
    if (reset) begin
      image_1292 <= 4'h0;
    end else begin
      image_1292 <= 4'h6;
    end
    if (reset) begin
      image_1293 <= 4'h0;
    end else begin
      image_1293 <= 4'h6;
    end
    if (reset) begin
      image_1294 <= 4'h0;
    end else begin
      image_1294 <= 4'h6;
    end
    if (reset) begin
      image_1295 <= 4'h0;
    end else begin
      image_1295 <= 4'h6;
    end
    if (reset) begin
      image_1296 <= 4'h0;
    end else begin
      image_1296 <= 4'h6;
    end
    if (reset) begin
      image_1297 <= 4'h0;
    end else begin
      image_1297 <= 4'h6;
    end
    if (reset) begin
      image_1298 <= 4'h0;
    end else begin
      image_1298 <= 4'h6;
    end
    if (reset) begin
      image_1299 <= 4'h0;
    end else begin
      image_1299 <= 4'h6;
    end
    if (reset) begin
      image_1300 <= 4'h0;
    end else begin
      image_1300 <= 4'h6;
    end
    if (reset) begin
      image_1301 <= 4'h0;
    end else begin
      image_1301 <= 4'h6;
    end
    if (reset) begin
      image_1302 <= 4'h0;
    end else begin
      image_1302 <= 4'h6;
    end
    if (reset) begin
      image_1303 <= 4'h0;
    end else begin
      image_1303 <= 4'h6;
    end
    if (reset) begin
      image_1304 <= 4'h0;
    end else begin
      image_1304 <= 4'h6;
    end
    if (reset) begin
      image_1305 <= 4'h0;
    end else begin
      image_1305 <= 4'h5;
    end
    if (reset) begin
      image_1306 <= 4'h0;
    end else begin
      image_1306 <= 4'h4;
    end
    if (reset) begin
      image_1307 <= 4'h0;
    end else begin
      image_1307 <= 4'h4;
    end
    if (reset) begin
      image_1308 <= 4'h0;
    end else begin
      image_1308 <= 4'h4;
    end
    if (reset) begin
      image_1309 <= 4'h0;
    end else begin
      image_1309 <= 4'h5;
    end
    if (reset) begin
      image_1310 <= 4'h0;
    end else begin
      image_1310 <= 4'h4;
    end
    if (reset) begin
      image_1311 <= 4'h0;
    end else begin
      image_1311 <= 4'h4;
    end
    if (reset) begin
      image_1312 <= 4'h0;
    end else begin
      image_1312 <= 4'h4;
    end
    if (reset) begin
      image_1313 <= 4'h0;
    end else begin
      image_1313 <= 4'h4;
    end
    if (reset) begin
      image_1314 <= 4'h0;
    end else begin
      image_1314 <= 4'h4;
    end
    if (reset) begin
      image_1315 <= 4'h0;
    end else begin
      image_1315 <= 4'h4;
    end
    if (reset) begin
      image_1316 <= 4'h0;
    end else begin
      image_1316 <= 4'h4;
    end
    if (reset) begin
      image_1317 <= 4'h0;
    end else begin
      image_1317 <= 4'h5;
    end
    if (reset) begin
      image_1318 <= 4'h0;
    end else begin
      image_1318 <= 4'h6;
    end
    if (reset) begin
      image_1319 <= 4'h0;
    end else begin
      image_1319 <= 4'h6;
    end
    if (reset) begin
      image_1320 <= 4'h0;
    end else begin
      image_1320 <= 4'h6;
    end
    if (reset) begin
      image_1321 <= 4'h0;
    end else begin
      image_1321 <= 4'h6;
    end
    if (reset) begin
      image_1322 <= 4'h0;
    end else begin
      image_1322 <= 4'h6;
    end
    if (reset) begin
      image_1323 <= 4'h0;
    end else begin
      image_1323 <= 4'h6;
    end
    if (reset) begin
      image_1324 <= 4'h0;
    end else begin
      image_1324 <= 4'h6;
    end
    if (reset) begin
      image_1325 <= 4'h0;
    end else begin
      image_1325 <= 4'h6;
    end
    if (reset) begin
      image_1326 <= 4'h0;
    end else begin
      image_1326 <= 4'h6;
    end
    if (reset) begin
      image_1327 <= 4'h0;
    end else begin
      image_1327 <= 4'h6;
    end
    if (reset) begin
      image_1328 <= 4'h0;
    end else begin
      image_1328 <= 4'h6;
    end
    if (reset) begin
      image_1329 <= 4'h0;
    end else begin
      image_1329 <= 4'h6;
    end
    if (reset) begin
      image_1330 <= 4'h0;
    end else begin
      image_1330 <= 4'h6;
    end
    if (reset) begin
      image_1331 <= 4'h0;
    end else begin
      image_1331 <= 4'h6;
    end
    if (reset) begin
      image_1332 <= 4'h0;
    end else begin
      image_1332 <= 4'h6;
    end
    if (reset) begin
      image_1333 <= 4'h0;
    end else begin
      image_1333 <= 4'h6;
    end
    if (reset) begin
      image_1334 <= 4'h0;
    end else begin
      image_1334 <= 4'h6;
    end
    if (reset) begin
      image_1335 <= 4'h0;
    end else begin
      image_1335 <= 4'h6;
    end
    if (reset) begin
      image_1336 <= 4'h0;
    end else begin
      image_1336 <= 4'h6;
    end
    if (reset) begin
      image_1337 <= 4'h0;
    end else begin
      image_1337 <= 4'h6;
    end
    if (reset) begin
      image_1338 <= 4'h0;
    end else begin
      image_1338 <= 4'h6;
    end
    if (reset) begin
      image_1339 <= 4'h0;
    end else begin
      image_1339 <= 4'h6;
    end
    if (reset) begin
      image_1340 <= 4'h0;
    end else begin
      image_1340 <= 4'h4;
    end
    if (reset) begin
      image_1341 <= 4'h0;
    end else begin
      image_1341 <= 4'h1;
    end
    if (reset) begin
      image_1344 <= 4'h0;
    end else begin
      image_1344 <= 4'h3;
    end
    if (reset) begin
      image_1345 <= 4'h0;
    end else begin
      image_1345 <= 4'h5;
    end
    if (reset) begin
      image_1346 <= 4'h0;
    end else begin
      image_1346 <= 4'h5;
    end
    if (reset) begin
      image_1347 <= 4'h0;
    end else begin
      image_1347 <= 4'h5;
    end
    if (reset) begin
      image_1348 <= 4'h0;
    end else begin
      image_1348 <= 4'h5;
    end
    if (reset) begin
      image_1349 <= 4'h0;
    end else begin
      image_1349 <= 4'h6;
    end
    if (reset) begin
      image_1350 <= 4'h0;
    end else begin
      image_1350 <= 4'h6;
    end
    if (reset) begin
      image_1351 <= 4'h0;
    end else begin
      image_1351 <= 4'h6;
    end
    if (reset) begin
      image_1352 <= 4'h0;
    end else begin
      image_1352 <= 4'h6;
    end
    if (reset) begin
      image_1353 <= 4'h0;
    end else begin
      image_1353 <= 4'h6;
    end
    if (reset) begin
      image_1354 <= 4'h0;
    end else begin
      image_1354 <= 4'h6;
    end
    if (reset) begin
      image_1355 <= 4'h0;
    end else begin
      image_1355 <= 4'h6;
    end
    if (reset) begin
      image_1356 <= 4'h0;
    end else begin
      image_1356 <= 4'h6;
    end
    if (reset) begin
      image_1357 <= 4'h0;
    end else begin
      image_1357 <= 4'h6;
    end
    if (reset) begin
      image_1358 <= 4'h0;
    end else begin
      image_1358 <= 4'h6;
    end
    if (reset) begin
      image_1359 <= 4'h0;
    end else begin
      image_1359 <= 4'h6;
    end
    if (reset) begin
      image_1360 <= 4'h0;
    end else begin
      image_1360 <= 4'h6;
    end
    if (reset) begin
      image_1361 <= 4'h0;
    end else begin
      image_1361 <= 4'h6;
    end
    if (reset) begin
      image_1362 <= 4'h0;
    end else begin
      image_1362 <= 4'h6;
    end
    if (reset) begin
      image_1363 <= 4'h0;
    end else begin
      image_1363 <= 4'h6;
    end
    if (reset) begin
      image_1364 <= 4'h0;
    end else begin
      image_1364 <= 4'h6;
    end
    if (reset) begin
      image_1365 <= 4'h0;
    end else begin
      image_1365 <= 4'h6;
    end
    if (reset) begin
      image_1366 <= 4'h0;
    end else begin
      image_1366 <= 4'h6;
    end
    if (reset) begin
      image_1367 <= 4'h0;
    end else begin
      image_1367 <= 4'h6;
    end
    if (reset) begin
      image_1368 <= 4'h0;
    end else begin
      image_1368 <= 4'h6;
    end
    if (reset) begin
      image_1369 <= 4'h0;
    end else begin
      image_1369 <= 4'h6;
    end
    if (reset) begin
      image_1370 <= 4'h0;
    end else begin
      image_1370 <= 4'h6;
    end
    if (reset) begin
      image_1371 <= 4'h0;
    end else begin
      image_1371 <= 4'h6;
    end
    if (reset) begin
      image_1372 <= 4'h0;
    end else begin
      image_1372 <= 4'h6;
    end
    if (reset) begin
      image_1373 <= 4'h0;
    end else begin
      image_1373 <= 4'h6;
    end
    if (reset) begin
      image_1374 <= 4'h0;
    end else begin
      image_1374 <= 4'h6;
    end
    if (reset) begin
      image_1375 <= 4'h0;
    end else begin
      image_1375 <= 4'h6;
    end
    if (reset) begin
      image_1376 <= 4'h0;
    end else begin
      image_1376 <= 4'h6;
    end
    if (reset) begin
      image_1377 <= 4'h0;
    end else begin
      image_1377 <= 4'h6;
    end
    if (reset) begin
      image_1378 <= 4'h0;
    end else begin
      image_1378 <= 4'h6;
    end
    if (reset) begin
      image_1379 <= 4'h0;
    end else begin
      image_1379 <= 4'h6;
    end
    if (reset) begin
      image_1380 <= 4'h0;
    end else begin
      image_1380 <= 4'h6;
    end
    if (reset) begin
      image_1381 <= 4'h0;
    end else begin
      image_1381 <= 4'h6;
    end
    if (reset) begin
      image_1382 <= 4'h0;
    end else begin
      image_1382 <= 4'h6;
    end
    if (reset) begin
      image_1383 <= 4'h0;
    end else begin
      image_1383 <= 4'h6;
    end
    if (reset) begin
      image_1384 <= 4'h0;
    end else begin
      image_1384 <= 4'h6;
    end
    if (reset) begin
      image_1385 <= 4'h0;
    end else begin
      image_1385 <= 4'h6;
    end
    if (reset) begin
      image_1386 <= 4'h0;
    end else begin
      image_1386 <= 4'h6;
    end
    if (reset) begin
      image_1387 <= 4'h0;
    end else begin
      image_1387 <= 4'h6;
    end
    if (reset) begin
      image_1388 <= 4'h0;
    end else begin
      image_1388 <= 4'h6;
    end
    if (reset) begin
      image_1389 <= 4'h0;
    end else begin
      image_1389 <= 4'h6;
    end
    if (reset) begin
      image_1390 <= 4'h0;
    end else begin
      image_1390 <= 4'h6;
    end
    if (reset) begin
      image_1391 <= 4'h0;
    end else begin
      image_1391 <= 4'h6;
    end
    if (reset) begin
      image_1392 <= 4'h0;
    end else begin
      image_1392 <= 4'h6;
    end
    if (reset) begin
      image_1393 <= 4'h0;
    end else begin
      image_1393 <= 4'h6;
    end
    if (reset) begin
      image_1394 <= 4'h0;
    end else begin
      image_1394 <= 4'h5;
    end
    if (reset) begin
      image_1395 <= 4'h0;
    end else begin
      image_1395 <= 4'h5;
    end
    if (reset) begin
      image_1396 <= 4'h0;
    end else begin
      image_1396 <= 4'h5;
    end
    if (reset) begin
      image_1397 <= 4'h0;
    end else begin
      image_1397 <= 4'h5;
    end
    if (reset) begin
      image_1398 <= 4'h0;
    end else begin
      image_1398 <= 4'h5;
    end
    if (reset) begin
      image_1399 <= 4'h0;
    end else begin
      image_1399 <= 4'h6;
    end
    if (reset) begin
      image_1400 <= 4'h0;
    end else begin
      image_1400 <= 4'h6;
    end
    if (reset) begin
      image_1401 <= 4'h0;
    end else begin
      image_1401 <= 4'h6;
    end
    if (reset) begin
      image_1402 <= 4'h0;
    end else begin
      image_1402 <= 4'h6;
    end
    if (reset) begin
      image_1403 <= 4'h0;
    end else begin
      image_1403 <= 4'h6;
    end
    if (reset) begin
      image_1404 <= 4'h0;
    end else begin
      image_1404 <= 4'h6;
    end
    if (reset) begin
      image_1405 <= 4'h0;
    end else begin
      image_1405 <= 4'h4;
    end
    if (reset) begin
      image_1408 <= 4'h0;
    end else begin
      image_1408 <= 4'h3;
    end
    if (reset) begin
      image_1409 <= 4'h0;
    end else begin
      image_1409 <= 4'h5;
    end
    if (reset) begin
      image_1410 <= 4'h0;
    end else begin
      image_1410 <= 4'h5;
    end
    if (reset) begin
      image_1411 <= 4'h0;
    end else begin
      image_1411 <= 4'h5;
    end
    if (reset) begin
      image_1412 <= 4'h0;
    end else begin
      image_1412 <= 4'h5;
    end
    if (reset) begin
      image_1413 <= 4'h0;
    end else begin
      image_1413 <= 4'h6;
    end
    if (reset) begin
      image_1414 <= 4'h0;
    end else begin
      image_1414 <= 4'h6;
    end
    if (reset) begin
      image_1415 <= 4'h0;
    end else begin
      image_1415 <= 4'h6;
    end
    if (reset) begin
      image_1416 <= 4'h0;
    end else begin
      image_1416 <= 4'h6;
    end
    if (reset) begin
      image_1417 <= 4'h0;
    end else begin
      image_1417 <= 4'h6;
    end
    if (reset) begin
      image_1418 <= 4'h0;
    end else begin
      image_1418 <= 4'h6;
    end
    if (reset) begin
      image_1419 <= 4'h0;
    end else begin
      image_1419 <= 4'h6;
    end
    if (reset) begin
      image_1420 <= 4'h0;
    end else begin
      image_1420 <= 4'h6;
    end
    if (reset) begin
      image_1421 <= 4'h0;
    end else begin
      image_1421 <= 4'h6;
    end
    if (reset) begin
      image_1422 <= 4'h0;
    end else begin
      image_1422 <= 4'h6;
    end
    if (reset) begin
      image_1423 <= 4'h0;
    end else begin
      image_1423 <= 4'h6;
    end
    if (reset) begin
      image_1424 <= 4'h0;
    end else begin
      image_1424 <= 4'h6;
    end
    if (reset) begin
      image_1425 <= 4'h0;
    end else begin
      image_1425 <= 4'h6;
    end
    if (reset) begin
      image_1426 <= 4'h0;
    end else begin
      image_1426 <= 4'h6;
    end
    if (reset) begin
      image_1427 <= 4'h0;
    end else begin
      image_1427 <= 4'h6;
    end
    if (reset) begin
      image_1428 <= 4'h0;
    end else begin
      image_1428 <= 4'h6;
    end
    if (reset) begin
      image_1429 <= 4'h0;
    end else begin
      image_1429 <= 4'h6;
    end
    if (reset) begin
      image_1430 <= 4'h0;
    end else begin
      image_1430 <= 4'h6;
    end
    if (reset) begin
      image_1431 <= 4'h0;
    end else begin
      image_1431 <= 4'h6;
    end
    if (reset) begin
      image_1432 <= 4'h0;
    end else begin
      image_1432 <= 4'h6;
    end
    if (reset) begin
      image_1433 <= 4'h0;
    end else begin
      image_1433 <= 4'h6;
    end
    if (reset) begin
      image_1434 <= 4'h0;
    end else begin
      image_1434 <= 4'h6;
    end
    if (reset) begin
      image_1435 <= 4'h0;
    end else begin
      image_1435 <= 4'h6;
    end
    if (reset) begin
      image_1436 <= 4'h0;
    end else begin
      image_1436 <= 4'h6;
    end
    if (reset) begin
      image_1437 <= 4'h0;
    end else begin
      image_1437 <= 4'h6;
    end
    if (reset) begin
      image_1438 <= 4'h0;
    end else begin
      image_1438 <= 4'h6;
    end
    if (reset) begin
      image_1439 <= 4'h0;
    end else begin
      image_1439 <= 4'h6;
    end
    if (reset) begin
      image_1440 <= 4'h0;
    end else begin
      image_1440 <= 4'h6;
    end
    if (reset) begin
      image_1441 <= 4'h0;
    end else begin
      image_1441 <= 4'h6;
    end
    if (reset) begin
      image_1442 <= 4'h0;
    end else begin
      image_1442 <= 4'h6;
    end
    if (reset) begin
      image_1443 <= 4'h0;
    end else begin
      image_1443 <= 4'h6;
    end
    if (reset) begin
      image_1444 <= 4'h0;
    end else begin
      image_1444 <= 4'h6;
    end
    if (reset) begin
      image_1445 <= 4'h0;
    end else begin
      image_1445 <= 4'h6;
    end
    if (reset) begin
      image_1446 <= 4'h0;
    end else begin
      image_1446 <= 4'h6;
    end
    if (reset) begin
      image_1447 <= 4'h0;
    end else begin
      image_1447 <= 4'h6;
    end
    if (reset) begin
      image_1448 <= 4'h0;
    end else begin
      image_1448 <= 4'h5;
    end
    if (reset) begin
      image_1449 <= 4'h0;
    end else begin
      image_1449 <= 4'h5;
    end
    if (reset) begin
      image_1450 <= 4'h0;
    end else begin
      image_1450 <= 4'h4;
    end
    if (reset) begin
      image_1451 <= 4'h0;
    end else begin
      image_1451 <= 4'h4;
    end
    if (reset) begin
      image_1452 <= 4'h0;
    end else begin
      image_1452 <= 4'h5;
    end
    if (reset) begin
      image_1453 <= 4'h0;
    end else begin
      image_1453 <= 4'h4;
    end
    if (reset) begin
      image_1454 <= 4'h0;
    end else begin
      image_1454 <= 4'h4;
    end
    if (reset) begin
      image_1455 <= 4'h0;
    end else begin
      image_1455 <= 4'h4;
    end
    if (reset) begin
      image_1456 <= 4'h0;
    end else begin
      image_1456 <= 4'h5;
    end
    if (reset) begin
      image_1457 <= 4'h0;
    end else begin
      image_1457 <= 4'h5;
    end
    if (reset) begin
      image_1458 <= 4'h0;
    end else begin
      image_1458 <= 4'h5;
    end
    if (reset) begin
      image_1459 <= 4'h0;
    end else begin
      image_1459 <= 4'h5;
    end
    if (reset) begin
      image_1460 <= 4'h0;
    end else begin
      image_1460 <= 4'h5;
    end
    if (reset) begin
      image_1461 <= 4'h0;
    end else begin
      image_1461 <= 4'h5;
    end
    if (reset) begin
      image_1462 <= 4'h0;
    end else begin
      image_1462 <= 4'h5;
    end
    if (reset) begin
      image_1463 <= 4'h0;
    end else begin
      image_1463 <= 4'h5;
    end
    if (reset) begin
      image_1464 <= 4'h0;
    end else begin
      image_1464 <= 4'h5;
    end
    if (reset) begin
      image_1465 <= 4'h0;
    end else begin
      image_1465 <= 4'h4;
    end
    if (reset) begin
      image_1466 <= 4'h0;
    end else begin
      image_1466 <= 4'h4;
    end
    if (reset) begin
      image_1467 <= 4'h0;
    end else begin
      image_1467 <= 4'h4;
    end
    if (reset) begin
      image_1468 <= 4'h0;
    end else begin
      image_1468 <= 4'h5;
    end
    if (reset) begin
      image_1469 <= 4'h0;
    end else begin
      image_1469 <= 4'h4;
    end
    if (reset) begin
      image_1472 <= 4'h0;
    end else begin
      image_1472 <= 4'h3;
    end
    if (reset) begin
      image_1473 <= 4'h0;
    end else begin
      image_1473 <= 4'h5;
    end
    if (reset) begin
      image_1474 <= 4'h0;
    end else begin
      image_1474 <= 4'h5;
    end
    if (reset) begin
      image_1475 <= 4'h0;
    end else begin
      image_1475 <= 4'h5;
    end
    if (reset) begin
      image_1476 <= 4'h0;
    end else begin
      image_1476 <= 4'h5;
    end
    if (reset) begin
      image_1477 <= 4'h0;
    end else begin
      image_1477 <= 4'h6;
    end
    if (reset) begin
      image_1478 <= 4'h0;
    end else begin
      image_1478 <= 4'h6;
    end
    if (reset) begin
      image_1479 <= 4'h0;
    end else begin
      image_1479 <= 4'h6;
    end
    if (reset) begin
      image_1480 <= 4'h0;
    end else begin
      image_1480 <= 4'h6;
    end
    if (reset) begin
      image_1481 <= 4'h0;
    end else begin
      image_1481 <= 4'h6;
    end
    if (reset) begin
      image_1482 <= 4'h0;
    end else begin
      image_1482 <= 4'h6;
    end
    if (reset) begin
      image_1483 <= 4'h0;
    end else begin
      image_1483 <= 4'h6;
    end
    if (reset) begin
      image_1484 <= 4'h0;
    end else begin
      image_1484 <= 4'h6;
    end
    if (reset) begin
      image_1485 <= 4'h0;
    end else begin
      image_1485 <= 4'h6;
    end
    if (reset) begin
      image_1486 <= 4'h0;
    end else begin
      image_1486 <= 4'h6;
    end
    if (reset) begin
      image_1487 <= 4'h0;
    end else begin
      image_1487 <= 4'h6;
    end
    if (reset) begin
      image_1488 <= 4'h0;
    end else begin
      image_1488 <= 4'h6;
    end
    if (reset) begin
      image_1489 <= 4'h0;
    end else begin
      image_1489 <= 4'h6;
    end
    if (reset) begin
      image_1490 <= 4'h0;
    end else begin
      image_1490 <= 4'h6;
    end
    if (reset) begin
      image_1491 <= 4'h0;
    end else begin
      image_1491 <= 4'h6;
    end
    if (reset) begin
      image_1492 <= 4'h0;
    end else begin
      image_1492 <= 4'h6;
    end
    if (reset) begin
      image_1493 <= 4'h0;
    end else begin
      image_1493 <= 4'h6;
    end
    if (reset) begin
      image_1494 <= 4'h0;
    end else begin
      image_1494 <= 4'h6;
    end
    if (reset) begin
      image_1495 <= 4'h0;
    end else begin
      image_1495 <= 4'h6;
    end
    if (reset) begin
      image_1496 <= 4'h0;
    end else begin
      image_1496 <= 4'h6;
    end
    if (reset) begin
      image_1497 <= 4'h0;
    end else begin
      image_1497 <= 4'h6;
    end
    if (reset) begin
      image_1498 <= 4'h0;
    end else begin
      image_1498 <= 4'h6;
    end
    if (reset) begin
      image_1499 <= 4'h0;
    end else begin
      image_1499 <= 4'h6;
    end
    if (reset) begin
      image_1500 <= 4'h0;
    end else begin
      image_1500 <= 4'h6;
    end
    if (reset) begin
      image_1501 <= 4'h0;
    end else begin
      image_1501 <= 4'h6;
    end
    if (reset) begin
      image_1502 <= 4'h0;
    end else begin
      image_1502 <= 4'h6;
    end
    if (reset) begin
      image_1503 <= 4'h0;
    end else begin
      image_1503 <= 4'h6;
    end
    if (reset) begin
      image_1504 <= 4'h0;
    end else begin
      image_1504 <= 4'h6;
    end
    if (reset) begin
      image_1505 <= 4'h0;
    end else begin
      image_1505 <= 4'h6;
    end
    if (reset) begin
      image_1506 <= 4'h0;
    end else begin
      image_1506 <= 4'h5;
    end
    if (reset) begin
      image_1507 <= 4'h0;
    end else begin
      image_1507 <= 4'h5;
    end
    if (reset) begin
      image_1508 <= 4'h0;
    end else begin
      image_1508 <= 4'h4;
    end
    if (reset) begin
      image_1509 <= 4'h0;
    end else begin
      image_1509 <= 4'h4;
    end
    if (reset) begin
      image_1510 <= 4'h0;
    end else begin
      image_1510 <= 4'h4;
    end
    if (reset) begin
      image_1511 <= 4'h0;
    end else begin
      image_1511 <= 4'h5;
    end
    if (reset) begin
      image_1512 <= 4'h0;
    end else begin
      image_1512 <= 4'h5;
    end
    if (reset) begin
      image_1513 <= 4'h0;
    end else begin
      image_1513 <= 4'h6;
    end
    if (reset) begin
      image_1514 <= 4'h0;
    end else begin
      image_1514 <= 4'h6;
    end
    if (reset) begin
      image_1515 <= 4'h0;
    end else begin
      image_1515 <= 4'h6;
    end
    if (reset) begin
      image_1516 <= 4'h0;
    end else begin
      image_1516 <= 4'h6;
    end
    if (reset) begin
      image_1517 <= 4'h0;
    end else begin
      image_1517 <= 4'h6;
    end
    if (reset) begin
      image_1518 <= 4'h0;
    end else begin
      image_1518 <= 4'h6;
    end
    if (reset) begin
      image_1519 <= 4'h0;
    end else begin
      image_1519 <= 4'h6;
    end
    if (reset) begin
      image_1520 <= 4'h0;
    end else begin
      image_1520 <= 4'h6;
    end
    if (reset) begin
      image_1521 <= 4'h0;
    end else begin
      image_1521 <= 4'h6;
    end
    if (reset) begin
      image_1522 <= 4'h0;
    end else begin
      image_1522 <= 4'h6;
    end
    if (reset) begin
      image_1523 <= 4'h0;
    end else begin
      image_1523 <= 4'h6;
    end
    if (reset) begin
      image_1524 <= 4'h0;
    end else begin
      image_1524 <= 4'h6;
    end
    if (reset) begin
      image_1525 <= 4'h0;
    end else begin
      image_1525 <= 4'h6;
    end
    if (reset) begin
      image_1526 <= 4'h0;
    end else begin
      image_1526 <= 4'h6;
    end
    if (reset) begin
      image_1527 <= 4'h0;
    end else begin
      image_1527 <= 4'h6;
    end
    if (reset) begin
      image_1528 <= 4'h0;
    end else begin
      image_1528 <= 4'h6;
    end
    if (reset) begin
      image_1529 <= 4'h0;
    end else begin
      image_1529 <= 4'h6;
    end
    if (reset) begin
      image_1530 <= 4'h0;
    end else begin
      image_1530 <= 4'h6;
    end
    if (reset) begin
      image_1531 <= 4'h0;
    end else begin
      image_1531 <= 4'h6;
    end
    if (reset) begin
      image_1532 <= 4'h0;
    end else begin
      image_1532 <= 4'h5;
    end
    if (reset) begin
      image_1533 <= 4'h0;
    end else begin
      image_1533 <= 4'h2;
    end
    if (reset) begin
      image_1536 <= 4'h0;
    end else begin
      image_1536 <= 4'h3;
    end
    if (reset) begin
      image_1537 <= 4'h0;
    end else begin
      image_1537 <= 4'h5;
    end
    if (reset) begin
      image_1538 <= 4'h0;
    end else begin
      image_1538 <= 4'h5;
    end
    if (reset) begin
      image_1539 <= 4'h0;
    end else begin
      image_1539 <= 4'h5;
    end
    if (reset) begin
      image_1540 <= 4'h0;
    end else begin
      image_1540 <= 4'h5;
    end
    if (reset) begin
      image_1541 <= 4'h0;
    end else begin
      image_1541 <= 4'h6;
    end
    if (reset) begin
      image_1542 <= 4'h0;
    end else begin
      image_1542 <= 4'h6;
    end
    if (reset) begin
      image_1543 <= 4'h0;
    end else begin
      image_1543 <= 4'h6;
    end
    if (reset) begin
      image_1544 <= 4'h0;
    end else begin
      image_1544 <= 4'h6;
    end
    if (reset) begin
      image_1545 <= 4'h0;
    end else begin
      image_1545 <= 4'h6;
    end
    if (reset) begin
      image_1546 <= 4'h0;
    end else begin
      image_1546 <= 4'h6;
    end
    if (reset) begin
      image_1547 <= 4'h0;
    end else begin
      image_1547 <= 4'h6;
    end
    if (reset) begin
      image_1548 <= 4'h0;
    end else begin
      image_1548 <= 4'h6;
    end
    if (reset) begin
      image_1549 <= 4'h0;
    end else begin
      image_1549 <= 4'h6;
    end
    if (reset) begin
      image_1550 <= 4'h0;
    end else begin
      image_1550 <= 4'h6;
    end
    if (reset) begin
      image_1551 <= 4'h0;
    end else begin
      image_1551 <= 4'h6;
    end
    if (reset) begin
      image_1552 <= 4'h0;
    end else begin
      image_1552 <= 4'h6;
    end
    if (reset) begin
      image_1553 <= 4'h0;
    end else begin
      image_1553 <= 4'h6;
    end
    if (reset) begin
      image_1554 <= 4'h0;
    end else begin
      image_1554 <= 4'h6;
    end
    if (reset) begin
      image_1555 <= 4'h0;
    end else begin
      image_1555 <= 4'h6;
    end
    if (reset) begin
      image_1556 <= 4'h0;
    end else begin
      image_1556 <= 4'h6;
    end
    if (reset) begin
      image_1557 <= 4'h0;
    end else begin
      image_1557 <= 4'h6;
    end
    if (reset) begin
      image_1558 <= 4'h0;
    end else begin
      image_1558 <= 4'h6;
    end
    if (reset) begin
      image_1559 <= 4'h0;
    end else begin
      image_1559 <= 4'h6;
    end
    if (reset) begin
      image_1560 <= 4'h0;
    end else begin
      image_1560 <= 4'h6;
    end
    if (reset) begin
      image_1561 <= 4'h0;
    end else begin
      image_1561 <= 4'h6;
    end
    if (reset) begin
      image_1562 <= 4'h0;
    end else begin
      image_1562 <= 4'h6;
    end
    if (reset) begin
      image_1563 <= 4'h0;
    end else begin
      image_1563 <= 4'h6;
    end
    if (reset) begin
      image_1564 <= 4'h0;
    end else begin
      image_1564 <= 4'h6;
    end
    if (reset) begin
      image_1565 <= 4'h0;
    end else begin
      image_1565 <= 4'h6;
    end
    if (reset) begin
      image_1566 <= 4'h0;
    end else begin
      image_1566 <= 4'h5;
    end
    if (reset) begin
      image_1567 <= 4'h0;
    end else begin
      image_1567 <= 4'h4;
    end
    if (reset) begin
      image_1568 <= 4'h0;
    end else begin
      image_1568 <= 4'h4;
    end
    if (reset) begin
      image_1569 <= 4'h0;
    end else begin
      image_1569 <= 4'h5;
    end
    if (reset) begin
      image_1570 <= 4'h0;
    end else begin
      image_1570 <= 4'h5;
    end
    if (reset) begin
      image_1571 <= 4'h0;
    end else begin
      image_1571 <= 4'h6;
    end
    if (reset) begin
      image_1572 <= 4'h0;
    end else begin
      image_1572 <= 4'h6;
    end
    if (reset) begin
      image_1573 <= 4'h0;
    end else begin
      image_1573 <= 4'h6;
    end
    if (reset) begin
      image_1574 <= 4'h0;
    end else begin
      image_1574 <= 4'h6;
    end
    if (reset) begin
      image_1575 <= 4'h0;
    end else begin
      image_1575 <= 4'h6;
    end
    if (reset) begin
      image_1576 <= 4'h0;
    end else begin
      image_1576 <= 4'h6;
    end
    if (reset) begin
      image_1577 <= 4'h0;
    end else begin
      image_1577 <= 4'h6;
    end
    if (reset) begin
      image_1578 <= 4'h0;
    end else begin
      image_1578 <= 4'h6;
    end
    if (reset) begin
      image_1579 <= 4'h0;
    end else begin
      image_1579 <= 4'h6;
    end
    if (reset) begin
      image_1580 <= 4'h0;
    end else begin
      image_1580 <= 4'h6;
    end
    if (reset) begin
      image_1581 <= 4'h0;
    end else begin
      image_1581 <= 4'h5;
    end
    if (reset) begin
      image_1582 <= 4'h0;
    end else begin
      image_1582 <= 4'h5;
    end
    if (reset) begin
      image_1583 <= 4'h0;
    end else begin
      image_1583 <= 4'h4;
    end
    if (reset) begin
      image_1584 <= 4'h0;
    end else begin
      image_1584 <= 4'h4;
    end
    if (reset) begin
      image_1585 <= 4'h0;
    end else begin
      image_1585 <= 4'h4;
    end
    if (reset) begin
      image_1586 <= 4'h0;
    end else begin
      image_1586 <= 4'h4;
    end
    if (reset) begin
      image_1587 <= 4'h0;
    end else begin
      image_1587 <= 4'h4;
    end
    if (reset) begin
      image_1588 <= 4'h0;
    end else begin
      image_1588 <= 4'h4;
    end
    if (reset) begin
      image_1589 <= 4'h0;
    end else begin
      image_1589 <= 4'h4;
    end
    if (reset) begin
      image_1590 <= 4'h0;
    end else begin
      image_1590 <= 4'h4;
    end
    if (reset) begin
      image_1591 <= 4'h0;
    end else begin
      image_1591 <= 4'h4;
    end
    if (reset) begin
      image_1592 <= 4'h0;
    end else begin
      image_1592 <= 4'h5;
    end
    if (reset) begin
      image_1593 <= 4'h0;
    end else begin
      image_1593 <= 4'h6;
    end
    if (reset) begin
      image_1594 <= 4'h0;
    end else begin
      image_1594 <= 4'h6;
    end
    if (reset) begin
      image_1595 <= 4'h0;
    end else begin
      image_1595 <= 4'h6;
    end
    if (reset) begin
      image_1596 <= 4'h0;
    end else begin
      image_1596 <= 4'h6;
    end
    if (reset) begin
      image_1597 <= 4'h0;
    end else begin
      image_1597 <= 4'h3;
    end
    if (reset) begin
      image_1600 <= 4'h0;
    end else begin
      image_1600 <= 4'h3;
    end
    if (reset) begin
      image_1601 <= 4'h0;
    end else begin
      image_1601 <= 4'h5;
    end
    if (reset) begin
      image_1602 <= 4'h0;
    end else begin
      image_1602 <= 4'h5;
    end
    if (reset) begin
      image_1603 <= 4'h0;
    end else begin
      image_1603 <= 4'h5;
    end
    if (reset) begin
      image_1604 <= 4'h0;
    end else begin
      image_1604 <= 4'h5;
    end
    if (reset) begin
      image_1605 <= 4'h0;
    end else begin
      image_1605 <= 4'h6;
    end
    if (reset) begin
      image_1606 <= 4'h0;
    end else begin
      image_1606 <= 4'h6;
    end
    if (reset) begin
      image_1607 <= 4'h0;
    end else begin
      image_1607 <= 4'h6;
    end
    if (reset) begin
      image_1608 <= 4'h0;
    end else begin
      image_1608 <= 4'h6;
    end
    if (reset) begin
      image_1609 <= 4'h0;
    end else begin
      image_1609 <= 4'h6;
    end
    if (reset) begin
      image_1610 <= 4'h0;
    end else begin
      image_1610 <= 4'h6;
    end
    if (reset) begin
      image_1611 <= 4'h0;
    end else begin
      image_1611 <= 4'h6;
    end
    if (reset) begin
      image_1612 <= 4'h0;
    end else begin
      image_1612 <= 4'h6;
    end
    if (reset) begin
      image_1613 <= 4'h0;
    end else begin
      image_1613 <= 4'h6;
    end
    if (reset) begin
      image_1614 <= 4'h0;
    end else begin
      image_1614 <= 4'h6;
    end
    if (reset) begin
      image_1615 <= 4'h0;
    end else begin
      image_1615 <= 4'h6;
    end
    if (reset) begin
      image_1616 <= 4'h0;
    end else begin
      image_1616 <= 4'h6;
    end
    if (reset) begin
      image_1617 <= 4'h0;
    end else begin
      image_1617 <= 4'h6;
    end
    if (reset) begin
      image_1618 <= 4'h0;
    end else begin
      image_1618 <= 4'h6;
    end
    if (reset) begin
      image_1619 <= 4'h0;
    end else begin
      image_1619 <= 4'h6;
    end
    if (reset) begin
      image_1620 <= 4'h0;
    end else begin
      image_1620 <= 4'h6;
    end
    if (reset) begin
      image_1621 <= 4'h0;
    end else begin
      image_1621 <= 4'h6;
    end
    if (reset) begin
      image_1622 <= 4'h0;
    end else begin
      image_1622 <= 4'h6;
    end
    if (reset) begin
      image_1623 <= 4'h0;
    end else begin
      image_1623 <= 4'h6;
    end
    if (reset) begin
      image_1624 <= 4'h0;
    end else begin
      image_1624 <= 4'h6;
    end
    if (reset) begin
      image_1625 <= 4'h0;
    end else begin
      image_1625 <= 4'h6;
    end
    if (reset) begin
      image_1626 <= 4'h0;
    end else begin
      image_1626 <= 4'h5;
    end
    if (reset) begin
      image_1627 <= 4'h0;
    end else begin
      image_1627 <= 4'h4;
    end
    if (reset) begin
      image_1628 <= 4'h0;
    end else begin
      image_1628 <= 4'h4;
    end
    if (reset) begin
      image_1629 <= 4'h0;
    end else begin
      image_1629 <= 4'h5;
    end
    if (reset) begin
      image_1630 <= 4'h0;
    end else begin
      image_1630 <= 4'h6;
    end
    if (reset) begin
      image_1631 <= 4'h0;
    end else begin
      image_1631 <= 4'h6;
    end
    if (reset) begin
      image_1632 <= 4'h0;
    end else begin
      image_1632 <= 4'h6;
    end
    if (reset) begin
      image_1633 <= 4'h0;
    end else begin
      image_1633 <= 4'h6;
    end
    if (reset) begin
      image_1634 <= 4'h0;
    end else begin
      image_1634 <= 4'h6;
    end
    if (reset) begin
      image_1635 <= 4'h0;
    end else begin
      image_1635 <= 4'h6;
    end
    if (reset) begin
      image_1636 <= 4'h0;
    end else begin
      image_1636 <= 4'h6;
    end
    if (reset) begin
      image_1637 <= 4'h0;
    end else begin
      image_1637 <= 4'h6;
    end
    if (reset) begin
      image_1638 <= 4'h0;
    end else begin
      image_1638 <= 4'h5;
    end
    if (reset) begin
      image_1639 <= 4'h0;
    end else begin
      image_1639 <= 4'h5;
    end
    if (reset) begin
      image_1640 <= 4'h0;
    end else begin
      image_1640 <= 4'h4;
    end
    if (reset) begin
      image_1641 <= 4'h0;
    end else begin
      image_1641 <= 4'h4;
    end
    if (reset) begin
      image_1642 <= 4'h0;
    end else begin
      image_1642 <= 4'h4;
    end
    if (reset) begin
      image_1643 <= 4'h0;
    end else begin
      image_1643 <= 4'h3;
    end
    if (reset) begin
      image_1644 <= 4'h0;
    end else begin
      image_1644 <= 4'h4;
    end
    if (reset) begin
      image_1645 <= 4'h0;
    end else begin
      image_1645 <= 4'h4;
    end
    if (reset) begin
      image_1646 <= 4'h0;
    end else begin
      image_1646 <= 4'h5;
    end
    if (reset) begin
      image_1647 <= 4'h0;
    end else begin
      image_1647 <= 4'h5;
    end
    if (reset) begin
      image_1648 <= 4'h0;
    end else begin
      image_1648 <= 4'h5;
    end
    if (reset) begin
      image_1649 <= 4'h0;
    end else begin
      image_1649 <= 4'h6;
    end
    if (reset) begin
      image_1650 <= 4'h0;
    end else begin
      image_1650 <= 4'h6;
    end
    if (reset) begin
      image_1651 <= 4'h0;
    end else begin
      image_1651 <= 4'h6;
    end
    if (reset) begin
      image_1652 <= 4'h0;
    end else begin
      image_1652 <= 4'h6;
    end
    if (reset) begin
      image_1653 <= 4'h0;
    end else begin
      image_1653 <= 4'h6;
    end
    if (reset) begin
      image_1654 <= 4'h0;
    end else begin
      image_1654 <= 4'h6;
    end
    if (reset) begin
      image_1655 <= 4'h0;
    end else begin
      image_1655 <= 4'h6;
    end
    if (reset) begin
      image_1656 <= 4'h0;
    end else begin
      image_1656 <= 4'h4;
    end
    if (reset) begin
      image_1657 <= 4'h0;
    end else begin
      image_1657 <= 4'h5;
    end
    if (reset) begin
      image_1658 <= 4'h0;
    end else begin
      image_1658 <= 4'h6;
    end
    if (reset) begin
      image_1659 <= 4'h0;
    end else begin
      image_1659 <= 4'h6;
    end
    if (reset) begin
      image_1660 <= 4'h0;
    end else begin
      image_1660 <= 4'h3;
    end
    if (reset) begin
      image_1664 <= 4'h0;
    end else begin
      image_1664 <= 4'h2;
    end
    if (reset) begin
      image_1665 <= 4'h0;
    end else begin
      image_1665 <= 4'h5;
    end
    if (reset) begin
      image_1666 <= 4'h0;
    end else begin
      image_1666 <= 4'h5;
    end
    if (reset) begin
      image_1667 <= 4'h0;
    end else begin
      image_1667 <= 4'h5;
    end
    if (reset) begin
      image_1668 <= 4'h0;
    end else begin
      image_1668 <= 4'h5;
    end
    if (reset) begin
      image_1669 <= 4'h0;
    end else begin
      image_1669 <= 4'h6;
    end
    if (reset) begin
      image_1670 <= 4'h0;
    end else begin
      image_1670 <= 4'h6;
    end
    if (reset) begin
      image_1671 <= 4'h0;
    end else begin
      image_1671 <= 4'h6;
    end
    if (reset) begin
      image_1672 <= 4'h0;
    end else begin
      image_1672 <= 4'h6;
    end
    if (reset) begin
      image_1673 <= 4'h0;
    end else begin
      image_1673 <= 4'h6;
    end
    if (reset) begin
      image_1674 <= 4'h0;
    end else begin
      image_1674 <= 4'h6;
    end
    if (reset) begin
      image_1675 <= 4'h0;
    end else begin
      image_1675 <= 4'h6;
    end
    if (reset) begin
      image_1676 <= 4'h0;
    end else begin
      image_1676 <= 4'h6;
    end
    if (reset) begin
      image_1677 <= 4'h0;
    end else begin
      image_1677 <= 4'h6;
    end
    if (reset) begin
      image_1678 <= 4'h0;
    end else begin
      image_1678 <= 4'h6;
    end
    if (reset) begin
      image_1679 <= 4'h0;
    end else begin
      image_1679 <= 4'h6;
    end
    if (reset) begin
      image_1680 <= 4'h0;
    end else begin
      image_1680 <= 4'h6;
    end
    if (reset) begin
      image_1681 <= 4'h0;
    end else begin
      image_1681 <= 4'h6;
    end
    if (reset) begin
      image_1682 <= 4'h0;
    end else begin
      image_1682 <= 4'h6;
    end
    if (reset) begin
      image_1683 <= 4'h0;
    end else begin
      image_1683 <= 4'h6;
    end
    if (reset) begin
      image_1684 <= 4'h0;
    end else begin
      image_1684 <= 4'h6;
    end
    if (reset) begin
      image_1685 <= 4'h0;
    end else begin
      image_1685 <= 4'h6;
    end
    if (reset) begin
      image_1686 <= 4'h0;
    end else begin
      image_1686 <= 4'h6;
    end
    if (reset) begin
      image_1687 <= 4'h0;
    end else begin
      image_1687 <= 4'h5;
    end
    if (reset) begin
      image_1688 <= 4'h0;
    end else begin
      image_1688 <= 4'h4;
    end
    if (reset) begin
      image_1689 <= 4'h0;
    end else begin
      image_1689 <= 4'h4;
    end
    if (reset) begin
      image_1690 <= 4'h0;
    end else begin
      image_1690 <= 4'h5;
    end
    if (reset) begin
      image_1691 <= 4'h0;
    end else begin
      image_1691 <= 4'h6;
    end
    if (reset) begin
      image_1692 <= 4'h0;
    end else begin
      image_1692 <= 4'h6;
    end
    if (reset) begin
      image_1693 <= 4'h0;
    end else begin
      image_1693 <= 4'h6;
    end
    if (reset) begin
      image_1694 <= 4'h0;
    end else begin
      image_1694 <= 4'h6;
    end
    if (reset) begin
      image_1695 <= 4'h0;
    end else begin
      image_1695 <= 4'h6;
    end
    if (reset) begin
      image_1696 <= 4'h0;
    end else begin
      image_1696 <= 4'h6;
    end
    if (reset) begin
      image_1697 <= 4'h0;
    end else begin
      image_1697 <= 4'h5;
    end
    if (reset) begin
      image_1698 <= 4'h0;
    end else begin
      image_1698 <= 4'h4;
    end
    if (reset) begin
      image_1699 <= 4'h0;
    end else begin
      image_1699 <= 4'h3;
    end
    if (reset) begin
      image_1700 <= 4'h0;
    end else begin
      image_1700 <= 4'h3;
    end
    if (reset) begin
      image_1701 <= 4'h0;
    end else begin
      image_1701 <= 4'h3;
    end
    if (reset) begin
      image_1702 <= 4'h0;
    end else begin
      image_1702 <= 4'h3;
    end
    if (reset) begin
      image_1703 <= 4'h0;
    end else begin
      image_1703 <= 4'h5;
    end
    if (reset) begin
      image_1704 <= 4'h0;
    end else begin
      image_1704 <= 4'h5;
    end
    if (reset) begin
      image_1705 <= 4'h0;
    end else begin
      image_1705 <= 4'h5;
    end
    if (reset) begin
      image_1706 <= 4'h0;
    end else begin
      image_1706 <= 4'h5;
    end
    if (reset) begin
      image_1707 <= 4'h0;
    end else begin
      image_1707 <= 4'h5;
    end
    if (reset) begin
      image_1708 <= 4'h0;
    end else begin
      image_1708 <= 4'h5;
    end
    if (reset) begin
      image_1709 <= 4'h0;
    end else begin
      image_1709 <= 4'h5;
    end
    if (reset) begin
      image_1710 <= 4'h0;
    end else begin
      image_1710 <= 4'h5;
    end
    if (reset) begin
      image_1711 <= 4'h0;
    end else begin
      image_1711 <= 4'h5;
    end
    if (reset) begin
      image_1712 <= 4'h0;
    end else begin
      image_1712 <= 4'h5;
    end
    if (reset) begin
      image_1713 <= 4'h0;
    end else begin
      image_1713 <= 4'h5;
    end
    if (reset) begin
      image_1714 <= 4'h0;
    end else begin
      image_1714 <= 4'h6;
    end
    if (reset) begin
      image_1715 <= 4'h0;
    end else begin
      image_1715 <= 4'h6;
    end
    if (reset) begin
      image_1716 <= 4'h0;
    end else begin
      image_1716 <= 4'h6;
    end
    if (reset) begin
      image_1717 <= 4'h0;
    end else begin
      image_1717 <= 4'h6;
    end
    if (reset) begin
      image_1718 <= 4'h0;
    end else begin
      image_1718 <= 4'h6;
    end
    if (reset) begin
      image_1719 <= 4'h0;
    end else begin
      image_1719 <= 4'h6;
    end
    if (reset) begin
      image_1720 <= 4'h0;
    end else begin
      image_1720 <= 4'h4;
    end
    if (reset) begin
      image_1721 <= 4'h0;
    end else begin
      image_1721 <= 4'h6;
    end
    if (reset) begin
      image_1722 <= 4'h0;
    end else begin
      image_1722 <= 4'h5;
    end
    if (reset) begin
      image_1723 <= 4'h0;
    end else begin
      image_1723 <= 4'h2;
    end
    if (reset) begin
      image_1728 <= 4'h0;
    end else begin
      image_1728 <= 4'h1;
    end
    if (reset) begin
      image_1729 <= 4'h0;
    end else begin
      image_1729 <= 4'h5;
    end
    if (reset) begin
      image_1730 <= 4'h0;
    end else begin
      image_1730 <= 4'h5;
    end
    if (reset) begin
      image_1731 <= 4'h0;
    end else begin
      image_1731 <= 4'h5;
    end
    if (reset) begin
      image_1732 <= 4'h0;
    end else begin
      image_1732 <= 4'h5;
    end
    if (reset) begin
      image_1733 <= 4'h0;
    end else begin
      image_1733 <= 4'h6;
    end
    if (reset) begin
      image_1734 <= 4'h0;
    end else begin
      image_1734 <= 4'h6;
    end
    if (reset) begin
      image_1735 <= 4'h0;
    end else begin
      image_1735 <= 4'h6;
    end
    if (reset) begin
      image_1736 <= 4'h0;
    end else begin
      image_1736 <= 4'h6;
    end
    if (reset) begin
      image_1737 <= 4'h0;
    end else begin
      image_1737 <= 4'h6;
    end
    if (reset) begin
      image_1738 <= 4'h0;
    end else begin
      image_1738 <= 4'h6;
    end
    if (reset) begin
      image_1739 <= 4'h0;
    end else begin
      image_1739 <= 4'h6;
    end
    if (reset) begin
      image_1740 <= 4'h0;
    end else begin
      image_1740 <= 4'h6;
    end
    if (reset) begin
      image_1741 <= 4'h0;
    end else begin
      image_1741 <= 4'h6;
    end
    if (reset) begin
      image_1742 <= 4'h0;
    end else begin
      image_1742 <= 4'h6;
    end
    if (reset) begin
      image_1743 <= 4'h0;
    end else begin
      image_1743 <= 4'h6;
    end
    if (reset) begin
      image_1744 <= 4'h0;
    end else begin
      image_1744 <= 4'h6;
    end
    if (reset) begin
      image_1745 <= 4'h0;
    end else begin
      image_1745 <= 4'h6;
    end
    if (reset) begin
      image_1746 <= 4'h0;
    end else begin
      image_1746 <= 4'h6;
    end
    if (reset) begin
      image_1747 <= 4'h0;
    end else begin
      image_1747 <= 4'h6;
    end
    if (reset) begin
      image_1748 <= 4'h0;
    end else begin
      image_1748 <= 4'h6;
    end
    if (reset) begin
      image_1749 <= 4'h0;
    end else begin
      image_1749 <= 4'h5;
    end
    if (reset) begin
      image_1750 <= 4'h0;
    end else begin
      image_1750 <= 4'h3;
    end
    if (reset) begin
      image_1751 <= 4'h0;
    end else begin
      image_1751 <= 4'h5;
    end
    if (reset) begin
      image_1752 <= 4'h0;
    end else begin
      image_1752 <= 4'h6;
    end
    if (reset) begin
      image_1753 <= 4'h0;
    end else begin
      image_1753 <= 4'h6;
    end
    if (reset) begin
      image_1754 <= 4'h0;
    end else begin
      image_1754 <= 4'h6;
    end
    if (reset) begin
      image_1755 <= 4'h0;
    end else begin
      image_1755 <= 4'h6;
    end
    if (reset) begin
      image_1756 <= 4'h0;
    end else begin
      image_1756 <= 4'h6;
    end
    if (reset) begin
      image_1757 <= 4'h0;
    end else begin
      image_1757 <= 4'h5;
    end
    if (reset) begin
      image_1758 <= 4'h0;
    end else begin
      image_1758 <= 4'h4;
    end
    if (reset) begin
      image_1759 <= 4'h0;
    end else begin
      image_1759 <= 4'h3;
    end
    if (reset) begin
      image_1760 <= 4'h0;
    end else begin
      image_1760 <= 4'h3;
    end
    if (reset) begin
      image_1761 <= 4'h0;
    end else begin
      image_1761 <= 4'h3;
    end
    if (reset) begin
      image_1762 <= 4'h0;
    end else begin
      image_1762 <= 4'h4;
    end
    if (reset) begin
      image_1763 <= 4'h0;
    end else begin
      image_1763 <= 4'h4;
    end
    if (reset) begin
      image_1764 <= 4'h0;
    end else begin
      image_1764 <= 4'h4;
    end
    if (reset) begin
      image_1765 <= 4'h0;
    end else begin
      image_1765 <= 4'h4;
    end
    if (reset) begin
      image_1766 <= 4'h0;
    end else begin
      image_1766 <= 4'h4;
    end
    if (reset) begin
      image_1767 <= 4'h0;
    end else begin
      image_1767 <= 4'h4;
    end
    if (reset) begin
      image_1768 <= 4'h0;
    end else begin
      image_1768 <= 4'h5;
    end
    if (reset) begin
      image_1769 <= 4'h0;
    end else begin
      image_1769 <= 4'h5;
    end
    if (reset) begin
      image_1770 <= 4'h0;
    end else begin
      image_1770 <= 4'h5;
    end
    if (reset) begin
      image_1771 <= 4'h0;
    end else begin
      image_1771 <= 4'h5;
    end
    if (reset) begin
      image_1772 <= 4'h0;
    end else begin
      image_1772 <= 4'h5;
    end
    if (reset) begin
      image_1773 <= 4'h0;
    end else begin
      image_1773 <= 4'h5;
    end
    if (reset) begin
      image_1774 <= 4'h0;
    end else begin
      image_1774 <= 4'h5;
    end
    if (reset) begin
      image_1775 <= 4'h0;
    end else begin
      image_1775 <= 4'h5;
    end
    if (reset) begin
      image_1776 <= 4'h0;
    end else begin
      image_1776 <= 4'h5;
    end
    if (reset) begin
      image_1777 <= 4'h0;
    end else begin
      image_1777 <= 4'h5;
    end
    if (reset) begin
      image_1778 <= 4'h0;
    end else begin
      image_1778 <= 4'h5;
    end
    if (reset) begin
      image_1779 <= 4'h0;
    end else begin
      image_1779 <= 4'h6;
    end
    if (reset) begin
      image_1780 <= 4'h0;
    end else begin
      image_1780 <= 4'h6;
    end
    if (reset) begin
      image_1781 <= 4'h0;
    end else begin
      image_1781 <= 4'h6;
    end
    if (reset) begin
      image_1782 <= 4'h0;
    end else begin
      image_1782 <= 4'h6;
    end
    if (reset) begin
      image_1783 <= 4'h0;
    end else begin
      image_1783 <= 4'h3;
    end
    if (reset) begin
      image_1784 <= 4'h0;
    end else begin
      image_1784 <= 4'h6;
    end
    if (reset) begin
      image_1785 <= 4'h0;
    end else begin
      image_1785 <= 4'h6;
    end
    if (reset) begin
      image_1786 <= 4'h0;
    end else begin
      image_1786 <= 4'h3;
    end
    if (reset) begin
      image_1793 <= 4'h0;
    end else begin
      image_1793 <= 4'h5;
    end
    if (reset) begin
      image_1794 <= 4'h0;
    end else begin
      image_1794 <= 4'h5;
    end
    if (reset) begin
      image_1795 <= 4'h0;
    end else begin
      image_1795 <= 4'h5;
    end
    if (reset) begin
      image_1796 <= 4'h0;
    end else begin
      image_1796 <= 4'h5;
    end
    if (reset) begin
      image_1797 <= 4'h0;
    end else begin
      image_1797 <= 4'h6;
    end
    if (reset) begin
      image_1798 <= 4'h0;
    end else begin
      image_1798 <= 4'h6;
    end
    if (reset) begin
      image_1799 <= 4'h0;
    end else begin
      image_1799 <= 4'h6;
    end
    if (reset) begin
      image_1800 <= 4'h0;
    end else begin
      image_1800 <= 4'h6;
    end
    if (reset) begin
      image_1801 <= 4'h0;
    end else begin
      image_1801 <= 4'h6;
    end
    if (reset) begin
      image_1802 <= 4'h0;
    end else begin
      image_1802 <= 4'h6;
    end
    if (reset) begin
      image_1803 <= 4'h0;
    end else begin
      image_1803 <= 4'h6;
    end
    if (reset) begin
      image_1804 <= 4'h0;
    end else begin
      image_1804 <= 4'h6;
    end
    if (reset) begin
      image_1805 <= 4'h0;
    end else begin
      image_1805 <= 4'h6;
    end
    if (reset) begin
      image_1806 <= 4'h0;
    end else begin
      image_1806 <= 4'h6;
    end
    if (reset) begin
      image_1807 <= 4'h0;
    end else begin
      image_1807 <= 4'h6;
    end
    if (reset) begin
      image_1808 <= 4'h0;
    end else begin
      image_1808 <= 4'h6;
    end
    if (reset) begin
      image_1809 <= 4'h0;
    end else begin
      image_1809 <= 4'h6;
    end
    if (reset) begin
      image_1810 <= 4'h0;
    end else begin
      image_1810 <= 4'h6;
    end
    if (reset) begin
      image_1811 <= 4'h0;
    end else begin
      image_1811 <= 4'h6;
    end
    if (reset) begin
      image_1812 <= 4'h0;
    end else begin
      image_1812 <= 4'h6;
    end
    if (reset) begin
      image_1813 <= 4'h0;
    end else begin
      image_1813 <= 4'h3;
    end
    if (reset) begin
      image_1814 <= 4'h0;
    end else begin
      image_1814 <= 4'h5;
    end
    if (reset) begin
      image_1815 <= 4'h0;
    end else begin
      image_1815 <= 4'h6;
    end
    if (reset) begin
      image_1816 <= 4'h0;
    end else begin
      image_1816 <= 4'h6;
    end
    if (reset) begin
      image_1817 <= 4'h0;
    end else begin
      image_1817 <= 4'h6;
    end
    if (reset) begin
      image_1818 <= 4'h0;
    end else begin
      image_1818 <= 4'h5;
    end
    if (reset) begin
      image_1819 <= 4'h0;
    end else begin
      image_1819 <= 4'h3;
    end
    if (reset) begin
      image_1820 <= 4'h0;
    end else begin
      image_1820 <= 4'h2;
    end
    if (reset) begin
      image_1821 <= 4'h0;
    end else begin
      image_1821 <= 4'h3;
    end
    if (reset) begin
      image_1822 <= 4'h0;
    end else begin
      image_1822 <= 4'h3;
    end
    if (reset) begin
      image_1823 <= 4'h0;
    end else begin
      image_1823 <= 4'h3;
    end
    if (reset) begin
      image_1824 <= 4'h0;
    end else begin
      image_1824 <= 4'h4;
    end
    if (reset) begin
      image_1825 <= 4'h0;
    end else begin
      image_1825 <= 4'h4;
    end
    if (reset) begin
      image_1826 <= 4'h0;
    end else begin
      image_1826 <= 4'h4;
    end
    if (reset) begin
      image_1827 <= 4'h0;
    end else begin
      image_1827 <= 4'h4;
    end
    if (reset) begin
      image_1828 <= 4'h0;
    end else begin
      image_1828 <= 4'h4;
    end
    if (reset) begin
      image_1829 <= 4'h0;
    end else begin
      image_1829 <= 4'h4;
    end
    if (reset) begin
      image_1830 <= 4'h0;
    end else begin
      image_1830 <= 4'h4;
    end
    if (reset) begin
      image_1831 <= 4'h0;
    end else begin
      image_1831 <= 4'h4;
    end
    if (reset) begin
      image_1832 <= 4'h0;
    end else begin
      image_1832 <= 4'h5;
    end
    if (reset) begin
      image_1833 <= 4'h0;
    end else begin
      image_1833 <= 4'h5;
    end
    if (reset) begin
      image_1834 <= 4'h0;
    end else begin
      image_1834 <= 4'h5;
    end
    if (reset) begin
      image_1835 <= 4'h0;
    end else begin
      image_1835 <= 4'h5;
    end
    if (reset) begin
      image_1836 <= 4'h0;
    end else begin
      image_1836 <= 4'h5;
    end
    if (reset) begin
      image_1837 <= 4'h0;
    end else begin
      image_1837 <= 4'h5;
    end
    if (reset) begin
      image_1838 <= 4'h0;
    end else begin
      image_1838 <= 4'h5;
    end
    if (reset) begin
      image_1839 <= 4'h0;
    end else begin
      image_1839 <= 4'h5;
    end
    if (reset) begin
      image_1840 <= 4'h0;
    end else begin
      image_1840 <= 4'h5;
    end
    if (reset) begin
      image_1841 <= 4'h0;
    end else begin
      image_1841 <= 4'h5;
    end
    if (reset) begin
      image_1842 <= 4'h0;
    end else begin
      image_1842 <= 4'h5;
    end
    if (reset) begin
      image_1843 <= 4'h0;
    end else begin
      image_1843 <= 4'h6;
    end
    if (reset) begin
      image_1844 <= 4'h0;
    end else begin
      image_1844 <= 4'h6;
    end
    if (reset) begin
      image_1845 <= 4'h0;
    end else begin
      image_1845 <= 4'h6;
    end
    if (reset) begin
      image_1846 <= 4'h0;
    end else begin
      image_1846 <= 4'h5;
    end
    if (reset) begin
      image_1847 <= 4'h0;
    end else begin
      image_1847 <= 4'h5;
    end
    if (reset) begin
      image_1848 <= 4'h0;
    end else begin
      image_1848 <= 4'h6;
    end
    if (reset) begin
      image_1849 <= 4'h0;
    end else begin
      image_1849 <= 4'h6;
    end
    if (reset) begin
      image_1857 <= 4'h0;
    end else begin
      image_1857 <= 4'h4;
    end
    if (reset) begin
      image_1858 <= 4'h0;
    end else begin
      image_1858 <= 4'h5;
    end
    if (reset) begin
      image_1859 <= 4'h0;
    end else begin
      image_1859 <= 4'h5;
    end
    if (reset) begin
      image_1860 <= 4'h0;
    end else begin
      image_1860 <= 4'h5;
    end
    if (reset) begin
      image_1861 <= 4'h0;
    end else begin
      image_1861 <= 4'h6;
    end
    if (reset) begin
      image_1862 <= 4'h0;
    end else begin
      image_1862 <= 4'h6;
    end
    if (reset) begin
      image_1863 <= 4'h0;
    end else begin
      image_1863 <= 4'h6;
    end
    if (reset) begin
      image_1864 <= 4'h0;
    end else begin
      image_1864 <= 4'h6;
    end
    if (reset) begin
      image_1865 <= 4'h0;
    end else begin
      image_1865 <= 4'h6;
    end
    if (reset) begin
      image_1866 <= 4'h0;
    end else begin
      image_1866 <= 4'h6;
    end
    if (reset) begin
      image_1867 <= 4'h0;
    end else begin
      image_1867 <= 4'h6;
    end
    if (reset) begin
      image_1868 <= 4'h0;
    end else begin
      image_1868 <= 4'h6;
    end
    if (reset) begin
      image_1869 <= 4'h0;
    end else begin
      image_1869 <= 4'h6;
    end
    if (reset) begin
      image_1870 <= 4'h0;
    end else begin
      image_1870 <= 4'h6;
    end
    if (reset) begin
      image_1871 <= 4'h0;
    end else begin
      image_1871 <= 4'h6;
    end
    if (reset) begin
      image_1872 <= 4'h0;
    end else begin
      image_1872 <= 4'h6;
    end
    if (reset) begin
      image_1873 <= 4'h0;
    end else begin
      image_1873 <= 4'h6;
    end
    if (reset) begin
      image_1874 <= 4'h0;
    end else begin
      image_1874 <= 4'h6;
    end
    if (reset) begin
      image_1875 <= 4'h0;
    end else begin
      image_1875 <= 4'h6;
    end
    if (reset) begin
      image_1876 <= 4'h0;
    end else begin
      image_1876 <= 4'h6;
    end
    if (reset) begin
      image_1877 <= 4'h0;
    end else begin
      image_1877 <= 4'h4;
    end
    if (reset) begin
      image_1878 <= 4'h0;
    end else begin
      image_1878 <= 4'h5;
    end
    if (reset) begin
      image_1879 <= 4'h0;
    end else begin
      image_1879 <= 4'h6;
    end
    if (reset) begin
      image_1880 <= 4'h0;
    end else begin
      image_1880 <= 4'h6;
    end
    if (reset) begin
      image_1881 <= 4'h0;
    end else begin
      image_1881 <= 4'h3;
    end
    if (reset) begin
      image_1882 <= 4'h0;
    end else begin
      image_1882 <= 4'h3;
    end
    if (reset) begin
      image_1883 <= 4'h0;
    end else begin
      image_1883 <= 4'h3;
    end
    if (reset) begin
      image_1884 <= 4'h0;
    end else begin
      image_1884 <= 4'h3;
    end
    if (reset) begin
      image_1885 <= 4'h0;
    end else begin
      image_1885 <= 4'h3;
    end
    if (reset) begin
      image_1886 <= 4'h0;
    end else begin
      image_1886 <= 4'h3;
    end
    if (reset) begin
      image_1887 <= 4'h0;
    end else begin
      image_1887 <= 4'h3;
    end
    if (reset) begin
      image_1888 <= 4'h0;
    end else begin
      image_1888 <= 4'h4;
    end
    if (reset) begin
      image_1889 <= 4'h0;
    end else begin
      image_1889 <= 4'h4;
    end
    if (reset) begin
      image_1890 <= 4'h0;
    end else begin
      image_1890 <= 4'h4;
    end
    if (reset) begin
      image_1891 <= 4'h0;
    end else begin
      image_1891 <= 4'h4;
    end
    if (reset) begin
      image_1892 <= 4'h0;
    end else begin
      image_1892 <= 4'h4;
    end
    if (reset) begin
      image_1893 <= 4'h0;
    end else begin
      image_1893 <= 4'h4;
    end
    if (reset) begin
      image_1894 <= 4'h0;
    end else begin
      image_1894 <= 4'h4;
    end
    if (reset) begin
      image_1895 <= 4'h0;
    end else begin
      image_1895 <= 4'h4;
    end
    if (reset) begin
      image_1896 <= 4'h0;
    end else begin
      image_1896 <= 4'h5;
    end
    if (reset) begin
      image_1897 <= 4'h0;
    end else begin
      image_1897 <= 4'h5;
    end
    if (reset) begin
      image_1898 <= 4'h0;
    end else begin
      image_1898 <= 4'h5;
    end
    if (reset) begin
      image_1899 <= 4'h0;
    end else begin
      image_1899 <= 4'h5;
    end
    if (reset) begin
      image_1900 <= 4'h0;
    end else begin
      image_1900 <= 4'h5;
    end
    if (reset) begin
      image_1901 <= 4'h0;
    end else begin
      image_1901 <= 4'h5;
    end
    if (reset) begin
      image_1902 <= 4'h0;
    end else begin
      image_1902 <= 4'h5;
    end
    if (reset) begin
      image_1903 <= 4'h0;
    end else begin
      image_1903 <= 4'h5;
    end
    if (reset) begin
      image_1904 <= 4'h0;
    end else begin
      image_1904 <= 4'h5;
    end
    if (reset) begin
      image_1905 <= 4'h0;
    end else begin
      image_1905 <= 4'h5;
    end
    if (reset) begin
      image_1906 <= 4'h0;
    end else begin
      image_1906 <= 4'h5;
    end
    if (reset) begin
      image_1907 <= 4'h0;
    end else begin
      image_1907 <= 4'h6;
    end
    if (reset) begin
      image_1908 <= 4'h0;
    end else begin
      image_1908 <= 4'h6;
    end
    if (reset) begin
      image_1909 <= 4'h0;
    end else begin
      image_1909 <= 4'h6;
    end
    if (reset) begin
      image_1910 <= 4'h0;
    end else begin
      image_1910 <= 4'h5;
    end
    if (reset) begin
      image_1911 <= 4'h0;
    end else begin
      image_1911 <= 4'h5;
    end
    if (reset) begin
      image_1912 <= 4'h0;
    end else begin
      image_1912 <= 4'h6;
    end
    if (reset) begin
      image_1913 <= 4'h0;
    end else begin
      image_1913 <= 4'h6;
    end
    if (reset) begin
      image_1921 <= 4'h0;
    end else begin
      image_1921 <= 4'h4;
    end
    if (reset) begin
      image_1922 <= 4'h0;
    end else begin
      image_1922 <= 4'h5;
    end
    if (reset) begin
      image_1923 <= 4'h0;
    end else begin
      image_1923 <= 4'h5;
    end
    if (reset) begin
      image_1924 <= 4'h0;
    end else begin
      image_1924 <= 4'h5;
    end
    if (reset) begin
      image_1925 <= 4'h0;
    end else begin
      image_1925 <= 4'h5;
    end
    if (reset) begin
      image_1926 <= 4'h0;
    end else begin
      image_1926 <= 4'h6;
    end
    if (reset) begin
      image_1927 <= 4'h0;
    end else begin
      image_1927 <= 4'h6;
    end
    if (reset) begin
      image_1928 <= 4'h0;
    end else begin
      image_1928 <= 4'h6;
    end
    if (reset) begin
      image_1929 <= 4'h0;
    end else begin
      image_1929 <= 4'h6;
    end
    if (reset) begin
      image_1930 <= 4'h0;
    end else begin
      image_1930 <= 4'h6;
    end
    if (reset) begin
      image_1931 <= 4'h0;
    end else begin
      image_1931 <= 4'h6;
    end
    if (reset) begin
      image_1932 <= 4'h0;
    end else begin
      image_1932 <= 4'h6;
    end
    if (reset) begin
      image_1933 <= 4'h0;
    end else begin
      image_1933 <= 4'h6;
    end
    if (reset) begin
      image_1934 <= 4'h0;
    end else begin
      image_1934 <= 4'h6;
    end
    if (reset) begin
      image_1935 <= 4'h0;
    end else begin
      image_1935 <= 4'h6;
    end
    if (reset) begin
      image_1936 <= 4'h0;
    end else begin
      image_1936 <= 4'h6;
    end
    if (reset) begin
      image_1937 <= 4'h0;
    end else begin
      image_1937 <= 4'h6;
    end
    if (reset) begin
      image_1938 <= 4'h0;
    end else begin
      image_1938 <= 4'h6;
    end
    if (reset) begin
      image_1939 <= 4'h0;
    end else begin
      image_1939 <= 4'h6;
    end
    if (reset) begin
      image_1940 <= 4'h0;
    end else begin
      image_1940 <= 4'h6;
    end
    if (reset) begin
      image_1941 <= 4'h0;
    end else begin
      image_1941 <= 4'h5;
    end
    if (reset) begin
      image_1942 <= 4'h0;
    end else begin
      image_1942 <= 4'h5;
    end
    if (reset) begin
      image_1943 <= 4'h0;
    end else begin
      image_1943 <= 4'h6;
    end
    if (reset) begin
      image_1944 <= 4'h0;
    end else begin
      image_1944 <= 4'h4;
    end
    if (reset) begin
      image_1945 <= 4'h0;
    end else begin
      image_1945 <= 4'h3;
    end
    if (reset) begin
      image_1946 <= 4'h0;
    end else begin
      image_1946 <= 4'h3;
    end
    if (reset) begin
      image_1947 <= 4'h0;
    end else begin
      image_1947 <= 4'h3;
    end
    if (reset) begin
      image_1948 <= 4'h0;
    end else begin
      image_1948 <= 4'h3;
    end
    if (reset) begin
      image_1949 <= 4'h0;
    end else begin
      image_1949 <= 4'h3;
    end
    if (reset) begin
      image_1950 <= 4'h0;
    end else begin
      image_1950 <= 4'h3;
    end
    if (reset) begin
      image_1951 <= 4'h0;
    end else begin
      image_1951 <= 4'h4;
    end
    if (reset) begin
      image_1952 <= 4'h0;
    end else begin
      image_1952 <= 4'h4;
    end
    if (reset) begin
      image_1953 <= 4'h0;
    end else begin
      image_1953 <= 4'h4;
    end
    if (reset) begin
      image_1954 <= 4'h0;
    end else begin
      image_1954 <= 4'h4;
    end
    if (reset) begin
      image_1955 <= 4'h0;
    end else begin
      image_1955 <= 4'h4;
    end
    if (reset) begin
      image_1956 <= 4'h0;
    end else begin
      image_1956 <= 4'h4;
    end
    if (reset) begin
      image_1957 <= 4'h0;
    end else begin
      image_1957 <= 4'h4;
    end
    if (reset) begin
      image_1958 <= 4'h0;
    end else begin
      image_1958 <= 4'h4;
    end
    if (reset) begin
      image_1959 <= 4'h0;
    end else begin
      image_1959 <= 4'h5;
    end
    if (reset) begin
      image_1960 <= 4'h0;
    end else begin
      image_1960 <= 4'h5;
    end
    if (reset) begin
      image_1961 <= 4'h0;
    end else begin
      image_1961 <= 4'h5;
    end
    if (reset) begin
      image_1962 <= 4'h0;
    end else begin
      image_1962 <= 4'h5;
    end
    if (reset) begin
      image_1963 <= 4'h0;
    end else begin
      image_1963 <= 4'h5;
    end
    if (reset) begin
      image_1964 <= 4'h0;
    end else begin
      image_1964 <= 4'h5;
    end
    if (reset) begin
      image_1965 <= 4'h0;
    end else begin
      image_1965 <= 4'h5;
    end
    if (reset) begin
      image_1966 <= 4'h0;
    end else begin
      image_1966 <= 4'h5;
    end
    if (reset) begin
      image_1967 <= 4'h0;
    end else begin
      image_1967 <= 4'h5;
    end
    if (reset) begin
      image_1968 <= 4'h0;
    end else begin
      image_1968 <= 4'h5;
    end
    if (reset) begin
      image_1969 <= 4'h0;
    end else begin
      image_1969 <= 4'h5;
    end
    if (reset) begin
      image_1970 <= 4'h0;
    end else begin
      image_1970 <= 4'h6;
    end
    if (reset) begin
      image_1971 <= 4'h0;
    end else begin
      image_1971 <= 4'h6;
    end
    if (reset) begin
      image_1972 <= 4'h0;
    end else begin
      image_1972 <= 4'h6;
    end
    if (reset) begin
      image_1973 <= 4'h0;
    end else begin
      image_1973 <= 4'h6;
    end
    if (reset) begin
      image_1974 <= 4'h0;
    end else begin
      image_1974 <= 4'h5;
    end
    if (reset) begin
      image_1975 <= 4'h0;
    end else begin
      image_1975 <= 4'h5;
    end
    if (reset) begin
      image_1976 <= 4'h0;
    end else begin
      image_1976 <= 4'h6;
    end
    if (reset) begin
      image_1977 <= 4'h0;
    end else begin
      image_1977 <= 4'h6;
    end
    if (reset) begin
      image_1985 <= 4'h0;
    end else begin
      image_1985 <= 4'h3;
    end
    if (reset) begin
      image_1986 <= 4'h0;
    end else begin
      image_1986 <= 4'h5;
    end
    if (reset) begin
      image_1987 <= 4'h0;
    end else begin
      image_1987 <= 4'h5;
    end
    if (reset) begin
      image_1988 <= 4'h0;
    end else begin
      image_1988 <= 4'h5;
    end
    if (reset) begin
      image_1989 <= 4'h0;
    end else begin
      image_1989 <= 4'h5;
    end
    if (reset) begin
      image_1990 <= 4'h0;
    end else begin
      image_1990 <= 4'h6;
    end
    if (reset) begin
      image_1991 <= 4'h0;
    end else begin
      image_1991 <= 4'h6;
    end
    if (reset) begin
      image_1992 <= 4'h0;
    end else begin
      image_1992 <= 4'h6;
    end
    if (reset) begin
      image_1993 <= 4'h0;
    end else begin
      image_1993 <= 4'h6;
    end
    if (reset) begin
      image_1994 <= 4'h0;
    end else begin
      image_1994 <= 4'h6;
    end
    if (reset) begin
      image_1995 <= 4'h0;
    end else begin
      image_1995 <= 4'h6;
    end
    if (reset) begin
      image_1996 <= 4'h0;
    end else begin
      image_1996 <= 4'h6;
    end
    if (reset) begin
      image_1997 <= 4'h0;
    end else begin
      image_1997 <= 4'h6;
    end
    if (reset) begin
      image_1998 <= 4'h0;
    end else begin
      image_1998 <= 4'h6;
    end
    if (reset) begin
      image_1999 <= 4'h0;
    end else begin
      image_1999 <= 4'h6;
    end
    if (reset) begin
      image_2000 <= 4'h0;
    end else begin
      image_2000 <= 4'h6;
    end
    if (reset) begin
      image_2001 <= 4'h0;
    end else begin
      image_2001 <= 4'h6;
    end
    if (reset) begin
      image_2002 <= 4'h0;
    end else begin
      image_2002 <= 4'h6;
    end
    if (reset) begin
      image_2003 <= 4'h0;
    end else begin
      image_2003 <= 4'h6;
    end
    if (reset) begin
      image_2004 <= 4'h0;
    end else begin
      image_2004 <= 4'h6;
    end
    if (reset) begin
      image_2005 <= 4'h0;
    end else begin
      image_2005 <= 4'h5;
    end
    if (reset) begin
      image_2006 <= 4'h0;
    end else begin
      image_2006 <= 4'h4;
    end
    if (reset) begin
      image_2007 <= 4'h0;
    end else begin
      image_2007 <= 4'h6;
    end
    if (reset) begin
      image_2008 <= 4'h0;
    end else begin
      image_2008 <= 4'h2;
    end
    if (reset) begin
      image_2009 <= 4'h0;
    end else begin
      image_2009 <= 4'h3;
    end
    if (reset) begin
      image_2010 <= 4'h0;
    end else begin
      image_2010 <= 4'h3;
    end
    if (reset) begin
      image_2011 <= 4'h0;
    end else begin
      image_2011 <= 4'h3;
    end
    if (reset) begin
      image_2012 <= 4'h0;
    end else begin
      image_2012 <= 4'h3;
    end
    if (reset) begin
      image_2013 <= 4'h0;
    end else begin
      image_2013 <= 4'h3;
    end
    if (reset) begin
      image_2014 <= 4'h0;
    end else begin
      image_2014 <= 4'h3;
    end
    if (reset) begin
      image_2015 <= 4'h0;
    end else begin
      image_2015 <= 4'h4;
    end
    if (reset) begin
      image_2016 <= 4'h0;
    end else begin
      image_2016 <= 4'h4;
    end
    if (reset) begin
      image_2017 <= 4'h0;
    end else begin
      image_2017 <= 4'h4;
    end
    if (reset) begin
      image_2018 <= 4'h0;
    end else begin
      image_2018 <= 4'h4;
    end
    if (reset) begin
      image_2019 <= 4'h0;
    end else begin
      image_2019 <= 4'h4;
    end
    if (reset) begin
      image_2020 <= 4'h0;
    end else begin
      image_2020 <= 4'h4;
    end
    if (reset) begin
      image_2021 <= 4'h0;
    end else begin
      image_2021 <= 4'h4;
    end
    if (reset) begin
      image_2022 <= 4'h0;
    end else begin
      image_2022 <= 4'h4;
    end
    if (reset) begin
      image_2023 <= 4'h0;
    end else begin
      image_2023 <= 4'h5;
    end
    if (reset) begin
      image_2024 <= 4'h0;
    end else begin
      image_2024 <= 4'h5;
    end
    if (reset) begin
      image_2025 <= 4'h0;
    end else begin
      image_2025 <= 4'h5;
    end
    if (reset) begin
      image_2026 <= 4'h0;
    end else begin
      image_2026 <= 4'h5;
    end
    if (reset) begin
      image_2027 <= 4'h0;
    end else begin
      image_2027 <= 4'h5;
    end
    if (reset) begin
      image_2028 <= 4'h0;
    end else begin
      image_2028 <= 4'h5;
    end
    if (reset) begin
      image_2029 <= 4'h0;
    end else begin
      image_2029 <= 4'h5;
    end
    if (reset) begin
      image_2030 <= 4'h0;
    end else begin
      image_2030 <= 4'h5;
    end
    if (reset) begin
      image_2031 <= 4'h0;
    end else begin
      image_2031 <= 4'h5;
    end
    if (reset) begin
      image_2032 <= 4'h0;
    end else begin
      image_2032 <= 4'h5;
    end
    if (reset) begin
      image_2033 <= 4'h0;
    end else begin
      image_2033 <= 4'h5;
    end
    if (reset) begin
      image_2034 <= 4'h0;
    end else begin
      image_2034 <= 4'h6;
    end
    if (reset) begin
      image_2035 <= 4'h0;
    end else begin
      image_2035 <= 4'h6;
    end
    if (reset) begin
      image_2036 <= 4'h0;
    end else begin
      image_2036 <= 4'h6;
    end
    if (reset) begin
      image_2037 <= 4'h0;
    end else begin
      image_2037 <= 4'h6;
    end
    if (reset) begin
      image_2038 <= 4'h0;
    end else begin
      image_2038 <= 4'h5;
    end
    if (reset) begin
      image_2039 <= 4'h0;
    end else begin
      image_2039 <= 4'h5;
    end
    if (reset) begin
      image_2040 <= 4'h0;
    end else begin
      image_2040 <= 4'h6;
    end
    if (reset) begin
      image_2041 <= 4'h0;
    end else begin
      image_2041 <= 4'h6;
    end
    if (reset) begin
      image_2049 <= 4'h0;
    end else begin
      image_2049 <= 4'h2;
    end
    if (reset) begin
      image_2050 <= 4'h0;
    end else begin
      image_2050 <= 4'h5;
    end
    if (reset) begin
      image_2051 <= 4'h0;
    end else begin
      image_2051 <= 4'h5;
    end
    if (reset) begin
      image_2052 <= 4'h0;
    end else begin
      image_2052 <= 4'h5;
    end
    if (reset) begin
      image_2053 <= 4'h0;
    end else begin
      image_2053 <= 4'h5;
    end
    if (reset) begin
      image_2054 <= 4'h0;
    end else begin
      image_2054 <= 4'h5;
    end
    if (reset) begin
      image_2055 <= 4'h0;
    end else begin
      image_2055 <= 4'h6;
    end
    if (reset) begin
      image_2056 <= 4'h0;
    end else begin
      image_2056 <= 4'h6;
    end
    if (reset) begin
      image_2057 <= 4'h0;
    end else begin
      image_2057 <= 4'h6;
    end
    if (reset) begin
      image_2058 <= 4'h0;
    end else begin
      image_2058 <= 4'h6;
    end
    if (reset) begin
      image_2059 <= 4'h0;
    end else begin
      image_2059 <= 4'h6;
    end
    if (reset) begin
      image_2060 <= 4'h0;
    end else begin
      image_2060 <= 4'h6;
    end
    if (reset) begin
      image_2061 <= 4'h0;
    end else begin
      image_2061 <= 4'h6;
    end
    if (reset) begin
      image_2062 <= 4'h0;
    end else begin
      image_2062 <= 4'h6;
    end
    if (reset) begin
      image_2063 <= 4'h0;
    end else begin
      image_2063 <= 4'h6;
    end
    if (reset) begin
      image_2064 <= 4'h0;
    end else begin
      image_2064 <= 4'h6;
    end
    if (reset) begin
      image_2065 <= 4'h0;
    end else begin
      image_2065 <= 4'h6;
    end
    if (reset) begin
      image_2066 <= 4'h0;
    end else begin
      image_2066 <= 4'h6;
    end
    if (reset) begin
      image_2067 <= 4'h0;
    end else begin
      image_2067 <= 4'h6;
    end
    if (reset) begin
      image_2068 <= 4'h0;
    end else begin
      image_2068 <= 4'h6;
    end
    if (reset) begin
      image_2069 <= 4'h0;
    end else begin
      image_2069 <= 4'h6;
    end
    if (reset) begin
      image_2070 <= 4'h0;
    end else begin
      image_2070 <= 4'h3;
    end
    if (reset) begin
      image_2071 <= 4'h0;
    end else begin
      image_2071 <= 4'h6;
    end
    if (reset) begin
      image_2072 <= 4'h0;
    end else begin
      image_2072 <= 4'h5;
    end
    if (reset) begin
      image_2073 <= 4'h0;
    end else begin
      image_2073 <= 4'h2;
    end
    if (reset) begin
      image_2074 <= 4'h0;
    end else begin
      image_2074 <= 4'h3;
    end
    if (reset) begin
      image_2075 <= 4'h0;
    end else begin
      image_2075 <= 4'h3;
    end
    if (reset) begin
      image_2076 <= 4'h0;
    end else begin
      image_2076 <= 4'h3;
    end
    if (reset) begin
      image_2077 <= 4'h0;
    end else begin
      image_2077 <= 4'h3;
    end
    if (reset) begin
      image_2078 <= 4'h0;
    end else begin
      image_2078 <= 4'h4;
    end
    if (reset) begin
      image_2079 <= 4'h0;
    end else begin
      image_2079 <= 4'h4;
    end
    if (reset) begin
      image_2080 <= 4'h0;
    end else begin
      image_2080 <= 4'h4;
    end
    if (reset) begin
      image_2081 <= 4'h0;
    end else begin
      image_2081 <= 4'h4;
    end
    if (reset) begin
      image_2082 <= 4'h0;
    end else begin
      image_2082 <= 4'h4;
    end
    if (reset) begin
      image_2083 <= 4'h0;
    end else begin
      image_2083 <= 4'h4;
    end
    if (reset) begin
      image_2084 <= 4'h0;
    end else begin
      image_2084 <= 4'h4;
    end
    if (reset) begin
      image_2085 <= 4'h0;
    end else begin
      image_2085 <= 4'h4;
    end
    if (reset) begin
      image_2086 <= 4'h0;
    end else begin
      image_2086 <= 4'h5;
    end
    if (reset) begin
      image_2087 <= 4'h0;
    end else begin
      image_2087 <= 4'h5;
    end
    if (reset) begin
      image_2088 <= 4'h0;
    end else begin
      image_2088 <= 4'h5;
    end
    if (reset) begin
      image_2089 <= 4'h0;
    end else begin
      image_2089 <= 4'h5;
    end
    if (reset) begin
      image_2090 <= 4'h0;
    end else begin
      image_2090 <= 4'h5;
    end
    if (reset) begin
      image_2091 <= 4'h0;
    end else begin
      image_2091 <= 4'h5;
    end
    if (reset) begin
      image_2092 <= 4'h0;
    end else begin
      image_2092 <= 4'h5;
    end
    if (reset) begin
      image_2093 <= 4'h0;
    end else begin
      image_2093 <= 4'h5;
    end
    if (reset) begin
      image_2094 <= 4'h0;
    end else begin
      image_2094 <= 4'h5;
    end
    if (reset) begin
      image_2095 <= 4'h0;
    end else begin
      image_2095 <= 4'h5;
    end
    if (reset) begin
      image_2096 <= 4'h0;
    end else begin
      image_2096 <= 4'h5;
    end
    if (reset) begin
      image_2097 <= 4'h0;
    end else begin
      image_2097 <= 4'h6;
    end
    if (reset) begin
      image_2098 <= 4'h0;
    end else begin
      image_2098 <= 4'h6;
    end
    if (reset) begin
      image_2099 <= 4'h0;
    end else begin
      image_2099 <= 4'h6;
    end
    if (reset) begin
      image_2100 <= 4'h0;
    end else begin
      image_2100 <= 4'h6;
    end
    if (reset) begin
      image_2101 <= 4'h0;
    end else begin
      image_2101 <= 4'h6;
    end
    if (reset) begin
      image_2102 <= 4'h0;
    end else begin
      image_2102 <= 4'h5;
    end
    if (reset) begin
      image_2103 <= 4'h0;
    end else begin
      image_2103 <= 4'h5;
    end
    if (reset) begin
      image_2104 <= 4'h0;
    end else begin
      image_2104 <= 4'h6;
    end
    if (reset) begin
      image_2105 <= 4'h0;
    end else begin
      image_2105 <= 4'h6;
    end
    if (reset) begin
      image_2106 <= 4'h0;
    end else begin
      image_2106 <= 4'h1;
    end
    if (reset) begin
      image_2114 <= 4'h0;
    end else begin
      image_2114 <= 4'h4;
    end
    if (reset) begin
      image_2115 <= 4'h0;
    end else begin
      image_2115 <= 4'h5;
    end
    if (reset) begin
      image_2116 <= 4'h0;
    end else begin
      image_2116 <= 4'h5;
    end
    if (reset) begin
      image_2117 <= 4'h0;
    end else begin
      image_2117 <= 4'h5;
    end
    if (reset) begin
      image_2118 <= 4'h0;
    end else begin
      image_2118 <= 4'h5;
    end
    if (reset) begin
      image_2119 <= 4'h0;
    end else begin
      image_2119 <= 4'h6;
    end
    if (reset) begin
      image_2120 <= 4'h0;
    end else begin
      image_2120 <= 4'h6;
    end
    if (reset) begin
      image_2121 <= 4'h0;
    end else begin
      image_2121 <= 4'h6;
    end
    if (reset) begin
      image_2122 <= 4'h0;
    end else begin
      image_2122 <= 4'h6;
    end
    if (reset) begin
      image_2123 <= 4'h0;
    end else begin
      image_2123 <= 4'h6;
    end
    if (reset) begin
      image_2124 <= 4'h0;
    end else begin
      image_2124 <= 4'h6;
    end
    if (reset) begin
      image_2125 <= 4'h0;
    end else begin
      image_2125 <= 4'h6;
    end
    if (reset) begin
      image_2126 <= 4'h0;
    end else begin
      image_2126 <= 4'h6;
    end
    if (reset) begin
      image_2127 <= 4'h0;
    end else begin
      image_2127 <= 4'h6;
    end
    if (reset) begin
      image_2128 <= 4'h0;
    end else begin
      image_2128 <= 4'h6;
    end
    if (reset) begin
      image_2129 <= 4'h0;
    end else begin
      image_2129 <= 4'h6;
    end
    if (reset) begin
      image_2130 <= 4'h0;
    end else begin
      image_2130 <= 4'h6;
    end
    if (reset) begin
      image_2131 <= 4'h0;
    end else begin
      image_2131 <= 4'h6;
    end
    if (reset) begin
      image_2132 <= 4'h0;
    end else begin
      image_2132 <= 4'h6;
    end
    if (reset) begin
      image_2133 <= 4'h0;
    end else begin
      image_2133 <= 4'h6;
    end
    if (reset) begin
      image_2134 <= 4'h0;
    end else begin
      image_2134 <= 4'h5;
    end
    if (reset) begin
      image_2135 <= 4'h0;
    end else begin
      image_2135 <= 4'h5;
    end
    if (reset) begin
      image_2136 <= 4'h0;
    end else begin
      image_2136 <= 4'h6;
    end
    if (reset) begin
      image_2137 <= 4'h0;
    end else begin
      image_2137 <= 4'h5;
    end
    if (reset) begin
      image_2138 <= 4'h0;
    end else begin
      image_2138 <= 4'h3;
    end
    if (reset) begin
      image_2139 <= 4'h0;
    end else begin
      image_2139 <= 4'h2;
    end
    if (reset) begin
      image_2140 <= 4'h0;
    end else begin
      image_2140 <= 4'h4;
    end
    if (reset) begin
      image_2141 <= 4'h0;
    end else begin
      image_2141 <= 4'h4;
    end
    if (reset) begin
      image_2142 <= 4'h0;
    end else begin
      image_2142 <= 4'h4;
    end
    if (reset) begin
      image_2143 <= 4'h0;
    end else begin
      image_2143 <= 4'h4;
    end
    if (reset) begin
      image_2144 <= 4'h0;
    end else begin
      image_2144 <= 4'h4;
    end
    if (reset) begin
      image_2145 <= 4'h0;
    end else begin
      image_2145 <= 4'h4;
    end
    if (reset) begin
      image_2146 <= 4'h0;
    end else begin
      image_2146 <= 4'h4;
    end
    if (reset) begin
      image_2147 <= 4'h0;
    end else begin
      image_2147 <= 4'h4;
    end
    if (reset) begin
      image_2148 <= 4'h0;
    end else begin
      image_2148 <= 4'h4;
    end
    if (reset) begin
      image_2149 <= 4'h0;
    end else begin
      image_2149 <= 4'h5;
    end
    if (reset) begin
      image_2150 <= 4'h0;
    end else begin
      image_2150 <= 4'h5;
    end
    if (reset) begin
      image_2151 <= 4'h0;
    end else begin
      image_2151 <= 4'h5;
    end
    if (reset) begin
      image_2152 <= 4'h0;
    end else begin
      image_2152 <= 4'h5;
    end
    if (reset) begin
      image_2153 <= 4'h0;
    end else begin
      image_2153 <= 4'h5;
    end
    if (reset) begin
      image_2154 <= 4'h0;
    end else begin
      image_2154 <= 4'h5;
    end
    if (reset) begin
      image_2155 <= 4'h0;
    end else begin
      image_2155 <= 4'h5;
    end
    if (reset) begin
      image_2156 <= 4'h0;
    end else begin
      image_2156 <= 4'h5;
    end
    if (reset) begin
      image_2157 <= 4'h0;
    end else begin
      image_2157 <= 4'h5;
    end
    if (reset) begin
      image_2158 <= 4'h0;
    end else begin
      image_2158 <= 4'h5;
    end
    if (reset) begin
      image_2159 <= 4'h0;
    end else begin
      image_2159 <= 4'h5;
    end
    if (reset) begin
      image_2160 <= 4'h0;
    end else begin
      image_2160 <= 4'h6;
    end
    if (reset) begin
      image_2161 <= 4'h0;
    end else begin
      image_2161 <= 4'h6;
    end
    if (reset) begin
      image_2162 <= 4'h0;
    end else begin
      image_2162 <= 4'h6;
    end
    if (reset) begin
      image_2163 <= 4'h0;
    end else begin
      image_2163 <= 4'h6;
    end
    if (reset) begin
      image_2164 <= 4'h0;
    end else begin
      image_2164 <= 4'h6;
    end
    if (reset) begin
      image_2165 <= 4'h0;
    end else begin
      image_2165 <= 4'h6;
    end
    if (reset) begin
      image_2166 <= 4'h0;
    end else begin
      image_2166 <= 4'h6;
    end
    if (reset) begin
      image_2167 <= 4'h0;
    end else begin
      image_2167 <= 4'h4;
    end
    if (reset) begin
      image_2168 <= 4'h0;
    end else begin
      image_2168 <= 4'h6;
    end
    if (reset) begin
      image_2169 <= 4'h0;
    end else begin
      image_2169 <= 4'h6;
    end
    if (reset) begin
      image_2170 <= 4'h0;
    end else begin
      image_2170 <= 4'h1;
    end
    if (reset) begin
      image_2177 <= 4'h0;
    end else begin
      image_2177 <= 4'h1;
    end
    if (reset) begin
      image_2178 <= 4'h0;
    end else begin
      image_2178 <= 4'h3;
    end
    if (reset) begin
      image_2179 <= 4'h0;
    end else begin
      image_2179 <= 4'h5;
    end
    if (reset) begin
      image_2180 <= 4'h0;
    end else begin
      image_2180 <= 4'h5;
    end
    if (reset) begin
      image_2181 <= 4'h0;
    end else begin
      image_2181 <= 4'h5;
    end
    if (reset) begin
      image_2182 <= 4'h0;
    end else begin
      image_2182 <= 4'h5;
    end
    if (reset) begin
      image_2183 <= 4'h0;
    end else begin
      image_2183 <= 4'h5;
    end
    if (reset) begin
      image_2184 <= 4'h0;
    end else begin
      image_2184 <= 4'h6;
    end
    if (reset) begin
      image_2185 <= 4'h0;
    end else begin
      image_2185 <= 4'h6;
    end
    if (reset) begin
      image_2186 <= 4'h0;
    end else begin
      image_2186 <= 4'h6;
    end
    if (reset) begin
      image_2187 <= 4'h0;
    end else begin
      image_2187 <= 4'h6;
    end
    if (reset) begin
      image_2188 <= 4'h0;
    end else begin
      image_2188 <= 4'h6;
    end
    if (reset) begin
      image_2189 <= 4'h0;
    end else begin
      image_2189 <= 4'h6;
    end
    if (reset) begin
      image_2190 <= 4'h0;
    end else begin
      image_2190 <= 4'h6;
    end
    if (reset) begin
      image_2191 <= 4'h0;
    end else begin
      image_2191 <= 4'h6;
    end
    if (reset) begin
      image_2192 <= 4'h0;
    end else begin
      image_2192 <= 4'h6;
    end
    if (reset) begin
      image_2193 <= 4'h0;
    end else begin
      image_2193 <= 4'h6;
    end
    if (reset) begin
      image_2194 <= 4'h0;
    end else begin
      image_2194 <= 4'h6;
    end
    if (reset) begin
      image_2195 <= 4'h0;
    end else begin
      image_2195 <= 4'h6;
    end
    if (reset) begin
      image_2196 <= 4'h0;
    end else begin
      image_2196 <= 4'h6;
    end
    if (reset) begin
      image_2197 <= 4'h0;
    end else begin
      image_2197 <= 4'h6;
    end
    if (reset) begin
      image_2198 <= 4'h0;
    end else begin
      image_2198 <= 4'h6;
    end
    if (reset) begin
      image_2199 <= 4'h0;
    end else begin
      image_2199 <= 4'h4;
    end
    if (reset) begin
      image_2200 <= 4'h0;
    end else begin
      image_2200 <= 4'h6;
    end
    if (reset) begin
      image_2201 <= 4'h0;
    end else begin
      image_2201 <= 4'h6;
    end
    if (reset) begin
      image_2202 <= 4'h0;
    end else begin
      image_2202 <= 4'h6;
    end
    if (reset) begin
      image_2203 <= 4'h0;
    end else begin
      image_2203 <= 4'h5;
    end
    if (reset) begin
      image_2204 <= 4'h0;
    end else begin
      image_2204 <= 4'h3;
    end
    if (reset) begin
      image_2205 <= 4'h0;
    end else begin
      image_2205 <= 4'h4;
    end
    if (reset) begin
      image_2206 <= 4'h0;
    end else begin
      image_2206 <= 4'h4;
    end
    if (reset) begin
      image_2207 <= 4'h0;
    end else begin
      image_2207 <= 4'h4;
    end
    if (reset) begin
      image_2208 <= 4'h0;
    end else begin
      image_2208 <= 4'h4;
    end
    if (reset) begin
      image_2209 <= 4'h0;
    end else begin
      image_2209 <= 4'h4;
    end
    if (reset) begin
      image_2210 <= 4'h0;
    end else begin
      image_2210 <= 4'h4;
    end
    if (reset) begin
      image_2211 <= 4'h0;
    end else begin
      image_2211 <= 4'h4;
    end
    if (reset) begin
      image_2212 <= 4'h0;
    end else begin
      image_2212 <= 4'h5;
    end
    if (reset) begin
      image_2213 <= 4'h0;
    end else begin
      image_2213 <= 4'h5;
    end
    if (reset) begin
      image_2214 <= 4'h0;
    end else begin
      image_2214 <= 4'h5;
    end
    if (reset) begin
      image_2215 <= 4'h0;
    end else begin
      image_2215 <= 4'h5;
    end
    if (reset) begin
      image_2216 <= 4'h0;
    end else begin
      image_2216 <= 4'h5;
    end
    if (reset) begin
      image_2217 <= 4'h0;
    end else begin
      image_2217 <= 4'h5;
    end
    if (reset) begin
      image_2218 <= 4'h0;
    end else begin
      image_2218 <= 4'h5;
    end
    if (reset) begin
      image_2219 <= 4'h0;
    end else begin
      image_2219 <= 4'h5;
    end
    if (reset) begin
      image_2220 <= 4'h0;
    end else begin
      image_2220 <= 4'h5;
    end
    if (reset) begin
      image_2221 <= 4'h0;
    end else begin
      image_2221 <= 4'h5;
    end
    if (reset) begin
      image_2222 <= 4'h0;
    end else begin
      image_2222 <= 4'h5;
    end
    if (reset) begin
      image_2223 <= 4'h0;
    end else begin
      image_2223 <= 4'h6;
    end
    if (reset) begin
      image_2224 <= 4'h0;
    end else begin
      image_2224 <= 4'h6;
    end
    if (reset) begin
      image_2225 <= 4'h0;
    end else begin
      image_2225 <= 4'h6;
    end
    if (reset) begin
      image_2226 <= 4'h0;
    end else begin
      image_2226 <= 4'h6;
    end
    if (reset) begin
      image_2227 <= 4'h0;
    end else begin
      image_2227 <= 4'h6;
    end
    if (reset) begin
      image_2228 <= 4'h0;
    end else begin
      image_2228 <= 4'h6;
    end
    if (reset) begin
      image_2229 <= 4'h0;
    end else begin
      image_2229 <= 4'h6;
    end
    if (reset) begin
      image_2230 <= 4'h0;
    end else begin
      image_2230 <= 4'h6;
    end
    if (reset) begin
      image_2231 <= 4'h0;
    end else begin
      image_2231 <= 4'h4;
    end
    if (reset) begin
      image_2232 <= 4'h0;
    end else begin
      image_2232 <= 4'h6;
    end
    if (reset) begin
      image_2233 <= 4'h0;
    end else begin
      image_2233 <= 4'h6;
    end
    if (reset) begin
      image_2234 <= 4'h0;
    end else begin
      image_2234 <= 4'h2;
    end
    if (reset) begin
      image_2243 <= 4'h0;
    end else begin
      image_2243 <= 4'h5;
    end
    if (reset) begin
      image_2244 <= 4'h0;
    end else begin
      image_2244 <= 4'h5;
    end
    if (reset) begin
      image_2245 <= 4'h0;
    end else begin
      image_2245 <= 4'h5;
    end
    if (reset) begin
      image_2246 <= 4'h0;
    end else begin
      image_2246 <= 4'h5;
    end
    if (reset) begin
      image_2247 <= 4'h0;
    end else begin
      image_2247 <= 4'h5;
    end
    if (reset) begin
      image_2248 <= 4'h0;
    end else begin
      image_2248 <= 4'h6;
    end
    if (reset) begin
      image_2249 <= 4'h0;
    end else begin
      image_2249 <= 4'h6;
    end
    if (reset) begin
      image_2250 <= 4'h0;
    end else begin
      image_2250 <= 4'h6;
    end
    if (reset) begin
      image_2251 <= 4'h0;
    end else begin
      image_2251 <= 4'h6;
    end
    if (reset) begin
      image_2252 <= 4'h0;
    end else begin
      image_2252 <= 4'h6;
    end
    if (reset) begin
      image_2253 <= 4'h0;
    end else begin
      image_2253 <= 4'h6;
    end
    if (reset) begin
      image_2254 <= 4'h0;
    end else begin
      image_2254 <= 4'h6;
    end
    if (reset) begin
      image_2255 <= 4'h0;
    end else begin
      image_2255 <= 4'h6;
    end
    if (reset) begin
      image_2256 <= 4'h0;
    end else begin
      image_2256 <= 4'h6;
    end
    if (reset) begin
      image_2257 <= 4'h0;
    end else begin
      image_2257 <= 4'h6;
    end
    if (reset) begin
      image_2258 <= 4'h0;
    end else begin
      image_2258 <= 4'h6;
    end
    if (reset) begin
      image_2259 <= 4'h0;
    end else begin
      image_2259 <= 4'h6;
    end
    if (reset) begin
      image_2260 <= 4'h0;
    end else begin
      image_2260 <= 4'h6;
    end
    if (reset) begin
      image_2261 <= 4'h0;
    end else begin
      image_2261 <= 4'h6;
    end
    if (reset) begin
      image_2262 <= 4'h0;
    end else begin
      image_2262 <= 4'h6;
    end
    if (reset) begin
      image_2263 <= 4'h0;
    end else begin
      image_2263 <= 4'h6;
    end
    if (reset) begin
      image_2264 <= 4'h0;
    end else begin
      image_2264 <= 4'h4;
    end
    if (reset) begin
      image_2265 <= 4'h0;
    end else begin
      image_2265 <= 4'h5;
    end
    if (reset) begin
      image_2266 <= 4'h0;
    end else begin
      image_2266 <= 4'h6;
    end
    if (reset) begin
      image_2267 <= 4'h0;
    end else begin
      image_2267 <= 4'h6;
    end
    if (reset) begin
      image_2268 <= 4'h0;
    end else begin
      image_2268 <= 4'h6;
    end
    if (reset) begin
      image_2269 <= 4'h0;
    end else begin
      image_2269 <= 4'h2;
    end
    if (reset) begin
      image_2270 <= 4'h0;
    end else begin
      image_2270 <= 4'h4;
    end
    if (reset) begin
      image_2271 <= 4'h0;
    end else begin
      image_2271 <= 4'h4;
    end
    if (reset) begin
      image_2272 <= 4'h0;
    end else begin
      image_2272 <= 4'h4;
    end
    if (reset) begin
      image_2273 <= 4'h0;
    end else begin
      image_2273 <= 4'h4;
    end
    if (reset) begin
      image_2274 <= 4'h0;
    end else begin
      image_2274 <= 4'h5;
    end
    if (reset) begin
      image_2275 <= 4'h0;
    end else begin
      image_2275 <= 4'h5;
    end
    if (reset) begin
      image_2276 <= 4'h0;
    end else begin
      image_2276 <= 4'h5;
    end
    if (reset) begin
      image_2277 <= 4'h0;
    end else begin
      image_2277 <= 4'h5;
    end
    if (reset) begin
      image_2278 <= 4'h0;
    end else begin
      image_2278 <= 4'h5;
    end
    if (reset) begin
      image_2279 <= 4'h0;
    end else begin
      image_2279 <= 4'h5;
    end
    if (reset) begin
      image_2280 <= 4'h0;
    end else begin
      image_2280 <= 4'h5;
    end
    if (reset) begin
      image_2281 <= 4'h0;
    end else begin
      image_2281 <= 4'h5;
    end
    if (reset) begin
      image_2282 <= 4'h0;
    end else begin
      image_2282 <= 4'h5;
    end
    if (reset) begin
      image_2283 <= 4'h0;
    end else begin
      image_2283 <= 4'h5;
    end
    if (reset) begin
      image_2284 <= 4'h0;
    end else begin
      image_2284 <= 4'h5;
    end
    if (reset) begin
      image_2285 <= 4'h0;
    end else begin
      image_2285 <= 4'h5;
    end
    if (reset) begin
      image_2286 <= 4'h0;
    end else begin
      image_2286 <= 4'h6;
    end
    if (reset) begin
      image_2287 <= 4'h0;
    end else begin
      image_2287 <= 4'h6;
    end
    if (reset) begin
      image_2288 <= 4'h0;
    end else begin
      image_2288 <= 4'h6;
    end
    if (reset) begin
      image_2289 <= 4'h0;
    end else begin
      image_2289 <= 4'h6;
    end
    if (reset) begin
      image_2290 <= 4'h0;
    end else begin
      image_2290 <= 4'h6;
    end
    if (reset) begin
      image_2291 <= 4'h0;
    end else begin
      image_2291 <= 4'h6;
    end
    if (reset) begin
      image_2292 <= 4'h0;
    end else begin
      image_2292 <= 4'h6;
    end
    if (reset) begin
      image_2293 <= 4'h0;
    end else begin
      image_2293 <= 4'h6;
    end
    if (reset) begin
      image_2294 <= 4'h0;
    end else begin
      image_2294 <= 4'h6;
    end
    if (reset) begin
      image_2295 <= 4'h0;
    end else begin
      image_2295 <= 4'h3;
    end
    if (reset) begin
      image_2296 <= 4'h0;
    end else begin
      image_2296 <= 4'h6;
    end
    if (reset) begin
      image_2297 <= 4'h0;
    end else begin
      image_2297 <= 4'h6;
    end
    if (reset) begin
      image_2298 <= 4'h0;
    end else begin
      image_2298 <= 4'h2;
    end
    if (reset) begin
      image_2307 <= 4'h0;
    end else begin
      image_2307 <= 4'h2;
    end
    if (reset) begin
      image_2308 <= 4'h0;
    end else begin
      image_2308 <= 4'h5;
    end
    if (reset) begin
      image_2309 <= 4'h0;
    end else begin
      image_2309 <= 4'h5;
    end
    if (reset) begin
      image_2310 <= 4'h0;
    end else begin
      image_2310 <= 4'h5;
    end
    if (reset) begin
      image_2311 <= 4'h0;
    end else begin
      image_2311 <= 4'h5;
    end
    if (reset) begin
      image_2312 <= 4'h0;
    end else begin
      image_2312 <= 4'h5;
    end
    if (reset) begin
      image_2313 <= 4'h0;
    end else begin
      image_2313 <= 4'h6;
    end
    if (reset) begin
      image_2314 <= 4'h0;
    end else begin
      image_2314 <= 4'h6;
    end
    if (reset) begin
      image_2315 <= 4'h0;
    end else begin
      image_2315 <= 4'h6;
    end
    if (reset) begin
      image_2316 <= 4'h0;
    end else begin
      image_2316 <= 4'h6;
    end
    if (reset) begin
      image_2317 <= 4'h0;
    end else begin
      image_2317 <= 4'h6;
    end
    if (reset) begin
      image_2318 <= 4'h0;
    end else begin
      image_2318 <= 4'h6;
    end
    if (reset) begin
      image_2319 <= 4'h0;
    end else begin
      image_2319 <= 4'h6;
    end
    if (reset) begin
      image_2320 <= 4'h0;
    end else begin
      image_2320 <= 4'h6;
    end
    if (reset) begin
      image_2321 <= 4'h0;
    end else begin
      image_2321 <= 4'h6;
    end
    if (reset) begin
      image_2322 <= 4'h0;
    end else begin
      image_2322 <= 4'h6;
    end
    if (reset) begin
      image_2323 <= 4'h0;
    end else begin
      image_2323 <= 4'h6;
    end
    if (reset) begin
      image_2324 <= 4'h0;
    end else begin
      image_2324 <= 4'h6;
    end
    if (reset) begin
      image_2325 <= 4'h0;
    end else begin
      image_2325 <= 4'h6;
    end
    if (reset) begin
      image_2326 <= 4'h0;
    end else begin
      image_2326 <= 4'h6;
    end
    if (reset) begin
      image_2327 <= 4'h0;
    end else begin
      image_2327 <= 4'h6;
    end
    if (reset) begin
      image_2328 <= 4'h0;
    end else begin
      image_2328 <= 4'h6;
    end
    if (reset) begin
      image_2329 <= 4'h0;
    end else begin
      image_2329 <= 4'h4;
    end
    if (reset) begin
      image_2330 <= 4'h0;
    end else begin
      image_2330 <= 4'h5;
    end
    if (reset) begin
      image_2331 <= 4'h0;
    end else begin
      image_2331 <= 4'h6;
    end
    if (reset) begin
      image_2332 <= 4'h0;
    end else begin
      image_2332 <= 4'h6;
    end
    if (reset) begin
      image_2333 <= 4'h0;
    end else begin
      image_2333 <= 4'h5;
    end
    if (reset) begin
      image_2334 <= 4'h0;
    end else begin
      image_2334 <= 4'h2;
    end
    if (reset) begin
      image_2335 <= 4'h0;
    end else begin
      image_2335 <= 4'h4;
    end
    if (reset) begin
      image_2336 <= 4'h0;
    end else begin
      image_2336 <= 4'h5;
    end
    if (reset) begin
      image_2337 <= 4'h0;
    end else begin
      image_2337 <= 4'h5;
    end
    if (reset) begin
      image_2338 <= 4'h0;
    end else begin
      image_2338 <= 4'h5;
    end
    if (reset) begin
      image_2339 <= 4'h0;
    end else begin
      image_2339 <= 4'h5;
    end
    if (reset) begin
      image_2340 <= 4'h0;
    end else begin
      image_2340 <= 4'h5;
    end
    if (reset) begin
      image_2341 <= 4'h0;
    end else begin
      image_2341 <= 4'h5;
    end
    if (reset) begin
      image_2342 <= 4'h0;
    end else begin
      image_2342 <= 4'h5;
    end
    if (reset) begin
      image_2343 <= 4'h0;
    end else begin
      image_2343 <= 4'h5;
    end
    if (reset) begin
      image_2344 <= 4'h0;
    end else begin
      image_2344 <= 4'h5;
    end
    if (reset) begin
      image_2345 <= 4'h0;
    end else begin
      image_2345 <= 4'h5;
    end
    if (reset) begin
      image_2346 <= 4'h0;
    end else begin
      image_2346 <= 4'h5;
    end
    if (reset) begin
      image_2347 <= 4'h0;
    end else begin
      image_2347 <= 4'h5;
    end
    if (reset) begin
      image_2348 <= 4'h0;
    end else begin
      image_2348 <= 4'h6;
    end
    if (reset) begin
      image_2349 <= 4'h0;
    end else begin
      image_2349 <= 4'h6;
    end
    if (reset) begin
      image_2350 <= 4'h0;
    end else begin
      image_2350 <= 4'h6;
    end
    if (reset) begin
      image_2351 <= 4'h0;
    end else begin
      image_2351 <= 4'h6;
    end
    if (reset) begin
      image_2352 <= 4'h0;
    end else begin
      image_2352 <= 4'h6;
    end
    if (reset) begin
      image_2353 <= 4'h0;
    end else begin
      image_2353 <= 4'h6;
    end
    if (reset) begin
      image_2354 <= 4'h0;
    end else begin
      image_2354 <= 4'h6;
    end
    if (reset) begin
      image_2355 <= 4'h0;
    end else begin
      image_2355 <= 4'h6;
    end
    if (reset) begin
      image_2356 <= 4'h0;
    end else begin
      image_2356 <= 4'h6;
    end
    if (reset) begin
      image_2357 <= 4'h0;
    end else begin
      image_2357 <= 4'h6;
    end
    if (reset) begin
      image_2358 <= 4'h0;
    end else begin
      image_2358 <= 4'h6;
    end
    if (reset) begin
      image_2359 <= 4'h0;
    end else begin
      image_2359 <= 4'h3;
    end
    if (reset) begin
      image_2360 <= 4'h0;
    end else begin
      image_2360 <= 4'h6;
    end
    if (reset) begin
      image_2361 <= 4'h0;
    end else begin
      image_2361 <= 4'h6;
    end
    if (reset) begin
      image_2362 <= 4'h0;
    end else begin
      image_2362 <= 4'h2;
    end
    if (reset) begin
      image_2372 <= 4'h0;
    end else begin
      image_2372 <= 4'h3;
    end
    if (reset) begin
      image_2373 <= 4'h0;
    end else begin
      image_2373 <= 4'h5;
    end
    if (reset) begin
      image_2374 <= 4'h0;
    end else begin
      image_2374 <= 4'h5;
    end
    if (reset) begin
      image_2375 <= 4'h0;
    end else begin
      image_2375 <= 4'h5;
    end
    if (reset) begin
      image_2376 <= 4'h0;
    end else begin
      image_2376 <= 4'h5;
    end
    if (reset) begin
      image_2377 <= 4'h0;
    end else begin
      image_2377 <= 4'h5;
    end
    if (reset) begin
      image_2378 <= 4'h0;
    end else begin
      image_2378 <= 4'h6;
    end
    if (reset) begin
      image_2379 <= 4'h0;
    end else begin
      image_2379 <= 4'h6;
    end
    if (reset) begin
      image_2380 <= 4'h0;
    end else begin
      image_2380 <= 4'h6;
    end
    if (reset) begin
      image_2381 <= 4'h0;
    end else begin
      image_2381 <= 4'h6;
    end
    if (reset) begin
      image_2382 <= 4'h0;
    end else begin
      image_2382 <= 4'h6;
    end
    if (reset) begin
      image_2383 <= 4'h0;
    end else begin
      image_2383 <= 4'h6;
    end
    if (reset) begin
      image_2384 <= 4'h0;
    end else begin
      image_2384 <= 4'h6;
    end
    if (reset) begin
      image_2385 <= 4'h0;
    end else begin
      image_2385 <= 4'h6;
    end
    if (reset) begin
      image_2386 <= 4'h0;
    end else begin
      image_2386 <= 4'h6;
    end
    if (reset) begin
      image_2387 <= 4'h0;
    end else begin
      image_2387 <= 4'h6;
    end
    if (reset) begin
      image_2388 <= 4'h0;
    end else begin
      image_2388 <= 4'h6;
    end
    if (reset) begin
      image_2389 <= 4'h0;
    end else begin
      image_2389 <= 4'h6;
    end
    if (reset) begin
      image_2390 <= 4'h0;
    end else begin
      image_2390 <= 4'h6;
    end
    if (reset) begin
      image_2391 <= 4'h0;
    end else begin
      image_2391 <= 4'h6;
    end
    if (reset) begin
      image_2392 <= 4'h0;
    end else begin
      image_2392 <= 4'h6;
    end
    if (reset) begin
      image_2393 <= 4'h0;
    end else begin
      image_2393 <= 4'h6;
    end
    if (reset) begin
      image_2394 <= 4'h0;
    end else begin
      image_2394 <= 4'h4;
    end
    if (reset) begin
      image_2395 <= 4'h0;
    end else begin
      image_2395 <= 4'h5;
    end
    if (reset) begin
      image_2396 <= 4'h0;
    end else begin
      image_2396 <= 4'h6;
    end
    if (reset) begin
      image_2397 <= 4'h0;
    end else begin
      image_2397 <= 4'h6;
    end
    if (reset) begin
      image_2398 <= 4'h0;
    end else begin
      image_2398 <= 4'h5;
    end
    if (reset) begin
      image_2399 <= 4'h0;
    end else begin
      image_2399 <= 4'h3;
    end
    if (reset) begin
      image_2400 <= 4'h0;
    end else begin
      image_2400 <= 4'h5;
    end
    if (reset) begin
      image_2401 <= 4'h0;
    end else begin
      image_2401 <= 4'h5;
    end
    if (reset) begin
      image_2402 <= 4'h0;
    end else begin
      image_2402 <= 4'h5;
    end
    if (reset) begin
      image_2403 <= 4'h0;
    end else begin
      image_2403 <= 4'h5;
    end
    if (reset) begin
      image_2404 <= 4'h0;
    end else begin
      image_2404 <= 4'h5;
    end
    if (reset) begin
      image_2405 <= 4'h0;
    end else begin
      image_2405 <= 4'h5;
    end
    if (reset) begin
      image_2406 <= 4'h0;
    end else begin
      image_2406 <= 4'h5;
    end
    if (reset) begin
      image_2407 <= 4'h0;
    end else begin
      image_2407 <= 4'h5;
    end
    if (reset) begin
      image_2408 <= 4'h0;
    end else begin
      image_2408 <= 4'h5;
    end
    if (reset) begin
      image_2409 <= 4'h0;
    end else begin
      image_2409 <= 4'h5;
    end
    if (reset) begin
      image_2410 <= 4'h0;
    end else begin
      image_2410 <= 4'h6;
    end
    if (reset) begin
      image_2411 <= 4'h0;
    end else begin
      image_2411 <= 4'h6;
    end
    if (reset) begin
      image_2412 <= 4'h0;
    end else begin
      image_2412 <= 4'h6;
    end
    if (reset) begin
      image_2413 <= 4'h0;
    end else begin
      image_2413 <= 4'h6;
    end
    if (reset) begin
      image_2414 <= 4'h0;
    end else begin
      image_2414 <= 4'h6;
    end
    if (reset) begin
      image_2415 <= 4'h0;
    end else begin
      image_2415 <= 4'h6;
    end
    if (reset) begin
      image_2416 <= 4'h0;
    end else begin
      image_2416 <= 4'h6;
    end
    if (reset) begin
      image_2417 <= 4'h0;
    end else begin
      image_2417 <= 4'h6;
    end
    if (reset) begin
      image_2418 <= 4'h0;
    end else begin
      image_2418 <= 4'h6;
    end
    if (reset) begin
      image_2419 <= 4'h0;
    end else begin
      image_2419 <= 4'h6;
    end
    if (reset) begin
      image_2420 <= 4'h0;
    end else begin
      image_2420 <= 4'h6;
    end
    if (reset) begin
      image_2421 <= 4'h0;
    end else begin
      image_2421 <= 4'h6;
    end
    if (reset) begin
      image_2422 <= 4'h0;
    end else begin
      image_2422 <= 4'h6;
    end
    if (reset) begin
      image_2423 <= 4'h0;
    end else begin
      image_2423 <= 4'h4;
    end
    if (reset) begin
      image_2424 <= 4'h0;
    end else begin
      image_2424 <= 4'h6;
    end
    if (reset) begin
      image_2425 <= 4'h0;
    end else begin
      image_2425 <= 4'h6;
    end
    if (reset) begin
      image_2426 <= 4'h0;
    end else begin
      image_2426 <= 4'h2;
    end
    if (reset) begin
      image_2437 <= 4'h0;
    end else begin
      image_2437 <= 4'h4;
    end
    if (reset) begin
      image_2438 <= 4'h0;
    end else begin
      image_2438 <= 4'h5;
    end
    if (reset) begin
      image_2439 <= 4'h0;
    end else begin
      image_2439 <= 4'h5;
    end
    if (reset) begin
      image_2440 <= 4'h0;
    end else begin
      image_2440 <= 4'h5;
    end
    if (reset) begin
      image_2441 <= 4'h0;
    end else begin
      image_2441 <= 4'h5;
    end
    if (reset) begin
      image_2442 <= 4'h0;
    end else begin
      image_2442 <= 4'h5;
    end
    if (reset) begin
      image_2443 <= 4'h0;
    end else begin
      image_2443 <= 4'h6;
    end
    if (reset) begin
      image_2444 <= 4'h0;
    end else begin
      image_2444 <= 4'h6;
    end
    if (reset) begin
      image_2445 <= 4'h0;
    end else begin
      image_2445 <= 4'h6;
    end
    if (reset) begin
      image_2446 <= 4'h0;
    end else begin
      image_2446 <= 4'h6;
    end
    if (reset) begin
      image_2447 <= 4'h0;
    end else begin
      image_2447 <= 4'h6;
    end
    if (reset) begin
      image_2448 <= 4'h0;
    end else begin
      image_2448 <= 4'h6;
    end
    if (reset) begin
      image_2449 <= 4'h0;
    end else begin
      image_2449 <= 4'h6;
    end
    if (reset) begin
      image_2450 <= 4'h0;
    end else begin
      image_2450 <= 4'h6;
    end
    if (reset) begin
      image_2451 <= 4'h0;
    end else begin
      image_2451 <= 4'h6;
    end
    if (reset) begin
      image_2452 <= 4'h0;
    end else begin
      image_2452 <= 4'h6;
    end
    if (reset) begin
      image_2453 <= 4'h0;
    end else begin
      image_2453 <= 4'h6;
    end
    if (reset) begin
      image_2454 <= 4'h0;
    end else begin
      image_2454 <= 4'h6;
    end
    if (reset) begin
      image_2455 <= 4'h0;
    end else begin
      image_2455 <= 4'h6;
    end
    if (reset) begin
      image_2456 <= 4'h0;
    end else begin
      image_2456 <= 4'h6;
    end
    if (reset) begin
      image_2457 <= 4'h0;
    end else begin
      image_2457 <= 4'h6;
    end
    if (reset) begin
      image_2458 <= 4'h0;
    end else begin
      image_2458 <= 4'h6;
    end
    if (reset) begin
      image_2459 <= 4'h0;
    end else begin
      image_2459 <= 4'h5;
    end
    if (reset) begin
      image_2460 <= 4'h0;
    end else begin
      image_2460 <= 4'h4;
    end
    if (reset) begin
      image_2461 <= 4'h0;
    end else begin
      image_2461 <= 4'h6;
    end
    if (reset) begin
      image_2462 <= 4'h0;
    end else begin
      image_2462 <= 4'h6;
    end
    if (reset) begin
      image_2463 <= 4'h0;
    end else begin
      image_2463 <= 4'h6;
    end
    if (reset) begin
      image_2464 <= 4'h0;
    end else begin
      image_2464 <= 4'h4;
    end
    if (reset) begin
      image_2465 <= 4'h0;
    end else begin
      image_2465 <= 4'h3;
    end
    if (reset) begin
      image_2466 <= 4'h0;
    end else begin
      image_2466 <= 4'h5;
    end
    if (reset) begin
      image_2467 <= 4'h0;
    end else begin
      image_2467 <= 4'h5;
    end
    if (reset) begin
      image_2468 <= 4'h0;
    end else begin
      image_2468 <= 4'h5;
    end
    if (reset) begin
      image_2469 <= 4'h0;
    end else begin
      image_2469 <= 4'h5;
    end
    if (reset) begin
      image_2470 <= 4'h0;
    end else begin
      image_2470 <= 4'h5;
    end
    if (reset) begin
      image_2471 <= 4'h0;
    end else begin
      image_2471 <= 4'h5;
    end
    if (reset) begin
      image_2472 <= 4'h0;
    end else begin
      image_2472 <= 4'h6;
    end
    if (reset) begin
      image_2473 <= 4'h0;
    end else begin
      image_2473 <= 4'h6;
    end
    if (reset) begin
      image_2474 <= 4'h0;
    end else begin
      image_2474 <= 4'h6;
    end
    if (reset) begin
      image_2475 <= 4'h0;
    end else begin
      image_2475 <= 4'h6;
    end
    if (reset) begin
      image_2476 <= 4'h0;
    end else begin
      image_2476 <= 4'h6;
    end
    if (reset) begin
      image_2477 <= 4'h0;
    end else begin
      image_2477 <= 4'h6;
    end
    if (reset) begin
      image_2478 <= 4'h0;
    end else begin
      image_2478 <= 4'h6;
    end
    if (reset) begin
      image_2479 <= 4'h0;
    end else begin
      image_2479 <= 4'h6;
    end
    if (reset) begin
      image_2480 <= 4'h0;
    end else begin
      image_2480 <= 4'h6;
    end
    if (reset) begin
      image_2481 <= 4'h0;
    end else begin
      image_2481 <= 4'h6;
    end
    if (reset) begin
      image_2482 <= 4'h0;
    end else begin
      image_2482 <= 4'h6;
    end
    if (reset) begin
      image_2483 <= 4'h0;
    end else begin
      image_2483 <= 4'h6;
    end
    if (reset) begin
      image_2484 <= 4'h0;
    end else begin
      image_2484 <= 4'h6;
    end
    if (reset) begin
      image_2485 <= 4'h0;
    end else begin
      image_2485 <= 4'h6;
    end
    if (reset) begin
      image_2486 <= 4'h0;
    end else begin
      image_2486 <= 4'h6;
    end
    if (reset) begin
      image_2487 <= 4'h0;
    end else begin
      image_2487 <= 4'h4;
    end
    if (reset) begin
      image_2488 <= 4'h0;
    end else begin
      image_2488 <= 4'h6;
    end
    if (reset) begin
      image_2489 <= 4'h0;
    end else begin
      image_2489 <= 4'h6;
    end
    if (reset) begin
      image_2490 <= 4'h0;
    end else begin
      image_2490 <= 4'h2;
    end
    if (reset) begin
      image_2502 <= 4'h0;
    end else begin
      image_2502 <= 4'h4;
    end
    if (reset) begin
      image_2503 <= 4'h0;
    end else begin
      image_2503 <= 4'h5;
    end
    if (reset) begin
      image_2504 <= 4'h0;
    end else begin
      image_2504 <= 4'h5;
    end
    if (reset) begin
      image_2505 <= 4'h0;
    end else begin
      image_2505 <= 4'h5;
    end
    if (reset) begin
      image_2506 <= 4'h0;
    end else begin
      image_2506 <= 4'h5;
    end
    if (reset) begin
      image_2507 <= 4'h0;
    end else begin
      image_2507 <= 4'h5;
    end
    if (reset) begin
      image_2508 <= 4'h0;
    end else begin
      image_2508 <= 4'h6;
    end
    if (reset) begin
      image_2509 <= 4'h0;
    end else begin
      image_2509 <= 4'h6;
    end
    if (reset) begin
      image_2510 <= 4'h0;
    end else begin
      image_2510 <= 4'h6;
    end
    if (reset) begin
      image_2511 <= 4'h0;
    end else begin
      image_2511 <= 4'h6;
    end
    if (reset) begin
      image_2512 <= 4'h0;
    end else begin
      image_2512 <= 4'h6;
    end
    if (reset) begin
      image_2513 <= 4'h0;
    end else begin
      image_2513 <= 4'h6;
    end
    if (reset) begin
      image_2514 <= 4'h0;
    end else begin
      image_2514 <= 4'h6;
    end
    if (reset) begin
      image_2515 <= 4'h0;
    end else begin
      image_2515 <= 4'h6;
    end
    if (reset) begin
      image_2516 <= 4'h0;
    end else begin
      image_2516 <= 4'h6;
    end
    if (reset) begin
      image_2517 <= 4'h0;
    end else begin
      image_2517 <= 4'h6;
    end
    if (reset) begin
      image_2518 <= 4'h0;
    end else begin
      image_2518 <= 4'h6;
    end
    if (reset) begin
      image_2519 <= 4'h0;
    end else begin
      image_2519 <= 4'h6;
    end
    if (reset) begin
      image_2520 <= 4'h0;
    end else begin
      image_2520 <= 4'h6;
    end
    if (reset) begin
      image_2521 <= 4'h0;
    end else begin
      image_2521 <= 4'h6;
    end
    if (reset) begin
      image_2522 <= 4'h0;
    end else begin
      image_2522 <= 4'h6;
    end
    if (reset) begin
      image_2523 <= 4'h0;
    end else begin
      image_2523 <= 4'h6;
    end
    if (reset) begin
      image_2524 <= 4'h0;
    end else begin
      image_2524 <= 4'h5;
    end
    if (reset) begin
      image_2525 <= 4'h0;
    end else begin
      image_2525 <= 4'h4;
    end
    if (reset) begin
      image_2526 <= 4'h0;
    end else begin
      image_2526 <= 4'h6;
    end
    if (reset) begin
      image_2527 <= 4'h0;
    end else begin
      image_2527 <= 4'h6;
    end
    if (reset) begin
      image_2528 <= 4'h0;
    end else begin
      image_2528 <= 4'h6;
    end
    if (reset) begin
      image_2529 <= 4'h0;
    end else begin
      image_2529 <= 4'h6;
    end
    if (reset) begin
      image_2530 <= 4'h0;
    end else begin
      image_2530 <= 4'h4;
    end
    if (reset) begin
      image_2531 <= 4'h0;
    end else begin
      image_2531 <= 4'h4;
    end
    if (reset) begin
      image_2532 <= 4'h0;
    end else begin
      image_2532 <= 4'h5;
    end
    if (reset) begin
      image_2533 <= 4'h0;
    end else begin
      image_2533 <= 4'h6;
    end
    if (reset) begin
      image_2534 <= 4'h0;
    end else begin
      image_2534 <= 4'h6;
    end
    if (reset) begin
      image_2535 <= 4'h0;
    end else begin
      image_2535 <= 4'h6;
    end
    if (reset) begin
      image_2536 <= 4'h0;
    end else begin
      image_2536 <= 4'h6;
    end
    if (reset) begin
      image_2537 <= 4'h0;
    end else begin
      image_2537 <= 4'h6;
    end
    if (reset) begin
      image_2538 <= 4'h0;
    end else begin
      image_2538 <= 4'h6;
    end
    if (reset) begin
      image_2539 <= 4'h0;
    end else begin
      image_2539 <= 4'h6;
    end
    if (reset) begin
      image_2540 <= 4'h0;
    end else begin
      image_2540 <= 4'h6;
    end
    if (reset) begin
      image_2541 <= 4'h0;
    end else begin
      image_2541 <= 4'h6;
    end
    if (reset) begin
      image_2542 <= 4'h0;
    end else begin
      image_2542 <= 4'h6;
    end
    if (reset) begin
      image_2543 <= 4'h0;
    end else begin
      image_2543 <= 4'h6;
    end
    if (reset) begin
      image_2544 <= 4'h0;
    end else begin
      image_2544 <= 4'h6;
    end
    if (reset) begin
      image_2545 <= 4'h0;
    end else begin
      image_2545 <= 4'h6;
    end
    if (reset) begin
      image_2546 <= 4'h0;
    end else begin
      image_2546 <= 4'h6;
    end
    if (reset) begin
      image_2547 <= 4'h0;
    end else begin
      image_2547 <= 4'h6;
    end
    if (reset) begin
      image_2548 <= 4'h0;
    end else begin
      image_2548 <= 4'h6;
    end
    if (reset) begin
      image_2549 <= 4'h0;
    end else begin
      image_2549 <= 4'h6;
    end
    if (reset) begin
      image_2550 <= 4'h0;
    end else begin
      image_2550 <= 4'h6;
    end
    if (reset) begin
      image_2551 <= 4'h0;
    end else begin
      image_2551 <= 4'h3;
    end
    if (reset) begin
      image_2552 <= 4'h0;
    end else begin
      image_2552 <= 4'h6;
    end
    if (reset) begin
      image_2553 <= 4'h0;
    end else begin
      image_2553 <= 4'h6;
    end
    if (reset) begin
      image_2554 <= 4'h0;
    end else begin
      image_2554 <= 4'h2;
    end
    if (reset) begin
      image_2567 <= 4'h0;
    end else begin
      image_2567 <= 4'h4;
    end
    if (reset) begin
      image_2568 <= 4'h0;
    end else begin
      image_2568 <= 4'h5;
    end
    if (reset) begin
      image_2569 <= 4'h0;
    end else begin
      image_2569 <= 4'h5;
    end
    if (reset) begin
      image_2570 <= 4'h0;
    end else begin
      image_2570 <= 4'h5;
    end
    if (reset) begin
      image_2571 <= 4'h0;
    end else begin
      image_2571 <= 4'h5;
    end
    if (reset) begin
      image_2572 <= 4'h0;
    end else begin
      image_2572 <= 4'h5;
    end
    if (reset) begin
      image_2573 <= 4'h0;
    end else begin
      image_2573 <= 4'h6;
    end
    if (reset) begin
      image_2574 <= 4'h0;
    end else begin
      image_2574 <= 4'h6;
    end
    if (reset) begin
      image_2575 <= 4'h0;
    end else begin
      image_2575 <= 4'h6;
    end
    if (reset) begin
      image_2576 <= 4'h0;
    end else begin
      image_2576 <= 4'h6;
    end
    if (reset) begin
      image_2577 <= 4'h0;
    end else begin
      image_2577 <= 4'h6;
    end
    if (reset) begin
      image_2578 <= 4'h0;
    end else begin
      image_2578 <= 4'h6;
    end
    if (reset) begin
      image_2579 <= 4'h0;
    end else begin
      image_2579 <= 4'h6;
    end
    if (reset) begin
      image_2580 <= 4'h0;
    end else begin
      image_2580 <= 4'h6;
    end
    if (reset) begin
      image_2581 <= 4'h0;
    end else begin
      image_2581 <= 4'h6;
    end
    if (reset) begin
      image_2582 <= 4'h0;
    end else begin
      image_2582 <= 4'h6;
    end
    if (reset) begin
      image_2583 <= 4'h0;
    end else begin
      image_2583 <= 4'h6;
    end
    if (reset) begin
      image_2584 <= 4'h0;
    end else begin
      image_2584 <= 4'h6;
    end
    if (reset) begin
      image_2585 <= 4'h0;
    end else begin
      image_2585 <= 4'h6;
    end
    if (reset) begin
      image_2586 <= 4'h0;
    end else begin
      image_2586 <= 4'h6;
    end
    if (reset) begin
      image_2587 <= 4'h0;
    end else begin
      image_2587 <= 4'h6;
    end
    if (reset) begin
      image_2588 <= 4'h0;
    end else begin
      image_2588 <= 4'h6;
    end
    if (reset) begin
      image_2589 <= 4'h0;
    end else begin
      image_2589 <= 4'h6;
    end
    if (reset) begin
      image_2590 <= 4'h0;
    end else begin
      image_2590 <= 4'h4;
    end
    if (reset) begin
      image_2591 <= 4'h0;
    end else begin
      image_2591 <= 4'h4;
    end
    if (reset) begin
      image_2592 <= 4'h0;
    end else begin
      image_2592 <= 4'h6;
    end
    if (reset) begin
      image_2593 <= 4'h0;
    end else begin
      image_2593 <= 4'h6;
    end
    if (reset) begin
      image_2594 <= 4'h0;
    end else begin
      image_2594 <= 4'h6;
    end
    if (reset) begin
      image_2595 <= 4'h0;
    end else begin
      image_2595 <= 4'h6;
    end
    if (reset) begin
      image_2596 <= 4'h0;
    end else begin
      image_2596 <= 4'h5;
    end
    if (reset) begin
      image_2597 <= 4'h0;
    end else begin
      image_2597 <= 4'h4;
    end
    if (reset) begin
      image_2598 <= 4'h0;
    end else begin
      image_2598 <= 4'h5;
    end
    if (reset) begin
      image_2599 <= 4'h0;
    end else begin
      image_2599 <= 4'h6;
    end
    if (reset) begin
      image_2600 <= 4'h0;
    end else begin
      image_2600 <= 4'h6;
    end
    if (reset) begin
      image_2601 <= 4'h0;
    end else begin
      image_2601 <= 4'h6;
    end
    if (reset) begin
      image_2602 <= 4'h0;
    end else begin
      image_2602 <= 4'h6;
    end
    if (reset) begin
      image_2603 <= 4'h0;
    end else begin
      image_2603 <= 4'h6;
    end
    if (reset) begin
      image_2604 <= 4'h0;
    end else begin
      image_2604 <= 4'h6;
    end
    if (reset) begin
      image_2605 <= 4'h0;
    end else begin
      image_2605 <= 4'h6;
    end
    if (reset) begin
      image_2606 <= 4'h0;
    end else begin
      image_2606 <= 4'h6;
    end
    if (reset) begin
      image_2607 <= 4'h0;
    end else begin
      image_2607 <= 4'h6;
    end
    if (reset) begin
      image_2608 <= 4'h0;
    end else begin
      image_2608 <= 4'h6;
    end
    if (reset) begin
      image_2609 <= 4'h0;
    end else begin
      image_2609 <= 4'h6;
    end
    if (reset) begin
      image_2610 <= 4'h0;
    end else begin
      image_2610 <= 4'h6;
    end
    if (reset) begin
      image_2611 <= 4'h0;
    end else begin
      image_2611 <= 4'h6;
    end
    if (reset) begin
      image_2612 <= 4'h0;
    end else begin
      image_2612 <= 4'h6;
    end
    if (reset) begin
      image_2613 <= 4'h0;
    end else begin
      image_2613 <= 4'h5;
    end
    if (reset) begin
      image_2614 <= 4'h0;
    end else begin
      image_2614 <= 4'h4;
    end
    if (reset) begin
      image_2615 <= 4'h0;
    end else begin
      image_2615 <= 4'h6;
    end
    if (reset) begin
      image_2616 <= 4'h0;
    end else begin
      image_2616 <= 4'h6;
    end
    if (reset) begin
      image_2617 <= 4'h0;
    end else begin
      image_2617 <= 4'h6;
    end
    if (reset) begin
      image_2618 <= 4'h0;
    end else begin
      image_2618 <= 4'h2;
    end
    if (reset) begin
      image_2632 <= 4'h0;
    end else begin
      image_2632 <= 4'h3;
    end
    if (reset) begin
      image_2633 <= 4'h0;
    end else begin
      image_2633 <= 4'h5;
    end
    if (reset) begin
      image_2634 <= 4'h0;
    end else begin
      image_2634 <= 4'h5;
    end
    if (reset) begin
      image_2635 <= 4'h0;
    end else begin
      image_2635 <= 4'h5;
    end
    if (reset) begin
      image_2636 <= 4'h0;
    end else begin
      image_2636 <= 4'h5;
    end
    if (reset) begin
      image_2637 <= 4'h0;
    end else begin
      image_2637 <= 4'h5;
    end
    if (reset) begin
      image_2638 <= 4'h0;
    end else begin
      image_2638 <= 4'h5;
    end
    if (reset) begin
      image_2639 <= 4'h0;
    end else begin
      image_2639 <= 4'h6;
    end
    if (reset) begin
      image_2640 <= 4'h0;
    end else begin
      image_2640 <= 4'h6;
    end
    if (reset) begin
      image_2641 <= 4'h0;
    end else begin
      image_2641 <= 4'h6;
    end
    if (reset) begin
      image_2642 <= 4'h0;
    end else begin
      image_2642 <= 4'h6;
    end
    if (reset) begin
      image_2643 <= 4'h0;
    end else begin
      image_2643 <= 4'h6;
    end
    if (reset) begin
      image_2644 <= 4'h0;
    end else begin
      image_2644 <= 4'h6;
    end
    if (reset) begin
      image_2645 <= 4'h0;
    end else begin
      image_2645 <= 4'h6;
    end
    if (reset) begin
      image_2646 <= 4'h0;
    end else begin
      image_2646 <= 4'h6;
    end
    if (reset) begin
      image_2647 <= 4'h0;
    end else begin
      image_2647 <= 4'h6;
    end
    if (reset) begin
      image_2648 <= 4'h0;
    end else begin
      image_2648 <= 4'h6;
    end
    if (reset) begin
      image_2649 <= 4'h0;
    end else begin
      image_2649 <= 4'h6;
    end
    if (reset) begin
      image_2650 <= 4'h0;
    end else begin
      image_2650 <= 4'h6;
    end
    if (reset) begin
      image_2651 <= 4'h0;
    end else begin
      image_2651 <= 4'h6;
    end
    if (reset) begin
      image_2652 <= 4'h0;
    end else begin
      image_2652 <= 4'h6;
    end
    if (reset) begin
      image_2653 <= 4'h0;
    end else begin
      image_2653 <= 4'h6;
    end
    if (reset) begin
      image_2654 <= 4'h0;
    end else begin
      image_2654 <= 4'h6;
    end
    if (reset) begin
      image_2655 <= 4'h0;
    end else begin
      image_2655 <= 4'h6;
    end
    if (reset) begin
      image_2656 <= 4'h0;
    end else begin
      image_2656 <= 4'h4;
    end
    if (reset) begin
      image_2657 <= 4'h0;
    end else begin
      image_2657 <= 4'h4;
    end
    if (reset) begin
      image_2658 <= 4'h0;
    end else begin
      image_2658 <= 4'h6;
    end
    if (reset) begin
      image_2659 <= 4'h0;
    end else begin
      image_2659 <= 4'h6;
    end
    if (reset) begin
      image_2660 <= 4'h0;
    end else begin
      image_2660 <= 4'h6;
    end
    if (reset) begin
      image_2661 <= 4'h0;
    end else begin
      image_2661 <= 4'h6;
    end
    if (reset) begin
      image_2662 <= 4'h0;
    end else begin
      image_2662 <= 4'h5;
    end
    if (reset) begin
      image_2663 <= 4'h0;
    end else begin
      image_2663 <= 4'h4;
    end
    if (reset) begin
      image_2664 <= 4'h0;
    end else begin
      image_2664 <= 4'h4;
    end
    if (reset) begin
      image_2665 <= 4'h0;
    end else begin
      image_2665 <= 4'h5;
    end
    if (reset) begin
      image_2666 <= 4'h0;
    end else begin
      image_2666 <= 4'h5;
    end
    if (reset) begin
      image_2667 <= 4'h0;
    end else begin
      image_2667 <= 4'h6;
    end
    if (reset) begin
      image_2668 <= 4'h0;
    end else begin
      image_2668 <= 4'h6;
    end
    if (reset) begin
      image_2669 <= 4'h0;
    end else begin
      image_2669 <= 4'h6;
    end
    if (reset) begin
      image_2670 <= 4'h0;
    end else begin
      image_2670 <= 4'h6;
    end
    if (reset) begin
      image_2671 <= 4'h0;
    end else begin
      image_2671 <= 4'h6;
    end
    if (reset) begin
      image_2672 <= 4'h0;
    end else begin
      image_2672 <= 4'h6;
    end
    if (reset) begin
      image_2673 <= 4'h0;
    end else begin
      image_2673 <= 4'h5;
    end
    if (reset) begin
      image_2674 <= 4'h0;
    end else begin
      image_2674 <= 4'h5;
    end
    if (reset) begin
      image_2675 <= 4'h0;
    end else begin
      image_2675 <= 4'h4;
    end
    if (reset) begin
      image_2676 <= 4'h0;
    end else begin
      image_2676 <= 4'h4;
    end
    if (reset) begin
      image_2677 <= 4'h0;
    end else begin
      image_2677 <= 4'h5;
    end
    if (reset) begin
      image_2678 <= 4'h0;
    end else begin
      image_2678 <= 4'h6;
    end
    if (reset) begin
      image_2679 <= 4'h0;
    end else begin
      image_2679 <= 4'h6;
    end
    if (reset) begin
      image_2680 <= 4'h0;
    end else begin
      image_2680 <= 4'h6;
    end
    if (reset) begin
      image_2681 <= 4'h0;
    end else begin
      image_2681 <= 4'h5;
    end
    if (reset) begin
      image_2682 <= 4'h0;
    end else begin
      image_2682 <= 4'h1;
    end
    if (reset) begin
      image_2697 <= 4'h0;
    end else begin
      image_2697 <= 4'h2;
    end
    if (reset) begin
      image_2698 <= 4'h0;
    end else begin
      image_2698 <= 4'h4;
    end
    if (reset) begin
      image_2699 <= 4'h0;
    end else begin
      image_2699 <= 4'h5;
    end
    if (reset) begin
      image_2700 <= 4'h0;
    end else begin
      image_2700 <= 4'h5;
    end
    if (reset) begin
      image_2701 <= 4'h0;
    end else begin
      image_2701 <= 4'h5;
    end
    if (reset) begin
      image_2702 <= 4'h0;
    end else begin
      image_2702 <= 4'h5;
    end
    if (reset) begin
      image_2703 <= 4'h0;
    end else begin
      image_2703 <= 4'h5;
    end
    if (reset) begin
      image_2704 <= 4'h0;
    end else begin
      image_2704 <= 4'h6;
    end
    if (reset) begin
      image_2705 <= 4'h0;
    end else begin
      image_2705 <= 4'h6;
    end
    if (reset) begin
      image_2706 <= 4'h0;
    end else begin
      image_2706 <= 4'h6;
    end
    if (reset) begin
      image_2707 <= 4'h0;
    end else begin
      image_2707 <= 4'h6;
    end
    if (reset) begin
      image_2708 <= 4'h0;
    end else begin
      image_2708 <= 4'h6;
    end
    if (reset) begin
      image_2709 <= 4'h0;
    end else begin
      image_2709 <= 4'h6;
    end
    if (reset) begin
      image_2710 <= 4'h0;
    end else begin
      image_2710 <= 4'h6;
    end
    if (reset) begin
      image_2711 <= 4'h0;
    end else begin
      image_2711 <= 4'h6;
    end
    if (reset) begin
      image_2712 <= 4'h0;
    end else begin
      image_2712 <= 4'h6;
    end
    if (reset) begin
      image_2713 <= 4'h0;
    end else begin
      image_2713 <= 4'h6;
    end
    if (reset) begin
      image_2714 <= 4'h0;
    end else begin
      image_2714 <= 4'h6;
    end
    if (reset) begin
      image_2715 <= 4'h0;
    end else begin
      image_2715 <= 4'h6;
    end
    if (reset) begin
      image_2716 <= 4'h0;
    end else begin
      image_2716 <= 4'h6;
    end
    if (reset) begin
      image_2717 <= 4'h0;
    end else begin
      image_2717 <= 4'h6;
    end
    if (reset) begin
      image_2718 <= 4'h0;
    end else begin
      image_2718 <= 4'h6;
    end
    if (reset) begin
      image_2719 <= 4'h0;
    end else begin
      image_2719 <= 4'h6;
    end
    if (reset) begin
      image_2720 <= 4'h0;
    end else begin
      image_2720 <= 4'h6;
    end
    if (reset) begin
      image_2721 <= 4'h0;
    end else begin
      image_2721 <= 4'h6;
    end
    if (reset) begin
      image_2722 <= 4'h0;
    end else begin
      image_2722 <= 4'h4;
    end
    if (reset) begin
      image_2723 <= 4'h0;
    end else begin
      image_2723 <= 4'h4;
    end
    if (reset) begin
      image_2724 <= 4'h0;
    end else begin
      image_2724 <= 4'h5;
    end
    if (reset) begin
      image_2725 <= 4'h0;
    end else begin
      image_2725 <= 4'h6;
    end
    if (reset) begin
      image_2726 <= 4'h0;
    end else begin
      image_2726 <= 4'h6;
    end
    if (reset) begin
      image_2727 <= 4'h0;
    end else begin
      image_2727 <= 4'h6;
    end
    if (reset) begin
      image_2728 <= 4'h0;
    end else begin
      image_2728 <= 4'h6;
    end
    if (reset) begin
      image_2729 <= 4'h0;
    end else begin
      image_2729 <= 4'h6;
    end
    if (reset) begin
      image_2730 <= 4'h0;
    end else begin
      image_2730 <= 4'h5;
    end
    if (reset) begin
      image_2731 <= 4'h0;
    end else begin
      image_2731 <= 4'h5;
    end
    if (reset) begin
      image_2732 <= 4'h0;
    end else begin
      image_2732 <= 4'h4;
    end
    if (reset) begin
      image_2733 <= 4'h0;
    end else begin
      image_2733 <= 4'h4;
    end
    if (reset) begin
      image_2734 <= 4'h0;
    end else begin
      image_2734 <= 4'h4;
    end
    if (reset) begin
      image_2735 <= 4'h0;
    end else begin
      image_2735 <= 4'h5;
    end
    if (reset) begin
      image_2736 <= 4'h0;
    end else begin
      image_2736 <= 4'h5;
    end
    if (reset) begin
      image_2737 <= 4'h0;
    end else begin
      image_2737 <= 4'h5;
    end
    if (reset) begin
      image_2738 <= 4'h0;
    end else begin
      image_2738 <= 4'h6;
    end
    if (reset) begin
      image_2739 <= 4'h0;
    end else begin
      image_2739 <= 4'h6;
    end
    if (reset) begin
      image_2740 <= 4'h0;
    end else begin
      image_2740 <= 4'h6;
    end
    if (reset) begin
      image_2741 <= 4'h0;
    end else begin
      image_2741 <= 4'h6;
    end
    if (reset) begin
      image_2742 <= 4'h0;
    end else begin
      image_2742 <= 4'h6;
    end
    if (reset) begin
      image_2743 <= 4'h0;
    end else begin
      image_2743 <= 4'h6;
    end
    if (reset) begin
      image_2744 <= 4'h0;
    end else begin
      image_2744 <= 4'h6;
    end
    if (reset) begin
      image_2745 <= 4'h0;
    end else begin
      image_2745 <= 4'h4;
    end
    if (reset) begin
      image_2763 <= 4'h0;
    end else begin
      image_2763 <= 4'h3;
    end
    if (reset) begin
      image_2764 <= 4'h0;
    end else begin
      image_2764 <= 4'h5;
    end
    if (reset) begin
      image_2765 <= 4'h0;
    end else begin
      image_2765 <= 4'h5;
    end
    if (reset) begin
      image_2766 <= 4'h0;
    end else begin
      image_2766 <= 4'h5;
    end
    if (reset) begin
      image_2767 <= 4'h0;
    end else begin
      image_2767 <= 4'h5;
    end
    if (reset) begin
      image_2768 <= 4'h0;
    end else begin
      image_2768 <= 4'h5;
    end
    if (reset) begin
      image_2769 <= 4'h0;
    end else begin
      image_2769 <= 4'h5;
    end
    if (reset) begin
      image_2770 <= 4'h0;
    end else begin
      image_2770 <= 4'h6;
    end
    if (reset) begin
      image_2771 <= 4'h0;
    end else begin
      image_2771 <= 4'h6;
    end
    if (reset) begin
      image_2772 <= 4'h0;
    end else begin
      image_2772 <= 4'h6;
    end
    if (reset) begin
      image_2773 <= 4'h0;
    end else begin
      image_2773 <= 4'h6;
    end
    if (reset) begin
      image_2774 <= 4'h0;
    end else begin
      image_2774 <= 4'h6;
    end
    if (reset) begin
      image_2775 <= 4'h0;
    end else begin
      image_2775 <= 4'h6;
    end
    if (reset) begin
      image_2776 <= 4'h0;
    end else begin
      image_2776 <= 4'h6;
    end
    if (reset) begin
      image_2777 <= 4'h0;
    end else begin
      image_2777 <= 4'h6;
    end
    if (reset) begin
      image_2778 <= 4'h0;
    end else begin
      image_2778 <= 4'h6;
    end
    if (reset) begin
      image_2779 <= 4'h0;
    end else begin
      image_2779 <= 4'h6;
    end
    if (reset) begin
      image_2780 <= 4'h0;
    end else begin
      image_2780 <= 4'h6;
    end
    if (reset) begin
      image_2781 <= 4'h0;
    end else begin
      image_2781 <= 4'h6;
    end
    if (reset) begin
      image_2782 <= 4'h0;
    end else begin
      image_2782 <= 4'h6;
    end
    if (reset) begin
      image_2783 <= 4'h0;
    end else begin
      image_2783 <= 4'h6;
    end
    if (reset) begin
      image_2784 <= 4'h0;
    end else begin
      image_2784 <= 4'h6;
    end
    if (reset) begin
      image_2785 <= 4'h0;
    end else begin
      image_2785 <= 4'h6;
    end
    if (reset) begin
      image_2786 <= 4'h0;
    end else begin
      image_2786 <= 4'h6;
    end
    if (reset) begin
      image_2787 <= 4'h0;
    end else begin
      image_2787 <= 4'h6;
    end
    if (reset) begin
      image_2788 <= 4'h0;
    end else begin
      image_2788 <= 4'h5;
    end
    if (reset) begin
      image_2789 <= 4'h0;
    end else begin
      image_2789 <= 4'h4;
    end
    if (reset) begin
      image_2790 <= 4'h0;
    end else begin
      image_2790 <= 4'h4;
    end
    if (reset) begin
      image_2791 <= 4'h0;
    end else begin
      image_2791 <= 4'h5;
    end
    if (reset) begin
      image_2792 <= 4'h0;
    end else begin
      image_2792 <= 4'h6;
    end
    if (reset) begin
      image_2793 <= 4'h0;
    end else begin
      image_2793 <= 4'h6;
    end
    if (reset) begin
      image_2794 <= 4'h0;
    end else begin
      image_2794 <= 4'h6;
    end
    if (reset) begin
      image_2795 <= 4'h0;
    end else begin
      image_2795 <= 4'h6;
    end
    if (reset) begin
      image_2796 <= 4'h0;
    end else begin
      image_2796 <= 4'h6;
    end
    if (reset) begin
      image_2797 <= 4'h0;
    end else begin
      image_2797 <= 4'h6;
    end
    if (reset) begin
      image_2798 <= 4'h0;
    end else begin
      image_2798 <= 4'h6;
    end
    if (reset) begin
      image_2799 <= 4'h0;
    end else begin
      image_2799 <= 4'h6;
    end
    if (reset) begin
      image_2800 <= 4'h0;
    end else begin
      image_2800 <= 4'h6;
    end
    if (reset) begin
      image_2801 <= 4'h0;
    end else begin
      image_2801 <= 4'h6;
    end
    if (reset) begin
      image_2802 <= 4'h0;
    end else begin
      image_2802 <= 4'h6;
    end
    if (reset) begin
      image_2803 <= 4'h0;
    end else begin
      image_2803 <= 4'h6;
    end
    if (reset) begin
      image_2804 <= 4'h0;
    end else begin
      image_2804 <= 4'h6;
    end
    if (reset) begin
      image_2805 <= 4'h0;
    end else begin
      image_2805 <= 4'h5;
    end
    if (reset) begin
      image_2806 <= 4'h0;
    end else begin
      image_2806 <= 4'h5;
    end
    if (reset) begin
      image_2807 <= 4'h0;
    end else begin
      image_2807 <= 4'h4;
    end
    if (reset) begin
      image_2808 <= 4'h0;
    end else begin
      image_2808 <= 4'h2;
    end
    if (reset) begin
      image_2828 <= 4'h0;
    end else begin
      image_2828 <= 4'h1;
    end
    if (reset) begin
      image_2829 <= 4'h0;
    end else begin
      image_2829 <= 4'h3;
    end
    if (reset) begin
      image_2830 <= 4'h0;
    end else begin
      image_2830 <= 4'h4;
    end
    if (reset) begin
      image_2831 <= 4'h0;
    end else begin
      image_2831 <= 4'h5;
    end
    if (reset) begin
      image_2832 <= 4'h0;
    end else begin
      image_2832 <= 4'h5;
    end
    if (reset) begin
      image_2833 <= 4'h0;
    end else begin
      image_2833 <= 4'h5;
    end
    if (reset) begin
      image_2834 <= 4'h0;
    end else begin
      image_2834 <= 4'h5;
    end
    if (reset) begin
      image_2835 <= 4'h0;
    end else begin
      image_2835 <= 4'h5;
    end
    if (reset) begin
      image_2836 <= 4'h0;
    end else begin
      image_2836 <= 4'h6;
    end
    if (reset) begin
      image_2837 <= 4'h0;
    end else begin
      image_2837 <= 4'h6;
    end
    if (reset) begin
      image_2838 <= 4'h0;
    end else begin
      image_2838 <= 4'h6;
    end
    if (reset) begin
      image_2839 <= 4'h0;
    end else begin
      image_2839 <= 4'h6;
    end
    if (reset) begin
      image_2840 <= 4'h0;
    end else begin
      image_2840 <= 4'h6;
    end
    if (reset) begin
      image_2841 <= 4'h0;
    end else begin
      image_2841 <= 4'h6;
    end
    if (reset) begin
      image_2842 <= 4'h0;
    end else begin
      image_2842 <= 4'h6;
    end
    if (reset) begin
      image_2843 <= 4'h0;
    end else begin
      image_2843 <= 4'h6;
    end
    if (reset) begin
      image_2844 <= 4'h0;
    end else begin
      image_2844 <= 4'h6;
    end
    if (reset) begin
      image_2845 <= 4'h0;
    end else begin
      image_2845 <= 4'h6;
    end
    if (reset) begin
      image_2846 <= 4'h0;
    end else begin
      image_2846 <= 4'h6;
    end
    if (reset) begin
      image_2847 <= 4'h0;
    end else begin
      image_2847 <= 4'h6;
    end
    if (reset) begin
      image_2848 <= 4'h0;
    end else begin
      image_2848 <= 4'h6;
    end
    if (reset) begin
      image_2849 <= 4'h0;
    end else begin
      image_2849 <= 4'h6;
    end
    if (reset) begin
      image_2850 <= 4'h0;
    end else begin
      image_2850 <= 4'h6;
    end
    if (reset) begin
      image_2851 <= 4'h0;
    end else begin
      image_2851 <= 4'h6;
    end
    if (reset) begin
      image_2852 <= 4'h0;
    end else begin
      image_2852 <= 4'h6;
    end
    if (reset) begin
      image_2853 <= 4'h0;
    end else begin
      image_2853 <= 4'h6;
    end
    if (reset) begin
      image_2854 <= 4'h0;
    end else begin
      image_2854 <= 4'h6;
    end
    if (reset) begin
      image_2855 <= 4'h0;
    end else begin
      image_2855 <= 4'h5;
    end
    if (reset) begin
      image_2856 <= 4'h0;
    end else begin
      image_2856 <= 4'h4;
    end
    if (reset) begin
      image_2857 <= 4'h0;
    end else begin
      image_2857 <= 4'h4;
    end
    if (reset) begin
      image_2858 <= 4'h0;
    end else begin
      image_2858 <= 4'h4;
    end
    if (reset) begin
      image_2859 <= 4'h0;
    end else begin
      image_2859 <= 4'h4;
    end
    if (reset) begin
      image_2860 <= 4'h0;
    end else begin
      image_2860 <= 4'h4;
    end
    if (reset) begin
      image_2861 <= 4'h0;
    end else begin
      image_2861 <= 4'h4;
    end
    if (reset) begin
      image_2862 <= 4'h0;
    end else begin
      image_2862 <= 4'h4;
    end
    if (reset) begin
      image_2863 <= 4'h0;
    end else begin
      image_2863 <= 4'h4;
    end
    if (reset) begin
      image_2864 <= 4'h0;
    end else begin
      image_2864 <= 4'h4;
    end
    if (reset) begin
      image_2865 <= 4'h0;
    end else begin
      image_2865 <= 4'h4;
    end
    if (reset) begin
      image_2866 <= 4'h0;
    end else begin
      image_2866 <= 4'h4;
    end
    if (reset) begin
      image_2867 <= 4'h0;
    end else begin
      image_2867 <= 4'h4;
    end
    if (reset) begin
      image_2868 <= 4'h0;
    end else begin
      image_2868 <= 4'h5;
    end
    if (reset) begin
      image_2869 <= 4'h0;
    end else begin
      image_2869 <= 4'h5;
    end
    if (reset) begin
      image_2870 <= 4'h0;
    end else begin
      image_2870 <= 4'h5;
    end
    if (reset) begin
      image_2871 <= 4'h0;
    end else begin
      image_2871 <= 4'h3;
    end
    if (reset) begin
      image_2895 <= 4'h0;
    end else begin
      image_2895 <= 4'h1;
    end
    if (reset) begin
      image_2896 <= 4'h0;
    end else begin
      image_2896 <= 4'h3;
    end
    if (reset) begin
      image_2897 <= 4'h0;
    end else begin
      image_2897 <= 4'h4;
    end
    if (reset) begin
      image_2898 <= 4'h0;
    end else begin
      image_2898 <= 4'h4;
    end
    if (reset) begin
      image_2899 <= 4'h0;
    end else begin
      image_2899 <= 4'h4;
    end
    if (reset) begin
      image_2900 <= 4'h0;
    end else begin
      image_2900 <= 4'h5;
    end
    if (reset) begin
      image_2901 <= 4'h0;
    end else begin
      image_2901 <= 4'h5;
    end
    if (reset) begin
      image_2902 <= 4'h0;
    end else begin
      image_2902 <= 4'h6;
    end
    if (reset) begin
      image_2903 <= 4'h0;
    end else begin
      image_2903 <= 4'h6;
    end
    if (reset) begin
      image_2904 <= 4'h0;
    end else begin
      image_2904 <= 4'h6;
    end
    if (reset) begin
      image_2905 <= 4'h0;
    end else begin
      image_2905 <= 4'h6;
    end
    if (reset) begin
      image_2906 <= 4'h0;
    end else begin
      image_2906 <= 4'h6;
    end
    if (reset) begin
      image_2907 <= 4'h0;
    end else begin
      image_2907 <= 4'h6;
    end
    if (reset) begin
      image_2908 <= 4'h0;
    end else begin
      image_2908 <= 4'h6;
    end
    if (reset) begin
      image_2909 <= 4'h0;
    end else begin
      image_2909 <= 4'h6;
    end
    if (reset) begin
      image_2910 <= 4'h0;
    end else begin
      image_2910 <= 4'h6;
    end
    if (reset) begin
      image_2911 <= 4'h0;
    end else begin
      image_2911 <= 4'h6;
    end
    if (reset) begin
      image_2912 <= 4'h0;
    end else begin
      image_2912 <= 4'h6;
    end
    if (reset) begin
      image_2913 <= 4'h0;
    end else begin
      image_2913 <= 4'h6;
    end
    if (reset) begin
      image_2914 <= 4'h0;
    end else begin
      image_2914 <= 4'h6;
    end
    if (reset) begin
      image_2915 <= 4'h0;
    end else begin
      image_2915 <= 4'h6;
    end
    if (reset) begin
      image_2916 <= 4'h0;
    end else begin
      image_2916 <= 4'h6;
    end
    if (reset) begin
      image_2917 <= 4'h0;
    end else begin
      image_2917 <= 4'h6;
    end
    if (reset) begin
      image_2918 <= 4'h0;
    end else begin
      image_2918 <= 4'h6;
    end
    if (reset) begin
      image_2919 <= 4'h0;
    end else begin
      image_2919 <= 4'h6;
    end
    if (reset) begin
      image_2920 <= 4'h0;
    end else begin
      image_2920 <= 4'h6;
    end
    if (reset) begin
      image_2921 <= 4'h0;
    end else begin
      image_2921 <= 4'h6;
    end
    if (reset) begin
      image_2922 <= 4'h0;
    end else begin
      image_2922 <= 4'h6;
    end
    if (reset) begin
      image_2923 <= 4'h0;
    end else begin
      image_2923 <= 4'h6;
    end
    if (reset) begin
      image_2924 <= 4'h0;
    end else begin
      image_2924 <= 4'h6;
    end
    if (reset) begin
      image_2925 <= 4'h0;
    end else begin
      image_2925 <= 4'h6;
    end
    if (reset) begin
      image_2926 <= 4'h0;
    end else begin
      image_2926 <= 4'h6;
    end
    if (reset) begin
      image_2927 <= 4'h0;
    end else begin
      image_2927 <= 4'h6;
    end
    if (reset) begin
      image_2928 <= 4'h0;
    end else begin
      image_2928 <= 4'h6;
    end
    if (reset) begin
      image_2929 <= 4'h0;
    end else begin
      image_2929 <= 4'h6;
    end
    if (reset) begin
      image_2930 <= 4'h0;
    end else begin
      image_2930 <= 4'h6;
    end
    if (reset) begin
      image_2931 <= 4'h0;
    end else begin
      image_2931 <= 4'h6;
    end
    if (reset) begin
      image_2932 <= 4'h0;
    end else begin
      image_2932 <= 4'h6;
    end
    if (reset) begin
      image_2933 <= 4'h0;
    end else begin
      image_2933 <= 4'h4;
    end
    if (reset) begin
      image_2934 <= 4'h0;
    end else begin
      image_2934 <= 4'h2;
    end
    if (reset) begin
      image_2965 <= 4'h0;
    end else begin
      image_2965 <= 4'h2;
    end
    if (reset) begin
      image_2966 <= 4'h0;
    end else begin
      image_2966 <= 4'h3;
    end
    if (reset) begin
      image_2967 <= 4'h0;
    end else begin
      image_2967 <= 4'h4;
    end
    if (reset) begin
      image_2968 <= 4'h0;
    end else begin
      image_2968 <= 4'h4;
    end
    if (reset) begin
      image_2969 <= 4'h0;
    end else begin
      image_2969 <= 4'h5;
    end
    if (reset) begin
      image_2970 <= 4'h0;
    end else begin
      image_2970 <= 4'h6;
    end
    if (reset) begin
      image_2971 <= 4'h0;
    end else begin
      image_2971 <= 4'h6;
    end
    if (reset) begin
      image_2972 <= 4'h0;
    end else begin
      image_2972 <= 4'h6;
    end
    if (reset) begin
      image_2973 <= 4'h0;
    end else begin
      image_2973 <= 4'h6;
    end
    if (reset) begin
      image_2974 <= 4'h0;
    end else begin
      image_2974 <= 4'h6;
    end
    if (reset) begin
      image_2975 <= 4'h0;
    end else begin
      image_2975 <= 4'h6;
    end
    if (reset) begin
      image_2976 <= 4'h0;
    end else begin
      image_2976 <= 4'h6;
    end
    if (reset) begin
      image_2977 <= 4'h0;
    end else begin
      image_2977 <= 4'h6;
    end
    if (reset) begin
      image_2978 <= 4'h0;
    end else begin
      image_2978 <= 4'h6;
    end
    if (reset) begin
      image_2979 <= 4'h0;
    end else begin
      image_2979 <= 4'h6;
    end
    if (reset) begin
      image_2980 <= 4'h0;
    end else begin
      image_2980 <= 4'h6;
    end
    if (reset) begin
      image_2981 <= 4'h0;
    end else begin
      image_2981 <= 4'h6;
    end
    if (reset) begin
      image_2982 <= 4'h0;
    end else begin
      image_2982 <= 4'h6;
    end
    if (reset) begin
      image_2983 <= 4'h0;
    end else begin
      image_2983 <= 4'h6;
    end
    if (reset) begin
      image_2984 <= 4'h0;
    end else begin
      image_2984 <= 4'h6;
    end
    if (reset) begin
      image_2985 <= 4'h0;
    end else begin
      image_2985 <= 4'h6;
    end
    if (reset) begin
      image_2986 <= 4'h0;
    end else begin
      image_2986 <= 4'h6;
    end
    if (reset) begin
      image_2987 <= 4'h0;
    end else begin
      image_2987 <= 4'h6;
    end
    if (reset) begin
      image_2988 <= 4'h0;
    end else begin
      image_2988 <= 4'h6;
    end
    if (reset) begin
      image_2989 <= 4'h0;
    end else begin
      image_2989 <= 4'h6;
    end
    if (reset) begin
      image_2990 <= 4'h0;
    end else begin
      image_2990 <= 4'h6;
    end
    if (reset) begin
      image_2991 <= 4'h0;
    end else begin
      image_2991 <= 4'h6;
    end
    if (reset) begin
      image_2992 <= 4'h0;
    end else begin
      image_2992 <= 4'h6;
    end
    if (reset) begin
      image_2993 <= 4'h0;
    end else begin
      image_2993 <= 4'h5;
    end
    if (reset) begin
      image_2994 <= 4'h0;
    end else begin
      image_2994 <= 4'h5;
    end
    if (reset) begin
      image_2995 <= 4'h0;
    end else begin
      image_2995 <= 4'h4;
    end
    if (reset) begin
      image_2996 <= 4'h0;
    end else begin
      image_2996 <= 4'h2;
    end
    if (reset) begin
      image_3035 <= 4'h0;
    end else begin
      image_3035 <= 4'h1;
    end
    if (reset) begin
      image_3036 <= 4'h0;
    end else begin
      image_3036 <= 4'h2;
    end
    if (reset) begin
      image_3037 <= 4'h0;
    end else begin
      image_3037 <= 4'h3;
    end
    if (reset) begin
      image_3038 <= 4'h0;
    end else begin
      image_3038 <= 4'h4;
    end
    if (reset) begin
      image_3039 <= 4'h0;
    end else begin
      image_3039 <= 4'h4;
    end
    if (reset) begin
      image_3040 <= 4'h0;
    end else begin
      image_3040 <= 4'h4;
    end
    if (reset) begin
      image_3041 <= 4'h0;
    end else begin
      image_3041 <= 4'h5;
    end
    if (reset) begin
      image_3042 <= 4'h0;
    end else begin
      image_3042 <= 4'h5;
    end
    if (reset) begin
      image_3043 <= 4'h0;
    end else begin
      image_3043 <= 4'h5;
    end
    if (reset) begin
      image_3044 <= 4'h0;
    end else begin
      image_3044 <= 4'h5;
    end
    if (reset) begin
      image_3045 <= 4'h0;
    end else begin
      image_3045 <= 4'h5;
    end
    if (reset) begin
      image_3046 <= 4'h0;
    end else begin
      image_3046 <= 4'h5;
    end
    if (reset) begin
      image_3047 <= 4'h0;
    end else begin
      image_3047 <= 4'h5;
    end
    if (reset) begin
      image_3048 <= 4'h0;
    end else begin
      image_3048 <= 4'h5;
    end
    if (reset) begin
      image_3049 <= 4'h0;
    end else begin
      image_3049 <= 4'h5;
    end
    if (reset) begin
      image_3050 <= 4'h0;
    end else begin
      image_3050 <= 4'h5;
    end
    if (reset) begin
      image_3051 <= 4'h0;
    end else begin
      image_3051 <= 4'h5;
    end
    if (reset) begin
      image_3052 <= 4'h0;
    end else begin
      image_3052 <= 4'h5;
    end
    if (reset) begin
      image_3053 <= 4'h0;
    end else begin
      image_3053 <= 4'h4;
    end
    if (reset) begin
      image_3054 <= 4'h0;
    end else begin
      image_3054 <= 4'h4;
    end
    if (reset) begin
      image_3055 <= 4'h0;
    end else begin
      image_3055 <= 4'h2;
    end
    if (reset) begin
      image_3056 <= 4'h0;
    end else begin
      image_3056 <= 4'h1;
    end
    if (reset) begin
      kernelCounter <= 4'h0;
    end else if (kernelCountReset) begin
      kernelCounter <= 4'h0;
    end else begin
      kernelCounter <= _T_15;
    end
    if (reset) begin
      imageCounterX <= 2'h0;
    end else if (imageCounterXReset) begin
      imageCounterX <= 2'h0;
    end else begin
      imageCounterX <= _T_19;
    end
    if (reset) begin
      imageCounterY <= 2'h0;
    end else if (imageCounterXReset) begin
      if (_T_20) begin
        imageCounterY <= 2'h0;
      end else begin
        imageCounterY <= _T_22;
      end
    end
    if (reset) begin
      pixelIndex <= 32'h0;
    end else if (kernelCountReset) begin
      if (_T_282) begin
        pixelIndex <= 32'h0;
      end else begin
        pixelIndex <= _T_280;
      end
    end
  end
endmodule
