module VideoBuffer(
  input         clock,
  input         reset,
  input  [3:0]  io_pixelVal_in_0,
  input  [3:0]  io_pixelVal_in_1,
  input  [3:0]  io_pixelVal_in_2,
  input  [3:0]  io_pixelVal_in_3,
  input  [3:0]  io_pixelVal_in_4,
  input  [3:0]  io_pixelVal_in_5,
  input  [3:0]  io_pixelVal_in_6,
  input  [3:0]  io_pixelVal_in_7,
  input         io_valid_in,
  input  [10:0] io_rowIndex,
  input  [10:0] io_colIndex,
  output [3:0]  io_pixelVal_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] _T = io_rowIndex * 11'h10; // @[VideoBuffer.scala 29:46]
  wire [15:0] _GEN_1922 = {{5'd0}, io_colIndex}; // @[VideoBuffer.scala 29:61]
  wire [15:0] _T_2 = _T + _GEN_1922; // @[VideoBuffer.scala 29:61]
  reg [31:0] pixelIndex; // @[VideoBuffer.scala 31:33]
  wire [31:0] _T_26 = pixelIndex + 32'h7; // @[VideoBuffer.scala 35:42]
  wire [31:0] _T_23 = pixelIndex + 32'h6; // @[VideoBuffer.scala 35:42]
  wire [31:0] _T_20 = pixelIndex + 32'h5; // @[VideoBuffer.scala 35:42]
  wire [31:0] _T_17 = pixelIndex + 32'h4; // @[VideoBuffer.scala 35:42]
  wire [31:0] _T_14 = pixelIndex + 32'h3; // @[VideoBuffer.scala 35:42]
  wire [31:0] _T_11 = pixelIndex + 32'h2; // @[VideoBuffer.scala 35:42]
  wire [31:0] _T_8 = pixelIndex + 32'h1; // @[VideoBuffer.scala 35:42]
  wire [32:0] _T_4 = {{1'd0}, pixelIndex}; // @[VideoBuffer.scala 35:42]
  wire [3:0] _GEN_192 = 8'h0 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_384 = 8'h0 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_192; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_576 = 8'h0 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_384; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_768 = 8'h0 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_576; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_960 = 8'h0 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_768; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1152 = 8'h0 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_960; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1344 = 8'h0 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1152; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1536 = 8'h0 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1344; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_0 = io_valid_in ? _GEN_1536 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_193 = 8'h1 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_385 = 8'h1 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_193; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_577 = 8'h1 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_385; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_769 = 8'h1 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_577; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_961 = 8'h1 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_769; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1153 = 8'h1 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_961; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1345 = 8'h1 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1153; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1537 = 8'h1 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1345; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1 = io_valid_in ? _GEN_1537 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1 = 8'h1 == _T_2[7:0] ? image_1 : image_0; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_194 = 8'h2 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_386 = 8'h2 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_194; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_578 = 8'h2 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_386; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_770 = 8'h2 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_578; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_962 = 8'h2 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_770; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1154 = 8'h2 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_962; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1346 = 8'h2 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1154; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1538 = 8'h2 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1346; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2 = io_valid_in ? _GEN_1538 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2 = 8'h2 == _T_2[7:0] ? image_2 : _GEN_1; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_195 = 8'h3 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_387 = 8'h3 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_195; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_579 = 8'h3 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_387; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_771 = 8'h3 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_579; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_963 = 8'h3 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_771; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1155 = 8'h3 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_963; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1347 = 8'h3 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1155; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1539 = 8'h3 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1347; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3 = io_valid_in ? _GEN_1539 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3 = 8'h3 == _T_2[7:0] ? image_3 : _GEN_2; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_196 = 8'h4 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_388 = 8'h4 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_196; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_580 = 8'h4 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_388; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_772 = 8'h4 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_580; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_964 = 8'h4 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_772; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1156 = 8'h4 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_964; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1348 = 8'h4 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1156; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1540 = 8'h4 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1348; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_4 = io_valid_in ? _GEN_1540 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_4 = 8'h4 == _T_2[7:0] ? image_4 : _GEN_3; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_197 = 8'h5 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_389 = 8'h5 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_197; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_581 = 8'h5 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_389; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_773 = 8'h5 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_581; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_965 = 8'h5 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_773; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1157 = 8'h5 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_965; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1349 = 8'h5 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1157; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1541 = 8'h5 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1349; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_5 = io_valid_in ? _GEN_1541 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_5 = 8'h5 == _T_2[7:0] ? image_5 : _GEN_4; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_198 = 8'h6 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_390 = 8'h6 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_198; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_582 = 8'h6 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_390; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_774 = 8'h6 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_582; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_966 = 8'h6 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_774; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1158 = 8'h6 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_966; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1350 = 8'h6 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1158; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1542 = 8'h6 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1350; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_6 = io_valid_in ? _GEN_1542 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_6 = 8'h6 == _T_2[7:0] ? image_6 : _GEN_5; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_199 = 8'h7 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_391 = 8'h7 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_199; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_583 = 8'h7 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_391; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_775 = 8'h7 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_583; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_967 = 8'h7 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_775; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1159 = 8'h7 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_967; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1351 = 8'h7 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1159; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1543 = 8'h7 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1351; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_7 = io_valid_in ? _GEN_1543 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_7 = 8'h7 == _T_2[7:0] ? image_7 : _GEN_6; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_200 = 8'h8 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_392 = 8'h8 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_200; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_584 = 8'h8 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_392; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_776 = 8'h8 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_584; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_968 = 8'h8 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_776; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1160 = 8'h8 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_968; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1352 = 8'h8 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1160; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1544 = 8'h8 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1352; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_8 = io_valid_in ? _GEN_1544 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_8 = 8'h8 == _T_2[7:0] ? image_8 : _GEN_7; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_201 = 8'h9 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_393 = 8'h9 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_201; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_585 = 8'h9 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_393; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_777 = 8'h9 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_585; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_969 = 8'h9 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_777; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1161 = 8'h9 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_969; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1353 = 8'h9 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1161; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1545 = 8'h9 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1353; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_9 = io_valid_in ? _GEN_1545 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_9 = 8'h9 == _T_2[7:0] ? image_9 : _GEN_8; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_202 = 8'ha == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_394 = 8'ha == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_202; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_586 = 8'ha == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_394; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_778 = 8'ha == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_586; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_970 = 8'ha == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_778; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1162 = 8'ha == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_970; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1354 = 8'ha == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1162; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1546 = 8'ha == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1354; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_10 = io_valid_in ? _GEN_1546 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_10 = 8'ha == _T_2[7:0] ? image_10 : _GEN_9; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_203 = 8'hb == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_395 = 8'hb == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_203; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_587 = 8'hb == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_395; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_779 = 8'hb == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_587; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_971 = 8'hb == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_779; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1163 = 8'hb == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_971; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1355 = 8'hb == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1163; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1547 = 8'hb == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1355; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_11 = io_valid_in ? _GEN_1547 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_11 = 8'hb == _T_2[7:0] ? image_11 : _GEN_10; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_204 = 8'hc == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_396 = 8'hc == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_204; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_588 = 8'hc == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_396; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_780 = 8'hc == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_588; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_972 = 8'hc == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_780; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1164 = 8'hc == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_972; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1356 = 8'hc == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1164; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1548 = 8'hc == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1356; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_12 = io_valid_in ? _GEN_1548 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_12 = 8'hc == _T_2[7:0] ? image_12 : _GEN_11; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_205 = 8'hd == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_397 = 8'hd == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_205; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_589 = 8'hd == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_397; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_781 = 8'hd == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_589; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_973 = 8'hd == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_781; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1165 = 8'hd == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_973; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1357 = 8'hd == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1165; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1549 = 8'hd == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1357; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_13 = io_valid_in ? _GEN_1549 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_13 = 8'hd == _T_2[7:0] ? image_13 : _GEN_12; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_206 = 8'he == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_398 = 8'he == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_206; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_590 = 8'he == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_398; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_782 = 8'he == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_590; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_974 = 8'he == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_782; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1166 = 8'he == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_974; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1358 = 8'he == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1166; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1550 = 8'he == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1358; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_14 = io_valid_in ? _GEN_1550 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_14 = 8'he == _T_2[7:0] ? image_14 : _GEN_13; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_207 = 8'hf == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_399 = 8'hf == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_207; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_591 = 8'hf == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_399; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_783 = 8'hf == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_591; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_975 = 8'hf == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_783; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1167 = 8'hf == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_975; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1359 = 8'hf == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1167; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1551 = 8'hf == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1359; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_15 = io_valid_in ? _GEN_1551 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_15 = 8'hf == _T_2[7:0] ? image_15 : _GEN_14; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_208 = 8'h10 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_400 = 8'h10 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_208; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_592 = 8'h10 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_400; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_784 = 8'h10 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_592; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_976 = 8'h10 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_784; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1168 = 8'h10 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_976; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1360 = 8'h10 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1168; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1552 = 8'h10 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1360; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_16 = io_valid_in ? _GEN_1552 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_16 = 8'h10 == _T_2[7:0] ? image_16 : _GEN_15; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_209 = 8'h11 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_401 = 8'h11 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_209; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_593 = 8'h11 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_401; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_785 = 8'h11 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_593; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_977 = 8'h11 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_785; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1169 = 8'h11 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_977; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1361 = 8'h11 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1169; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1553 = 8'h11 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1361; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_17 = io_valid_in ? _GEN_1553 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_17 = 8'h11 == _T_2[7:0] ? image_17 : _GEN_16; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_210 = 8'h12 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_402 = 8'h12 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_210; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_594 = 8'h12 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_402; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_786 = 8'h12 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_594; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_978 = 8'h12 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_786; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1170 = 8'h12 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_978; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1362 = 8'h12 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1170; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1554 = 8'h12 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1362; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_18 = io_valid_in ? _GEN_1554 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_18 = 8'h12 == _T_2[7:0] ? image_18 : _GEN_17; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_211 = 8'h13 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_403 = 8'h13 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_211; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_595 = 8'h13 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_403; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_787 = 8'h13 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_595; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_979 = 8'h13 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_787; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1171 = 8'h13 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_979; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1363 = 8'h13 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1171; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1555 = 8'h13 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1363; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_19 = io_valid_in ? _GEN_1555 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_19 = 8'h13 == _T_2[7:0] ? image_19 : _GEN_18; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_212 = 8'h14 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_404 = 8'h14 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_212; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_596 = 8'h14 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_404; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_788 = 8'h14 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_596; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_980 = 8'h14 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_788; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1172 = 8'h14 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_980; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1364 = 8'h14 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1172; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1556 = 8'h14 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1364; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_20 = io_valid_in ? _GEN_1556 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_20 = 8'h14 == _T_2[7:0] ? image_20 : _GEN_19; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_213 = 8'h15 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_405 = 8'h15 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_213; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_597 = 8'h15 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_405; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_789 = 8'h15 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_597; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_981 = 8'h15 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_789; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1173 = 8'h15 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_981; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1365 = 8'h15 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1173; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1557 = 8'h15 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1365; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_21 = io_valid_in ? _GEN_1557 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_21 = 8'h15 == _T_2[7:0] ? image_21 : _GEN_20; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_214 = 8'h16 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_406 = 8'h16 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_214; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_598 = 8'h16 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_406; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_790 = 8'h16 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_598; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_982 = 8'h16 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_790; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1174 = 8'h16 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_982; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1366 = 8'h16 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1174; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1558 = 8'h16 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1366; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_22 = io_valid_in ? _GEN_1558 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_22 = 8'h16 == _T_2[7:0] ? image_22 : _GEN_21; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_215 = 8'h17 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_407 = 8'h17 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_215; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_599 = 8'h17 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_407; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_791 = 8'h17 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_599; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_983 = 8'h17 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_791; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1175 = 8'h17 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_983; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1367 = 8'h17 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1175; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1559 = 8'h17 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1367; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_23 = io_valid_in ? _GEN_1559 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_23 = 8'h17 == _T_2[7:0] ? image_23 : _GEN_22; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_216 = 8'h18 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_408 = 8'h18 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_216; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_600 = 8'h18 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_408; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_792 = 8'h18 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_600; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_984 = 8'h18 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_792; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1176 = 8'h18 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_984; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1368 = 8'h18 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1176; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1560 = 8'h18 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1368; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_24 = io_valid_in ? _GEN_1560 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_24 = 8'h18 == _T_2[7:0] ? image_24 : _GEN_23; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_217 = 8'h19 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_409 = 8'h19 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_217; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_601 = 8'h19 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_409; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_793 = 8'h19 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_601; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_985 = 8'h19 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_793; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1177 = 8'h19 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_985; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1369 = 8'h19 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1177; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1561 = 8'h19 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1369; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_25 = io_valid_in ? _GEN_1561 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_25 = 8'h19 == _T_2[7:0] ? image_25 : _GEN_24; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_218 = 8'h1a == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_410 = 8'h1a == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_218; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_602 = 8'h1a == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_410; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_794 = 8'h1a == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_602; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_986 = 8'h1a == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_794; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1178 = 8'h1a == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_986; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1370 = 8'h1a == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1178; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1562 = 8'h1a == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1370; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_26 = io_valid_in ? _GEN_1562 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_26 = 8'h1a == _T_2[7:0] ? image_26 : _GEN_25; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_219 = 8'h1b == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_411 = 8'h1b == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_219; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_603 = 8'h1b == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_411; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_795 = 8'h1b == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_603; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_987 = 8'h1b == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_795; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1179 = 8'h1b == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_987; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1371 = 8'h1b == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1179; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1563 = 8'h1b == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1371; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_27 = io_valid_in ? _GEN_1563 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_27 = 8'h1b == _T_2[7:0] ? image_27 : _GEN_26; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_220 = 8'h1c == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_412 = 8'h1c == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_220; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_604 = 8'h1c == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_412; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_796 = 8'h1c == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_604; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_988 = 8'h1c == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_796; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1180 = 8'h1c == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_988; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1372 = 8'h1c == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1180; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1564 = 8'h1c == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1372; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_28 = io_valid_in ? _GEN_1564 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_28 = 8'h1c == _T_2[7:0] ? image_28 : _GEN_27; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_221 = 8'h1d == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_413 = 8'h1d == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_221; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_605 = 8'h1d == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_413; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_797 = 8'h1d == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_605; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_989 = 8'h1d == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_797; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1181 = 8'h1d == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_989; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1373 = 8'h1d == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1181; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1565 = 8'h1d == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1373; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_29 = io_valid_in ? _GEN_1565 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_29 = 8'h1d == _T_2[7:0] ? image_29 : _GEN_28; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_222 = 8'h1e == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_414 = 8'h1e == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_222; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_606 = 8'h1e == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_414; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_798 = 8'h1e == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_606; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_990 = 8'h1e == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_798; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1182 = 8'h1e == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_990; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1374 = 8'h1e == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1182; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1566 = 8'h1e == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1374; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_30 = io_valid_in ? _GEN_1566 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_30 = 8'h1e == _T_2[7:0] ? image_30 : _GEN_29; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_223 = 8'h1f == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_415 = 8'h1f == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_223; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_607 = 8'h1f == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_415; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_799 = 8'h1f == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_607; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_991 = 8'h1f == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_799; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1183 = 8'h1f == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_991; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1375 = 8'h1f == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1183; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1567 = 8'h1f == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1375; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_31 = io_valid_in ? _GEN_1567 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_31 = 8'h1f == _T_2[7:0] ? image_31 : _GEN_30; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_224 = 8'h20 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_416 = 8'h20 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_224; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_608 = 8'h20 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_416; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_800 = 8'h20 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_608; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_992 = 8'h20 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_800; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1184 = 8'h20 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_992; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1376 = 8'h20 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1184; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1568 = 8'h20 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1376; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_32 = io_valid_in ? _GEN_1568 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_32 = 8'h20 == _T_2[7:0] ? image_32 : _GEN_31; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_225 = 8'h21 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_417 = 8'h21 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_225; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_609 = 8'h21 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_417; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_801 = 8'h21 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_609; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_993 = 8'h21 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_801; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1185 = 8'h21 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_993; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1377 = 8'h21 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1185; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1569 = 8'h21 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1377; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_33 = io_valid_in ? _GEN_1569 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_33 = 8'h21 == _T_2[7:0] ? image_33 : _GEN_32; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_226 = 8'h22 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_418 = 8'h22 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_226; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_610 = 8'h22 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_418; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_802 = 8'h22 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_610; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_994 = 8'h22 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_802; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1186 = 8'h22 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_994; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1378 = 8'h22 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1186; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1570 = 8'h22 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1378; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_34 = io_valid_in ? _GEN_1570 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_34 = 8'h22 == _T_2[7:0] ? image_34 : _GEN_33; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_227 = 8'h23 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_419 = 8'h23 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_227; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_611 = 8'h23 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_419; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_803 = 8'h23 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_611; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_995 = 8'h23 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_803; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1187 = 8'h23 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_995; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1379 = 8'h23 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1187; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1571 = 8'h23 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1379; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_35 = io_valid_in ? _GEN_1571 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_35 = 8'h23 == _T_2[7:0] ? image_35 : _GEN_34; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_228 = 8'h24 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_420 = 8'h24 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_228; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_612 = 8'h24 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_420; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_804 = 8'h24 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_612; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_996 = 8'h24 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_804; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1188 = 8'h24 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_996; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1380 = 8'h24 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1188; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1572 = 8'h24 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1380; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_36 = io_valid_in ? _GEN_1572 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_36 = 8'h24 == _T_2[7:0] ? image_36 : _GEN_35; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_229 = 8'h25 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_421 = 8'h25 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_229; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_613 = 8'h25 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_421; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_805 = 8'h25 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_613; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_997 = 8'h25 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_805; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1189 = 8'h25 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_997; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1381 = 8'h25 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1189; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1573 = 8'h25 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1381; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_37 = io_valid_in ? _GEN_1573 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_37 = 8'h25 == _T_2[7:0] ? image_37 : _GEN_36; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_230 = 8'h26 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_422 = 8'h26 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_230; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_614 = 8'h26 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_422; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_806 = 8'h26 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_614; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_998 = 8'h26 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_806; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1190 = 8'h26 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_998; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1382 = 8'h26 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1190; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1574 = 8'h26 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1382; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_38 = io_valid_in ? _GEN_1574 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_38 = 8'h26 == _T_2[7:0] ? image_38 : _GEN_37; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_231 = 8'h27 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_423 = 8'h27 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_231; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_615 = 8'h27 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_423; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_807 = 8'h27 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_615; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_999 = 8'h27 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_807; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1191 = 8'h27 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_999; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1383 = 8'h27 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1191; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1575 = 8'h27 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1383; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_39 = io_valid_in ? _GEN_1575 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_39 = 8'h27 == _T_2[7:0] ? image_39 : _GEN_38; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_232 = 8'h28 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_424 = 8'h28 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_232; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_616 = 8'h28 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_424; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_808 = 8'h28 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_616; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1000 = 8'h28 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_808; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1192 = 8'h28 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1000; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1384 = 8'h28 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1192; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1576 = 8'h28 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1384; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_40 = io_valid_in ? _GEN_1576 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_40 = 8'h28 == _T_2[7:0] ? image_40 : _GEN_39; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_233 = 8'h29 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_425 = 8'h29 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_233; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_617 = 8'h29 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_425; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_809 = 8'h29 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_617; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1001 = 8'h29 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_809; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1193 = 8'h29 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1001; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1385 = 8'h29 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1193; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1577 = 8'h29 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1385; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_41 = io_valid_in ? _GEN_1577 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_41 = 8'h29 == _T_2[7:0] ? image_41 : _GEN_40; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_234 = 8'h2a == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_426 = 8'h2a == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_234; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_618 = 8'h2a == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_426; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_810 = 8'h2a == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_618; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1002 = 8'h2a == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_810; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1194 = 8'h2a == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1002; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1386 = 8'h2a == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1194; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1578 = 8'h2a == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1386; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_42 = io_valid_in ? _GEN_1578 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_42 = 8'h2a == _T_2[7:0] ? image_42 : _GEN_41; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_235 = 8'h2b == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_427 = 8'h2b == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_235; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_619 = 8'h2b == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_427; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_811 = 8'h2b == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_619; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1003 = 8'h2b == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_811; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1195 = 8'h2b == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1003; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1387 = 8'h2b == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1195; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1579 = 8'h2b == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1387; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_43 = io_valid_in ? _GEN_1579 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_43 = 8'h2b == _T_2[7:0] ? image_43 : _GEN_42; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_236 = 8'h2c == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_428 = 8'h2c == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_236; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_620 = 8'h2c == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_428; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_812 = 8'h2c == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_620; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1004 = 8'h2c == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_812; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1196 = 8'h2c == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1004; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1388 = 8'h2c == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1196; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1580 = 8'h2c == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1388; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_44 = io_valid_in ? _GEN_1580 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_44 = 8'h2c == _T_2[7:0] ? image_44 : _GEN_43; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_237 = 8'h2d == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_429 = 8'h2d == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_237; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_621 = 8'h2d == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_429; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_813 = 8'h2d == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_621; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1005 = 8'h2d == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_813; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1197 = 8'h2d == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1005; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1389 = 8'h2d == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1197; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1581 = 8'h2d == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1389; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_45 = io_valid_in ? _GEN_1581 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_45 = 8'h2d == _T_2[7:0] ? image_45 : _GEN_44; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_238 = 8'h2e == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_430 = 8'h2e == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_238; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_622 = 8'h2e == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_430; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_814 = 8'h2e == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_622; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1006 = 8'h2e == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_814; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1198 = 8'h2e == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1006; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1390 = 8'h2e == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1198; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1582 = 8'h2e == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1390; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_46 = io_valid_in ? _GEN_1582 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_46 = 8'h2e == _T_2[7:0] ? image_46 : _GEN_45; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_239 = 8'h2f == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_431 = 8'h2f == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_239; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_623 = 8'h2f == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_431; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_815 = 8'h2f == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_623; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1007 = 8'h2f == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_815; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1199 = 8'h2f == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1007; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1391 = 8'h2f == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1199; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1583 = 8'h2f == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1391; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_47 = io_valid_in ? _GEN_1583 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_47 = 8'h2f == _T_2[7:0] ? image_47 : _GEN_46; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_240 = 8'h30 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_432 = 8'h30 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_240; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_624 = 8'h30 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_432; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_816 = 8'h30 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_624; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1008 = 8'h30 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_816; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1200 = 8'h30 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1008; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1392 = 8'h30 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1200; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1584 = 8'h30 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1392; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_48 = io_valid_in ? _GEN_1584 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_48 = 8'h30 == _T_2[7:0] ? image_48 : _GEN_47; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_241 = 8'h31 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_433 = 8'h31 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_241; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_625 = 8'h31 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_433; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_817 = 8'h31 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_625; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1009 = 8'h31 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_817; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1201 = 8'h31 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1009; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1393 = 8'h31 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1201; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1585 = 8'h31 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1393; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_49 = io_valid_in ? _GEN_1585 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_49 = 8'h31 == _T_2[7:0] ? image_49 : _GEN_48; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_242 = 8'h32 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_434 = 8'h32 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_242; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_626 = 8'h32 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_434; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_818 = 8'h32 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_626; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1010 = 8'h32 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_818; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1202 = 8'h32 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1010; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1394 = 8'h32 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1202; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1586 = 8'h32 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1394; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_50 = io_valid_in ? _GEN_1586 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_50 = 8'h32 == _T_2[7:0] ? image_50 : _GEN_49; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_243 = 8'h33 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_435 = 8'h33 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_243; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_627 = 8'h33 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_435; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_819 = 8'h33 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_627; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1011 = 8'h33 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_819; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1203 = 8'h33 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1011; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1395 = 8'h33 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1203; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1587 = 8'h33 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1395; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_51 = io_valid_in ? _GEN_1587 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_51 = 8'h33 == _T_2[7:0] ? image_51 : _GEN_50; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_244 = 8'h34 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_436 = 8'h34 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_244; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_628 = 8'h34 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_436; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_820 = 8'h34 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_628; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1012 = 8'h34 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_820; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1204 = 8'h34 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1012; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1396 = 8'h34 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1204; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1588 = 8'h34 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1396; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_52 = io_valid_in ? _GEN_1588 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_52 = 8'h34 == _T_2[7:0] ? image_52 : _GEN_51; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_245 = 8'h35 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_437 = 8'h35 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_245; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_629 = 8'h35 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_437; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_821 = 8'h35 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_629; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1013 = 8'h35 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_821; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1205 = 8'h35 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1013; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1397 = 8'h35 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1205; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1589 = 8'h35 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1397; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_53 = io_valid_in ? _GEN_1589 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_53 = 8'h35 == _T_2[7:0] ? image_53 : _GEN_52; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_246 = 8'h36 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_438 = 8'h36 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_246; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_630 = 8'h36 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_438; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_822 = 8'h36 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_630; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1014 = 8'h36 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_822; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1206 = 8'h36 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1014; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1398 = 8'h36 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1206; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1590 = 8'h36 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1398; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_54 = io_valid_in ? _GEN_1590 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_54 = 8'h36 == _T_2[7:0] ? image_54 : _GEN_53; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_247 = 8'h37 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_439 = 8'h37 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_247; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_631 = 8'h37 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_439; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_823 = 8'h37 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_631; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1015 = 8'h37 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_823; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1207 = 8'h37 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1015; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1399 = 8'h37 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1207; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1591 = 8'h37 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1399; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_55 = io_valid_in ? _GEN_1591 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_55 = 8'h37 == _T_2[7:0] ? image_55 : _GEN_54; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_248 = 8'h38 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_440 = 8'h38 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_248; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_632 = 8'h38 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_440; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_824 = 8'h38 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_632; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1016 = 8'h38 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_824; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1208 = 8'h38 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1016; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1400 = 8'h38 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1208; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1592 = 8'h38 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1400; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_56 = io_valid_in ? _GEN_1592 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_56 = 8'h38 == _T_2[7:0] ? image_56 : _GEN_55; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_249 = 8'h39 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_441 = 8'h39 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_249; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_633 = 8'h39 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_441; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_825 = 8'h39 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_633; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1017 = 8'h39 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_825; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1209 = 8'h39 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1017; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1401 = 8'h39 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1209; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1593 = 8'h39 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1401; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_57 = io_valid_in ? _GEN_1593 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_57 = 8'h39 == _T_2[7:0] ? image_57 : _GEN_56; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_250 = 8'h3a == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_442 = 8'h3a == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_250; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_634 = 8'h3a == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_442; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_826 = 8'h3a == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_634; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1018 = 8'h3a == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_826; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1210 = 8'h3a == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1018; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1402 = 8'h3a == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1210; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1594 = 8'h3a == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1402; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_58 = io_valid_in ? _GEN_1594 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_58 = 8'h3a == _T_2[7:0] ? image_58 : _GEN_57; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_251 = 8'h3b == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_443 = 8'h3b == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_251; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_635 = 8'h3b == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_443; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_827 = 8'h3b == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_635; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1019 = 8'h3b == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_827; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1211 = 8'h3b == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1019; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1403 = 8'h3b == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1211; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1595 = 8'h3b == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1403; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_59 = io_valid_in ? _GEN_1595 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_59 = 8'h3b == _T_2[7:0] ? image_59 : _GEN_58; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_252 = 8'h3c == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_444 = 8'h3c == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_252; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_636 = 8'h3c == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_444; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_828 = 8'h3c == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_636; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1020 = 8'h3c == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_828; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1212 = 8'h3c == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1020; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1404 = 8'h3c == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1212; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1596 = 8'h3c == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1404; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_60 = io_valid_in ? _GEN_1596 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_60 = 8'h3c == _T_2[7:0] ? image_60 : _GEN_59; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_253 = 8'h3d == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_445 = 8'h3d == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_253; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_637 = 8'h3d == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_445; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_829 = 8'h3d == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_637; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1021 = 8'h3d == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_829; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1213 = 8'h3d == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1021; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1405 = 8'h3d == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1213; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1597 = 8'h3d == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1405; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_61 = io_valid_in ? _GEN_1597 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_61 = 8'h3d == _T_2[7:0] ? image_61 : _GEN_60; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_254 = 8'h3e == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_446 = 8'h3e == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_254; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_638 = 8'h3e == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_446; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_830 = 8'h3e == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_638; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1022 = 8'h3e == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_830; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1214 = 8'h3e == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1022; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1406 = 8'h3e == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1214; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1598 = 8'h3e == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1406; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_62 = io_valid_in ? _GEN_1598 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_62 = 8'h3e == _T_2[7:0] ? image_62 : _GEN_61; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_255 = 8'h3f == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_447 = 8'h3f == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_255; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_639 = 8'h3f == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_447; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_831 = 8'h3f == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_639; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1023 = 8'h3f == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_831; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1215 = 8'h3f == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1023; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1407 = 8'h3f == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1215; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1599 = 8'h3f == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1407; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_63 = io_valid_in ? _GEN_1599 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_63 = 8'h3f == _T_2[7:0] ? image_63 : _GEN_62; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_256 = 8'h40 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_448 = 8'h40 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_256; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_640 = 8'h40 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_448; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_832 = 8'h40 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_640; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1024 = 8'h40 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_832; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1216 = 8'h40 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1024; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1408 = 8'h40 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1216; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1600 = 8'h40 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1408; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_64 = io_valid_in ? _GEN_1600 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_64 = 8'h40 == _T_2[7:0] ? image_64 : _GEN_63; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_257 = 8'h41 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_449 = 8'h41 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_257; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_641 = 8'h41 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_449; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_833 = 8'h41 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_641; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1025 = 8'h41 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_833; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1217 = 8'h41 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1025; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1409 = 8'h41 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1217; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1601 = 8'h41 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1409; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_65 = io_valid_in ? _GEN_1601 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_65 = 8'h41 == _T_2[7:0] ? image_65 : _GEN_64; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_258 = 8'h42 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_450 = 8'h42 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_258; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_642 = 8'h42 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_450; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_834 = 8'h42 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_642; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1026 = 8'h42 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_834; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1218 = 8'h42 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1026; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1410 = 8'h42 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1218; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1602 = 8'h42 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1410; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_66 = io_valid_in ? _GEN_1602 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_66 = 8'h42 == _T_2[7:0] ? image_66 : _GEN_65; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_259 = 8'h43 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_451 = 8'h43 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_259; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_643 = 8'h43 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_451; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_835 = 8'h43 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_643; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1027 = 8'h43 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_835; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1219 = 8'h43 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1027; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1411 = 8'h43 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1219; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1603 = 8'h43 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1411; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_67 = io_valid_in ? _GEN_1603 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_67 = 8'h43 == _T_2[7:0] ? image_67 : _GEN_66; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_260 = 8'h44 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_452 = 8'h44 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_260; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_644 = 8'h44 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_452; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_836 = 8'h44 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_644; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1028 = 8'h44 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_836; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1220 = 8'h44 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1028; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1412 = 8'h44 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1220; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1604 = 8'h44 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1412; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_68 = io_valid_in ? _GEN_1604 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_68 = 8'h44 == _T_2[7:0] ? image_68 : _GEN_67; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_261 = 8'h45 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_453 = 8'h45 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_261; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_645 = 8'h45 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_453; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_837 = 8'h45 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_645; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1029 = 8'h45 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_837; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1221 = 8'h45 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1029; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1413 = 8'h45 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1221; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1605 = 8'h45 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1413; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_69 = io_valid_in ? _GEN_1605 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_69 = 8'h45 == _T_2[7:0] ? image_69 : _GEN_68; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_262 = 8'h46 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_454 = 8'h46 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_262; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_646 = 8'h46 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_454; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_838 = 8'h46 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_646; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1030 = 8'h46 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_838; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1222 = 8'h46 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1030; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1414 = 8'h46 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1222; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1606 = 8'h46 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1414; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_70 = io_valid_in ? _GEN_1606 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_70 = 8'h46 == _T_2[7:0] ? image_70 : _GEN_69; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_263 = 8'h47 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_455 = 8'h47 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_263; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_647 = 8'h47 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_455; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_839 = 8'h47 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_647; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1031 = 8'h47 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_839; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1223 = 8'h47 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1031; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1415 = 8'h47 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1223; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1607 = 8'h47 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1415; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_71 = io_valid_in ? _GEN_1607 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_71 = 8'h47 == _T_2[7:0] ? image_71 : _GEN_70; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_264 = 8'h48 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_456 = 8'h48 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_264; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_648 = 8'h48 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_456; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_840 = 8'h48 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_648; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1032 = 8'h48 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_840; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1224 = 8'h48 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1032; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1416 = 8'h48 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1224; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1608 = 8'h48 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1416; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_72 = io_valid_in ? _GEN_1608 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_72 = 8'h48 == _T_2[7:0] ? image_72 : _GEN_71; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_265 = 8'h49 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_457 = 8'h49 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_265; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_649 = 8'h49 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_457; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_841 = 8'h49 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_649; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1033 = 8'h49 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_841; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1225 = 8'h49 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1033; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1417 = 8'h49 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1225; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1609 = 8'h49 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1417; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_73 = io_valid_in ? _GEN_1609 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_73 = 8'h49 == _T_2[7:0] ? image_73 : _GEN_72; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_266 = 8'h4a == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_458 = 8'h4a == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_266; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_650 = 8'h4a == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_458; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_842 = 8'h4a == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_650; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1034 = 8'h4a == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_842; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1226 = 8'h4a == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1034; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1418 = 8'h4a == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1226; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1610 = 8'h4a == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1418; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_74 = io_valid_in ? _GEN_1610 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_74 = 8'h4a == _T_2[7:0] ? image_74 : _GEN_73; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_267 = 8'h4b == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_459 = 8'h4b == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_267; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_651 = 8'h4b == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_459; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_843 = 8'h4b == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_651; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1035 = 8'h4b == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_843; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1227 = 8'h4b == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1035; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1419 = 8'h4b == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1227; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1611 = 8'h4b == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1419; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_75 = io_valid_in ? _GEN_1611 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_75 = 8'h4b == _T_2[7:0] ? image_75 : _GEN_74; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_268 = 8'h4c == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_460 = 8'h4c == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_268; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_652 = 8'h4c == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_460; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_844 = 8'h4c == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_652; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1036 = 8'h4c == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_844; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1228 = 8'h4c == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1036; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1420 = 8'h4c == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1228; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1612 = 8'h4c == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1420; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_76 = io_valid_in ? _GEN_1612 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_76 = 8'h4c == _T_2[7:0] ? image_76 : _GEN_75; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_269 = 8'h4d == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_461 = 8'h4d == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_269; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_653 = 8'h4d == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_461; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_845 = 8'h4d == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_653; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1037 = 8'h4d == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_845; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1229 = 8'h4d == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1037; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1421 = 8'h4d == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1229; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1613 = 8'h4d == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1421; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_77 = io_valid_in ? _GEN_1613 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_77 = 8'h4d == _T_2[7:0] ? image_77 : _GEN_76; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_270 = 8'h4e == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_462 = 8'h4e == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_270; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_654 = 8'h4e == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_462; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_846 = 8'h4e == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_654; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1038 = 8'h4e == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_846; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1230 = 8'h4e == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1038; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1422 = 8'h4e == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1230; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1614 = 8'h4e == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1422; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_78 = io_valid_in ? _GEN_1614 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_78 = 8'h4e == _T_2[7:0] ? image_78 : _GEN_77; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_271 = 8'h4f == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_463 = 8'h4f == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_271; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_655 = 8'h4f == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_463; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_847 = 8'h4f == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_655; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1039 = 8'h4f == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_847; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1231 = 8'h4f == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1039; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1423 = 8'h4f == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1231; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1615 = 8'h4f == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1423; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_79 = io_valid_in ? _GEN_1615 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_79 = 8'h4f == _T_2[7:0] ? image_79 : _GEN_78; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_272 = 8'h50 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_464 = 8'h50 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_272; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_656 = 8'h50 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_464; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_848 = 8'h50 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_656; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1040 = 8'h50 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_848; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1232 = 8'h50 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1040; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1424 = 8'h50 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1232; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1616 = 8'h50 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1424; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_80 = io_valid_in ? _GEN_1616 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_80 = 8'h50 == _T_2[7:0] ? image_80 : _GEN_79; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_273 = 8'h51 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_465 = 8'h51 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_273; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_657 = 8'h51 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_465; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_849 = 8'h51 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_657; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1041 = 8'h51 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_849; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1233 = 8'h51 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1041; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1425 = 8'h51 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1233; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1617 = 8'h51 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1425; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_81 = io_valid_in ? _GEN_1617 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_81 = 8'h51 == _T_2[7:0] ? image_81 : _GEN_80; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_274 = 8'h52 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_466 = 8'h52 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_274; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_658 = 8'h52 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_466; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_850 = 8'h52 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_658; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1042 = 8'h52 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_850; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1234 = 8'h52 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1042; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1426 = 8'h52 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1234; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1618 = 8'h52 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1426; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_82 = io_valid_in ? _GEN_1618 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_82 = 8'h52 == _T_2[7:0] ? image_82 : _GEN_81; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_275 = 8'h53 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_467 = 8'h53 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_275; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_659 = 8'h53 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_467; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_851 = 8'h53 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_659; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1043 = 8'h53 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_851; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1235 = 8'h53 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1043; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1427 = 8'h53 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1235; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1619 = 8'h53 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1427; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_83 = io_valid_in ? _GEN_1619 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_83 = 8'h53 == _T_2[7:0] ? image_83 : _GEN_82; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_276 = 8'h54 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_468 = 8'h54 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_276; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_660 = 8'h54 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_468; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_852 = 8'h54 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_660; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1044 = 8'h54 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_852; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1236 = 8'h54 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1044; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1428 = 8'h54 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1236; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1620 = 8'h54 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1428; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_84 = io_valid_in ? _GEN_1620 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_84 = 8'h54 == _T_2[7:0] ? image_84 : _GEN_83; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_277 = 8'h55 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_469 = 8'h55 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_277; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_661 = 8'h55 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_469; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_853 = 8'h55 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_661; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1045 = 8'h55 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_853; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1237 = 8'h55 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1045; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1429 = 8'h55 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1237; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1621 = 8'h55 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1429; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_85 = io_valid_in ? _GEN_1621 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_85 = 8'h55 == _T_2[7:0] ? image_85 : _GEN_84; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_278 = 8'h56 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_470 = 8'h56 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_278; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_662 = 8'h56 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_470; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_854 = 8'h56 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_662; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1046 = 8'h56 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_854; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1238 = 8'h56 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1046; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1430 = 8'h56 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1238; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1622 = 8'h56 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1430; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_86 = io_valid_in ? _GEN_1622 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_86 = 8'h56 == _T_2[7:0] ? image_86 : _GEN_85; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_279 = 8'h57 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_471 = 8'h57 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_279; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_663 = 8'h57 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_471; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_855 = 8'h57 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_663; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1047 = 8'h57 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_855; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1239 = 8'h57 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1047; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1431 = 8'h57 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1239; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1623 = 8'h57 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1431; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_87 = io_valid_in ? _GEN_1623 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_87 = 8'h57 == _T_2[7:0] ? image_87 : _GEN_86; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_280 = 8'h58 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_472 = 8'h58 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_280; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_664 = 8'h58 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_472; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_856 = 8'h58 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_664; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1048 = 8'h58 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_856; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1240 = 8'h58 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1048; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1432 = 8'h58 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1240; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1624 = 8'h58 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1432; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_88 = io_valid_in ? _GEN_1624 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_88 = 8'h58 == _T_2[7:0] ? image_88 : _GEN_87; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_281 = 8'h59 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_473 = 8'h59 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_281; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_665 = 8'h59 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_473; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_857 = 8'h59 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_665; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1049 = 8'h59 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_857; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1241 = 8'h59 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1049; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1433 = 8'h59 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1241; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1625 = 8'h59 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1433; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_89 = io_valid_in ? _GEN_1625 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_89 = 8'h59 == _T_2[7:0] ? image_89 : _GEN_88; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_282 = 8'h5a == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_474 = 8'h5a == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_282; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_666 = 8'h5a == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_474; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_858 = 8'h5a == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_666; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1050 = 8'h5a == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_858; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1242 = 8'h5a == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1050; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1434 = 8'h5a == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1242; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1626 = 8'h5a == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1434; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_90 = io_valid_in ? _GEN_1626 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_90 = 8'h5a == _T_2[7:0] ? image_90 : _GEN_89; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_283 = 8'h5b == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_475 = 8'h5b == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_283; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_667 = 8'h5b == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_475; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_859 = 8'h5b == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_667; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1051 = 8'h5b == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_859; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1243 = 8'h5b == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1051; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1435 = 8'h5b == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1243; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1627 = 8'h5b == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1435; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_91 = io_valid_in ? _GEN_1627 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_91 = 8'h5b == _T_2[7:0] ? image_91 : _GEN_90; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_284 = 8'h5c == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_476 = 8'h5c == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_284; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_668 = 8'h5c == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_476; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_860 = 8'h5c == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_668; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1052 = 8'h5c == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_860; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1244 = 8'h5c == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1052; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1436 = 8'h5c == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1244; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1628 = 8'h5c == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1436; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_92 = io_valid_in ? _GEN_1628 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_92 = 8'h5c == _T_2[7:0] ? image_92 : _GEN_91; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_285 = 8'h5d == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_477 = 8'h5d == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_285; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_669 = 8'h5d == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_477; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_861 = 8'h5d == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_669; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1053 = 8'h5d == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_861; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1245 = 8'h5d == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1053; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1437 = 8'h5d == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1245; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1629 = 8'h5d == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1437; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_93 = io_valid_in ? _GEN_1629 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_93 = 8'h5d == _T_2[7:0] ? image_93 : _GEN_92; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_286 = 8'h5e == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_478 = 8'h5e == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_286; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_670 = 8'h5e == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_478; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_862 = 8'h5e == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_670; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1054 = 8'h5e == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_862; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1246 = 8'h5e == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1054; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1438 = 8'h5e == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1246; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1630 = 8'h5e == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1438; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_94 = io_valid_in ? _GEN_1630 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_94 = 8'h5e == _T_2[7:0] ? image_94 : _GEN_93; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_287 = 8'h5f == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_479 = 8'h5f == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_287; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_671 = 8'h5f == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_479; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_863 = 8'h5f == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_671; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1055 = 8'h5f == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_863; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1247 = 8'h5f == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1055; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1439 = 8'h5f == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1247; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1631 = 8'h5f == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1439; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_95 = io_valid_in ? _GEN_1631 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_95 = 8'h5f == _T_2[7:0] ? image_95 : _GEN_94; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_288 = 8'h60 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_480 = 8'h60 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_288; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_672 = 8'h60 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_480; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_864 = 8'h60 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_672; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1056 = 8'h60 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_864; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1248 = 8'h60 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1056; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1440 = 8'h60 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1248; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1632 = 8'h60 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1440; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_96 = io_valid_in ? _GEN_1632 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_96 = 8'h60 == _T_2[7:0] ? image_96 : _GEN_95; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_289 = 8'h61 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_481 = 8'h61 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_289; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_673 = 8'h61 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_481; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_865 = 8'h61 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_673; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1057 = 8'h61 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_865; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1249 = 8'h61 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1057; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1441 = 8'h61 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1249; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1633 = 8'h61 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1441; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_97 = io_valid_in ? _GEN_1633 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_97 = 8'h61 == _T_2[7:0] ? image_97 : _GEN_96; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_290 = 8'h62 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_482 = 8'h62 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_290; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_674 = 8'h62 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_482; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_866 = 8'h62 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_674; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1058 = 8'h62 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_866; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1250 = 8'h62 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1058; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1442 = 8'h62 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1250; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1634 = 8'h62 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1442; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_98 = io_valid_in ? _GEN_1634 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_98 = 8'h62 == _T_2[7:0] ? image_98 : _GEN_97; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_291 = 8'h63 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_483 = 8'h63 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_291; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_675 = 8'h63 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_483; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_867 = 8'h63 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_675; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1059 = 8'h63 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_867; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1251 = 8'h63 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1059; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1443 = 8'h63 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1251; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1635 = 8'h63 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1443; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_99 = io_valid_in ? _GEN_1635 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_99 = 8'h63 == _T_2[7:0] ? image_99 : _GEN_98; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_292 = 8'h64 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_484 = 8'h64 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_292; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_676 = 8'h64 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_484; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_868 = 8'h64 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_676; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1060 = 8'h64 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_868; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1252 = 8'h64 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1060; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1444 = 8'h64 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1252; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1636 = 8'h64 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1444; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_100 = io_valid_in ? _GEN_1636 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_100 = 8'h64 == _T_2[7:0] ? image_100 : _GEN_99; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_293 = 8'h65 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_485 = 8'h65 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_293; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_677 = 8'h65 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_485; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_869 = 8'h65 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_677; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1061 = 8'h65 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_869; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1253 = 8'h65 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1061; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1445 = 8'h65 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1253; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1637 = 8'h65 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1445; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_101 = io_valid_in ? _GEN_1637 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_101 = 8'h65 == _T_2[7:0] ? image_101 : _GEN_100; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_294 = 8'h66 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_486 = 8'h66 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_294; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_678 = 8'h66 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_486; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_870 = 8'h66 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_678; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1062 = 8'h66 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_870; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1254 = 8'h66 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1062; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1446 = 8'h66 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1254; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1638 = 8'h66 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1446; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_102 = io_valid_in ? _GEN_1638 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_102 = 8'h66 == _T_2[7:0] ? image_102 : _GEN_101; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_295 = 8'h67 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_487 = 8'h67 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_295; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_679 = 8'h67 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_487; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_871 = 8'h67 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_679; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1063 = 8'h67 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_871; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1255 = 8'h67 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1063; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1447 = 8'h67 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1255; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1639 = 8'h67 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1447; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_103 = io_valid_in ? _GEN_1639 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_103 = 8'h67 == _T_2[7:0] ? image_103 : _GEN_102; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_296 = 8'h68 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_488 = 8'h68 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_296; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_680 = 8'h68 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_488; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_872 = 8'h68 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_680; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1064 = 8'h68 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_872; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1256 = 8'h68 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1064; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1448 = 8'h68 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1256; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1640 = 8'h68 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1448; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_104 = io_valid_in ? _GEN_1640 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_104 = 8'h68 == _T_2[7:0] ? image_104 : _GEN_103; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_297 = 8'h69 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_489 = 8'h69 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_297; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_681 = 8'h69 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_489; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_873 = 8'h69 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_681; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1065 = 8'h69 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_873; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1257 = 8'h69 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1065; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1449 = 8'h69 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1257; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1641 = 8'h69 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1449; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_105 = io_valid_in ? _GEN_1641 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_105 = 8'h69 == _T_2[7:0] ? image_105 : _GEN_104; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_298 = 8'h6a == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_490 = 8'h6a == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_298; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_682 = 8'h6a == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_490; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_874 = 8'h6a == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_682; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1066 = 8'h6a == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_874; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1258 = 8'h6a == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1066; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1450 = 8'h6a == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1258; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1642 = 8'h6a == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1450; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_106 = io_valid_in ? _GEN_1642 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_106 = 8'h6a == _T_2[7:0] ? image_106 : _GEN_105; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_299 = 8'h6b == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_491 = 8'h6b == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_299; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_683 = 8'h6b == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_491; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_875 = 8'h6b == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_683; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1067 = 8'h6b == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_875; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1259 = 8'h6b == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1067; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1451 = 8'h6b == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1259; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1643 = 8'h6b == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1451; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_107 = io_valid_in ? _GEN_1643 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_107 = 8'h6b == _T_2[7:0] ? image_107 : _GEN_106; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_300 = 8'h6c == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_492 = 8'h6c == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_300; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_684 = 8'h6c == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_492; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_876 = 8'h6c == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_684; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1068 = 8'h6c == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_876; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1260 = 8'h6c == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1068; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1452 = 8'h6c == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1260; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1644 = 8'h6c == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1452; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_108 = io_valid_in ? _GEN_1644 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_108 = 8'h6c == _T_2[7:0] ? image_108 : _GEN_107; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_301 = 8'h6d == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_493 = 8'h6d == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_301; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_685 = 8'h6d == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_493; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_877 = 8'h6d == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_685; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1069 = 8'h6d == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_877; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1261 = 8'h6d == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1069; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1453 = 8'h6d == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1261; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1645 = 8'h6d == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1453; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_109 = io_valid_in ? _GEN_1645 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_109 = 8'h6d == _T_2[7:0] ? image_109 : _GEN_108; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_302 = 8'h6e == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_494 = 8'h6e == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_302; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_686 = 8'h6e == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_494; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_878 = 8'h6e == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_686; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1070 = 8'h6e == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_878; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1262 = 8'h6e == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1070; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1454 = 8'h6e == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1262; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1646 = 8'h6e == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1454; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_110 = io_valid_in ? _GEN_1646 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_110 = 8'h6e == _T_2[7:0] ? image_110 : _GEN_109; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_303 = 8'h6f == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_495 = 8'h6f == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_303; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_687 = 8'h6f == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_495; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_879 = 8'h6f == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_687; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1071 = 8'h6f == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_879; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1263 = 8'h6f == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1071; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1455 = 8'h6f == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1263; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1647 = 8'h6f == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1455; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_111 = io_valid_in ? _GEN_1647 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_111 = 8'h6f == _T_2[7:0] ? image_111 : _GEN_110; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_304 = 8'h70 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_496 = 8'h70 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_304; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_688 = 8'h70 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_496; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_880 = 8'h70 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_688; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1072 = 8'h70 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_880; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1264 = 8'h70 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1072; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1456 = 8'h70 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1264; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1648 = 8'h70 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1456; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_112 = io_valid_in ? _GEN_1648 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_112 = 8'h70 == _T_2[7:0] ? image_112 : _GEN_111; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_305 = 8'h71 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_497 = 8'h71 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_305; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_689 = 8'h71 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_497; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_881 = 8'h71 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_689; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1073 = 8'h71 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_881; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1265 = 8'h71 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1073; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1457 = 8'h71 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1265; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1649 = 8'h71 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1457; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_113 = io_valid_in ? _GEN_1649 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_113 = 8'h71 == _T_2[7:0] ? image_113 : _GEN_112; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_306 = 8'h72 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_498 = 8'h72 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_306; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_690 = 8'h72 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_498; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_882 = 8'h72 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_690; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1074 = 8'h72 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_882; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1266 = 8'h72 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1074; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1458 = 8'h72 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1266; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1650 = 8'h72 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1458; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_114 = io_valid_in ? _GEN_1650 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_114 = 8'h72 == _T_2[7:0] ? image_114 : _GEN_113; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_307 = 8'h73 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_499 = 8'h73 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_307; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_691 = 8'h73 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_499; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_883 = 8'h73 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_691; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1075 = 8'h73 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_883; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1267 = 8'h73 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1075; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1459 = 8'h73 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1267; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1651 = 8'h73 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1459; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_115 = io_valid_in ? _GEN_1651 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_115 = 8'h73 == _T_2[7:0] ? image_115 : _GEN_114; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_308 = 8'h74 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_500 = 8'h74 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_308; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_692 = 8'h74 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_500; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_884 = 8'h74 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_692; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1076 = 8'h74 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_884; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1268 = 8'h74 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1076; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1460 = 8'h74 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1268; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1652 = 8'h74 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1460; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_116 = io_valid_in ? _GEN_1652 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_116 = 8'h74 == _T_2[7:0] ? image_116 : _GEN_115; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_309 = 8'h75 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_501 = 8'h75 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_309; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_693 = 8'h75 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_501; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_885 = 8'h75 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_693; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1077 = 8'h75 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_885; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1269 = 8'h75 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1077; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1461 = 8'h75 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1269; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1653 = 8'h75 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1461; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_117 = io_valid_in ? _GEN_1653 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_117 = 8'h75 == _T_2[7:0] ? image_117 : _GEN_116; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_310 = 8'h76 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_502 = 8'h76 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_310; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_694 = 8'h76 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_502; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_886 = 8'h76 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_694; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1078 = 8'h76 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_886; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1270 = 8'h76 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1078; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1462 = 8'h76 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1270; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1654 = 8'h76 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1462; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_118 = io_valid_in ? _GEN_1654 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_118 = 8'h76 == _T_2[7:0] ? image_118 : _GEN_117; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_311 = 8'h77 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_503 = 8'h77 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_311; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_695 = 8'h77 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_503; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_887 = 8'h77 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_695; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1079 = 8'h77 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_887; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1271 = 8'h77 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1079; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1463 = 8'h77 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1271; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1655 = 8'h77 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1463; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_119 = io_valid_in ? _GEN_1655 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_119 = 8'h77 == _T_2[7:0] ? image_119 : _GEN_118; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_312 = 8'h78 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_504 = 8'h78 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_312; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_696 = 8'h78 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_504; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_888 = 8'h78 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_696; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1080 = 8'h78 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_888; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1272 = 8'h78 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1080; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1464 = 8'h78 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1272; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1656 = 8'h78 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1464; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_120 = io_valid_in ? _GEN_1656 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_120 = 8'h78 == _T_2[7:0] ? image_120 : _GEN_119; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_313 = 8'h79 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_505 = 8'h79 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_313; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_697 = 8'h79 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_505; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_889 = 8'h79 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_697; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1081 = 8'h79 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_889; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1273 = 8'h79 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1081; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1465 = 8'h79 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1273; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1657 = 8'h79 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1465; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_121 = io_valid_in ? _GEN_1657 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_121 = 8'h79 == _T_2[7:0] ? image_121 : _GEN_120; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_314 = 8'h7a == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_506 = 8'h7a == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_314; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_698 = 8'h7a == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_506; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_890 = 8'h7a == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_698; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1082 = 8'h7a == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_890; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1274 = 8'h7a == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1082; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1466 = 8'h7a == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1274; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1658 = 8'h7a == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1466; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_122 = io_valid_in ? _GEN_1658 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_122 = 8'h7a == _T_2[7:0] ? image_122 : _GEN_121; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_315 = 8'h7b == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_507 = 8'h7b == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_315; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_699 = 8'h7b == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_507; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_891 = 8'h7b == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_699; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1083 = 8'h7b == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_891; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1275 = 8'h7b == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1083; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1467 = 8'h7b == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1275; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1659 = 8'h7b == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1467; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_123 = io_valid_in ? _GEN_1659 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_123 = 8'h7b == _T_2[7:0] ? image_123 : _GEN_122; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_316 = 8'h7c == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_508 = 8'h7c == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_316; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_700 = 8'h7c == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_508; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_892 = 8'h7c == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_700; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1084 = 8'h7c == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_892; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1276 = 8'h7c == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1084; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1468 = 8'h7c == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1276; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1660 = 8'h7c == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1468; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_124 = io_valid_in ? _GEN_1660 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_124 = 8'h7c == _T_2[7:0] ? image_124 : _GEN_123; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_317 = 8'h7d == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_509 = 8'h7d == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_317; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_701 = 8'h7d == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_509; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_893 = 8'h7d == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_701; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1085 = 8'h7d == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_893; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1277 = 8'h7d == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1085; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1469 = 8'h7d == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1277; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1661 = 8'h7d == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1469; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_125 = io_valid_in ? _GEN_1661 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_125 = 8'h7d == _T_2[7:0] ? image_125 : _GEN_124; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_318 = 8'h7e == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_510 = 8'h7e == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_318; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_702 = 8'h7e == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_510; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_894 = 8'h7e == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_702; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1086 = 8'h7e == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_894; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1278 = 8'h7e == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1086; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1470 = 8'h7e == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1278; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1662 = 8'h7e == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1470; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_126 = io_valid_in ? _GEN_1662 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_126 = 8'h7e == _T_2[7:0] ? image_126 : _GEN_125; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_319 = 8'h7f == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_511 = 8'h7f == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_319; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_703 = 8'h7f == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_511; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_895 = 8'h7f == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_703; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1087 = 8'h7f == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_895; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1279 = 8'h7f == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1087; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1471 = 8'h7f == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1279; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1663 = 8'h7f == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1471; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_127 = io_valid_in ? _GEN_1663 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_127 = 8'h7f == _T_2[7:0] ? image_127 : _GEN_126; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_320 = 8'h80 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_512 = 8'h80 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_320; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_704 = 8'h80 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_512; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_896 = 8'h80 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_704; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1088 = 8'h80 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_896; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1280 = 8'h80 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1088; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1472 = 8'h80 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1280; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1664 = 8'h80 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1472; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_128 = io_valid_in ? _GEN_1664 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_128 = 8'h80 == _T_2[7:0] ? image_128 : _GEN_127; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_321 = 8'h81 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_513 = 8'h81 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_321; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_705 = 8'h81 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_513; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_897 = 8'h81 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_705; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1089 = 8'h81 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_897; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1281 = 8'h81 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1089; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1473 = 8'h81 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1281; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1665 = 8'h81 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1473; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_129 = io_valid_in ? _GEN_1665 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_129 = 8'h81 == _T_2[7:0] ? image_129 : _GEN_128; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_322 = 8'h82 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_514 = 8'h82 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_322; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_706 = 8'h82 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_514; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_898 = 8'h82 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_706; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1090 = 8'h82 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_898; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1282 = 8'h82 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1090; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1474 = 8'h82 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1282; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1666 = 8'h82 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1474; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_130 = io_valid_in ? _GEN_1666 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_130 = 8'h82 == _T_2[7:0] ? image_130 : _GEN_129; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_323 = 8'h83 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_515 = 8'h83 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_323; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_707 = 8'h83 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_515; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_899 = 8'h83 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_707; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1091 = 8'h83 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_899; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1283 = 8'h83 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1091; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1475 = 8'h83 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1283; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1667 = 8'h83 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1475; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_131 = io_valid_in ? _GEN_1667 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_131 = 8'h83 == _T_2[7:0] ? image_131 : _GEN_130; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_324 = 8'h84 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_516 = 8'h84 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_324; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_708 = 8'h84 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_516; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_900 = 8'h84 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_708; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1092 = 8'h84 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_900; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1284 = 8'h84 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1092; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1476 = 8'h84 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1284; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1668 = 8'h84 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1476; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_132 = io_valid_in ? _GEN_1668 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_132 = 8'h84 == _T_2[7:0] ? image_132 : _GEN_131; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_325 = 8'h85 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_517 = 8'h85 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_325; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_709 = 8'h85 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_517; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_901 = 8'h85 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_709; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1093 = 8'h85 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_901; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1285 = 8'h85 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1093; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1477 = 8'h85 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1285; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1669 = 8'h85 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1477; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_133 = io_valid_in ? _GEN_1669 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_133 = 8'h85 == _T_2[7:0] ? image_133 : _GEN_132; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_326 = 8'h86 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_518 = 8'h86 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_326; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_710 = 8'h86 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_518; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_902 = 8'h86 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_710; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1094 = 8'h86 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_902; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1286 = 8'h86 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1094; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1478 = 8'h86 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1286; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1670 = 8'h86 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1478; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_134 = io_valid_in ? _GEN_1670 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_134 = 8'h86 == _T_2[7:0] ? image_134 : _GEN_133; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_327 = 8'h87 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_519 = 8'h87 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_327; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_711 = 8'h87 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_519; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_903 = 8'h87 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_711; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1095 = 8'h87 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_903; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1287 = 8'h87 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1095; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1479 = 8'h87 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1287; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1671 = 8'h87 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1479; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_135 = io_valid_in ? _GEN_1671 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_135 = 8'h87 == _T_2[7:0] ? image_135 : _GEN_134; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_328 = 8'h88 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_520 = 8'h88 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_328; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_712 = 8'h88 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_520; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_904 = 8'h88 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_712; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1096 = 8'h88 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_904; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1288 = 8'h88 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1096; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1480 = 8'h88 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1288; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1672 = 8'h88 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1480; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_136 = io_valid_in ? _GEN_1672 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_136 = 8'h88 == _T_2[7:0] ? image_136 : _GEN_135; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_329 = 8'h89 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_521 = 8'h89 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_329; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_713 = 8'h89 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_521; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_905 = 8'h89 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_713; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1097 = 8'h89 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_905; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1289 = 8'h89 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1097; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1481 = 8'h89 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1289; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1673 = 8'h89 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1481; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_137 = io_valid_in ? _GEN_1673 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_137 = 8'h89 == _T_2[7:0] ? image_137 : _GEN_136; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_330 = 8'h8a == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_522 = 8'h8a == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_330; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_714 = 8'h8a == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_522; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_906 = 8'h8a == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_714; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1098 = 8'h8a == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_906; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1290 = 8'h8a == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1098; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1482 = 8'h8a == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1290; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1674 = 8'h8a == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1482; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_138 = io_valid_in ? _GEN_1674 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_138 = 8'h8a == _T_2[7:0] ? image_138 : _GEN_137; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_331 = 8'h8b == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_523 = 8'h8b == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_331; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_715 = 8'h8b == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_523; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_907 = 8'h8b == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_715; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1099 = 8'h8b == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_907; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1291 = 8'h8b == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1099; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1483 = 8'h8b == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1291; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1675 = 8'h8b == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1483; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_139 = io_valid_in ? _GEN_1675 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_139 = 8'h8b == _T_2[7:0] ? image_139 : _GEN_138; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_332 = 8'h8c == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_524 = 8'h8c == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_332; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_716 = 8'h8c == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_524; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_908 = 8'h8c == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_716; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1100 = 8'h8c == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_908; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1292 = 8'h8c == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1100; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1484 = 8'h8c == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1292; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1676 = 8'h8c == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1484; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_140 = io_valid_in ? _GEN_1676 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_140 = 8'h8c == _T_2[7:0] ? image_140 : _GEN_139; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_333 = 8'h8d == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_525 = 8'h8d == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_333; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_717 = 8'h8d == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_525; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_909 = 8'h8d == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_717; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1101 = 8'h8d == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_909; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1293 = 8'h8d == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1101; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1485 = 8'h8d == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1293; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1677 = 8'h8d == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1485; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_141 = io_valid_in ? _GEN_1677 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_141 = 8'h8d == _T_2[7:0] ? image_141 : _GEN_140; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_334 = 8'h8e == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_526 = 8'h8e == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_334; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_718 = 8'h8e == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_526; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_910 = 8'h8e == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_718; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1102 = 8'h8e == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_910; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1294 = 8'h8e == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1102; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1486 = 8'h8e == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1294; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1678 = 8'h8e == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1486; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_142 = io_valid_in ? _GEN_1678 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_142 = 8'h8e == _T_2[7:0] ? image_142 : _GEN_141; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_335 = 8'h8f == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_527 = 8'h8f == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_335; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_719 = 8'h8f == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_527; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_911 = 8'h8f == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_719; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1103 = 8'h8f == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_911; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1295 = 8'h8f == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1103; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1487 = 8'h8f == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1295; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1679 = 8'h8f == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1487; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_143 = io_valid_in ? _GEN_1679 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_143 = 8'h8f == _T_2[7:0] ? image_143 : _GEN_142; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_336 = 8'h90 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_528 = 8'h90 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_336; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_720 = 8'h90 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_528; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_912 = 8'h90 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_720; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1104 = 8'h90 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_912; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1296 = 8'h90 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1104; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1488 = 8'h90 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1296; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1680 = 8'h90 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1488; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_144 = io_valid_in ? _GEN_1680 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_144 = 8'h90 == _T_2[7:0] ? image_144 : _GEN_143; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_337 = 8'h91 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_529 = 8'h91 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_337; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_721 = 8'h91 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_529; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_913 = 8'h91 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_721; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1105 = 8'h91 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_913; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1297 = 8'h91 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1105; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1489 = 8'h91 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1297; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1681 = 8'h91 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1489; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_145 = io_valid_in ? _GEN_1681 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_145 = 8'h91 == _T_2[7:0] ? image_145 : _GEN_144; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_338 = 8'h92 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_530 = 8'h92 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_338; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_722 = 8'h92 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_530; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_914 = 8'h92 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_722; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1106 = 8'h92 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_914; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1298 = 8'h92 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1106; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1490 = 8'h92 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1298; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1682 = 8'h92 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1490; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_146 = io_valid_in ? _GEN_1682 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_146 = 8'h92 == _T_2[7:0] ? image_146 : _GEN_145; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_339 = 8'h93 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_531 = 8'h93 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_339; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_723 = 8'h93 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_531; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_915 = 8'h93 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_723; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1107 = 8'h93 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_915; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1299 = 8'h93 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1107; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1491 = 8'h93 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1299; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1683 = 8'h93 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1491; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_147 = io_valid_in ? _GEN_1683 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_147 = 8'h93 == _T_2[7:0] ? image_147 : _GEN_146; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_340 = 8'h94 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_532 = 8'h94 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_340; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_724 = 8'h94 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_532; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_916 = 8'h94 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_724; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1108 = 8'h94 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_916; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1300 = 8'h94 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1108; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1492 = 8'h94 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1300; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1684 = 8'h94 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1492; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_148 = io_valid_in ? _GEN_1684 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_148 = 8'h94 == _T_2[7:0] ? image_148 : _GEN_147; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_341 = 8'h95 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_533 = 8'h95 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_341; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_725 = 8'h95 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_533; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_917 = 8'h95 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_725; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1109 = 8'h95 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_917; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1301 = 8'h95 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1109; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1493 = 8'h95 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1301; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1685 = 8'h95 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1493; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_149 = io_valid_in ? _GEN_1685 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_149 = 8'h95 == _T_2[7:0] ? image_149 : _GEN_148; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_342 = 8'h96 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_534 = 8'h96 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_342; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_726 = 8'h96 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_534; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_918 = 8'h96 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_726; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1110 = 8'h96 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_918; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1302 = 8'h96 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1110; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1494 = 8'h96 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1302; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1686 = 8'h96 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1494; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_150 = io_valid_in ? _GEN_1686 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_150 = 8'h96 == _T_2[7:0] ? image_150 : _GEN_149; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_343 = 8'h97 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_535 = 8'h97 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_343; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_727 = 8'h97 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_535; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_919 = 8'h97 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_727; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1111 = 8'h97 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_919; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1303 = 8'h97 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1111; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1495 = 8'h97 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1303; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1687 = 8'h97 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1495; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_151 = io_valid_in ? _GEN_1687 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_151 = 8'h97 == _T_2[7:0] ? image_151 : _GEN_150; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_344 = 8'h98 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_536 = 8'h98 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_344; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_728 = 8'h98 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_536; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_920 = 8'h98 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_728; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1112 = 8'h98 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_920; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1304 = 8'h98 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1112; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1496 = 8'h98 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1304; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1688 = 8'h98 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1496; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_152 = io_valid_in ? _GEN_1688 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_152 = 8'h98 == _T_2[7:0] ? image_152 : _GEN_151; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_345 = 8'h99 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_537 = 8'h99 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_345; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_729 = 8'h99 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_537; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_921 = 8'h99 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_729; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1113 = 8'h99 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_921; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1305 = 8'h99 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1113; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1497 = 8'h99 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1305; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1689 = 8'h99 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1497; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_153 = io_valid_in ? _GEN_1689 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_153 = 8'h99 == _T_2[7:0] ? image_153 : _GEN_152; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_346 = 8'h9a == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_538 = 8'h9a == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_346; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_730 = 8'h9a == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_538; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_922 = 8'h9a == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_730; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1114 = 8'h9a == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_922; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1306 = 8'h9a == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1114; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1498 = 8'h9a == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1306; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1690 = 8'h9a == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1498; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_154 = io_valid_in ? _GEN_1690 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_154 = 8'h9a == _T_2[7:0] ? image_154 : _GEN_153; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_347 = 8'h9b == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_539 = 8'h9b == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_347; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_731 = 8'h9b == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_539; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_923 = 8'h9b == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_731; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1115 = 8'h9b == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_923; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1307 = 8'h9b == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1115; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1499 = 8'h9b == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1307; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1691 = 8'h9b == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1499; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_155 = io_valid_in ? _GEN_1691 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_155 = 8'h9b == _T_2[7:0] ? image_155 : _GEN_154; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_348 = 8'h9c == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_540 = 8'h9c == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_348; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_732 = 8'h9c == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_540; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_924 = 8'h9c == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_732; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1116 = 8'h9c == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_924; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1308 = 8'h9c == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1116; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1500 = 8'h9c == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1308; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1692 = 8'h9c == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1500; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_156 = io_valid_in ? _GEN_1692 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_156 = 8'h9c == _T_2[7:0] ? image_156 : _GEN_155; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_349 = 8'h9d == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_541 = 8'h9d == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_349; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_733 = 8'h9d == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_541; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_925 = 8'h9d == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_733; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1117 = 8'h9d == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_925; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1309 = 8'h9d == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1117; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1501 = 8'h9d == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1309; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1693 = 8'h9d == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1501; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_157 = io_valid_in ? _GEN_1693 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_157 = 8'h9d == _T_2[7:0] ? image_157 : _GEN_156; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_350 = 8'h9e == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_542 = 8'h9e == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_350; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_734 = 8'h9e == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_542; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_926 = 8'h9e == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_734; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1118 = 8'h9e == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_926; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1310 = 8'h9e == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1118; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1502 = 8'h9e == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1310; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1694 = 8'h9e == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1502; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_158 = io_valid_in ? _GEN_1694 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_158 = 8'h9e == _T_2[7:0] ? image_158 : _GEN_157; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_351 = 8'h9f == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_543 = 8'h9f == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_351; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_735 = 8'h9f == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_543; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_927 = 8'h9f == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_735; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1119 = 8'h9f == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_927; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1311 = 8'h9f == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1119; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1503 = 8'h9f == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1311; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1695 = 8'h9f == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1503; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_159 = io_valid_in ? _GEN_1695 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_159 = 8'h9f == _T_2[7:0] ? image_159 : _GEN_158; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_352 = 8'ha0 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_544 = 8'ha0 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_352; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_736 = 8'ha0 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_544; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_928 = 8'ha0 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_736; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1120 = 8'ha0 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_928; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1312 = 8'ha0 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1120; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1504 = 8'ha0 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1312; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1696 = 8'ha0 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1504; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_160 = io_valid_in ? _GEN_1696 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_160 = 8'ha0 == _T_2[7:0] ? image_160 : _GEN_159; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_353 = 8'ha1 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_545 = 8'ha1 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_353; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_737 = 8'ha1 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_545; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_929 = 8'ha1 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_737; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1121 = 8'ha1 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_929; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1313 = 8'ha1 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1121; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1505 = 8'ha1 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1313; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1697 = 8'ha1 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1505; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_161 = io_valid_in ? _GEN_1697 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_161 = 8'ha1 == _T_2[7:0] ? image_161 : _GEN_160; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_354 = 8'ha2 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_546 = 8'ha2 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_354; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_738 = 8'ha2 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_546; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_930 = 8'ha2 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_738; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1122 = 8'ha2 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_930; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1314 = 8'ha2 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1122; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1506 = 8'ha2 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1314; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1698 = 8'ha2 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1506; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_162 = io_valid_in ? _GEN_1698 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_162 = 8'ha2 == _T_2[7:0] ? image_162 : _GEN_161; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_355 = 8'ha3 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_547 = 8'ha3 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_355; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_739 = 8'ha3 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_547; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_931 = 8'ha3 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_739; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1123 = 8'ha3 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_931; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1315 = 8'ha3 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1123; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1507 = 8'ha3 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1315; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1699 = 8'ha3 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1507; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_163 = io_valid_in ? _GEN_1699 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_163 = 8'ha3 == _T_2[7:0] ? image_163 : _GEN_162; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_356 = 8'ha4 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_548 = 8'ha4 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_356; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_740 = 8'ha4 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_548; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_932 = 8'ha4 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_740; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1124 = 8'ha4 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_932; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1316 = 8'ha4 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1124; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1508 = 8'ha4 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1316; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1700 = 8'ha4 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1508; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_164 = io_valid_in ? _GEN_1700 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_164 = 8'ha4 == _T_2[7:0] ? image_164 : _GEN_163; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_357 = 8'ha5 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_549 = 8'ha5 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_357; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_741 = 8'ha5 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_549; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_933 = 8'ha5 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_741; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1125 = 8'ha5 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_933; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1317 = 8'ha5 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1125; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1509 = 8'ha5 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1317; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1701 = 8'ha5 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1509; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_165 = io_valid_in ? _GEN_1701 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_165 = 8'ha5 == _T_2[7:0] ? image_165 : _GEN_164; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_358 = 8'ha6 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_550 = 8'ha6 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_358; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_742 = 8'ha6 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_550; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_934 = 8'ha6 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_742; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1126 = 8'ha6 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_934; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1318 = 8'ha6 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1126; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1510 = 8'ha6 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1318; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1702 = 8'ha6 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1510; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_166 = io_valid_in ? _GEN_1702 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_166 = 8'ha6 == _T_2[7:0] ? image_166 : _GEN_165; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_359 = 8'ha7 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_551 = 8'ha7 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_359; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_743 = 8'ha7 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_551; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_935 = 8'ha7 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_743; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1127 = 8'ha7 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_935; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1319 = 8'ha7 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1127; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1511 = 8'ha7 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1319; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1703 = 8'ha7 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1511; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_167 = io_valid_in ? _GEN_1703 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_167 = 8'ha7 == _T_2[7:0] ? image_167 : _GEN_166; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_360 = 8'ha8 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_552 = 8'ha8 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_360; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_744 = 8'ha8 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_552; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_936 = 8'ha8 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_744; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1128 = 8'ha8 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_936; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1320 = 8'ha8 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1128; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1512 = 8'ha8 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1320; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1704 = 8'ha8 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1512; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_168 = io_valid_in ? _GEN_1704 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_168 = 8'ha8 == _T_2[7:0] ? image_168 : _GEN_167; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_361 = 8'ha9 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_553 = 8'ha9 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_361; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_745 = 8'ha9 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_553; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_937 = 8'ha9 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_745; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1129 = 8'ha9 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_937; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1321 = 8'ha9 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1129; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1513 = 8'ha9 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1321; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1705 = 8'ha9 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1513; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_169 = io_valid_in ? _GEN_1705 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_169 = 8'ha9 == _T_2[7:0] ? image_169 : _GEN_168; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_362 = 8'haa == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_554 = 8'haa == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_362; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_746 = 8'haa == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_554; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_938 = 8'haa == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_746; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1130 = 8'haa == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_938; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1322 = 8'haa == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1130; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1514 = 8'haa == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1322; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1706 = 8'haa == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1514; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_170 = io_valid_in ? _GEN_1706 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_170 = 8'haa == _T_2[7:0] ? image_170 : _GEN_169; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_363 = 8'hab == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_555 = 8'hab == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_363; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_747 = 8'hab == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_555; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_939 = 8'hab == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_747; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1131 = 8'hab == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_939; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1323 = 8'hab == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1131; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1515 = 8'hab == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1323; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1707 = 8'hab == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1515; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_171 = io_valid_in ? _GEN_1707 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_171 = 8'hab == _T_2[7:0] ? image_171 : _GEN_170; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_364 = 8'hac == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_556 = 8'hac == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_364; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_748 = 8'hac == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_556; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_940 = 8'hac == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_748; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1132 = 8'hac == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_940; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1324 = 8'hac == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1132; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1516 = 8'hac == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1324; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1708 = 8'hac == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1516; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_172 = io_valid_in ? _GEN_1708 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_172 = 8'hac == _T_2[7:0] ? image_172 : _GEN_171; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_365 = 8'had == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_557 = 8'had == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_365; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_749 = 8'had == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_557; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_941 = 8'had == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_749; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1133 = 8'had == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_941; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1325 = 8'had == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1133; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1517 = 8'had == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1325; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1709 = 8'had == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1517; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_173 = io_valid_in ? _GEN_1709 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_173 = 8'had == _T_2[7:0] ? image_173 : _GEN_172; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_366 = 8'hae == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_558 = 8'hae == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_366; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_750 = 8'hae == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_558; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_942 = 8'hae == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_750; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1134 = 8'hae == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_942; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1326 = 8'hae == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1134; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1518 = 8'hae == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1326; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1710 = 8'hae == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1518; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_174 = io_valid_in ? _GEN_1710 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_174 = 8'hae == _T_2[7:0] ? image_174 : _GEN_173; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_367 = 8'haf == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_559 = 8'haf == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_367; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_751 = 8'haf == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_559; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_943 = 8'haf == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_751; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1135 = 8'haf == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_943; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1327 = 8'haf == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1135; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1519 = 8'haf == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1327; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1711 = 8'haf == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1519; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_175 = io_valid_in ? _GEN_1711 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_175 = 8'haf == _T_2[7:0] ? image_175 : _GEN_174; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_368 = 8'hb0 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_560 = 8'hb0 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_368; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_752 = 8'hb0 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_560; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_944 = 8'hb0 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_752; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1136 = 8'hb0 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_944; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1328 = 8'hb0 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1136; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1520 = 8'hb0 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1328; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1712 = 8'hb0 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1520; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_176 = io_valid_in ? _GEN_1712 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_176 = 8'hb0 == _T_2[7:0] ? image_176 : _GEN_175; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_369 = 8'hb1 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_561 = 8'hb1 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_369; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_753 = 8'hb1 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_561; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_945 = 8'hb1 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_753; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1137 = 8'hb1 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_945; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1329 = 8'hb1 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1137; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1521 = 8'hb1 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1329; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1713 = 8'hb1 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1521; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_177 = io_valid_in ? _GEN_1713 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_177 = 8'hb1 == _T_2[7:0] ? image_177 : _GEN_176; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_370 = 8'hb2 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_562 = 8'hb2 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_370; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_754 = 8'hb2 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_562; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_946 = 8'hb2 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_754; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1138 = 8'hb2 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_946; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1330 = 8'hb2 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1138; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1522 = 8'hb2 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1330; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1714 = 8'hb2 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1522; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_178 = io_valid_in ? _GEN_1714 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_178 = 8'hb2 == _T_2[7:0] ? image_178 : _GEN_177; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_371 = 8'hb3 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_563 = 8'hb3 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_371; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_755 = 8'hb3 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_563; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_947 = 8'hb3 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_755; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1139 = 8'hb3 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_947; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1331 = 8'hb3 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1139; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1523 = 8'hb3 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1331; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1715 = 8'hb3 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1523; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_179 = io_valid_in ? _GEN_1715 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_179 = 8'hb3 == _T_2[7:0] ? image_179 : _GEN_178; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_372 = 8'hb4 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_564 = 8'hb4 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_372; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_756 = 8'hb4 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_564; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_948 = 8'hb4 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_756; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1140 = 8'hb4 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_948; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1332 = 8'hb4 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1140; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1524 = 8'hb4 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1332; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1716 = 8'hb4 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1524; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_180 = io_valid_in ? _GEN_1716 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_180 = 8'hb4 == _T_2[7:0] ? image_180 : _GEN_179; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_373 = 8'hb5 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_565 = 8'hb5 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_373; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_757 = 8'hb5 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_565; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_949 = 8'hb5 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_757; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1141 = 8'hb5 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_949; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1333 = 8'hb5 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1141; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1525 = 8'hb5 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1333; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1717 = 8'hb5 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1525; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_181 = io_valid_in ? _GEN_1717 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_181 = 8'hb5 == _T_2[7:0] ? image_181 : _GEN_180; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_374 = 8'hb6 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_566 = 8'hb6 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_374; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_758 = 8'hb6 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_566; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_950 = 8'hb6 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_758; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1142 = 8'hb6 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_950; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1334 = 8'hb6 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1142; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1526 = 8'hb6 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1334; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1718 = 8'hb6 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1526; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_182 = io_valid_in ? _GEN_1718 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_182 = 8'hb6 == _T_2[7:0] ? image_182 : _GEN_181; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_375 = 8'hb7 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_567 = 8'hb7 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_375; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_759 = 8'hb7 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_567; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_951 = 8'hb7 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_759; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1143 = 8'hb7 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_951; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1335 = 8'hb7 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1143; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1527 = 8'hb7 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1335; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1719 = 8'hb7 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1527; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_183 = io_valid_in ? _GEN_1719 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_183 = 8'hb7 == _T_2[7:0] ? image_183 : _GEN_182; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_376 = 8'hb8 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_568 = 8'hb8 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_376; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_760 = 8'hb8 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_568; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_952 = 8'hb8 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_760; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1144 = 8'hb8 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_952; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1336 = 8'hb8 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1144; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1528 = 8'hb8 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1336; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1720 = 8'hb8 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1528; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_184 = io_valid_in ? _GEN_1720 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_184 = 8'hb8 == _T_2[7:0] ? image_184 : _GEN_183; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_377 = 8'hb9 == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_569 = 8'hb9 == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_377; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_761 = 8'hb9 == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_569; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_953 = 8'hb9 == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_761; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1145 = 8'hb9 == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_953; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1337 = 8'hb9 == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1145; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1529 = 8'hb9 == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1337; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1721 = 8'hb9 == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1529; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_185 = io_valid_in ? _GEN_1721 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_185 = 8'hb9 == _T_2[7:0] ? image_185 : _GEN_184; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_378 = 8'hba == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_570 = 8'hba == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_378; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_762 = 8'hba == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_570; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_954 = 8'hba == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_762; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1146 = 8'hba == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_954; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1338 = 8'hba == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1146; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1530 = 8'hba == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1338; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1722 = 8'hba == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1530; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_186 = io_valid_in ? _GEN_1722 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_186 = 8'hba == _T_2[7:0] ? image_186 : _GEN_185; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_379 = 8'hbb == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_571 = 8'hbb == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_379; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_763 = 8'hbb == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_571; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_955 = 8'hbb == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_763; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1147 = 8'hbb == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_955; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1339 = 8'hbb == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1147; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1531 = 8'hbb == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1339; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1723 = 8'hbb == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1531; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_187 = io_valid_in ? _GEN_1723 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_187 = 8'hbb == _T_2[7:0] ? image_187 : _GEN_186; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_380 = 8'hbc == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_572 = 8'hbc == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_380; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_764 = 8'hbc == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_572; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_956 = 8'hbc == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_764; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1148 = 8'hbc == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_956; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1340 = 8'hbc == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1148; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1532 = 8'hbc == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1340; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1724 = 8'hbc == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1532; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_188 = io_valid_in ? _GEN_1724 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_188 = 8'hbc == _T_2[7:0] ? image_188 : _GEN_187; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_381 = 8'hbd == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_573 = 8'hbd == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_381; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_765 = 8'hbd == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_573; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_957 = 8'hbd == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_765; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1149 = 8'hbd == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_957; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1341 = 8'hbd == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1149; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1533 = 8'hbd == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1341; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1725 = 8'hbd == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1533; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_189 = io_valid_in ? _GEN_1725 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_189 = 8'hbd == _T_2[7:0] ? image_189 : _GEN_188; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_382 = 8'hbe == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_574 = 8'hbe == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_382; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_766 = 8'hbe == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_574; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_958 = 8'hbe == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_766; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1150 = 8'hbe == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_958; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1342 = 8'hbe == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1150; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1534 = 8'hbe == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1342; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1726 = 8'hbe == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1534; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_190 = io_valid_in ? _GEN_1726 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_190 = 8'hbe == _T_2[7:0] ? image_190 : _GEN_189; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_383 = 8'hbf == _T_4[7:0] ? io_pixelVal_in_0 : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_575 = 8'hbf == _T_8[7:0] ? io_pixelVal_in_1 : _GEN_383; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_767 = 8'hbf == _T_11[7:0] ? io_pixelVal_in_2 : _GEN_575; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_959 = 8'hbf == _T_14[7:0] ? io_pixelVal_in_3 : _GEN_767; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1151 = 8'hbf == _T_17[7:0] ? io_pixelVal_in_4 : _GEN_959; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1343 = 8'hbf == _T_20[7:0] ? io_pixelVal_in_5 : _GEN_1151; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1535 = 8'hbf == _T_23[7:0] ? io_pixelVal_in_6 : _GEN_1343; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_1727 = 8'hbf == _T_26[7:0] ? io_pixelVal_in_7 : _GEN_1535; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_191 = io_valid_in ? _GEN_1727 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [31:0] _T_29 = pixelIndex + 32'h8; // @[VideoBuffer.scala 37:42]
  wire [8:0] _T_30 = 5'h10 * 5'hc; // @[VideoBuffer.scala 38:42]
  wire [31:0] _GEN_1923 = {{23'd0}, _T_30}; // @[VideoBuffer.scala 38:25]
  wire  _T_31 = pixelIndex == _GEN_1923; // @[VideoBuffer.scala 38:25]
  assign io_pixelVal_out = 8'hbf == _T_2[7:0] ? image_191 : _GEN_190; // @[VideoBuffer.scala 29:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pixelIndex = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      pixelIndex <= 32'h0;
    end else if (io_valid_in) begin
      if (_T_31) begin
        pixelIndex <= 32'h0;
      end else begin
        pixelIndex <= _T_29;
      end
    end
  end
endmodule
