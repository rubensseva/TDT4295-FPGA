module VideoBuffer(
  input         clock,
  input         reset,
  input  [15:0] io_pixelVal_in_0,
  input  [15:0] io_pixelVal_in_1,
  input  [15:0] io_pixelVal_in_2,
  input  [15:0] io_pixelVal_in_3,
  input  [15:0] io_pixelVal_in_4,
  input  [15:0] io_pixelVal_in_5,
  input  [15:0] io_pixelVal_in_6,
  input  [15:0] io_pixelVal_in_7,
  input  [15:0] io_pixelVal_in_8,
  input  [15:0] io_pixelVal_in_9,
  input  [15:0] io_pixelVal_in_10,
  input  [15:0] io_pixelVal_in_11,
  input  [15:0] io_pixelVal_in_12,
  input  [15:0] io_pixelVal_in_13,
  input  [15:0] io_pixelVal_in_14,
  input  [15:0] io_pixelVal_in_15,
  input  [15:0] io_pixelVal_in_16,
  input  [15:0] io_pixelVal_in_17,
  input         io_valid_in,
  input  [10:0] io_rowIndex,
  input  [10:0] io_colIndex,
  output [15:0] io_pixelVal_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [13:0] _T = io_rowIndex * 11'h6; // @[VideoBuffer.scala 29:46]
  wire [13:0] _GEN_962 = {{3'd0}, io_colIndex}; // @[VideoBuffer.scala 29:61]
  wire [13:0] _T_2 = _T + _GEN_962; // @[VideoBuffer.scala 29:61]
  reg [31:0] pixelIndex; // @[VideoBuffer.scala 31:33]
  wire [31:0] _T_56 = pixelIndex + 32'h11; // @[VideoBuffer.scala 35:42]
  wire [31:0] _T_53 = pixelIndex + 32'h10; // @[VideoBuffer.scala 35:42]
  wire [31:0] _T_50 = pixelIndex + 32'hf; // @[VideoBuffer.scala 35:42]
  wire [31:0] _T_47 = pixelIndex + 32'he; // @[VideoBuffer.scala 35:42]
  wire [31:0] _T_44 = pixelIndex + 32'hd; // @[VideoBuffer.scala 35:42]
  wire [31:0] _T_41 = pixelIndex + 32'hc; // @[VideoBuffer.scala 35:42]
  wire [31:0] _T_38 = pixelIndex + 32'hb; // @[VideoBuffer.scala 35:42]
  wire [31:0] _T_35 = pixelIndex + 32'ha; // @[VideoBuffer.scala 35:42]
  wire [31:0] _T_32 = pixelIndex + 32'h9; // @[VideoBuffer.scala 35:42]
  wire [31:0] _T_29 = pixelIndex + 32'h8; // @[VideoBuffer.scala 35:42]
  wire [31:0] _T_26 = pixelIndex + 32'h7; // @[VideoBuffer.scala 35:42]
  wire [31:0] _T_23 = pixelIndex + 32'h6; // @[VideoBuffer.scala 35:42]
  wire [31:0] _T_20 = pixelIndex + 32'h5; // @[VideoBuffer.scala 35:42]
  wire [31:0] _T_17 = pixelIndex + 32'h4; // @[VideoBuffer.scala 35:42]
  wire [31:0] _T_14 = pixelIndex + 32'h3; // @[VideoBuffer.scala 35:42]
  wire [31:0] _T_11 = pixelIndex + 32'h2; // @[VideoBuffer.scala 35:42]
  wire [31:0] _T_8 = pixelIndex + 32'h1; // @[VideoBuffer.scala 35:42]
  wire [32:0] _T_4 = {{1'd0}, pixelIndex}; // @[VideoBuffer.scala 35:42]
  wire [3:0] _GEN_48 = 6'h0 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_96 = 6'h0 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_48; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_144 = 6'h0 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_96; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_192 = 6'h0 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_144; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_240 = 6'h0 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_192; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_288 = 6'h0 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_240; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_336 = 6'h0 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_288; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_384 = 6'h0 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_336; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_432 = 6'h0 == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_384; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_480 = 6'h0 == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_432; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_528 = 6'h0 == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_480; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_576 = 6'h0 == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_528; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_624 = 6'h0 == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_576; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_672 = 6'h0 == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_624; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_720 = 6'h0 == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_672; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_768 = 6'h0 == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_720; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_816 = 6'h0 == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_768; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_864 = 6'h0 == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_816; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_0 = io_valid_in ? _GEN_864 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_49 = 6'h1 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_97 = 6'h1 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_49; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_145 = 6'h1 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_97; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_193 = 6'h1 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_145; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_241 = 6'h1 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_193; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_289 = 6'h1 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_241; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_337 = 6'h1 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_289; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_385 = 6'h1 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_337; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_433 = 6'h1 == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_385; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_481 = 6'h1 == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_433; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_529 = 6'h1 == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_481; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_577 = 6'h1 == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_529; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_625 = 6'h1 == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_577; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_673 = 6'h1 == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_625; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_721 = 6'h1 == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_673; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_769 = 6'h1 == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_721; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_817 = 6'h1 == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_769; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_865 = 6'h1 == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_817; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1 = io_valid_in ? _GEN_865 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1 = 6'h1 == _T_2[5:0] ? image_1 : image_0; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_50 = 6'h2 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_98 = 6'h2 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_50; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_146 = 6'h2 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_98; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_194 = 6'h2 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_146; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_242 = 6'h2 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_194; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_290 = 6'h2 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_242; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_338 = 6'h2 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_290; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_386 = 6'h2 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_338; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_434 = 6'h2 == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_386; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_482 = 6'h2 == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_434; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_530 = 6'h2 == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_482; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_578 = 6'h2 == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_530; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_626 = 6'h2 == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_578; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_674 = 6'h2 == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_626; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_722 = 6'h2 == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_674; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_770 = 6'h2 == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_722; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_818 = 6'h2 == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_770; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_866 = 6'h2 == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_818; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2 = io_valid_in ? _GEN_866 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2 = 6'h2 == _T_2[5:0] ? image_2 : _GEN_1; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_51 = 6'h3 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_99 = 6'h3 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_51; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_147 = 6'h3 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_99; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_195 = 6'h3 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_147; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_243 = 6'h3 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_195; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_291 = 6'h3 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_243; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_339 = 6'h3 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_291; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_387 = 6'h3 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_339; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_435 = 6'h3 == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_387; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_483 = 6'h3 == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_435; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_531 = 6'h3 == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_483; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_579 = 6'h3 == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_531; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_627 = 6'h3 == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_579; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_675 = 6'h3 == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_627; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_723 = 6'h3 == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_675; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_771 = 6'h3 == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_723; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_819 = 6'h3 == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_771; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_867 = 6'h3 == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_819; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3 = io_valid_in ? _GEN_867 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3 = 6'h3 == _T_2[5:0] ? image_3 : _GEN_2; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_52 = 6'h4 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_100 = 6'h4 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_52; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_148 = 6'h4 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_100; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_196 = 6'h4 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_148; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_244 = 6'h4 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_196; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_292 = 6'h4 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_244; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_340 = 6'h4 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_292; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_388 = 6'h4 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_340; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_436 = 6'h4 == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_388; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_484 = 6'h4 == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_436; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_532 = 6'h4 == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_484; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_580 = 6'h4 == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_532; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_628 = 6'h4 == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_580; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_676 = 6'h4 == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_628; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_724 = 6'h4 == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_676; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_772 = 6'h4 == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_724; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_820 = 6'h4 == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_772; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_868 = 6'h4 == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_820; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_4 = io_valid_in ? _GEN_868 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_4 = 6'h4 == _T_2[5:0] ? image_4 : _GEN_3; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_53 = 6'h5 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_101 = 6'h5 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_53; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_149 = 6'h5 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_101; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_197 = 6'h5 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_149; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_245 = 6'h5 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_197; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_293 = 6'h5 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_245; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_341 = 6'h5 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_293; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_389 = 6'h5 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_341; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_437 = 6'h5 == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_389; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_485 = 6'h5 == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_437; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_533 = 6'h5 == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_485; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_581 = 6'h5 == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_533; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_629 = 6'h5 == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_581; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_677 = 6'h5 == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_629; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_725 = 6'h5 == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_677; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_773 = 6'h5 == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_725; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_821 = 6'h5 == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_773; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_869 = 6'h5 == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_821; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_5 = io_valid_in ? _GEN_869 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_5 = 6'h5 == _T_2[5:0] ? image_5 : _GEN_4; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_54 = 6'h6 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_102 = 6'h6 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_54; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_150 = 6'h6 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_102; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_198 = 6'h6 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_150; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_246 = 6'h6 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_198; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_294 = 6'h6 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_246; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_342 = 6'h6 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_294; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_390 = 6'h6 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_342; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_438 = 6'h6 == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_390; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_486 = 6'h6 == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_438; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_534 = 6'h6 == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_486; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_582 = 6'h6 == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_534; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_630 = 6'h6 == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_582; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_678 = 6'h6 == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_630; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_726 = 6'h6 == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_678; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_774 = 6'h6 == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_726; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_822 = 6'h6 == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_774; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_870 = 6'h6 == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_822; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_6 = io_valid_in ? _GEN_870 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_6 = 6'h6 == _T_2[5:0] ? image_6 : _GEN_5; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_55 = 6'h7 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_103 = 6'h7 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_55; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_151 = 6'h7 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_103; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_199 = 6'h7 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_151; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_247 = 6'h7 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_199; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_295 = 6'h7 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_247; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_343 = 6'h7 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_295; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_391 = 6'h7 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_343; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_439 = 6'h7 == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_391; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_487 = 6'h7 == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_439; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_535 = 6'h7 == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_487; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_583 = 6'h7 == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_535; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_631 = 6'h7 == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_583; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_679 = 6'h7 == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_631; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_727 = 6'h7 == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_679; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_775 = 6'h7 == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_727; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_823 = 6'h7 == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_775; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_871 = 6'h7 == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_823; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_7 = io_valid_in ? _GEN_871 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_7 = 6'h7 == _T_2[5:0] ? image_7 : _GEN_6; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_56 = 6'h8 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_104 = 6'h8 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_56; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_152 = 6'h8 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_104; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_200 = 6'h8 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_152; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_248 = 6'h8 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_200; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_296 = 6'h8 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_248; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_344 = 6'h8 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_296; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_392 = 6'h8 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_344; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_440 = 6'h8 == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_392; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_488 = 6'h8 == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_440; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_536 = 6'h8 == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_488; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_584 = 6'h8 == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_536; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_632 = 6'h8 == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_584; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_680 = 6'h8 == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_632; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_728 = 6'h8 == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_680; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_776 = 6'h8 == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_728; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_824 = 6'h8 == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_776; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_872 = 6'h8 == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_824; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_8 = io_valid_in ? _GEN_872 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_8 = 6'h8 == _T_2[5:0] ? image_8 : _GEN_7; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_57 = 6'h9 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_105 = 6'h9 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_57; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_153 = 6'h9 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_105; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_201 = 6'h9 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_153; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_249 = 6'h9 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_201; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_297 = 6'h9 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_249; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_345 = 6'h9 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_297; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_393 = 6'h9 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_345; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_441 = 6'h9 == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_393; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_489 = 6'h9 == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_441; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_537 = 6'h9 == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_489; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_585 = 6'h9 == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_537; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_633 = 6'h9 == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_585; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_681 = 6'h9 == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_633; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_729 = 6'h9 == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_681; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_777 = 6'h9 == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_729; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_825 = 6'h9 == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_777; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_873 = 6'h9 == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_825; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_9 = io_valid_in ? _GEN_873 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_9 = 6'h9 == _T_2[5:0] ? image_9 : _GEN_8; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_58 = 6'ha == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_106 = 6'ha == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_58; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_154 = 6'ha == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_106; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_202 = 6'ha == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_154; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_250 = 6'ha == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_202; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_298 = 6'ha == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_250; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_346 = 6'ha == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_298; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_394 = 6'ha == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_346; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_442 = 6'ha == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_394; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_490 = 6'ha == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_442; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_538 = 6'ha == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_490; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_586 = 6'ha == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_538; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_634 = 6'ha == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_586; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_682 = 6'ha == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_634; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_730 = 6'ha == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_682; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_778 = 6'ha == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_730; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_826 = 6'ha == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_778; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_874 = 6'ha == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_826; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_10 = io_valid_in ? _GEN_874 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_10 = 6'ha == _T_2[5:0] ? image_10 : _GEN_9; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_59 = 6'hb == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_107 = 6'hb == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_59; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_155 = 6'hb == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_107; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_203 = 6'hb == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_155; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_251 = 6'hb == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_203; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_299 = 6'hb == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_251; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_347 = 6'hb == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_299; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_395 = 6'hb == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_347; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_443 = 6'hb == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_395; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_491 = 6'hb == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_443; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_539 = 6'hb == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_491; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_587 = 6'hb == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_539; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_635 = 6'hb == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_587; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_683 = 6'hb == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_635; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_731 = 6'hb == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_683; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_779 = 6'hb == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_731; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_827 = 6'hb == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_779; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_875 = 6'hb == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_827; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_11 = io_valid_in ? _GEN_875 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_11 = 6'hb == _T_2[5:0] ? image_11 : _GEN_10; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_60 = 6'hc == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_108 = 6'hc == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_60; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_156 = 6'hc == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_108; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_204 = 6'hc == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_156; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_252 = 6'hc == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_204; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_300 = 6'hc == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_252; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_348 = 6'hc == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_300; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_396 = 6'hc == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_348; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_444 = 6'hc == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_396; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_492 = 6'hc == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_444; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_540 = 6'hc == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_492; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_588 = 6'hc == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_540; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_636 = 6'hc == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_588; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_684 = 6'hc == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_636; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_732 = 6'hc == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_684; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_780 = 6'hc == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_732; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_828 = 6'hc == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_780; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_876 = 6'hc == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_828; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_12 = io_valid_in ? _GEN_876 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_12 = 6'hc == _T_2[5:0] ? image_12 : _GEN_11; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_61 = 6'hd == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_109 = 6'hd == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_61; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_157 = 6'hd == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_109; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_205 = 6'hd == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_157; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_253 = 6'hd == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_205; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_301 = 6'hd == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_253; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_349 = 6'hd == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_301; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_397 = 6'hd == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_349; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_445 = 6'hd == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_397; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_493 = 6'hd == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_445; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_541 = 6'hd == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_493; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_589 = 6'hd == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_541; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_637 = 6'hd == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_589; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_685 = 6'hd == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_637; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_733 = 6'hd == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_685; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_781 = 6'hd == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_733; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_829 = 6'hd == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_781; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_877 = 6'hd == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_829; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_13 = io_valid_in ? _GEN_877 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_13 = 6'hd == _T_2[5:0] ? image_13 : _GEN_12; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_62 = 6'he == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_110 = 6'he == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_62; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_158 = 6'he == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_110; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_206 = 6'he == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_158; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_254 = 6'he == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_206; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_302 = 6'he == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_254; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_350 = 6'he == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_302; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_398 = 6'he == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_350; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_446 = 6'he == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_398; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_494 = 6'he == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_446; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_542 = 6'he == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_494; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_590 = 6'he == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_542; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_638 = 6'he == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_590; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_686 = 6'he == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_638; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_734 = 6'he == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_686; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_782 = 6'he == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_734; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_830 = 6'he == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_782; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_878 = 6'he == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_830; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_14 = io_valid_in ? _GEN_878 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_14 = 6'he == _T_2[5:0] ? image_14 : _GEN_13; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_63 = 6'hf == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_111 = 6'hf == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_63; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_159 = 6'hf == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_111; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_207 = 6'hf == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_159; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_255 = 6'hf == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_207; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_303 = 6'hf == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_255; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_351 = 6'hf == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_303; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_399 = 6'hf == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_351; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_447 = 6'hf == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_399; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_495 = 6'hf == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_447; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_543 = 6'hf == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_495; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_591 = 6'hf == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_543; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_639 = 6'hf == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_591; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_687 = 6'hf == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_639; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_735 = 6'hf == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_687; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_783 = 6'hf == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_735; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_831 = 6'hf == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_783; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_879 = 6'hf == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_831; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_15 = io_valid_in ? _GEN_879 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_15 = 6'hf == _T_2[5:0] ? image_15 : _GEN_14; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_64 = 6'h10 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_112 = 6'h10 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_64; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_160 = 6'h10 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_112; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_208 = 6'h10 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_160; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_256 = 6'h10 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_208; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_304 = 6'h10 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_256; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_352 = 6'h10 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_304; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_400 = 6'h10 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_352; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_448 = 6'h10 == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_400; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_496 = 6'h10 == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_448; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_544 = 6'h10 == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_496; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_592 = 6'h10 == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_544; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_640 = 6'h10 == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_592; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_688 = 6'h10 == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_640; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_736 = 6'h10 == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_688; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_784 = 6'h10 == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_736; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_832 = 6'h10 == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_784; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_880 = 6'h10 == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_832; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_16 = io_valid_in ? _GEN_880 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_16 = 6'h10 == _T_2[5:0] ? image_16 : _GEN_15; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_65 = 6'h11 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_113 = 6'h11 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_65; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_161 = 6'h11 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_113; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_209 = 6'h11 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_161; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_257 = 6'h11 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_209; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_305 = 6'h11 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_257; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_353 = 6'h11 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_305; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_401 = 6'h11 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_353; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_449 = 6'h11 == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_401; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_497 = 6'h11 == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_449; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_545 = 6'h11 == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_497; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_593 = 6'h11 == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_545; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_641 = 6'h11 == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_593; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_689 = 6'h11 == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_641; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_737 = 6'h11 == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_689; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_785 = 6'h11 == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_737; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_833 = 6'h11 == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_785; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_881 = 6'h11 == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_833; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_17 = io_valid_in ? _GEN_881 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_17 = 6'h11 == _T_2[5:0] ? image_17 : _GEN_16; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_66 = 6'h12 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'hf; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_114 = 6'h12 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_66; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_162 = 6'h12 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_114; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_210 = 6'h12 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_162; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_258 = 6'h12 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_210; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_306 = 6'h12 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_258; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_354 = 6'h12 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_306; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_402 = 6'h12 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_354; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_450 = 6'h12 == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_402; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_498 = 6'h12 == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_450; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_546 = 6'h12 == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_498; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_594 = 6'h12 == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_546; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_642 = 6'h12 == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_594; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_690 = 6'h12 == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_642; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_738 = 6'h12 == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_690; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_786 = 6'h12 == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_738; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_834 = 6'h12 == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_786; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_882 = 6'h12 == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_834; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_18 = io_valid_in ? _GEN_882 : 4'hf; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_18 = 6'h12 == _T_2[5:0] ? image_18 : _GEN_17; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_67 = 6'h13 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'hf; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_115 = 6'h13 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_67; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_163 = 6'h13 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_115; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_211 = 6'h13 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_163; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_259 = 6'h13 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_211; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_307 = 6'h13 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_259; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_355 = 6'h13 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_307; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_403 = 6'h13 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_355; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_451 = 6'h13 == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_403; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_499 = 6'h13 == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_451; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_547 = 6'h13 == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_499; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_595 = 6'h13 == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_547; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_643 = 6'h13 == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_595; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_691 = 6'h13 == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_643; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_739 = 6'h13 == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_691; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_787 = 6'h13 == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_739; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_835 = 6'h13 == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_787; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_883 = 6'h13 == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_835; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_19 = io_valid_in ? _GEN_883 : 4'hf; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_19 = 6'h13 == _T_2[5:0] ? image_19 : _GEN_18; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_68 = 6'h14 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'hf; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_116 = 6'h14 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_68; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_164 = 6'h14 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_116; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_212 = 6'h14 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_164; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_260 = 6'h14 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_212; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_308 = 6'h14 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_260; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_356 = 6'h14 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_308; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_404 = 6'h14 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_356; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_452 = 6'h14 == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_404; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_500 = 6'h14 == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_452; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_548 = 6'h14 == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_500; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_596 = 6'h14 == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_548; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_644 = 6'h14 == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_596; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_692 = 6'h14 == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_644; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_740 = 6'h14 == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_692; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_788 = 6'h14 == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_740; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_836 = 6'h14 == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_788; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_884 = 6'h14 == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_836; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_20 = io_valid_in ? _GEN_884 : 4'hf; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_20 = 6'h14 == _T_2[5:0] ? image_20 : _GEN_19; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_69 = 6'h15 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_117 = 6'h15 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_69; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_165 = 6'h15 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_117; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_213 = 6'h15 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_165; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_261 = 6'h15 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_213; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_309 = 6'h15 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_261; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_357 = 6'h15 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_309; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_405 = 6'h15 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_357; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_453 = 6'h15 == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_405; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_501 = 6'h15 == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_453; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_549 = 6'h15 == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_501; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_597 = 6'h15 == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_549; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_645 = 6'h15 == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_597; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_693 = 6'h15 == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_645; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_741 = 6'h15 == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_693; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_789 = 6'h15 == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_741; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_837 = 6'h15 == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_789; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_885 = 6'h15 == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_837; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_21 = io_valid_in ? _GEN_885 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_21 = 6'h15 == _T_2[5:0] ? image_21 : _GEN_20; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_70 = 6'h16 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_118 = 6'h16 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_70; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_166 = 6'h16 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_118; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_214 = 6'h16 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_166; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_262 = 6'h16 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_214; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_310 = 6'h16 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_262; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_358 = 6'h16 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_310; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_406 = 6'h16 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_358; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_454 = 6'h16 == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_406; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_502 = 6'h16 == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_454; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_550 = 6'h16 == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_502; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_598 = 6'h16 == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_550; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_646 = 6'h16 == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_598; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_694 = 6'h16 == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_646; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_742 = 6'h16 == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_694; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_790 = 6'h16 == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_742; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_838 = 6'h16 == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_790; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_886 = 6'h16 == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_838; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_22 = io_valid_in ? _GEN_886 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_22 = 6'h16 == _T_2[5:0] ? image_22 : _GEN_21; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_71 = 6'h17 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_119 = 6'h17 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_71; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_167 = 6'h17 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_119; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_215 = 6'h17 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_167; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_263 = 6'h17 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_215; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_311 = 6'h17 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_263; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_359 = 6'h17 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_311; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_407 = 6'h17 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_359; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_455 = 6'h17 == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_407; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_503 = 6'h17 == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_455; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_551 = 6'h17 == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_503; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_599 = 6'h17 == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_551; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_647 = 6'h17 == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_599; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_695 = 6'h17 == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_647; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_743 = 6'h17 == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_695; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_791 = 6'h17 == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_743; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_839 = 6'h17 == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_791; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_887 = 6'h17 == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_839; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_23 = io_valid_in ? _GEN_887 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_23 = 6'h17 == _T_2[5:0] ? image_23 : _GEN_22; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_72 = 6'h18 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_120 = 6'h18 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_72; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_168 = 6'h18 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_120; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_216 = 6'h18 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_168; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_264 = 6'h18 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_216; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_312 = 6'h18 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_264; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_360 = 6'h18 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_312; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_408 = 6'h18 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_360; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_456 = 6'h18 == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_408; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_504 = 6'h18 == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_456; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_552 = 6'h18 == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_504; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_600 = 6'h18 == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_552; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_648 = 6'h18 == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_600; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_696 = 6'h18 == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_648; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_744 = 6'h18 == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_696; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_792 = 6'h18 == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_744; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_840 = 6'h18 == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_792; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_888 = 6'h18 == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_840; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_24 = io_valid_in ? _GEN_888 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_24 = 6'h18 == _T_2[5:0] ? image_24 : _GEN_23; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_73 = 6'h19 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_121 = 6'h19 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_73; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_169 = 6'h19 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_121; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_217 = 6'h19 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_169; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_265 = 6'h19 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_217; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_313 = 6'h19 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_265; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_361 = 6'h19 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_313; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_409 = 6'h19 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_361; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_457 = 6'h19 == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_409; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_505 = 6'h19 == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_457; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_553 = 6'h19 == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_505; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_601 = 6'h19 == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_553; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_649 = 6'h19 == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_601; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_697 = 6'h19 == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_649; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_745 = 6'h19 == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_697; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_793 = 6'h19 == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_745; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_841 = 6'h19 == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_793; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_889 = 6'h19 == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_841; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_25 = io_valid_in ? _GEN_889 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_25 = 6'h19 == _T_2[5:0] ? image_25 : _GEN_24; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_74 = 6'h1a == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'hf; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_122 = 6'h1a == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_74; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_170 = 6'h1a == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_122; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_218 = 6'h1a == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_170; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_266 = 6'h1a == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_218; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_314 = 6'h1a == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_266; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_362 = 6'h1a == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_314; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_410 = 6'h1a == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_362; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_458 = 6'h1a == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_410; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_506 = 6'h1a == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_458; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_554 = 6'h1a == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_506; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_602 = 6'h1a == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_554; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_650 = 6'h1a == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_602; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_698 = 6'h1a == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_650; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_746 = 6'h1a == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_698; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_794 = 6'h1a == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_746; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_842 = 6'h1a == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_794; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_890 = 6'h1a == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_842; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_26 = io_valid_in ? _GEN_890 : 4'hf; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_26 = 6'h1a == _T_2[5:0] ? image_26 : _GEN_25; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_75 = 6'h1b == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'hf; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_123 = 6'h1b == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_75; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_171 = 6'h1b == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_123; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_219 = 6'h1b == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_171; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_267 = 6'h1b == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_219; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_315 = 6'h1b == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_267; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_363 = 6'h1b == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_315; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_411 = 6'h1b == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_363; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_459 = 6'h1b == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_411; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_507 = 6'h1b == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_459; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_555 = 6'h1b == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_507; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_603 = 6'h1b == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_555; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_651 = 6'h1b == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_603; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_699 = 6'h1b == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_651; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_747 = 6'h1b == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_699; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_795 = 6'h1b == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_747; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_843 = 6'h1b == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_795; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_891 = 6'h1b == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_843; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_27 = io_valid_in ? _GEN_891 : 4'hf; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_27 = 6'h1b == _T_2[5:0] ? image_27 : _GEN_26; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_76 = 6'h1c == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'hf; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_124 = 6'h1c == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_76; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_172 = 6'h1c == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_124; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_220 = 6'h1c == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_172; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_268 = 6'h1c == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_220; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_316 = 6'h1c == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_268; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_364 = 6'h1c == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_316; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_412 = 6'h1c == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_364; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_460 = 6'h1c == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_412; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_508 = 6'h1c == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_460; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_556 = 6'h1c == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_508; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_604 = 6'h1c == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_556; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_652 = 6'h1c == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_604; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_700 = 6'h1c == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_652; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_748 = 6'h1c == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_700; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_796 = 6'h1c == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_748; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_844 = 6'h1c == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_796; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_892 = 6'h1c == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_844; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_28 = io_valid_in ? _GEN_892 : 4'hf; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_28 = 6'h1c == _T_2[5:0] ? image_28 : _GEN_27; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_77 = 6'h1d == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_125 = 6'h1d == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_77; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_173 = 6'h1d == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_125; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_221 = 6'h1d == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_173; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_269 = 6'h1d == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_221; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_317 = 6'h1d == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_269; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_365 = 6'h1d == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_317; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_413 = 6'h1d == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_365; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_461 = 6'h1d == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_413; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_509 = 6'h1d == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_461; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_557 = 6'h1d == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_509; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_605 = 6'h1d == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_557; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_653 = 6'h1d == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_605; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_701 = 6'h1d == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_653; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_749 = 6'h1d == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_701; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_797 = 6'h1d == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_749; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_845 = 6'h1d == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_797; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_893 = 6'h1d == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_845; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_29 = io_valid_in ? _GEN_893 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_29 = 6'h1d == _T_2[5:0] ? image_29 : _GEN_28; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_78 = 6'h1e == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_126 = 6'h1e == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_78; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_174 = 6'h1e == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_126; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_222 = 6'h1e == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_174; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_270 = 6'h1e == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_222; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_318 = 6'h1e == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_270; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_366 = 6'h1e == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_318; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_414 = 6'h1e == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_366; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_462 = 6'h1e == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_414; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_510 = 6'h1e == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_462; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_558 = 6'h1e == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_510; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_606 = 6'h1e == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_558; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_654 = 6'h1e == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_606; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_702 = 6'h1e == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_654; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_750 = 6'h1e == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_702; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_798 = 6'h1e == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_750; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_846 = 6'h1e == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_798; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_894 = 6'h1e == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_846; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_30 = io_valid_in ? _GEN_894 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_30 = 6'h1e == _T_2[5:0] ? image_30 : _GEN_29; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_79 = 6'h1f == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_127 = 6'h1f == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_79; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_175 = 6'h1f == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_127; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_223 = 6'h1f == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_175; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_271 = 6'h1f == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_223; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_319 = 6'h1f == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_271; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_367 = 6'h1f == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_319; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_415 = 6'h1f == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_367; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_463 = 6'h1f == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_415; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_511 = 6'h1f == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_463; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_559 = 6'h1f == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_511; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_607 = 6'h1f == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_559; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_655 = 6'h1f == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_607; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_703 = 6'h1f == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_655; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_751 = 6'h1f == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_703; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_799 = 6'h1f == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_751; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_847 = 6'h1f == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_799; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_895 = 6'h1f == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_847; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_31 = io_valid_in ? _GEN_895 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_31 = 6'h1f == _T_2[5:0] ? image_31 : _GEN_30; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_80 = 6'h20 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_128 = 6'h20 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_80; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_176 = 6'h20 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_128; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_224 = 6'h20 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_176; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_272 = 6'h20 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_224; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_320 = 6'h20 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_272; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_368 = 6'h20 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_320; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_416 = 6'h20 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_368; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_464 = 6'h20 == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_416; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_512 = 6'h20 == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_464; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_560 = 6'h20 == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_512; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_608 = 6'h20 == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_560; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_656 = 6'h20 == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_608; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_704 = 6'h20 == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_656; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_752 = 6'h20 == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_704; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_800 = 6'h20 == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_752; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_848 = 6'h20 == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_800; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_896 = 6'h20 == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_848; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_32 = io_valid_in ? _GEN_896 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_32 = 6'h20 == _T_2[5:0] ? image_32 : _GEN_31; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_81 = 6'h21 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_129 = 6'h21 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_81; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_177 = 6'h21 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_129; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_225 = 6'h21 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_177; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_273 = 6'h21 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_225; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_321 = 6'h21 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_273; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_369 = 6'h21 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_321; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_417 = 6'h21 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_369; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_465 = 6'h21 == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_417; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_513 = 6'h21 == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_465; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_561 = 6'h21 == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_513; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_609 = 6'h21 == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_561; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_657 = 6'h21 == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_609; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_705 = 6'h21 == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_657; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_753 = 6'h21 == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_705; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_801 = 6'h21 == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_753; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_849 = 6'h21 == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_801; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_897 = 6'h21 == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_849; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_33 = io_valid_in ? _GEN_897 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_33 = 6'h21 == _T_2[5:0] ? image_33 : _GEN_32; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_82 = 6'h22 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'hf; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_130 = 6'h22 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_82; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_178 = 6'h22 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_130; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_226 = 6'h22 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_178; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_274 = 6'h22 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_226; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_322 = 6'h22 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_274; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_370 = 6'h22 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_322; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_418 = 6'h22 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_370; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_466 = 6'h22 == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_418; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_514 = 6'h22 == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_466; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_562 = 6'h22 == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_514; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_610 = 6'h22 == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_562; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_658 = 6'h22 == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_610; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_706 = 6'h22 == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_658; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_754 = 6'h22 == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_706; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_802 = 6'h22 == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_754; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_850 = 6'h22 == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_802; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_898 = 6'h22 == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_850; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_34 = io_valid_in ? _GEN_898 : 4'hf; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_34 = 6'h22 == _T_2[5:0] ? image_34 : _GEN_33; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_83 = 6'h23 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'hf; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_131 = 6'h23 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_83; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_179 = 6'h23 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_131; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_227 = 6'h23 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_179; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_275 = 6'h23 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_227; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_323 = 6'h23 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_275; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_371 = 6'h23 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_323; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_419 = 6'h23 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_371; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_467 = 6'h23 == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_419; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_515 = 6'h23 == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_467; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_563 = 6'h23 == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_515; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_611 = 6'h23 == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_563; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_659 = 6'h23 == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_611; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_707 = 6'h23 == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_659; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_755 = 6'h23 == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_707; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_803 = 6'h23 == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_755; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_851 = 6'h23 == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_803; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_899 = 6'h23 == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_851; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_35 = io_valid_in ? _GEN_899 : 4'hf; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_35 = 6'h23 == _T_2[5:0] ? image_35 : _GEN_34; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_84 = 6'h24 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'hf; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_132 = 6'h24 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_84; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_180 = 6'h24 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_132; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_228 = 6'h24 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_180; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_276 = 6'h24 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_228; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_324 = 6'h24 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_276; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_372 = 6'h24 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_324; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_420 = 6'h24 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_372; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_468 = 6'h24 == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_420; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_516 = 6'h24 == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_468; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_564 = 6'h24 == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_516; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_612 = 6'h24 == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_564; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_660 = 6'h24 == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_612; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_708 = 6'h24 == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_660; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_756 = 6'h24 == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_708; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_804 = 6'h24 == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_756; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_852 = 6'h24 == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_804; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_900 = 6'h24 == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_852; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_36 = io_valid_in ? _GEN_900 : 4'hf; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_36 = 6'h24 == _T_2[5:0] ? image_36 : _GEN_35; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_85 = 6'h25 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_133 = 6'h25 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_85; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_181 = 6'h25 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_133; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_229 = 6'h25 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_181; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_277 = 6'h25 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_229; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_325 = 6'h25 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_277; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_373 = 6'h25 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_325; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_421 = 6'h25 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_373; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_469 = 6'h25 == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_421; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_517 = 6'h25 == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_469; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_565 = 6'h25 == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_517; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_613 = 6'h25 == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_565; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_661 = 6'h25 == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_613; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_709 = 6'h25 == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_661; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_757 = 6'h25 == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_709; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_805 = 6'h25 == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_757; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_853 = 6'h25 == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_805; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_901 = 6'h25 == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_853; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_37 = io_valid_in ? _GEN_901 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_37 = 6'h25 == _T_2[5:0] ? image_37 : _GEN_36; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_86 = 6'h26 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_134 = 6'h26 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_86; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_182 = 6'h26 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_134; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_230 = 6'h26 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_182; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_278 = 6'h26 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_230; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_326 = 6'h26 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_278; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_374 = 6'h26 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_326; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_422 = 6'h26 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_374; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_470 = 6'h26 == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_422; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_518 = 6'h26 == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_470; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_566 = 6'h26 == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_518; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_614 = 6'h26 == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_566; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_662 = 6'h26 == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_614; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_710 = 6'h26 == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_662; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_758 = 6'h26 == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_710; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_806 = 6'h26 == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_758; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_854 = 6'h26 == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_806; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_902 = 6'h26 == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_854; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_38 = io_valid_in ? _GEN_902 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_38 = 6'h26 == _T_2[5:0] ? image_38 : _GEN_37; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_87 = 6'h27 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_135 = 6'h27 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_87; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_183 = 6'h27 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_135; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_231 = 6'h27 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_183; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_279 = 6'h27 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_231; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_327 = 6'h27 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_279; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_375 = 6'h27 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_327; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_423 = 6'h27 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_375; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_471 = 6'h27 == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_423; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_519 = 6'h27 == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_471; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_567 = 6'h27 == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_519; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_615 = 6'h27 == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_567; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_663 = 6'h27 == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_615; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_711 = 6'h27 == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_663; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_759 = 6'h27 == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_711; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_807 = 6'h27 == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_759; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_855 = 6'h27 == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_807; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_903 = 6'h27 == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_855; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_39 = io_valid_in ? _GEN_903 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_39 = 6'h27 == _T_2[5:0] ? image_39 : _GEN_38; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_88 = 6'h28 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_136 = 6'h28 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_88; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_184 = 6'h28 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_136; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_232 = 6'h28 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_184; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_280 = 6'h28 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_232; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_328 = 6'h28 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_280; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_376 = 6'h28 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_328; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_424 = 6'h28 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_376; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_472 = 6'h28 == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_424; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_520 = 6'h28 == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_472; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_568 = 6'h28 == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_520; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_616 = 6'h28 == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_568; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_664 = 6'h28 == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_616; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_712 = 6'h28 == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_664; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_760 = 6'h28 == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_712; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_808 = 6'h28 == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_760; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_856 = 6'h28 == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_808; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_904 = 6'h28 == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_856; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_40 = io_valid_in ? _GEN_904 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_40 = 6'h28 == _T_2[5:0] ? image_40 : _GEN_39; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_89 = 6'h29 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_137 = 6'h29 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_89; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_185 = 6'h29 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_137; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_233 = 6'h29 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_185; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_281 = 6'h29 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_233; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_329 = 6'h29 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_281; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_377 = 6'h29 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_329; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_425 = 6'h29 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_377; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_473 = 6'h29 == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_425; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_521 = 6'h29 == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_473; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_569 = 6'h29 == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_521; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_617 = 6'h29 == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_569; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_665 = 6'h29 == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_617; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_713 = 6'h29 == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_665; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_761 = 6'h29 == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_713; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_809 = 6'h29 == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_761; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_857 = 6'h29 == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_809; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_905 = 6'h29 == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_857; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_41 = io_valid_in ? _GEN_905 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_41 = 6'h29 == _T_2[5:0] ? image_41 : _GEN_40; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_90 = 6'h2a == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_138 = 6'h2a == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_90; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_186 = 6'h2a == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_138; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_234 = 6'h2a == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_186; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_282 = 6'h2a == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_234; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_330 = 6'h2a == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_282; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_378 = 6'h2a == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_330; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_426 = 6'h2a == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_378; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_474 = 6'h2a == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_426; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_522 = 6'h2a == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_474; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_570 = 6'h2a == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_522; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_618 = 6'h2a == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_570; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_666 = 6'h2a == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_618; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_714 = 6'h2a == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_666; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_762 = 6'h2a == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_714; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_810 = 6'h2a == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_762; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_858 = 6'h2a == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_810; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_906 = 6'h2a == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_858; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_42 = io_valid_in ? _GEN_906 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_42 = 6'h2a == _T_2[5:0] ? image_42 : _GEN_41; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_91 = 6'h2b == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_139 = 6'h2b == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_91; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_187 = 6'h2b == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_139; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_235 = 6'h2b == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_187; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_283 = 6'h2b == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_235; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_331 = 6'h2b == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_283; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_379 = 6'h2b == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_331; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_427 = 6'h2b == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_379; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_475 = 6'h2b == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_427; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_523 = 6'h2b == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_475; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_571 = 6'h2b == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_523; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_619 = 6'h2b == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_571; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_667 = 6'h2b == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_619; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_715 = 6'h2b == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_667; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_763 = 6'h2b == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_715; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_811 = 6'h2b == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_763; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_859 = 6'h2b == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_811; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_907 = 6'h2b == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_859; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_43 = io_valid_in ? _GEN_907 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_43 = 6'h2b == _T_2[5:0] ? image_43 : _GEN_42; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_92 = 6'h2c == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_140 = 6'h2c == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_92; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_188 = 6'h2c == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_140; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_236 = 6'h2c == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_188; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_284 = 6'h2c == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_236; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_332 = 6'h2c == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_284; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_380 = 6'h2c == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_332; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_428 = 6'h2c == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_380; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_476 = 6'h2c == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_428; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_524 = 6'h2c == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_476; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_572 = 6'h2c == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_524; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_620 = 6'h2c == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_572; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_668 = 6'h2c == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_620; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_716 = 6'h2c == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_668; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_764 = 6'h2c == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_716; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_812 = 6'h2c == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_764; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_860 = 6'h2c == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_812; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_908 = 6'h2c == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_860; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_44 = io_valid_in ? _GEN_908 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_44 = 6'h2c == _T_2[5:0] ? image_44 : _GEN_43; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_93 = 6'h2d == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_141 = 6'h2d == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_93; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_189 = 6'h2d == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_141; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_237 = 6'h2d == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_189; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_285 = 6'h2d == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_237; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_333 = 6'h2d == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_285; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_381 = 6'h2d == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_333; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_429 = 6'h2d == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_381; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_477 = 6'h2d == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_429; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_525 = 6'h2d == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_477; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_573 = 6'h2d == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_525; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_621 = 6'h2d == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_573; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_669 = 6'h2d == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_621; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_717 = 6'h2d == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_669; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_765 = 6'h2d == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_717; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_813 = 6'h2d == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_765; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_861 = 6'h2d == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_813; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_909 = 6'h2d == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_861; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_45 = io_valid_in ? _GEN_909 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_45 = 6'h2d == _T_2[5:0] ? image_45 : _GEN_44; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_94 = 6'h2e == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_142 = 6'h2e == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_94; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_190 = 6'h2e == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_142; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_238 = 6'h2e == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_190; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_286 = 6'h2e == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_238; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_334 = 6'h2e == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_286; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_382 = 6'h2e == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_334; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_430 = 6'h2e == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_382; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_478 = 6'h2e == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_430; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_526 = 6'h2e == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_478; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_574 = 6'h2e == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_526; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_622 = 6'h2e == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_574; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_670 = 6'h2e == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_622; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_718 = 6'h2e == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_670; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_766 = 6'h2e == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_718; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_814 = 6'h2e == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_766; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_862 = 6'h2e == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_814; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_910 = 6'h2e == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_862; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_46 = io_valid_in ? _GEN_910 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_46 = 6'h2e == _T_2[5:0] ? image_46 : _GEN_45; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_95 = 6'h2f == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_143 = 6'h2f == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_95; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_191 = 6'h2f == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_143; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_239 = 6'h2f == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_191; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_287 = 6'h2f == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_239; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_335 = 6'h2f == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_287; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_383 = 6'h2f == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_335; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_431 = 6'h2f == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_383; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_479 = 6'h2f == _T_29[5:0] ? io_pixelVal_in_8[3:0] : _GEN_431; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_527 = 6'h2f == _T_32[5:0] ? io_pixelVal_in_9[3:0] : _GEN_479; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_575 = 6'h2f == _T_35[5:0] ? io_pixelVal_in_10[3:0] : _GEN_527; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_623 = 6'h2f == _T_38[5:0] ? io_pixelVal_in_11[3:0] : _GEN_575; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_671 = 6'h2f == _T_41[5:0] ? io_pixelVal_in_12[3:0] : _GEN_623; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_719 = 6'h2f == _T_44[5:0] ? io_pixelVal_in_13[3:0] : _GEN_671; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_767 = 6'h2f == _T_47[5:0] ? io_pixelVal_in_14[3:0] : _GEN_719; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_815 = 6'h2f == _T_50[5:0] ? io_pixelVal_in_15[3:0] : _GEN_767; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_863 = 6'h2f == _T_53[5:0] ? io_pixelVal_in_16[3:0] : _GEN_815; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_911 = 6'h2f == _T_56[5:0] ? io_pixelVal_in_17[3:0] : _GEN_863; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_47 = io_valid_in ? _GEN_911 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_47 = 6'h2f == _T_2[5:0] ? image_47 : _GEN_46; // @[VideoBuffer.scala 29:25]
  wire [31:0] _T_59 = pixelIndex + 32'h12; // @[VideoBuffer.scala 37:42]
  wire [5:0] _T_60 = 3'h6 * 3'h6; // @[VideoBuffer.scala 38:42]
  wire [31:0] _GEN_963 = {{26'd0}, _T_60}; // @[VideoBuffer.scala 38:25]
  wire  _T_61 = pixelIndex == _GEN_963; // @[VideoBuffer.scala 38:25]
  assign io_pixelVal_out = {{12'd0}, _GEN_47}; // @[VideoBuffer.scala 29:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pixelIndex = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      pixelIndex <= 32'h0;
    end else if (io_valid_in) begin
      if (_T_61) begin
        pixelIndex <= 32'h0;
      end else begin
        pixelIndex <= _T_59;
      end
    end
  end
endmodule
