module VideoBuffer(
  input         clock,
  input         reset,
  input  [15:0] io_pixelVal_in_0,
  input  [15:0] io_pixelVal_in_1,
  input  [15:0] io_pixelVal_in_2,
  input  [15:0] io_pixelVal_in_3,
  input  [15:0] io_pixelVal_in_4,
  input  [15:0] io_pixelVal_in_5,
  input  [15:0] io_pixelVal_in_6,
  input  [15:0] io_pixelVal_in_7,
  input         io_valid_in,
  input  [10:0] io_rowIndex,
  input  [10:0] io_colIndex,
  output [15:0] io_pixelVal_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [14:0] _T = io_rowIndex * 11'h8; // @[VideoBuffer.scala 29:46]
  wire [14:0] _GEN_482 = {{4'd0}, io_colIndex}; // @[VideoBuffer.scala 29:61]
  wire [14:0] _T_2 = _T + _GEN_482; // @[VideoBuffer.scala 29:61]
  reg [31:0] pixelIndex; // @[VideoBuffer.scala 31:33]
  wire [31:0] _T_26 = pixelIndex + 32'h7; // @[VideoBuffer.scala 35:42]
  wire [31:0] _T_23 = pixelIndex + 32'h6; // @[VideoBuffer.scala 35:42]
  wire [31:0] _T_20 = pixelIndex + 32'h5; // @[VideoBuffer.scala 35:42]
  wire [31:0] _T_17 = pixelIndex + 32'h4; // @[VideoBuffer.scala 35:42]
  wire [31:0] _T_14 = pixelIndex + 32'h3; // @[VideoBuffer.scala 35:42]
  wire [31:0] _T_11 = pixelIndex + 32'h2; // @[VideoBuffer.scala 35:42]
  wire [31:0] _T_8 = pixelIndex + 32'h1; // @[VideoBuffer.scala 35:42]
  wire [32:0] _T_4 = {{1'd0}, pixelIndex}; // @[VideoBuffer.scala 35:42]
  wire [3:0] _GEN_48 = 6'h0 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_96 = 6'h0 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_48; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_144 = 6'h0 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_96; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_192 = 6'h0 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_144; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_240 = 6'h0 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_192; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_288 = 6'h0 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_240; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_336 = 6'h0 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_288; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_384 = 6'h0 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_336; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_0 = io_valid_in ? _GEN_384 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_49 = 6'h1 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_97 = 6'h1 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_49; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_145 = 6'h1 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_97; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_193 = 6'h1 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_145; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_241 = 6'h1 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_193; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_289 = 6'h1 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_241; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_337 = 6'h1 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_289; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_385 = 6'h1 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_337; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_1 = io_valid_in ? _GEN_385 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_1 = 6'h1 == _T_2[5:0] ? image_1 : image_0; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_50 = 6'h2 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_98 = 6'h2 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_50; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_146 = 6'h2 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_98; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_194 = 6'h2 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_146; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_242 = 6'h2 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_194; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_290 = 6'h2 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_242; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_338 = 6'h2 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_290; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_386 = 6'h2 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_338; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_2 = io_valid_in ? _GEN_386 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_2 = 6'h2 == _T_2[5:0] ? image_2 : _GEN_1; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_51 = 6'h3 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_99 = 6'h3 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_51; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_147 = 6'h3 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_99; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_195 = 6'h3 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_147; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_243 = 6'h3 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_195; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_291 = 6'h3 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_243; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_339 = 6'h3 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_291; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_387 = 6'h3 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_339; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_3 = io_valid_in ? _GEN_387 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_3 = 6'h3 == _T_2[5:0] ? image_3 : _GEN_2; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_52 = 6'h4 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_100 = 6'h4 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_52; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_148 = 6'h4 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_100; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_196 = 6'h4 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_148; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_244 = 6'h4 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_196; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_292 = 6'h4 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_244; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_340 = 6'h4 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_292; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_388 = 6'h4 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_340; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_4 = io_valid_in ? _GEN_388 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_4 = 6'h4 == _T_2[5:0] ? image_4 : _GEN_3; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_53 = 6'h5 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_101 = 6'h5 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_53; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_149 = 6'h5 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_101; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_197 = 6'h5 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_149; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_245 = 6'h5 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_197; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_293 = 6'h5 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_245; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_341 = 6'h5 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_293; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_389 = 6'h5 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_341; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_5 = io_valid_in ? _GEN_389 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_5 = 6'h5 == _T_2[5:0] ? image_5 : _GEN_4; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_54 = 6'h6 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_102 = 6'h6 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_54; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_150 = 6'h6 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_102; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_198 = 6'h6 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_150; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_246 = 6'h6 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_198; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_294 = 6'h6 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_246; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_342 = 6'h6 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_294; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_390 = 6'h6 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_342; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_6 = io_valid_in ? _GEN_390 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_6 = 6'h6 == _T_2[5:0] ? image_6 : _GEN_5; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_55 = 6'h7 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_103 = 6'h7 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_55; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_151 = 6'h7 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_103; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_199 = 6'h7 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_151; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_247 = 6'h7 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_199; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_295 = 6'h7 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_247; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_343 = 6'h7 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_295; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_391 = 6'h7 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_343; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_7 = io_valid_in ? _GEN_391 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_7 = 6'h7 == _T_2[5:0] ? image_7 : _GEN_6; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_56 = 6'h8 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_104 = 6'h8 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_56; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_152 = 6'h8 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_104; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_200 = 6'h8 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_152; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_248 = 6'h8 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_200; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_296 = 6'h8 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_248; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_344 = 6'h8 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_296; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_392 = 6'h8 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_344; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_8 = io_valid_in ? _GEN_392 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_8 = 6'h8 == _T_2[5:0] ? image_8 : _GEN_7; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_57 = 6'h9 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_105 = 6'h9 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_57; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_153 = 6'h9 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_105; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_201 = 6'h9 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_153; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_249 = 6'h9 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_201; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_297 = 6'h9 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_249; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_345 = 6'h9 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_297; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_393 = 6'h9 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_345; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_9 = io_valid_in ? _GEN_393 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_9 = 6'h9 == _T_2[5:0] ? image_9 : _GEN_8; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_58 = 6'ha == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_106 = 6'ha == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_58; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_154 = 6'ha == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_106; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_202 = 6'ha == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_154; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_250 = 6'ha == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_202; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_298 = 6'ha == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_250; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_346 = 6'ha == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_298; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_394 = 6'ha == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_346; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_10 = io_valid_in ? _GEN_394 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_10 = 6'ha == _T_2[5:0] ? image_10 : _GEN_9; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_59 = 6'hb == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_107 = 6'hb == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_59; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_155 = 6'hb == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_107; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_203 = 6'hb == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_155; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_251 = 6'hb == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_203; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_299 = 6'hb == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_251; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_347 = 6'hb == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_299; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_395 = 6'hb == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_347; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_11 = io_valid_in ? _GEN_395 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_11 = 6'hb == _T_2[5:0] ? image_11 : _GEN_10; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_60 = 6'hc == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_108 = 6'hc == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_60; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_156 = 6'hc == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_108; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_204 = 6'hc == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_156; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_252 = 6'hc == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_204; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_300 = 6'hc == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_252; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_348 = 6'hc == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_300; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_396 = 6'hc == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_348; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_12 = io_valid_in ? _GEN_396 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_12 = 6'hc == _T_2[5:0] ? image_12 : _GEN_11; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_61 = 6'hd == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_109 = 6'hd == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_61; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_157 = 6'hd == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_109; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_205 = 6'hd == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_157; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_253 = 6'hd == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_205; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_301 = 6'hd == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_253; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_349 = 6'hd == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_301; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_397 = 6'hd == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_349; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_13 = io_valid_in ? _GEN_397 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_13 = 6'hd == _T_2[5:0] ? image_13 : _GEN_12; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_62 = 6'he == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_110 = 6'he == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_62; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_158 = 6'he == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_110; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_206 = 6'he == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_158; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_254 = 6'he == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_206; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_302 = 6'he == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_254; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_350 = 6'he == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_302; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_398 = 6'he == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_350; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_14 = io_valid_in ? _GEN_398 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_14 = 6'he == _T_2[5:0] ? image_14 : _GEN_13; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_63 = 6'hf == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_111 = 6'hf == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_63; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_159 = 6'hf == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_111; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_207 = 6'hf == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_159; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_255 = 6'hf == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_207; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_303 = 6'hf == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_255; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_351 = 6'hf == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_303; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_399 = 6'hf == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_351; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_15 = io_valid_in ? _GEN_399 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_15 = 6'hf == _T_2[5:0] ? image_15 : _GEN_14; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_64 = 6'h10 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_112 = 6'h10 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_64; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_160 = 6'h10 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_112; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_208 = 6'h10 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_160; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_256 = 6'h10 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_208; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_304 = 6'h10 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_256; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_352 = 6'h10 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_304; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_400 = 6'h10 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_352; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_16 = io_valid_in ? _GEN_400 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_16 = 6'h10 == _T_2[5:0] ? image_16 : _GEN_15; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_65 = 6'h11 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_113 = 6'h11 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_65; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_161 = 6'h11 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_113; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_209 = 6'h11 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_161; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_257 = 6'h11 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_209; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_305 = 6'h11 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_257; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_353 = 6'h11 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_305; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_401 = 6'h11 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_353; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_17 = io_valid_in ? _GEN_401 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_17 = 6'h11 == _T_2[5:0] ? image_17 : _GEN_16; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_66 = 6'h12 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'hf; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_114 = 6'h12 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_66; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_162 = 6'h12 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_114; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_210 = 6'h12 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_162; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_258 = 6'h12 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_210; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_306 = 6'h12 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_258; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_354 = 6'h12 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_306; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_402 = 6'h12 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_354; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_18 = io_valid_in ? _GEN_402 : 4'hf; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_18 = 6'h12 == _T_2[5:0] ? image_18 : _GEN_17; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_67 = 6'h13 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'hf; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_115 = 6'h13 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_67; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_163 = 6'h13 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_115; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_211 = 6'h13 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_163; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_259 = 6'h13 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_211; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_307 = 6'h13 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_259; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_355 = 6'h13 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_307; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_403 = 6'h13 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_355; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_19 = io_valid_in ? _GEN_403 : 4'hf; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_19 = 6'h13 == _T_2[5:0] ? image_19 : _GEN_18; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_68 = 6'h14 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'hf; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_116 = 6'h14 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_68; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_164 = 6'h14 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_116; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_212 = 6'h14 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_164; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_260 = 6'h14 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_212; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_308 = 6'h14 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_260; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_356 = 6'h14 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_308; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_404 = 6'h14 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_356; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_20 = io_valid_in ? _GEN_404 : 4'hf; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_20 = 6'h14 == _T_2[5:0] ? image_20 : _GEN_19; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_69 = 6'h15 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_117 = 6'h15 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_69; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_165 = 6'h15 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_117; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_213 = 6'h15 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_165; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_261 = 6'h15 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_213; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_309 = 6'h15 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_261; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_357 = 6'h15 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_309; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_405 = 6'h15 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_357; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_21 = io_valid_in ? _GEN_405 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_21 = 6'h15 == _T_2[5:0] ? image_21 : _GEN_20; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_70 = 6'h16 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_118 = 6'h16 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_70; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_166 = 6'h16 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_118; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_214 = 6'h16 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_166; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_262 = 6'h16 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_214; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_310 = 6'h16 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_262; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_358 = 6'h16 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_310; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_406 = 6'h16 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_358; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_22 = io_valid_in ? _GEN_406 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_22 = 6'h16 == _T_2[5:0] ? image_22 : _GEN_21; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_71 = 6'h17 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_119 = 6'h17 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_71; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_167 = 6'h17 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_119; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_215 = 6'h17 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_167; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_263 = 6'h17 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_215; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_311 = 6'h17 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_263; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_359 = 6'h17 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_311; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_407 = 6'h17 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_359; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_23 = io_valid_in ? _GEN_407 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_23 = 6'h17 == _T_2[5:0] ? image_23 : _GEN_22; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_72 = 6'h18 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_120 = 6'h18 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_72; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_168 = 6'h18 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_120; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_216 = 6'h18 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_168; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_264 = 6'h18 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_216; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_312 = 6'h18 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_264; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_360 = 6'h18 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_312; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_408 = 6'h18 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_360; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_24 = io_valid_in ? _GEN_408 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_24 = 6'h18 == _T_2[5:0] ? image_24 : _GEN_23; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_73 = 6'h19 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_121 = 6'h19 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_73; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_169 = 6'h19 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_121; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_217 = 6'h19 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_169; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_265 = 6'h19 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_217; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_313 = 6'h19 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_265; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_361 = 6'h19 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_313; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_409 = 6'h19 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_361; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_25 = io_valid_in ? _GEN_409 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_25 = 6'h19 == _T_2[5:0] ? image_25 : _GEN_24; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_74 = 6'h1a == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'hf; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_122 = 6'h1a == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_74; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_170 = 6'h1a == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_122; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_218 = 6'h1a == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_170; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_266 = 6'h1a == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_218; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_314 = 6'h1a == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_266; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_362 = 6'h1a == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_314; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_410 = 6'h1a == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_362; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_26 = io_valid_in ? _GEN_410 : 4'hf; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_26 = 6'h1a == _T_2[5:0] ? image_26 : _GEN_25; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_75 = 6'h1b == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'hf; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_123 = 6'h1b == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_75; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_171 = 6'h1b == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_123; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_219 = 6'h1b == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_171; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_267 = 6'h1b == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_219; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_315 = 6'h1b == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_267; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_363 = 6'h1b == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_315; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_411 = 6'h1b == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_363; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_27 = io_valid_in ? _GEN_411 : 4'hf; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_27 = 6'h1b == _T_2[5:0] ? image_27 : _GEN_26; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_76 = 6'h1c == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'hf; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_124 = 6'h1c == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_76; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_172 = 6'h1c == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_124; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_220 = 6'h1c == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_172; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_268 = 6'h1c == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_220; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_316 = 6'h1c == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_268; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_364 = 6'h1c == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_316; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_412 = 6'h1c == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_364; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_28 = io_valid_in ? _GEN_412 : 4'hf; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_28 = 6'h1c == _T_2[5:0] ? image_28 : _GEN_27; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_77 = 6'h1d == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_125 = 6'h1d == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_77; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_173 = 6'h1d == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_125; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_221 = 6'h1d == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_173; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_269 = 6'h1d == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_221; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_317 = 6'h1d == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_269; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_365 = 6'h1d == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_317; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_413 = 6'h1d == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_365; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_29 = io_valid_in ? _GEN_413 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_29 = 6'h1d == _T_2[5:0] ? image_29 : _GEN_28; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_78 = 6'h1e == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_126 = 6'h1e == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_78; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_174 = 6'h1e == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_126; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_222 = 6'h1e == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_174; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_270 = 6'h1e == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_222; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_318 = 6'h1e == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_270; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_366 = 6'h1e == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_318; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_414 = 6'h1e == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_366; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_30 = io_valid_in ? _GEN_414 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_30 = 6'h1e == _T_2[5:0] ? image_30 : _GEN_29; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_79 = 6'h1f == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_127 = 6'h1f == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_79; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_175 = 6'h1f == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_127; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_223 = 6'h1f == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_175; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_271 = 6'h1f == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_223; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_319 = 6'h1f == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_271; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_367 = 6'h1f == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_319; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_415 = 6'h1f == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_367; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_31 = io_valid_in ? _GEN_415 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_31 = 6'h1f == _T_2[5:0] ? image_31 : _GEN_30; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_80 = 6'h20 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_128 = 6'h20 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_80; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_176 = 6'h20 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_128; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_224 = 6'h20 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_176; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_272 = 6'h20 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_224; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_320 = 6'h20 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_272; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_368 = 6'h20 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_320; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_416 = 6'h20 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_368; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_32 = io_valid_in ? _GEN_416 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_32 = 6'h20 == _T_2[5:0] ? image_32 : _GEN_31; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_81 = 6'h21 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_129 = 6'h21 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_81; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_177 = 6'h21 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_129; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_225 = 6'h21 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_177; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_273 = 6'h21 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_225; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_321 = 6'h21 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_273; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_369 = 6'h21 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_321; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_417 = 6'h21 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_369; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_33 = io_valid_in ? _GEN_417 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_33 = 6'h21 == _T_2[5:0] ? image_33 : _GEN_32; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_82 = 6'h22 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'hf; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_130 = 6'h22 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_82; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_178 = 6'h22 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_130; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_226 = 6'h22 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_178; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_274 = 6'h22 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_226; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_322 = 6'h22 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_274; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_370 = 6'h22 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_322; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_418 = 6'h22 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_370; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_34 = io_valid_in ? _GEN_418 : 4'hf; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_34 = 6'h22 == _T_2[5:0] ? image_34 : _GEN_33; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_83 = 6'h23 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'hf; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_131 = 6'h23 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_83; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_179 = 6'h23 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_131; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_227 = 6'h23 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_179; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_275 = 6'h23 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_227; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_323 = 6'h23 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_275; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_371 = 6'h23 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_323; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_419 = 6'h23 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_371; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_35 = io_valid_in ? _GEN_419 : 4'hf; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_35 = 6'h23 == _T_2[5:0] ? image_35 : _GEN_34; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_84 = 6'h24 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'hf; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_132 = 6'h24 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_84; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_180 = 6'h24 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_132; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_228 = 6'h24 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_180; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_276 = 6'h24 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_228; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_324 = 6'h24 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_276; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_372 = 6'h24 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_324; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_420 = 6'h24 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_372; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_36 = io_valid_in ? _GEN_420 : 4'hf; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_36 = 6'h24 == _T_2[5:0] ? image_36 : _GEN_35; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_85 = 6'h25 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_133 = 6'h25 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_85; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_181 = 6'h25 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_133; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_229 = 6'h25 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_181; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_277 = 6'h25 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_229; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_325 = 6'h25 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_277; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_373 = 6'h25 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_325; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_421 = 6'h25 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_373; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_37 = io_valid_in ? _GEN_421 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_37 = 6'h25 == _T_2[5:0] ? image_37 : _GEN_36; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_86 = 6'h26 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_134 = 6'h26 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_86; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_182 = 6'h26 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_134; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_230 = 6'h26 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_182; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_278 = 6'h26 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_230; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_326 = 6'h26 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_278; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_374 = 6'h26 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_326; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_422 = 6'h26 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_374; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_38 = io_valid_in ? _GEN_422 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_38 = 6'h26 == _T_2[5:0] ? image_38 : _GEN_37; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_87 = 6'h27 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_135 = 6'h27 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_87; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_183 = 6'h27 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_135; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_231 = 6'h27 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_183; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_279 = 6'h27 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_231; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_327 = 6'h27 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_279; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_375 = 6'h27 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_327; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_423 = 6'h27 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_375; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_39 = io_valid_in ? _GEN_423 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_39 = 6'h27 == _T_2[5:0] ? image_39 : _GEN_38; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_88 = 6'h28 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_136 = 6'h28 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_88; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_184 = 6'h28 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_136; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_232 = 6'h28 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_184; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_280 = 6'h28 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_232; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_328 = 6'h28 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_280; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_376 = 6'h28 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_328; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_424 = 6'h28 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_376; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_40 = io_valid_in ? _GEN_424 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_40 = 6'h28 == _T_2[5:0] ? image_40 : _GEN_39; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_89 = 6'h29 == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_137 = 6'h29 == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_89; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_185 = 6'h29 == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_137; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_233 = 6'h29 == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_185; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_281 = 6'h29 == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_233; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_329 = 6'h29 == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_281; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_377 = 6'h29 == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_329; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_425 = 6'h29 == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_377; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_41 = io_valid_in ? _GEN_425 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_41 = 6'h29 == _T_2[5:0] ? image_41 : _GEN_40; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_90 = 6'h2a == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_138 = 6'h2a == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_90; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_186 = 6'h2a == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_138; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_234 = 6'h2a == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_186; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_282 = 6'h2a == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_234; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_330 = 6'h2a == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_282; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_378 = 6'h2a == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_330; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_426 = 6'h2a == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_378; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_42 = io_valid_in ? _GEN_426 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_42 = 6'h2a == _T_2[5:0] ? image_42 : _GEN_41; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_91 = 6'h2b == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_139 = 6'h2b == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_91; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_187 = 6'h2b == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_139; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_235 = 6'h2b == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_187; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_283 = 6'h2b == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_235; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_331 = 6'h2b == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_283; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_379 = 6'h2b == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_331; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_427 = 6'h2b == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_379; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_43 = io_valid_in ? _GEN_427 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_43 = 6'h2b == _T_2[5:0] ? image_43 : _GEN_42; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_92 = 6'h2c == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_140 = 6'h2c == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_92; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_188 = 6'h2c == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_140; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_236 = 6'h2c == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_188; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_284 = 6'h2c == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_236; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_332 = 6'h2c == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_284; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_380 = 6'h2c == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_332; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_428 = 6'h2c == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_380; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_44 = io_valid_in ? _GEN_428 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_44 = 6'h2c == _T_2[5:0] ? image_44 : _GEN_43; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_93 = 6'h2d == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_141 = 6'h2d == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_93; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_189 = 6'h2d == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_141; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_237 = 6'h2d == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_189; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_285 = 6'h2d == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_237; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_333 = 6'h2d == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_285; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_381 = 6'h2d == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_333; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_429 = 6'h2d == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_381; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_45 = io_valid_in ? _GEN_429 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_45 = 6'h2d == _T_2[5:0] ? image_45 : _GEN_44; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_94 = 6'h2e == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_142 = 6'h2e == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_94; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_190 = 6'h2e == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_142; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_238 = 6'h2e == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_190; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_286 = 6'h2e == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_238; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_334 = 6'h2e == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_286; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_382 = 6'h2e == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_334; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_430 = 6'h2e == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_382; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_46 = io_valid_in ? _GEN_430 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_46 = 6'h2e == _T_2[5:0] ? image_46 : _GEN_45; // @[VideoBuffer.scala 29:25]
  wire [3:0] _GEN_95 = 6'h2f == _T_4[5:0] ? io_pixelVal_in_0[3:0] : 4'h0; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_143 = 6'h2f == _T_8[5:0] ? io_pixelVal_in_1[3:0] : _GEN_95; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_191 = 6'h2f == _T_11[5:0] ? io_pixelVal_in_2[3:0] : _GEN_143; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_239 = 6'h2f == _T_14[5:0] ? io_pixelVal_in_3[3:0] : _GEN_191; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_287 = 6'h2f == _T_17[5:0] ? io_pixelVal_in_4[3:0] : _GEN_239; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_335 = 6'h2f == _T_20[5:0] ? io_pixelVal_in_5[3:0] : _GEN_287; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_383 = 6'h2f == _T_23[5:0] ? io_pixelVal_in_6[3:0] : _GEN_335; // @[VideoBuffer.scala 35:49]
  wire [3:0] _GEN_431 = 6'h2f == _T_26[5:0] ? io_pixelVal_in_7[3:0] : _GEN_383; // @[VideoBuffer.scala 35:49]
  wire [3:0] image_47 = io_valid_in ? _GEN_431 : 4'h0; // @[VideoBuffer.scala 33:26]
  wire [3:0] _GEN_47 = 6'h2f == _T_2[5:0] ? image_47 : _GEN_46; // @[VideoBuffer.scala 29:25]
  wire [31:0] _T_29 = pixelIndex + 32'h8; // @[VideoBuffer.scala 37:42]
  wire [6:0] _T_30 = 4'h8 * 4'h6; // @[VideoBuffer.scala 38:42]
  wire [31:0] _GEN_483 = {{25'd0}, _T_30}; // @[VideoBuffer.scala 38:25]
  wire  _T_31 = pixelIndex == _GEN_483; // @[VideoBuffer.scala 38:25]
  assign io_pixelVal_out = {{12'd0}, _GEN_47}; // @[VideoBuffer.scala 29:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pixelIndex = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      pixelIndex <= 32'h0;
    end else if (io_valid_in) begin
      if (_T_31) begin
        pixelIndex <= 32'h0;
      end else begin
        pixelIndex <= _T_29;
      end
    end
  end
endmodule
