module DotProd(
  input        clock,
  input        reset,
  input  [7:0] io_dataInA,
  input  [7:0] io_dataInB,
  output [8:0] io_dataOut,
  output       io_outputValid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] countVal; // @[Counter.scala 29:33]
  wire  countReset = countVal == 4'h8; // @[Counter.scala 38:24]
  wire [3:0] _T_2 = countVal + 4'h1; // @[Counter.scala 39:22]
  reg [8:0] accumulator; // @[DotProd.scala 19:28]
  wire [15:0] product = $signed(io_dataInA) * $signed(io_dataInB); // @[DotProd.scala 20:35]
  wire [15:0] _GEN_5 = {{7{accumulator[8]}},accumulator}; // @[DotProd.scala 21:30]
  wire [15:0] _T_6 = $signed(_GEN_5) + $signed(product); // @[DotProd.scala 21:30]
  wire [15:0] _GEN_4 = countReset ? $signed(16'sh0) : $signed(_T_6); // @[DotProd.scala 25:20]
  assign io_dataOut = _T_6[8:0]; // @[DotProd.scala 23:14]
  assign io_outputValid = countVal == 4'h8; // @[DotProd.scala 26:20 DotProd.scala 29:20]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  countVal = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  accumulator = _RAND_1[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      countVal <= 4'h0;
    end else if (countReset) begin
      countVal <= 4'h0;
    end else begin
      countVal <= _T_2;
    end
    if (reset) begin
      accumulator <= 9'sh0;
    end else begin
      accumulator <= _GEN_4[8:0];
    end
  end
endmodule
module KernelConvolution(
  input        clock,
  input        reset,
  input  [4:0] io_kernelVal_in,
  input  [3:0] io_pixelVal_in_0,
  input  [3:0] io_pixelVal_in_1,
  input  [3:0] io_pixelVal_in_2,
  input  [3:0] io_pixelVal_in_3,
  input  [3:0] io_pixelVal_in_4,
  input  [3:0] io_pixelVal_in_5,
  input  [3:0] io_pixelVal_in_6,
  input  [3:0] io_pixelVal_in_7,
  output [8:0] io_pixelVal_out_0,
  output [8:0] io_pixelVal_out_1,
  output [8:0] io_pixelVal_out_2,
  output [8:0] io_pixelVal_out_3,
  output [8:0] io_pixelVal_out_4,
  output [8:0] io_pixelVal_out_5,
  output [8:0] io_pixelVal_out_6,
  output [8:0] io_pixelVal_out_7,
  output       io_valid_out
);
  wire  DotProd_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_1_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_1_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_1_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_1_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_1_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_1_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_2_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_2_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_2_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_2_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_2_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_2_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_3_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_3_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_3_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_3_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_3_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_3_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_4_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_4_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_4_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_4_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_4_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_4_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_5_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_5_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_5_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_5_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_5_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_5_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_6_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_6_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_6_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_6_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_6_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_6_io_outputValid; // @[KernelConvolution.scala 21:58]
  wire  DotProd_7_clock; // @[KernelConvolution.scala 21:58]
  wire  DotProd_7_reset; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_7_io_dataInA; // @[KernelConvolution.scala 21:58]
  wire [7:0] DotProd_7_io_dataInB; // @[KernelConvolution.scala 21:58]
  wire [8:0] DotProd_7_io_dataOut; // @[KernelConvolution.scala 21:58]
  wire  DotProd_7_io_outputValid; // @[KernelConvolution.scala 21:58]
  DotProd DotProd ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_clock),
    .reset(DotProd_reset),
    .io_dataInA(DotProd_io_dataInA),
    .io_dataInB(DotProd_io_dataInB),
    .io_dataOut(DotProd_io_dataOut),
    .io_outputValid(DotProd_io_outputValid)
  );
  DotProd DotProd_1 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_1_clock),
    .reset(DotProd_1_reset),
    .io_dataInA(DotProd_1_io_dataInA),
    .io_dataInB(DotProd_1_io_dataInB),
    .io_dataOut(DotProd_1_io_dataOut),
    .io_outputValid(DotProd_1_io_outputValid)
  );
  DotProd DotProd_2 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_2_clock),
    .reset(DotProd_2_reset),
    .io_dataInA(DotProd_2_io_dataInA),
    .io_dataInB(DotProd_2_io_dataInB),
    .io_dataOut(DotProd_2_io_dataOut),
    .io_outputValid(DotProd_2_io_outputValid)
  );
  DotProd DotProd_3 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_3_clock),
    .reset(DotProd_3_reset),
    .io_dataInA(DotProd_3_io_dataInA),
    .io_dataInB(DotProd_3_io_dataInB),
    .io_dataOut(DotProd_3_io_dataOut),
    .io_outputValid(DotProd_3_io_outputValid)
  );
  DotProd DotProd_4 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_4_clock),
    .reset(DotProd_4_reset),
    .io_dataInA(DotProd_4_io_dataInA),
    .io_dataInB(DotProd_4_io_dataInB),
    .io_dataOut(DotProd_4_io_dataOut),
    .io_outputValid(DotProd_4_io_outputValid)
  );
  DotProd DotProd_5 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_5_clock),
    .reset(DotProd_5_reset),
    .io_dataInA(DotProd_5_io_dataInA),
    .io_dataInB(DotProd_5_io_dataInB),
    .io_dataOut(DotProd_5_io_dataOut),
    .io_outputValid(DotProd_5_io_outputValid)
  );
  DotProd DotProd_6 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_6_clock),
    .reset(DotProd_6_reset),
    .io_dataInA(DotProd_6_io_dataInA),
    .io_dataInB(DotProd_6_io_dataInB),
    .io_dataOut(DotProd_6_io_dataOut),
    .io_outputValid(DotProd_6_io_outputValid)
  );
  DotProd DotProd_7 ( // @[KernelConvolution.scala 21:58]
    .clock(DotProd_7_clock),
    .reset(DotProd_7_reset),
    .io_dataInA(DotProd_7_io_dataInA),
    .io_dataInB(DotProd_7_io_dataInB),
    .io_dataOut(DotProd_7_io_dataOut),
    .io_outputValid(DotProd_7_io_outputValid)
  );
  assign io_pixelVal_out_0 = DotProd_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_1 = DotProd_1_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_2 = DotProd_2_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_3 = DotProd_3_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_4 = DotProd_4_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_5 = DotProd_5_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_6 = DotProd_6_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_pixelVal_out_7 = DotProd_7_io_dataOut; // @[KernelConvolution.scala 33:34]
  assign io_valid_out = DotProd_io_outputValid; // @[KernelConvolution.scala 35:30]
  assign DotProd_clock = clock;
  assign DotProd_reset = reset;
  assign DotProd_io_dataInA = {{4'd0}, io_pixelVal_in_0}; // @[KernelConvolution.scala 21:32]
  assign DotProd_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_1_clock = clock;
  assign DotProd_1_reset = reset;
  assign DotProd_1_io_dataInA = {{4'd0}, io_pixelVal_in_1}; // @[KernelConvolution.scala 21:32]
  assign DotProd_1_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_2_clock = clock;
  assign DotProd_2_reset = reset;
  assign DotProd_2_io_dataInA = {{4'd0}, io_pixelVal_in_2}; // @[KernelConvolution.scala 21:32]
  assign DotProd_2_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_3_clock = clock;
  assign DotProd_3_reset = reset;
  assign DotProd_3_io_dataInA = {{4'd0}, io_pixelVal_in_3}; // @[KernelConvolution.scala 21:32]
  assign DotProd_3_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_4_clock = clock;
  assign DotProd_4_reset = reset;
  assign DotProd_4_io_dataInA = {{4'd0}, io_pixelVal_in_4}; // @[KernelConvolution.scala 21:32]
  assign DotProd_4_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_5_clock = clock;
  assign DotProd_5_reset = reset;
  assign DotProd_5_io_dataInA = {{4'd0}, io_pixelVal_in_5}; // @[KernelConvolution.scala 21:32]
  assign DotProd_5_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_6_clock = clock;
  assign DotProd_6_reset = reset;
  assign DotProd_6_io_dataInA = {{4'd0}, io_pixelVal_in_6}; // @[KernelConvolution.scala 21:32]
  assign DotProd_6_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
  assign DotProd_7_clock = clock;
  assign DotProd_7_reset = reset;
  assign DotProd_7_io_dataInA = {{4'd0}, io_pixelVal_in_7}; // @[KernelConvolution.scala 21:32]
  assign DotProd_7_io_dataInB = {{3{io_kernelVal_in[4]}},io_kernelVal_in}; // @[KernelConvolution.scala 21:32]
endmodule
module Filter(
  input        clock,
  input        reset,
  input  [5:0] io_SPI_filterIndex,
  input        io_SPI_invert,
  input        io_SPI_distort,
  output [3:0] io_pixelVal_out_0_0,
  output [3:0] io_pixelVal_out_0_1,
  output [3:0] io_pixelVal_out_0_2,
  output [3:0] io_pixelVal_out_0_3,
  output [3:0] io_pixelVal_out_0_4,
  output [3:0] io_pixelVal_out_0_5,
  output [3:0] io_pixelVal_out_0_6,
  output [3:0] io_pixelVal_out_0_7,
  output [3:0] io_pixelVal_out_1_0,
  output [3:0] io_pixelVal_out_1_1,
  output [3:0] io_pixelVal_out_1_2,
  output [3:0] io_pixelVal_out_1_3,
  output [3:0] io_pixelVal_out_1_4,
  output [3:0] io_pixelVal_out_1_5,
  output [3:0] io_pixelVal_out_1_6,
  output [3:0] io_pixelVal_out_1_7,
  output [3:0] io_pixelVal_out_2_0,
  output [3:0] io_pixelVal_out_2_1,
  output [3:0] io_pixelVal_out_2_2,
  output [3:0] io_pixelVal_out_2_3,
  output [3:0] io_pixelVal_out_2_4,
  output [3:0] io_pixelVal_out_2_5,
  output [3:0] io_pixelVal_out_2_6,
  output [3:0] io_pixelVal_out_2_7,
  output       io_valid_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
`endif // RANDOMIZE_REG_INIT
  wire  KernelConvolution_clock; // @[Filter.scala 173:36]
  wire  KernelConvolution_reset; // @[Filter.scala 173:36]
  wire [4:0] KernelConvolution_io_kernelVal_in; // @[Filter.scala 173:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_0; // @[Filter.scala 173:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_1; // @[Filter.scala 173:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_2; // @[Filter.scala 173:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_3; // @[Filter.scala 173:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_4; // @[Filter.scala 173:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_5; // @[Filter.scala 173:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_6; // @[Filter.scala 173:36]
  wire [3:0] KernelConvolution_io_pixelVal_in_7; // @[Filter.scala 173:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_0; // @[Filter.scala 173:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_1; // @[Filter.scala 173:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_2; // @[Filter.scala 173:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_3; // @[Filter.scala 173:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_4; // @[Filter.scala 173:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_5; // @[Filter.scala 173:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_6; // @[Filter.scala 173:36]
  wire [8:0] KernelConvolution_io_pixelVal_out_7; // @[Filter.scala 173:36]
  wire  KernelConvolution_io_valid_out; // @[Filter.scala 173:36]
  wire  KernelConvolution_1_clock; // @[Filter.scala 174:36]
  wire  KernelConvolution_1_reset; // @[Filter.scala 174:36]
  wire [4:0] KernelConvolution_1_io_kernelVal_in; // @[Filter.scala 174:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_0; // @[Filter.scala 174:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_1; // @[Filter.scala 174:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_2; // @[Filter.scala 174:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_3; // @[Filter.scala 174:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_4; // @[Filter.scala 174:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_5; // @[Filter.scala 174:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_6; // @[Filter.scala 174:36]
  wire [3:0] KernelConvolution_1_io_pixelVal_in_7; // @[Filter.scala 174:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_0; // @[Filter.scala 174:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_1; // @[Filter.scala 174:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_2; // @[Filter.scala 174:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_3; // @[Filter.scala 174:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_4; // @[Filter.scala 174:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_5; // @[Filter.scala 174:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_6; // @[Filter.scala 174:36]
  wire [8:0] KernelConvolution_1_io_pixelVal_out_7; // @[Filter.scala 174:36]
  wire  KernelConvolution_1_io_valid_out; // @[Filter.scala 174:36]
  wire  KernelConvolution_2_clock; // @[Filter.scala 175:36]
  wire  KernelConvolution_2_reset; // @[Filter.scala 175:36]
  wire [4:0] KernelConvolution_2_io_kernelVal_in; // @[Filter.scala 175:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_0; // @[Filter.scala 175:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_1; // @[Filter.scala 175:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_2; // @[Filter.scala 175:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_3; // @[Filter.scala 175:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_4; // @[Filter.scala 175:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_5; // @[Filter.scala 175:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_6; // @[Filter.scala 175:36]
  wire [3:0] KernelConvolution_2_io_pixelVal_in_7; // @[Filter.scala 175:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_0; // @[Filter.scala 175:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_1; // @[Filter.scala 175:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_2; // @[Filter.scala 175:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_3; // @[Filter.scala 175:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_4; // @[Filter.scala 175:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_5; // @[Filter.scala 175:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_6; // @[Filter.scala 175:36]
  wire [8:0] KernelConvolution_2_io_pixelVal_out_7; // @[Filter.scala 175:36]
  wire  KernelConvolution_2_io_valid_out; // @[Filter.scala 175:36]
  reg [3:0] kernelCounter; // @[Counter.scala 29:33]
  wire  kernelCountReset = kernelCounter == 4'h8; // @[Counter.scala 38:24]
  wire [3:0] _T_17 = kernelCounter + 4'h1; // @[Counter.scala 39:22]
  wire  _GEN_27995 = 3'h0 == io_SPI_filterIndex[2:0]; // @[Filter.scala 181:41]
  wire  _GEN_27996 = 4'h4 == kernelCounter; // @[Filter.scala 181:41]
  wire [4:0] _GEN_7 = _GEN_27995 & _GEN_27996 ? $signed(5'sh1) : $signed(5'sh0); // @[Filter.scala 181:41]
  wire  _GEN_27998 = 4'h5 == kernelCounter; // @[Filter.scala 181:41]
  wire [4:0] _GEN_8 = _GEN_27995 & _GEN_27998 ? $signed(5'sh0) : $signed(_GEN_7); // @[Filter.scala 181:41]
  wire  _GEN_28000 = 4'h6 == kernelCounter; // @[Filter.scala 181:41]
  wire [4:0] _GEN_9 = _GEN_27995 & _GEN_28000 ? $signed(5'sh0) : $signed(_GEN_8); // @[Filter.scala 181:41]
  wire  _GEN_28002 = 4'h7 == kernelCounter; // @[Filter.scala 181:41]
  wire [4:0] _GEN_10 = _GEN_27995 & _GEN_28002 ? $signed(5'sh0) : $signed(_GEN_9); // @[Filter.scala 181:41]
  wire  _GEN_28004 = 4'h8 == kernelCounter; // @[Filter.scala 181:41]
  wire [4:0] _GEN_11 = _GEN_27995 & _GEN_28004 ? $signed(5'sh0) : $signed(_GEN_10); // @[Filter.scala 181:41]
  wire  _GEN_28005 = 3'h1 == io_SPI_filterIndex[2:0]; // @[Filter.scala 181:41]
  wire  _GEN_28006 = 4'h0 == kernelCounter; // @[Filter.scala 181:41]
  wire [4:0] _GEN_12 = _GEN_28005 & _GEN_28006 ? $signed(5'sh1) : $signed(_GEN_11); // @[Filter.scala 181:41]
  wire  _GEN_28008 = 4'h1 == kernelCounter; // @[Filter.scala 181:41]
  wire [4:0] _GEN_13 = _GEN_28005 & _GEN_28008 ? $signed(5'sh1) : $signed(_GEN_12); // @[Filter.scala 181:41]
  wire  _GEN_28010 = 4'h2 == kernelCounter; // @[Filter.scala 181:41]
  wire [4:0] _GEN_14 = _GEN_28005 & _GEN_28010 ? $signed(5'sh1) : $signed(_GEN_13); // @[Filter.scala 181:41]
  wire  _GEN_28012 = 4'h3 == kernelCounter; // @[Filter.scala 181:41]
  wire [4:0] _GEN_15 = _GEN_28005 & _GEN_28012 ? $signed(5'sh1) : $signed(_GEN_14); // @[Filter.scala 181:41]
  wire [4:0] _GEN_16 = _GEN_28005 & _GEN_27996 ? $signed(5'sh1) : $signed(_GEN_15); // @[Filter.scala 181:41]
  wire [4:0] _GEN_17 = _GEN_28005 & _GEN_27998 ? $signed(5'sh1) : $signed(_GEN_16); // @[Filter.scala 181:41]
  wire [4:0] _GEN_18 = _GEN_28005 & _GEN_28000 ? $signed(5'sh1) : $signed(_GEN_17); // @[Filter.scala 181:41]
  wire [4:0] _GEN_19 = _GEN_28005 & _GEN_28002 ? $signed(5'sh1) : $signed(_GEN_18); // @[Filter.scala 181:41]
  wire [4:0] _GEN_20 = _GEN_28005 & _GEN_28004 ? $signed(5'sh1) : $signed(_GEN_19); // @[Filter.scala 181:41]
  wire  _GEN_28023 = 3'h2 == io_SPI_filterIndex[2:0]; // @[Filter.scala 181:41]
  wire [4:0] _GEN_21 = _GEN_28023 & _GEN_28006 ? $signed(5'sh1) : $signed(_GEN_20); // @[Filter.scala 181:41]
  wire [4:0] _GEN_22 = _GEN_28023 & _GEN_28008 ? $signed(5'sh2) : $signed(_GEN_21); // @[Filter.scala 181:41]
  wire [4:0] _GEN_23 = _GEN_28023 & _GEN_28010 ? $signed(5'sh1) : $signed(_GEN_22); // @[Filter.scala 181:41]
  wire [4:0] _GEN_24 = _GEN_28023 & _GEN_28012 ? $signed(5'sh2) : $signed(_GEN_23); // @[Filter.scala 181:41]
  wire [4:0] _GEN_25 = _GEN_28023 & _GEN_27996 ? $signed(5'sh4) : $signed(_GEN_24); // @[Filter.scala 181:41]
  wire [4:0] _GEN_26 = _GEN_28023 & _GEN_27998 ? $signed(5'sh2) : $signed(_GEN_25); // @[Filter.scala 181:41]
  wire [4:0] _GEN_27 = _GEN_28023 & _GEN_28000 ? $signed(5'sh1) : $signed(_GEN_26); // @[Filter.scala 181:41]
  wire [4:0] _GEN_28 = _GEN_28023 & _GEN_28002 ? $signed(5'sh2) : $signed(_GEN_27); // @[Filter.scala 181:41]
  wire [4:0] _GEN_29 = _GEN_28023 & _GEN_28004 ? $signed(5'sh1) : $signed(_GEN_28); // @[Filter.scala 181:41]
  wire  _GEN_28041 = 3'h3 == io_SPI_filterIndex[2:0]; // @[Filter.scala 181:41]
  wire [4:0] _GEN_30 = _GEN_28041 & _GEN_28006 ? $signed(5'sh0) : $signed(_GEN_29); // @[Filter.scala 181:41]
  wire [4:0] _GEN_31 = _GEN_28041 & _GEN_28008 ? $signed(-5'sh1) : $signed(_GEN_30); // @[Filter.scala 181:41]
  wire [4:0] _GEN_32 = _GEN_28041 & _GEN_28010 ? $signed(5'sh0) : $signed(_GEN_31); // @[Filter.scala 181:41]
  wire [4:0] _GEN_33 = _GEN_28041 & _GEN_28012 ? $signed(-5'sh1) : $signed(_GEN_32); // @[Filter.scala 181:41]
  wire [4:0] _GEN_34 = _GEN_28041 & _GEN_27996 ? $signed(5'sh4) : $signed(_GEN_33); // @[Filter.scala 181:41]
  wire [4:0] _GEN_35 = _GEN_28041 & _GEN_27998 ? $signed(-5'sh1) : $signed(_GEN_34); // @[Filter.scala 181:41]
  wire [4:0] _GEN_36 = _GEN_28041 & _GEN_28000 ? $signed(5'sh0) : $signed(_GEN_35); // @[Filter.scala 181:41]
  wire [4:0] _GEN_37 = _GEN_28041 & _GEN_28002 ? $signed(-5'sh1) : $signed(_GEN_36); // @[Filter.scala 181:41]
  wire [4:0] _GEN_38 = _GEN_28041 & _GEN_28004 ? $signed(5'sh0) : $signed(_GEN_37); // @[Filter.scala 181:41]
  wire  _GEN_28059 = 3'h4 == io_SPI_filterIndex[2:0]; // @[Filter.scala 181:41]
  wire [4:0] _GEN_39 = _GEN_28059 & _GEN_28006 ? $signed(-5'sh1) : $signed(_GEN_38); // @[Filter.scala 181:41]
  wire [4:0] _GEN_40 = _GEN_28059 & _GEN_28008 ? $signed(-5'sh1) : $signed(_GEN_39); // @[Filter.scala 181:41]
  wire [4:0] _GEN_41 = _GEN_28059 & _GEN_28010 ? $signed(-5'sh1) : $signed(_GEN_40); // @[Filter.scala 181:41]
  wire [4:0] _GEN_42 = _GEN_28059 & _GEN_28012 ? $signed(-5'sh1) : $signed(_GEN_41); // @[Filter.scala 181:41]
  wire [4:0] _GEN_43 = _GEN_28059 & _GEN_27996 ? $signed(5'sh8) : $signed(_GEN_42); // @[Filter.scala 181:41]
  wire [4:0] _GEN_44 = _GEN_28059 & _GEN_27998 ? $signed(-5'sh1) : $signed(_GEN_43); // @[Filter.scala 181:41]
  wire [4:0] _GEN_45 = _GEN_28059 & _GEN_28000 ? $signed(-5'sh1) : $signed(_GEN_44); // @[Filter.scala 181:41]
  wire [4:0] _GEN_46 = _GEN_28059 & _GEN_28002 ? $signed(-5'sh1) : $signed(_GEN_45); // @[Filter.scala 181:41]
  wire [4:0] _GEN_47 = _GEN_28059 & _GEN_28004 ? $signed(-5'sh1) : $signed(_GEN_46); // @[Filter.scala 181:41]
  wire  _GEN_28077 = 3'h5 == io_SPI_filterIndex[2:0]; // @[Filter.scala 181:41]
  wire [4:0] _GEN_48 = _GEN_28077 & _GEN_28006 ? $signed(5'sh0) : $signed(_GEN_47); // @[Filter.scala 181:41]
  wire [4:0] _GEN_49 = _GEN_28077 & _GEN_28008 ? $signed(-5'sh1) : $signed(_GEN_48); // @[Filter.scala 181:41]
  wire [4:0] _GEN_50 = _GEN_28077 & _GEN_28010 ? $signed(5'sh0) : $signed(_GEN_49); // @[Filter.scala 181:41]
  wire [4:0] _GEN_51 = _GEN_28077 & _GEN_28012 ? $signed(-5'sh1) : $signed(_GEN_50); // @[Filter.scala 181:41]
  wire [4:0] _GEN_52 = _GEN_28077 & _GEN_27996 ? $signed(5'sh5) : $signed(_GEN_51); // @[Filter.scala 181:41]
  wire [4:0] _GEN_53 = _GEN_28077 & _GEN_27998 ? $signed(-5'sh1) : $signed(_GEN_52); // @[Filter.scala 181:41]
  wire [4:0] _GEN_54 = _GEN_28077 & _GEN_28000 ? $signed(5'sh0) : $signed(_GEN_53); // @[Filter.scala 181:41]
  wire [4:0] _GEN_55 = _GEN_28077 & _GEN_28002 ? $signed(-5'sh1) : $signed(_GEN_54); // @[Filter.scala 181:41]
  reg [1:0] imageCounterX; // @[Counter.scala 29:33]
  wire  imageCounterXReset = imageCounterX == 2'h2; // @[Counter.scala 38:24]
  wire [1:0] _T_23 = imageCounterX + 2'h1; // @[Counter.scala 39:22]
  reg [1:0] imageCounterY; // @[Counter.scala 29:33]
  wire  _T_24 = imageCounterY == 2'h2; // @[Counter.scala 38:24]
  wire [1:0] _T_26 = imageCounterY + 2'h1; // @[Counter.scala 39:22]
  reg [31:0] pixelIndex; // @[Filter.scala 186:31]
  wire [32:0] _T_27 = {{1'd0}, pixelIndex}; // @[Filter.scala 189:31]
  wire [31:0] _GEN_0 = _T_27[31:0] % 32'h20; // @[Filter.scala 189:38]
  wire [5:0] _T_29 = _GEN_0[5:0]; // @[Filter.scala 189:38]
  wire [5:0] _GEN_28295 = {{4'd0}, imageCounterX}; // @[Filter.scala 189:53]
  wire [5:0] _T_31 = _T_29 + _GEN_28295; // @[Filter.scala 189:53]
  wire [5:0] _T_33 = _T_31 - 6'h1; // @[Filter.scala 189:69]
  wire [31:0] _T_36 = _T_27[31:0] / 32'h20; // @[Filter.scala 190:38]
  wire [31:0] _GEN_28296 = {{30'd0}, imageCounterY}; // @[Filter.scala 190:53]
  wire [31:0] _T_38 = _T_36 + _GEN_28296; // @[Filter.scala 190:53]
  wire [31:0] _T_40 = _T_38 - 32'h1; // @[Filter.scala 190:69]
  wire [37:0] _T_41 = _T_40 * 32'h20; // @[Filter.scala 191:42]
  wire [37:0] _GEN_28297 = {{32'd0}, _T_33}; // @[Filter.scala 191:57]
  wire [37:0] _T_43 = _T_41 + _GEN_28297; // @[Filter.scala 191:57]
  wire [3:0] _GEN_174 = 10'h3 == _T_43[9:0] ? 4'h3 : 4'ha; // @[Filter.scala 191:62]
  wire [3:0] _GEN_175 = 10'h4 == _T_43[9:0] ? 4'ha : _GEN_174; // @[Filter.scala 191:62]
  wire [3:0] _GEN_176 = 10'h5 == _T_43[9:0] ? 4'ha : _GEN_175; // @[Filter.scala 191:62]
  wire [3:0] _GEN_177 = 10'h6 == _T_43[9:0] ? 4'ha : _GEN_176; // @[Filter.scala 191:62]
  wire [3:0] _GEN_178 = 10'h7 == _T_43[9:0] ? 4'ha : _GEN_177; // @[Filter.scala 191:62]
  wire [3:0] _GEN_179 = 10'h8 == _T_43[9:0] ? 4'ha : _GEN_178; // @[Filter.scala 191:62]
  wire [3:0] _GEN_180 = 10'h9 == _T_43[9:0] ? 4'ha : _GEN_179; // @[Filter.scala 191:62]
  wire [3:0] _GEN_181 = 10'ha == _T_43[9:0] ? 4'ha : _GEN_180; // @[Filter.scala 191:62]
  wire [3:0] _GEN_182 = 10'hb == _T_43[9:0] ? 4'ha : _GEN_181; // @[Filter.scala 191:62]
  wire [3:0] _GEN_183 = 10'hc == _T_43[9:0] ? 4'ha : _GEN_182; // @[Filter.scala 191:62]
  wire [3:0] _GEN_184 = 10'hd == _T_43[9:0] ? 4'ha : _GEN_183; // @[Filter.scala 191:62]
  wire [3:0] _GEN_185 = 10'he == _T_43[9:0] ? 4'ha : _GEN_184; // @[Filter.scala 191:62]
  wire [3:0] _GEN_186 = 10'hf == _T_43[9:0] ? 4'ha : _GEN_185; // @[Filter.scala 191:62]
  wire [3:0] _GEN_187 = 10'h10 == _T_43[9:0] ? 4'ha : _GEN_186; // @[Filter.scala 191:62]
  wire [3:0] _GEN_188 = 10'h11 == _T_43[9:0] ? 4'ha : _GEN_187; // @[Filter.scala 191:62]
  wire [3:0] _GEN_189 = 10'h12 == _T_43[9:0] ? 4'ha : _GEN_188; // @[Filter.scala 191:62]
  wire [3:0] _GEN_190 = 10'h13 == _T_43[9:0] ? 4'ha : _GEN_189; // @[Filter.scala 191:62]
  wire [3:0] _GEN_191 = 10'h14 == _T_43[9:0] ? 4'ha : _GEN_190; // @[Filter.scala 191:62]
  wire [3:0] _GEN_192 = 10'h15 == _T_43[9:0] ? 4'ha : _GEN_191; // @[Filter.scala 191:62]
  wire [3:0] _GEN_193 = 10'h16 == _T_43[9:0] ? 4'ha : _GEN_192; // @[Filter.scala 191:62]
  wire [3:0] _GEN_194 = 10'h17 == _T_43[9:0] ? 4'ha : _GEN_193; // @[Filter.scala 191:62]
  wire [3:0] _GEN_195 = 10'h18 == _T_43[9:0] ? 4'ha : _GEN_194; // @[Filter.scala 191:62]
  wire [3:0] _GEN_196 = 10'h19 == _T_43[9:0] ? 4'ha : _GEN_195; // @[Filter.scala 191:62]
  wire [3:0] _GEN_197 = 10'h1a == _T_43[9:0] ? 4'ha : _GEN_196; // @[Filter.scala 191:62]
  wire [3:0] _GEN_198 = 10'h1b == _T_43[9:0] ? 4'ha : _GEN_197; // @[Filter.scala 191:62]
  wire [3:0] _GEN_199 = 10'h1c == _T_43[9:0] ? 4'ha : _GEN_198; // @[Filter.scala 191:62]
  wire [3:0] _GEN_200 = 10'h1d == _T_43[9:0] ? 4'ha : _GEN_199; // @[Filter.scala 191:62]
  wire [3:0] _GEN_201 = 10'h1e == _T_43[9:0] ? 4'ha : _GEN_200; // @[Filter.scala 191:62]
  wire [3:0] _GEN_202 = 10'h1f == _T_43[9:0] ? 4'h0 : _GEN_201; // @[Filter.scala 191:62]
  wire [3:0] _GEN_203 = 10'h20 == _T_43[9:0] ? 4'ha : _GEN_202; // @[Filter.scala 191:62]
  wire [3:0] _GEN_204 = 10'h21 == _T_43[9:0] ? 4'ha : _GEN_203; // @[Filter.scala 191:62]
  wire [3:0] _GEN_205 = 10'h22 == _T_43[9:0] ? 4'ha : _GEN_204; // @[Filter.scala 191:62]
  wire [3:0] _GEN_206 = 10'h23 == _T_43[9:0] ? 4'h3 : _GEN_205; // @[Filter.scala 191:62]
  wire [3:0] _GEN_207 = 10'h24 == _T_43[9:0] ? 4'ha : _GEN_206; // @[Filter.scala 191:62]
  wire [3:0] _GEN_208 = 10'h25 == _T_43[9:0] ? 4'ha : _GEN_207; // @[Filter.scala 191:62]
  wire [3:0] _GEN_209 = 10'h26 == _T_43[9:0] ? 4'ha : _GEN_208; // @[Filter.scala 191:62]
  wire [3:0] _GEN_210 = 10'h27 == _T_43[9:0] ? 4'h1 : _GEN_209; // @[Filter.scala 191:62]
  wire [3:0] _GEN_211 = 10'h28 == _T_43[9:0] ? 4'h1 : _GEN_210; // @[Filter.scala 191:62]
  wire [3:0] _GEN_212 = 10'h29 == _T_43[9:0] ? 4'ha : _GEN_211; // @[Filter.scala 191:62]
  wire [3:0] _GEN_213 = 10'h2a == _T_43[9:0] ? 4'ha : _GEN_212; // @[Filter.scala 191:62]
  wire [3:0] _GEN_214 = 10'h2b == _T_43[9:0] ? 4'ha : _GEN_213; // @[Filter.scala 191:62]
  wire [3:0] _GEN_215 = 10'h2c == _T_43[9:0] ? 4'ha : _GEN_214; // @[Filter.scala 191:62]
  wire [3:0] _GEN_216 = 10'h2d == _T_43[9:0] ? 4'ha : _GEN_215; // @[Filter.scala 191:62]
  wire [3:0] _GEN_217 = 10'h2e == _T_43[9:0] ? 4'ha : _GEN_216; // @[Filter.scala 191:62]
  wire [3:0] _GEN_218 = 10'h2f == _T_43[9:0] ? 4'ha : _GEN_217; // @[Filter.scala 191:62]
  wire [3:0] _GEN_219 = 10'h30 == _T_43[9:0] ? 4'ha : _GEN_218; // @[Filter.scala 191:62]
  wire [3:0] _GEN_220 = 10'h31 == _T_43[9:0] ? 4'ha : _GEN_219; // @[Filter.scala 191:62]
  wire [3:0] _GEN_221 = 10'h32 == _T_43[9:0] ? 4'ha : _GEN_220; // @[Filter.scala 191:62]
  wire [3:0] _GEN_222 = 10'h33 == _T_43[9:0] ? 4'ha : _GEN_221; // @[Filter.scala 191:62]
  wire [3:0] _GEN_223 = 10'h34 == _T_43[9:0] ? 4'ha : _GEN_222; // @[Filter.scala 191:62]
  wire [3:0] _GEN_224 = 10'h35 == _T_43[9:0] ? 4'ha : _GEN_223; // @[Filter.scala 191:62]
  wire [3:0] _GEN_225 = 10'h36 == _T_43[9:0] ? 4'ha : _GEN_224; // @[Filter.scala 191:62]
  wire [3:0] _GEN_226 = 10'h37 == _T_43[9:0] ? 4'h1 : _GEN_225; // @[Filter.scala 191:62]
  wire [3:0] _GEN_227 = 10'h38 == _T_43[9:0] ? 4'h1 : _GEN_226; // @[Filter.scala 191:62]
  wire [3:0] _GEN_228 = 10'h39 == _T_43[9:0] ? 4'ha : _GEN_227; // @[Filter.scala 191:62]
  wire [3:0] _GEN_229 = 10'h3a == _T_43[9:0] ? 4'ha : _GEN_228; // @[Filter.scala 191:62]
  wire [3:0] _GEN_230 = 10'h3b == _T_43[9:0] ? 4'ha : _GEN_229; // @[Filter.scala 191:62]
  wire [3:0] _GEN_231 = 10'h3c == _T_43[9:0] ? 4'ha : _GEN_230; // @[Filter.scala 191:62]
  wire [3:0] _GEN_232 = 10'h3d == _T_43[9:0] ? 4'h3 : _GEN_231; // @[Filter.scala 191:62]
  wire [3:0] _GEN_233 = 10'h3e == _T_43[9:0] ? 4'ha : _GEN_232; // @[Filter.scala 191:62]
  wire [3:0] _GEN_234 = 10'h3f == _T_43[9:0] ? 4'h0 : _GEN_233; // @[Filter.scala 191:62]
  wire [3:0] _GEN_235 = 10'h40 == _T_43[9:0] ? 4'ha : _GEN_234; // @[Filter.scala 191:62]
  wire [3:0] _GEN_236 = 10'h41 == _T_43[9:0] ? 4'ha : _GEN_235; // @[Filter.scala 191:62]
  wire [3:0] _GEN_237 = 10'h42 == _T_43[9:0] ? 4'ha : _GEN_236; // @[Filter.scala 191:62]
  wire [3:0] _GEN_238 = 10'h43 == _T_43[9:0] ? 4'h2 : _GEN_237; // @[Filter.scala 191:62]
  wire [3:0] _GEN_239 = 10'h44 == _T_43[9:0] ? 4'h3 : _GEN_238; // @[Filter.scala 191:62]
  wire [3:0] _GEN_240 = 10'h45 == _T_43[9:0] ? 4'h0 : _GEN_239; // @[Filter.scala 191:62]
  wire [3:0] _GEN_241 = 10'h46 == _T_43[9:0] ? 4'h0 : _GEN_240; // @[Filter.scala 191:62]
  wire [3:0] _GEN_242 = 10'h47 == _T_43[9:0] ? 4'h0 : _GEN_241; // @[Filter.scala 191:62]
  wire [3:0] _GEN_243 = 10'h48 == _T_43[9:0] ? 4'h0 : _GEN_242; // @[Filter.scala 191:62]
  wire [3:0] _GEN_244 = 10'h49 == _T_43[9:0] ? 4'ha : _GEN_243; // @[Filter.scala 191:62]
  wire [3:0] _GEN_245 = 10'h4a == _T_43[9:0] ? 4'ha : _GEN_244; // @[Filter.scala 191:62]
  wire [3:0] _GEN_246 = 10'h4b == _T_43[9:0] ? 4'ha : _GEN_245; // @[Filter.scala 191:62]
  wire [3:0] _GEN_247 = 10'h4c == _T_43[9:0] ? 4'ha : _GEN_246; // @[Filter.scala 191:62]
  wire [3:0] _GEN_248 = 10'h4d == _T_43[9:0] ? 4'ha : _GEN_247; // @[Filter.scala 191:62]
  wire [3:0] _GEN_249 = 10'h4e == _T_43[9:0] ? 4'ha : _GEN_248; // @[Filter.scala 191:62]
  wire [3:0] _GEN_250 = 10'h4f == _T_43[9:0] ? 4'ha : _GEN_249; // @[Filter.scala 191:62]
  wire [3:0] _GEN_251 = 10'h50 == _T_43[9:0] ? 4'ha : _GEN_250; // @[Filter.scala 191:62]
  wire [3:0] _GEN_252 = 10'h51 == _T_43[9:0] ? 4'ha : _GEN_251; // @[Filter.scala 191:62]
  wire [3:0] _GEN_253 = 10'h52 == _T_43[9:0] ? 4'ha : _GEN_252; // @[Filter.scala 191:62]
  wire [3:0] _GEN_254 = 10'h53 == _T_43[9:0] ? 4'ha : _GEN_253; // @[Filter.scala 191:62]
  wire [3:0] _GEN_255 = 10'h54 == _T_43[9:0] ? 4'h1 : _GEN_254; // @[Filter.scala 191:62]
  wire [3:0] _GEN_256 = 10'h55 == _T_43[9:0] ? 4'h1 : _GEN_255; // @[Filter.scala 191:62]
  wire [3:0] _GEN_257 = 10'h56 == _T_43[9:0] ? 4'h1 : _GEN_256; // @[Filter.scala 191:62]
  wire [3:0] _GEN_258 = 10'h57 == _T_43[9:0] ? 4'h0 : _GEN_257; // @[Filter.scala 191:62]
  wire [3:0] _GEN_259 = 10'h58 == _T_43[9:0] ? 4'ha : _GEN_258; // @[Filter.scala 191:62]
  wire [3:0] _GEN_260 = 10'h59 == _T_43[9:0] ? 4'h0 : _GEN_259; // @[Filter.scala 191:62]
  wire [3:0] _GEN_261 = 10'h5a == _T_43[9:0] ? 4'ha : _GEN_260; // @[Filter.scala 191:62]
  wire [3:0] _GEN_262 = 10'h5b == _T_43[9:0] ? 4'ha : _GEN_261; // @[Filter.scala 191:62]
  wire [3:0] _GEN_263 = 10'h5c == _T_43[9:0] ? 4'ha : _GEN_262; // @[Filter.scala 191:62]
  wire [3:0] _GEN_264 = 10'h5d == _T_43[9:0] ? 4'h3 : _GEN_263; // @[Filter.scala 191:62]
  wire [3:0] _GEN_265 = 10'h5e == _T_43[9:0] ? 4'ha : _GEN_264; // @[Filter.scala 191:62]
  wire [3:0] _GEN_266 = 10'h5f == _T_43[9:0] ? 4'h0 : _GEN_265; // @[Filter.scala 191:62]
  wire [3:0] _GEN_267 = 10'h60 == _T_43[9:0] ? 4'ha : _GEN_266; // @[Filter.scala 191:62]
  wire [3:0] _GEN_268 = 10'h61 == _T_43[9:0] ? 4'ha : _GEN_267; // @[Filter.scala 191:62]
  wire [3:0] _GEN_269 = 10'h62 == _T_43[9:0] ? 4'ha : _GEN_268; // @[Filter.scala 191:62]
  wire [3:0] _GEN_270 = 10'h63 == _T_43[9:0] ? 4'ha : _GEN_269; // @[Filter.scala 191:62]
  wire [3:0] _GEN_271 = 10'h64 == _T_43[9:0] ? 4'h3 : _GEN_270; // @[Filter.scala 191:62]
  wire [3:0] _GEN_272 = 10'h65 == _T_43[9:0] ? 4'h0 : _GEN_271; // @[Filter.scala 191:62]
  wire [3:0] _GEN_273 = 10'h66 == _T_43[9:0] ? 4'ha : _GEN_272; // @[Filter.scala 191:62]
  wire [3:0] _GEN_274 = 10'h67 == _T_43[9:0] ? 4'ha : _GEN_273; // @[Filter.scala 191:62]
  wire [3:0] _GEN_275 = 10'h68 == _T_43[9:0] ? 4'ha : _GEN_274; // @[Filter.scala 191:62]
  wire [3:0] _GEN_276 = 10'h69 == _T_43[9:0] ? 4'h0 : _GEN_275; // @[Filter.scala 191:62]
  wire [3:0] _GEN_277 = 10'h6a == _T_43[9:0] ? 4'h1 : _GEN_276; // @[Filter.scala 191:62]
  wire [3:0] _GEN_278 = 10'h6b == _T_43[9:0] ? 4'h1 : _GEN_277; // @[Filter.scala 191:62]
  wire [3:0] _GEN_279 = 10'h6c == _T_43[9:0] ? 4'ha : _GEN_278; // @[Filter.scala 191:62]
  wire [3:0] _GEN_280 = 10'h6d == _T_43[9:0] ? 4'ha : _GEN_279; // @[Filter.scala 191:62]
  wire [3:0] _GEN_281 = 10'h6e == _T_43[9:0] ? 4'ha : _GEN_280; // @[Filter.scala 191:62]
  wire [3:0] _GEN_282 = 10'h6f == _T_43[9:0] ? 4'ha : _GEN_281; // @[Filter.scala 191:62]
  wire [3:0] _GEN_283 = 10'h70 == _T_43[9:0] ? 4'ha : _GEN_282; // @[Filter.scala 191:62]
  wire [3:0] _GEN_284 = 10'h71 == _T_43[9:0] ? 4'ha : _GEN_283; // @[Filter.scala 191:62]
  wire [3:0] _GEN_285 = 10'h72 == _T_43[9:0] ? 4'ha : _GEN_284; // @[Filter.scala 191:62]
  wire [3:0] _GEN_286 = 10'h73 == _T_43[9:0] ? 4'h1 : _GEN_285; // @[Filter.scala 191:62]
  wire [3:0] _GEN_287 = 10'h74 == _T_43[9:0] ? 4'h0 : _GEN_286; // @[Filter.scala 191:62]
  wire [3:0] _GEN_288 = 10'h75 == _T_43[9:0] ? 4'h0 : _GEN_287; // @[Filter.scala 191:62]
  wire [3:0] _GEN_289 = 10'h76 == _T_43[9:0] ? 4'h0 : _GEN_288; // @[Filter.scala 191:62]
  wire [3:0] _GEN_290 = 10'h77 == _T_43[9:0] ? 4'ha : _GEN_289; // @[Filter.scala 191:62]
  wire [3:0] _GEN_291 = 10'h78 == _T_43[9:0] ? 4'ha : _GEN_290; // @[Filter.scala 191:62]
  wire [3:0] _GEN_292 = 10'h79 == _T_43[9:0] ? 4'ha : _GEN_291; // @[Filter.scala 191:62]
  wire [3:0] _GEN_293 = 10'h7a == _T_43[9:0] ? 4'h0 : _GEN_292; // @[Filter.scala 191:62]
  wire [3:0] _GEN_294 = 10'h7b == _T_43[9:0] ? 4'ha : _GEN_293; // @[Filter.scala 191:62]
  wire [3:0] _GEN_295 = 10'h7c == _T_43[9:0] ? 4'ha : _GEN_294; // @[Filter.scala 191:62]
  wire [3:0] _GEN_296 = 10'h7d == _T_43[9:0] ? 4'h2 : _GEN_295; // @[Filter.scala 191:62]
  wire [3:0] _GEN_297 = 10'h7e == _T_43[9:0] ? 4'h3 : _GEN_296; // @[Filter.scala 191:62]
  wire [3:0] _GEN_298 = 10'h7f == _T_43[9:0] ? 4'h0 : _GEN_297; // @[Filter.scala 191:62]
  wire [3:0] _GEN_299 = 10'h80 == _T_43[9:0] ? 4'ha : _GEN_298; // @[Filter.scala 191:62]
  wire [3:0] _GEN_300 = 10'h81 == _T_43[9:0] ? 4'ha : _GEN_299; // @[Filter.scala 191:62]
  wire [3:0] _GEN_301 = 10'h82 == _T_43[9:0] ? 4'h1 : _GEN_300; // @[Filter.scala 191:62]
  wire [3:0] _GEN_302 = 10'h83 == _T_43[9:0] ? 4'h0 : _GEN_301; // @[Filter.scala 191:62]
  wire [3:0] _GEN_303 = 10'h84 == _T_43[9:0] ? 4'h2 : _GEN_302; // @[Filter.scala 191:62]
  wire [3:0] _GEN_304 = 10'h85 == _T_43[9:0] ? 4'h1 : _GEN_303; // @[Filter.scala 191:62]
  wire [3:0] _GEN_305 = 10'h86 == _T_43[9:0] ? 4'h1 : _GEN_304; // @[Filter.scala 191:62]
  wire [3:0] _GEN_306 = 10'h87 == _T_43[9:0] ? 4'ha : _GEN_305; // @[Filter.scala 191:62]
  wire [3:0] _GEN_307 = 10'h88 == _T_43[9:0] ? 4'ha : _GEN_306; // @[Filter.scala 191:62]
  wire [3:0] _GEN_308 = 10'h89 == _T_43[9:0] ? 4'h0 : _GEN_307; // @[Filter.scala 191:62]
  wire [3:0] _GEN_309 = 10'h8a == _T_43[9:0] ? 4'h0 : _GEN_308; // @[Filter.scala 191:62]
  wire [3:0] _GEN_310 = 10'h8b == _T_43[9:0] ? 4'h1 : _GEN_309; // @[Filter.scala 191:62]
  wire [3:0] _GEN_311 = 10'h8c == _T_43[9:0] ? 4'h1 : _GEN_310; // @[Filter.scala 191:62]
  wire [3:0] _GEN_312 = 10'h8d == _T_43[9:0] ? 4'h1 : _GEN_311; // @[Filter.scala 191:62]
  wire [3:0] _GEN_313 = 10'h8e == _T_43[9:0] ? 4'h1 : _GEN_312; // @[Filter.scala 191:62]
  wire [3:0] _GEN_314 = 10'h8f == _T_43[9:0] ? 4'h1 : _GEN_313; // @[Filter.scala 191:62]
  wire [3:0] _GEN_315 = 10'h90 == _T_43[9:0] ? 4'h1 : _GEN_314; // @[Filter.scala 191:62]
  wire [3:0] _GEN_316 = 10'h91 == _T_43[9:0] ? 4'h1 : _GEN_315; // @[Filter.scala 191:62]
  wire [3:0] _GEN_317 = 10'h92 == _T_43[9:0] ? 4'h1 : _GEN_316; // @[Filter.scala 191:62]
  wire [3:0] _GEN_318 = 10'h93 == _T_43[9:0] ? 4'h0 : _GEN_317; // @[Filter.scala 191:62]
  wire [3:0] _GEN_319 = 10'h94 == _T_43[9:0] ? 4'h0 : _GEN_318; // @[Filter.scala 191:62]
  wire [3:0] _GEN_320 = 10'h95 == _T_43[9:0] ? 4'ha : _GEN_319; // @[Filter.scala 191:62]
  wire [3:0] _GEN_321 = 10'h96 == _T_43[9:0] ? 4'ha : _GEN_320; // @[Filter.scala 191:62]
  wire [3:0] _GEN_322 = 10'h97 == _T_43[9:0] ? 4'ha : _GEN_321; // @[Filter.scala 191:62]
  wire [3:0] _GEN_323 = 10'h98 == _T_43[9:0] ? 4'h1 : _GEN_322; // @[Filter.scala 191:62]
  wire [3:0] _GEN_324 = 10'h99 == _T_43[9:0] ? 4'h0 : _GEN_323; // @[Filter.scala 191:62]
  wire [3:0] _GEN_325 = 10'h9a == _T_43[9:0] ? 4'h1 : _GEN_324; // @[Filter.scala 191:62]
  wire [3:0] _GEN_326 = 10'h9b == _T_43[9:0] ? 4'h1 : _GEN_325; // @[Filter.scala 191:62]
  wire [3:0] _GEN_327 = 10'h9c == _T_43[9:0] ? 4'ha : _GEN_326; // @[Filter.scala 191:62]
  wire [3:0] _GEN_328 = 10'h9d == _T_43[9:0] ? 4'ha : _GEN_327; // @[Filter.scala 191:62]
  wire [3:0] _GEN_329 = 10'h9e == _T_43[9:0] ? 4'h3 : _GEN_328; // @[Filter.scala 191:62]
  wire [3:0] _GEN_330 = 10'h9f == _T_43[9:0] ? 4'h0 : _GEN_329; // @[Filter.scala 191:62]
  wire [3:0] _GEN_331 = 10'ha0 == _T_43[9:0] ? 4'ha : _GEN_330; // @[Filter.scala 191:62]
  wire [3:0] _GEN_332 = 10'ha1 == _T_43[9:0] ? 4'h1 : _GEN_331; // @[Filter.scala 191:62]
  wire [3:0] _GEN_333 = 10'ha2 == _T_43[9:0] ? 4'h0 : _GEN_332; // @[Filter.scala 191:62]
  wire [3:0] _GEN_334 = 10'ha3 == _T_43[9:0] ? 4'h3 : _GEN_333; // @[Filter.scala 191:62]
  wire [3:0] _GEN_335 = 10'ha4 == _T_43[9:0] ? 4'ha : _GEN_334; // @[Filter.scala 191:62]
  wire [3:0] _GEN_336 = 10'ha5 == _T_43[9:0] ? 4'ha : _GEN_335; // @[Filter.scala 191:62]
  wire [3:0] _GEN_337 = 10'ha6 == _T_43[9:0] ? 4'ha : _GEN_336; // @[Filter.scala 191:62]
  wire [3:0] _GEN_338 = 10'ha7 == _T_43[9:0] ? 4'h0 : _GEN_337; // @[Filter.scala 191:62]
  wire [3:0] _GEN_339 = 10'ha8 == _T_43[9:0] ? 4'ha : _GEN_338; // @[Filter.scala 191:62]
  wire [3:0] _GEN_340 = 10'ha9 == _T_43[9:0] ? 4'h1 : _GEN_339; // @[Filter.scala 191:62]
  wire [3:0] _GEN_341 = 10'haa == _T_43[9:0] ? 4'h0 : _GEN_340; // @[Filter.scala 191:62]
  wire [3:0] _GEN_342 = 10'hab == _T_43[9:0] ? 4'h0 : _GEN_341; // @[Filter.scala 191:62]
  wire [3:0] _GEN_343 = 10'hac == _T_43[9:0] ? 4'h0 : _GEN_342; // @[Filter.scala 191:62]
  wire [3:0] _GEN_344 = 10'had == _T_43[9:0] ? 4'h0 : _GEN_343; // @[Filter.scala 191:62]
  wire [3:0] _GEN_345 = 10'hae == _T_43[9:0] ? 4'h0 : _GEN_344; // @[Filter.scala 191:62]
  wire [3:0] _GEN_346 = 10'haf == _T_43[9:0] ? 4'h0 : _GEN_345; // @[Filter.scala 191:62]
  wire [3:0] _GEN_347 = 10'hb0 == _T_43[9:0] ? 4'h0 : _GEN_346; // @[Filter.scala 191:62]
  wire [3:0] _GEN_348 = 10'hb1 == _T_43[9:0] ? 4'h0 : _GEN_347; // @[Filter.scala 191:62]
  wire [3:0] _GEN_349 = 10'hb2 == _T_43[9:0] ? 4'h0 : _GEN_348; // @[Filter.scala 191:62]
  wire [3:0] _GEN_350 = 10'hb3 == _T_43[9:0] ? 4'h0 : _GEN_349; // @[Filter.scala 191:62]
  wire [3:0] _GEN_351 = 10'hb4 == _T_43[9:0] ? 4'h1 : _GEN_350; // @[Filter.scala 191:62]
  wire [3:0] _GEN_352 = 10'hb5 == _T_43[9:0] ? 4'h1 : _GEN_351; // @[Filter.scala 191:62]
  wire [3:0] _GEN_353 = 10'hb6 == _T_43[9:0] ? 4'ha : _GEN_352; // @[Filter.scala 191:62]
  wire [3:0] _GEN_354 = 10'hb7 == _T_43[9:0] ? 4'h0 : _GEN_353; // @[Filter.scala 191:62]
  wire [3:0] _GEN_355 = 10'hb8 == _T_43[9:0] ? 4'ha : _GEN_354; // @[Filter.scala 191:62]
  wire [3:0] _GEN_356 = 10'hb9 == _T_43[9:0] ? 4'ha : _GEN_355; // @[Filter.scala 191:62]
  wire [3:0] _GEN_357 = 10'hba == _T_43[9:0] ? 4'ha : _GEN_356; // @[Filter.scala 191:62]
  wire [3:0] _GEN_358 = 10'hbb == _T_43[9:0] ? 4'h0 : _GEN_357; // @[Filter.scala 191:62]
  wire [3:0] _GEN_359 = 10'hbc == _T_43[9:0] ? 4'ha : _GEN_358; // @[Filter.scala 191:62]
  wire [3:0] _GEN_360 = 10'hbd == _T_43[9:0] ? 4'ha : _GEN_359; // @[Filter.scala 191:62]
  wire [3:0] _GEN_361 = 10'hbe == _T_43[9:0] ? 4'h3 : _GEN_360; // @[Filter.scala 191:62]
  wire [3:0] _GEN_362 = 10'hbf == _T_43[9:0] ? 4'h0 : _GEN_361; // @[Filter.scala 191:62]
  wire [3:0] _GEN_363 = 10'hc0 == _T_43[9:0] ? 4'ha : _GEN_362; // @[Filter.scala 191:62]
  wire [3:0] _GEN_364 = 10'hc1 == _T_43[9:0] ? 4'ha : _GEN_363; // @[Filter.scala 191:62]
  wire [3:0] _GEN_365 = 10'hc2 == _T_43[9:0] ? 4'h3 : _GEN_364; // @[Filter.scala 191:62]
  wire [3:0] _GEN_366 = 10'hc3 == _T_43[9:0] ? 4'h2 : _GEN_365; // @[Filter.scala 191:62]
  wire [3:0] _GEN_367 = 10'hc4 == _T_43[9:0] ? 4'h0 : _GEN_366; // @[Filter.scala 191:62]
  wire [3:0] _GEN_368 = 10'hc5 == _T_43[9:0] ? 4'h0 : _GEN_367; // @[Filter.scala 191:62]
  wire [3:0] _GEN_369 = 10'hc6 == _T_43[9:0] ? 4'h0 : _GEN_368; // @[Filter.scala 191:62]
  wire [3:0] _GEN_370 = 10'hc7 == _T_43[9:0] ? 4'ha : _GEN_369; // @[Filter.scala 191:62]
  wire [3:0] _GEN_371 = 10'hc8 == _T_43[9:0] ? 4'h1 : _GEN_370; // @[Filter.scala 191:62]
  wire [3:0] _GEN_372 = 10'hc9 == _T_43[9:0] ? 4'h0 : _GEN_371; // @[Filter.scala 191:62]
  wire [3:0] _GEN_373 = 10'hca == _T_43[9:0] ? 4'h0 : _GEN_372; // @[Filter.scala 191:62]
  wire [3:0] _GEN_374 = 10'hcb == _T_43[9:0] ? 4'h0 : _GEN_373; // @[Filter.scala 191:62]
  wire [3:0] _GEN_375 = 10'hcc == _T_43[9:0] ? 4'h0 : _GEN_374; // @[Filter.scala 191:62]
  wire [3:0] _GEN_376 = 10'hcd == _T_43[9:0] ? 4'h0 : _GEN_375; // @[Filter.scala 191:62]
  wire [3:0] _GEN_377 = 10'hce == _T_43[9:0] ? 4'h0 : _GEN_376; // @[Filter.scala 191:62]
  wire [3:0] _GEN_378 = 10'hcf == _T_43[9:0] ? 4'h0 : _GEN_377; // @[Filter.scala 191:62]
  wire [3:0] _GEN_379 = 10'hd0 == _T_43[9:0] ? 4'h0 : _GEN_378; // @[Filter.scala 191:62]
  wire [3:0] _GEN_380 = 10'hd1 == _T_43[9:0] ? 4'h0 : _GEN_379; // @[Filter.scala 191:62]
  wire [3:0] _GEN_381 = 10'hd2 == _T_43[9:0] ? 4'h0 : _GEN_380; // @[Filter.scala 191:62]
  wire [3:0] _GEN_382 = 10'hd3 == _T_43[9:0] ? 4'h0 : _GEN_381; // @[Filter.scala 191:62]
  wire [3:0] _GEN_383 = 10'hd4 == _T_43[9:0] ? 4'h0 : _GEN_382; // @[Filter.scala 191:62]
  wire [3:0] _GEN_384 = 10'hd5 == _T_43[9:0] ? 4'h0 : _GEN_383; // @[Filter.scala 191:62]
  wire [3:0] _GEN_385 = 10'hd6 == _T_43[9:0] ? 4'h1 : _GEN_384; // @[Filter.scala 191:62]
  wire [3:0] _GEN_386 = 10'hd7 == _T_43[9:0] ? 4'ha : _GEN_385; // @[Filter.scala 191:62]
  wire [3:0] _GEN_387 = 10'hd8 == _T_43[9:0] ? 4'h0 : _GEN_386; // @[Filter.scala 191:62]
  wire [3:0] _GEN_388 = 10'hd9 == _T_43[9:0] ? 4'ha : _GEN_387; // @[Filter.scala 191:62]
  wire [3:0] _GEN_389 = 10'hda == _T_43[9:0] ? 4'ha : _GEN_388; // @[Filter.scala 191:62]
  wire [3:0] _GEN_390 = 10'hdb == _T_43[9:0] ? 4'ha : _GEN_389; // @[Filter.scala 191:62]
  wire [3:0] _GEN_391 = 10'hdc == _T_43[9:0] ? 4'ha : _GEN_390; // @[Filter.scala 191:62]
  wire [3:0] _GEN_392 = 10'hdd == _T_43[9:0] ? 4'h3 : _GEN_391; // @[Filter.scala 191:62]
  wire [3:0] _GEN_393 = 10'hde == _T_43[9:0] ? 4'h2 : _GEN_392; // @[Filter.scala 191:62]
  wire [3:0] _GEN_394 = 10'hdf == _T_43[9:0] ? 4'h0 : _GEN_393; // @[Filter.scala 191:62]
  wire [3:0] _GEN_395 = 10'he0 == _T_43[9:0] ? 4'ha : _GEN_394; // @[Filter.scala 191:62]
  wire [3:0] _GEN_396 = 10'he1 == _T_43[9:0] ? 4'ha : _GEN_395; // @[Filter.scala 191:62]
  wire [3:0] _GEN_397 = 10'he2 == _T_43[9:0] ? 4'h3 : _GEN_396; // @[Filter.scala 191:62]
  wire [3:0] _GEN_398 = 10'he3 == _T_43[9:0] ? 4'ha : _GEN_397; // @[Filter.scala 191:62]
  wire [3:0] _GEN_399 = 10'he4 == _T_43[9:0] ? 4'ha : _GEN_398; // @[Filter.scala 191:62]
  wire [3:0] _GEN_400 = 10'he5 == _T_43[9:0] ? 4'ha : _GEN_399; // @[Filter.scala 191:62]
  wire [3:0] _GEN_401 = 10'he6 == _T_43[9:0] ? 4'ha : _GEN_400; // @[Filter.scala 191:62]
  wire [3:0] _GEN_402 = 10'he7 == _T_43[9:0] ? 4'h1 : _GEN_401; // @[Filter.scala 191:62]
  wire [3:0] _GEN_403 = 10'he8 == _T_43[9:0] ? 4'h1 : _GEN_402; // @[Filter.scala 191:62]
  wire [3:0] _GEN_404 = 10'he9 == _T_43[9:0] ? 4'h1 : _GEN_403; // @[Filter.scala 191:62]
  wire [3:0] _GEN_405 = 10'hea == _T_43[9:0] ? 4'h0 : _GEN_404; // @[Filter.scala 191:62]
  wire [3:0] _GEN_406 = 10'heb == _T_43[9:0] ? 4'h0 : _GEN_405; // @[Filter.scala 191:62]
  wire [3:0] _GEN_407 = 10'hec == _T_43[9:0] ? 4'h0 : _GEN_406; // @[Filter.scala 191:62]
  wire [3:0] _GEN_408 = 10'hed == _T_43[9:0] ? 4'h0 : _GEN_407; // @[Filter.scala 191:62]
  wire [3:0] _GEN_409 = 10'hee == _T_43[9:0] ? 4'h0 : _GEN_408; // @[Filter.scala 191:62]
  wire [3:0] _GEN_410 = 10'hef == _T_43[9:0] ? 4'h0 : _GEN_409; // @[Filter.scala 191:62]
  wire [3:0] _GEN_411 = 10'hf0 == _T_43[9:0] ? 4'h0 : _GEN_410; // @[Filter.scala 191:62]
  wire [3:0] _GEN_412 = 10'hf1 == _T_43[9:0] ? 4'h0 : _GEN_411; // @[Filter.scala 191:62]
  wire [3:0] _GEN_413 = 10'hf2 == _T_43[9:0] ? 4'h0 : _GEN_412; // @[Filter.scala 191:62]
  wire [3:0] _GEN_414 = 10'hf3 == _T_43[9:0] ? 4'h0 : _GEN_413; // @[Filter.scala 191:62]
  wire [3:0] _GEN_415 = 10'hf4 == _T_43[9:0] ? 4'h0 : _GEN_414; // @[Filter.scala 191:62]
  wire [3:0] _GEN_416 = 10'hf5 == _T_43[9:0] ? 4'h1 : _GEN_415; // @[Filter.scala 191:62]
  wire [3:0] _GEN_417 = 10'hf6 == _T_43[9:0] ? 4'h0 : _GEN_416; // @[Filter.scala 191:62]
  wire [3:0] _GEN_418 = 10'hf7 == _T_43[9:0] ? 4'h0 : _GEN_417; // @[Filter.scala 191:62]
  wire [3:0] _GEN_419 = 10'hf8 == _T_43[9:0] ? 4'h1 : _GEN_418; // @[Filter.scala 191:62]
  wire [3:0] _GEN_420 = 10'hf9 == _T_43[9:0] ? 4'h0 : _GEN_419; // @[Filter.scala 191:62]
  wire [3:0] _GEN_421 = 10'hfa == _T_43[9:0] ? 4'ha : _GEN_420; // @[Filter.scala 191:62]
  wire [3:0] _GEN_422 = 10'hfb == _T_43[9:0] ? 4'ha : _GEN_421; // @[Filter.scala 191:62]
  wire [3:0] _GEN_423 = 10'hfc == _T_43[9:0] ? 4'ha : _GEN_422; // @[Filter.scala 191:62]
  wire [3:0] _GEN_424 = 10'hfd == _T_43[9:0] ? 4'h3 : _GEN_423; // @[Filter.scala 191:62]
  wire [3:0] _GEN_425 = 10'hfe == _T_43[9:0] ? 4'ha : _GEN_424; // @[Filter.scala 191:62]
  wire [3:0] _GEN_426 = 10'hff == _T_43[9:0] ? 4'h0 : _GEN_425; // @[Filter.scala 191:62]
  wire [3:0] _GEN_427 = 10'h100 == _T_43[9:0] ? 4'ha : _GEN_426; // @[Filter.scala 191:62]
  wire [3:0] _GEN_428 = 10'h101 == _T_43[9:0] ? 4'h0 : _GEN_427; // @[Filter.scala 191:62]
  wire [3:0] _GEN_429 = 10'h102 == _T_43[9:0] ? 4'h3 : _GEN_428; // @[Filter.scala 191:62]
  wire [3:0] _GEN_430 = 10'h103 == _T_43[9:0] ? 4'ha : _GEN_429; // @[Filter.scala 191:62]
  wire [3:0] _GEN_431 = 10'h104 == _T_43[9:0] ? 4'ha : _GEN_430; // @[Filter.scala 191:62]
  wire [3:0] _GEN_432 = 10'h105 == _T_43[9:0] ? 4'ha : _GEN_431; // @[Filter.scala 191:62]
  wire [3:0] _GEN_433 = 10'h106 == _T_43[9:0] ? 4'ha : _GEN_432; // @[Filter.scala 191:62]
  wire [3:0] _GEN_434 = 10'h107 == _T_43[9:0] ? 4'ha : _GEN_433; // @[Filter.scala 191:62]
  wire [3:0] _GEN_435 = 10'h108 == _T_43[9:0] ? 4'h1 : _GEN_434; // @[Filter.scala 191:62]
  wire [3:0] _GEN_436 = 10'h109 == _T_43[9:0] ? 4'h0 : _GEN_435; // @[Filter.scala 191:62]
  wire [3:0] _GEN_437 = 10'h10a == _T_43[9:0] ? 4'h0 : _GEN_436; // @[Filter.scala 191:62]
  wire [3:0] _GEN_438 = 10'h10b == _T_43[9:0] ? 4'h0 : _GEN_437; // @[Filter.scala 191:62]
  wire [3:0] _GEN_439 = 10'h10c == _T_43[9:0] ? 4'h0 : _GEN_438; // @[Filter.scala 191:62]
  wire [3:0] _GEN_440 = 10'h10d == _T_43[9:0] ? 4'h0 : _GEN_439; // @[Filter.scala 191:62]
  wire [3:0] _GEN_441 = 10'h10e == _T_43[9:0] ? 4'h0 : _GEN_440; // @[Filter.scala 191:62]
  wire [3:0] _GEN_442 = 10'h10f == _T_43[9:0] ? 4'h0 : _GEN_441; // @[Filter.scala 191:62]
  wire [3:0] _GEN_443 = 10'h110 == _T_43[9:0] ? 4'h0 : _GEN_442; // @[Filter.scala 191:62]
  wire [3:0] _GEN_444 = 10'h111 == _T_43[9:0] ? 4'h0 : _GEN_443; // @[Filter.scala 191:62]
  wire [3:0] _GEN_445 = 10'h112 == _T_43[9:0] ? 4'h0 : _GEN_444; // @[Filter.scala 191:62]
  wire [3:0] _GEN_446 = 10'h113 == _T_43[9:0] ? 4'h0 : _GEN_445; // @[Filter.scala 191:62]
  wire [3:0] _GEN_447 = 10'h114 == _T_43[9:0] ? 4'h0 : _GEN_446; // @[Filter.scala 191:62]
  wire [3:0] _GEN_448 = 10'h115 == _T_43[9:0] ? 4'h0 : _GEN_447; // @[Filter.scala 191:62]
  wire [3:0] _GEN_449 = 10'h116 == _T_43[9:0] ? 4'h1 : _GEN_448; // @[Filter.scala 191:62]
  wire [3:0] _GEN_450 = 10'h117 == _T_43[9:0] ? 4'ha : _GEN_449; // @[Filter.scala 191:62]
  wire [3:0] _GEN_451 = 10'h118 == _T_43[9:0] ? 4'ha : _GEN_450; // @[Filter.scala 191:62]
  wire [3:0] _GEN_452 = 10'h119 == _T_43[9:0] ? 4'ha : _GEN_451; // @[Filter.scala 191:62]
  wire [3:0] _GEN_453 = 10'h11a == _T_43[9:0] ? 4'h0 : _GEN_452; // @[Filter.scala 191:62]
  wire [3:0] _GEN_454 = 10'h11b == _T_43[9:0] ? 4'ha : _GEN_453; // @[Filter.scala 191:62]
  wire [3:0] _GEN_455 = 10'h11c == _T_43[9:0] ? 4'ha : _GEN_454; // @[Filter.scala 191:62]
  wire [3:0] _GEN_456 = 10'h11d == _T_43[9:0] ? 4'h2 : _GEN_455; // @[Filter.scala 191:62]
  wire [3:0] _GEN_457 = 10'h11e == _T_43[9:0] ? 4'h3 : _GEN_456; // @[Filter.scala 191:62]
  wire [3:0] _GEN_458 = 10'h11f == _T_43[9:0] ? 4'h0 : _GEN_457; // @[Filter.scala 191:62]
  wire [3:0] _GEN_459 = 10'h120 == _T_43[9:0] ? 4'ha : _GEN_458; // @[Filter.scala 191:62]
  wire [3:0] _GEN_460 = 10'h121 == _T_43[9:0] ? 4'ha : _GEN_459; // @[Filter.scala 191:62]
  wire [3:0] _GEN_461 = 10'h122 == _T_43[9:0] ? 4'h3 : _GEN_460; // @[Filter.scala 191:62]
  wire [3:0] _GEN_462 = 10'h123 == _T_43[9:0] ? 4'ha : _GEN_461; // @[Filter.scala 191:62]
  wire [3:0] _GEN_463 = 10'h124 == _T_43[9:0] ? 4'ha : _GEN_462; // @[Filter.scala 191:62]
  wire [3:0] _GEN_464 = 10'h125 == _T_43[9:0] ? 4'ha : _GEN_463; // @[Filter.scala 191:62]
  wire [3:0] _GEN_465 = 10'h126 == _T_43[9:0] ? 4'ha : _GEN_464; // @[Filter.scala 191:62]
  wire [3:0] _GEN_466 = 10'h127 == _T_43[9:0] ? 4'h1 : _GEN_465; // @[Filter.scala 191:62]
  wire [3:0] _GEN_467 = 10'h128 == _T_43[9:0] ? 4'h0 : _GEN_466; // @[Filter.scala 191:62]
  wire [3:0] _GEN_468 = 10'h129 == _T_43[9:0] ? 4'ha : _GEN_467; // @[Filter.scala 191:62]
  wire [3:0] _GEN_469 = 10'h12a == _T_43[9:0] ? 4'ha : _GEN_468; // @[Filter.scala 191:62]
  wire [3:0] _GEN_470 = 10'h12b == _T_43[9:0] ? 4'h0 : _GEN_469; // @[Filter.scala 191:62]
  wire [3:0] _GEN_471 = 10'h12c == _T_43[9:0] ? 4'h0 : _GEN_470; // @[Filter.scala 191:62]
  wire [3:0] _GEN_472 = 10'h12d == _T_43[9:0] ? 4'h0 : _GEN_471; // @[Filter.scala 191:62]
  wire [3:0] _GEN_473 = 10'h12e == _T_43[9:0] ? 4'h0 : _GEN_472; // @[Filter.scala 191:62]
  wire [3:0] _GEN_474 = 10'h12f == _T_43[9:0] ? 4'h0 : _GEN_473; // @[Filter.scala 191:62]
  wire [3:0] _GEN_475 = 10'h130 == _T_43[9:0] ? 4'h0 : _GEN_474; // @[Filter.scala 191:62]
  wire [3:0] _GEN_476 = 10'h131 == _T_43[9:0] ? 4'h0 : _GEN_475; // @[Filter.scala 191:62]
  wire [3:0] _GEN_477 = 10'h132 == _T_43[9:0] ? 4'h0 : _GEN_476; // @[Filter.scala 191:62]
  wire [3:0] _GEN_478 = 10'h133 == _T_43[9:0] ? 4'h0 : _GEN_477; // @[Filter.scala 191:62]
  wire [3:0] _GEN_479 = 10'h134 == _T_43[9:0] ? 4'ha : _GEN_478; // @[Filter.scala 191:62]
  wire [3:0] _GEN_480 = 10'h135 == _T_43[9:0] ? 4'ha : _GEN_479; // @[Filter.scala 191:62]
  wire [3:0] _GEN_481 = 10'h136 == _T_43[9:0] ? 4'h0 : _GEN_480; // @[Filter.scala 191:62]
  wire [3:0] _GEN_482 = 10'h137 == _T_43[9:0] ? 4'h1 : _GEN_481; // @[Filter.scala 191:62]
  wire [3:0] _GEN_483 = 10'h138 == _T_43[9:0] ? 4'ha : _GEN_482; // @[Filter.scala 191:62]
  wire [3:0] _GEN_484 = 10'h139 == _T_43[9:0] ? 4'ha : _GEN_483; // @[Filter.scala 191:62]
  wire [3:0] _GEN_485 = 10'h13a == _T_43[9:0] ? 4'ha : _GEN_484; // @[Filter.scala 191:62]
  wire [3:0] _GEN_486 = 10'h13b == _T_43[9:0] ? 4'ha : _GEN_485; // @[Filter.scala 191:62]
  wire [3:0] _GEN_487 = 10'h13c == _T_43[9:0] ? 4'ha : _GEN_486; // @[Filter.scala 191:62]
  wire [3:0] _GEN_488 = 10'h13d == _T_43[9:0] ? 4'ha : _GEN_487; // @[Filter.scala 191:62]
  wire [3:0] _GEN_489 = 10'h13e == _T_43[9:0] ? 4'h3 : _GEN_488; // @[Filter.scala 191:62]
  wire [3:0] _GEN_490 = 10'h13f == _T_43[9:0] ? 4'h0 : _GEN_489; // @[Filter.scala 191:62]
  wire [3:0] _GEN_491 = 10'h140 == _T_43[9:0] ? 4'ha : _GEN_490; // @[Filter.scala 191:62]
  wire [3:0] _GEN_492 = 10'h141 == _T_43[9:0] ? 4'ha : _GEN_491; // @[Filter.scala 191:62]
  wire [3:0] _GEN_493 = 10'h142 == _T_43[9:0] ? 4'h2 : _GEN_492; // @[Filter.scala 191:62]
  wire [3:0] _GEN_494 = 10'h143 == _T_43[9:0] ? 4'h3 : _GEN_493; // @[Filter.scala 191:62]
  wire [3:0] _GEN_495 = 10'h144 == _T_43[9:0] ? 4'ha : _GEN_494; // @[Filter.scala 191:62]
  wire [3:0] _GEN_496 = 10'h145 == _T_43[9:0] ? 4'ha : _GEN_495; // @[Filter.scala 191:62]
  wire [3:0] _GEN_497 = 10'h146 == _T_43[9:0] ? 4'h1 : _GEN_496; // @[Filter.scala 191:62]
  wire [3:0] _GEN_498 = 10'h147 == _T_43[9:0] ? 4'h0 : _GEN_497; // @[Filter.scala 191:62]
  wire [3:0] _GEN_499 = 10'h148 == _T_43[9:0] ? 4'ha : _GEN_498; // @[Filter.scala 191:62]
  wire [3:0] _GEN_500 = 10'h149 == _T_43[9:0] ? 4'ha : _GEN_499; // @[Filter.scala 191:62]
  wire [3:0] _GEN_501 = 10'h14a == _T_43[9:0] ? 4'ha : _GEN_500; // @[Filter.scala 191:62]
  wire [3:0] _GEN_502 = 10'h14b == _T_43[9:0] ? 4'ha : _GEN_501; // @[Filter.scala 191:62]
  wire [3:0] _GEN_503 = 10'h14c == _T_43[9:0] ? 4'ha : _GEN_502; // @[Filter.scala 191:62]
  wire [3:0] _GEN_504 = 10'h14d == _T_43[9:0] ? 4'ha : _GEN_503; // @[Filter.scala 191:62]
  wire [3:0] _GEN_505 = 10'h14e == _T_43[9:0] ? 4'ha : _GEN_504; // @[Filter.scala 191:62]
  wire [3:0] _GEN_506 = 10'h14f == _T_43[9:0] ? 4'ha : _GEN_505; // @[Filter.scala 191:62]
  wire [3:0] _GEN_507 = 10'h150 == _T_43[9:0] ? 4'ha : _GEN_506; // @[Filter.scala 191:62]
  wire [3:0] _GEN_508 = 10'h151 == _T_43[9:0] ? 4'ha : _GEN_507; // @[Filter.scala 191:62]
  wire [3:0] _GEN_509 = 10'h152 == _T_43[9:0] ? 4'ha : _GEN_508; // @[Filter.scala 191:62]
  wire [3:0] _GEN_510 = 10'h153 == _T_43[9:0] ? 4'ha : _GEN_509; // @[Filter.scala 191:62]
  wire [3:0] _GEN_511 = 10'h154 == _T_43[9:0] ? 4'ha : _GEN_510; // @[Filter.scala 191:62]
  wire [3:0] _GEN_512 = 10'h155 == _T_43[9:0] ? 4'ha : _GEN_511; // @[Filter.scala 191:62]
  wire [3:0] _GEN_513 = 10'h156 == _T_43[9:0] ? 4'ha : _GEN_512; // @[Filter.scala 191:62]
  wire [3:0] _GEN_514 = 10'h157 == _T_43[9:0] ? 4'h0 : _GEN_513; // @[Filter.scala 191:62]
  wire [3:0] _GEN_515 = 10'h158 == _T_43[9:0] ? 4'ha : _GEN_514; // @[Filter.scala 191:62]
  wire [3:0] _GEN_516 = 10'h159 == _T_43[9:0] ? 4'ha : _GEN_515; // @[Filter.scala 191:62]
  wire [3:0] _GEN_517 = 10'h15a == _T_43[9:0] ? 4'ha : _GEN_516; // @[Filter.scala 191:62]
  wire [3:0] _GEN_518 = 10'h15b == _T_43[9:0] ? 4'ha : _GEN_517; // @[Filter.scala 191:62]
  wire [3:0] _GEN_519 = 10'h15c == _T_43[9:0] ? 4'ha : _GEN_518; // @[Filter.scala 191:62]
  wire [3:0] _GEN_520 = 10'h15d == _T_43[9:0] ? 4'h3 : _GEN_519; // @[Filter.scala 191:62]
  wire [3:0] _GEN_521 = 10'h15e == _T_43[9:0] ? 4'h2 : _GEN_520; // @[Filter.scala 191:62]
  wire [3:0] _GEN_522 = 10'h15f == _T_43[9:0] ? 4'h0 : _GEN_521; // @[Filter.scala 191:62]
  wire [3:0] _GEN_523 = 10'h160 == _T_43[9:0] ? 4'ha : _GEN_522; // @[Filter.scala 191:62]
  wire [3:0] _GEN_524 = 10'h161 == _T_43[9:0] ? 4'ha : _GEN_523; // @[Filter.scala 191:62]
  wire [3:0] _GEN_525 = 10'h162 == _T_43[9:0] ? 4'ha : _GEN_524; // @[Filter.scala 191:62]
  wire [3:0] _GEN_526 = 10'h163 == _T_43[9:0] ? 4'h2 : _GEN_525; // @[Filter.scala 191:62]
  wire [3:0] _GEN_527 = 10'h164 == _T_43[9:0] ? 4'h3 : _GEN_526; // @[Filter.scala 191:62]
  wire [3:0] _GEN_528 = 10'h165 == _T_43[9:0] ? 4'h1 : _GEN_527; // @[Filter.scala 191:62]
  wire [3:0] _GEN_529 = 10'h166 == _T_43[9:0] ? 4'h0 : _GEN_528; // @[Filter.scala 191:62]
  wire [3:0] _GEN_530 = 10'h167 == _T_43[9:0] ? 4'h0 : _GEN_529; // @[Filter.scala 191:62]
  wire [3:0] _GEN_531 = 10'h168 == _T_43[9:0] ? 4'h5 : _GEN_530; // @[Filter.scala 191:62]
  wire [3:0] _GEN_532 = 10'h169 == _T_43[9:0] ? 4'h3 : _GEN_531; // @[Filter.scala 191:62]
  wire [3:0] _GEN_533 = 10'h16a == _T_43[9:0] ? 4'h5 : _GEN_532; // @[Filter.scala 191:62]
  wire [3:0] _GEN_534 = 10'h16b == _T_43[9:0] ? 4'h5 : _GEN_533; // @[Filter.scala 191:62]
  wire [3:0] _GEN_535 = 10'h16c == _T_43[9:0] ? 4'ha : _GEN_534; // @[Filter.scala 191:62]
  wire [3:0] _GEN_536 = 10'h16d == _T_43[9:0] ? 4'ha : _GEN_535; // @[Filter.scala 191:62]
  wire [3:0] _GEN_537 = 10'h16e == _T_43[9:0] ? 4'ha : _GEN_536; // @[Filter.scala 191:62]
  wire [3:0] _GEN_538 = 10'h16f == _T_43[9:0] ? 4'ha : _GEN_537; // @[Filter.scala 191:62]
  wire [3:0] _GEN_539 = 10'h170 == _T_43[9:0] ? 4'ha : _GEN_538; // @[Filter.scala 191:62]
  wire [3:0] _GEN_540 = 10'h171 == _T_43[9:0] ? 4'ha : _GEN_539; // @[Filter.scala 191:62]
  wire [3:0] _GEN_541 = 10'h172 == _T_43[9:0] ? 4'ha : _GEN_540; // @[Filter.scala 191:62]
  wire [3:0] _GEN_542 = 10'h173 == _T_43[9:0] ? 4'ha : _GEN_541; // @[Filter.scala 191:62]
  wire [3:0] _GEN_543 = 10'h174 == _T_43[9:0] ? 4'ha : _GEN_542; // @[Filter.scala 191:62]
  wire [3:0] _GEN_544 = 10'h175 == _T_43[9:0] ? 4'ha : _GEN_543; // @[Filter.scala 191:62]
  wire [3:0] _GEN_545 = 10'h176 == _T_43[9:0] ? 4'h0 : _GEN_544; // @[Filter.scala 191:62]
  wire [3:0] _GEN_546 = 10'h177 == _T_43[9:0] ? 4'h0 : _GEN_545; // @[Filter.scala 191:62]
  wire [3:0] _GEN_547 = 10'h178 == _T_43[9:0] ? 4'h1 : _GEN_546; // @[Filter.scala 191:62]
  wire [3:0] _GEN_548 = 10'h179 == _T_43[9:0] ? 4'ha : _GEN_547; // @[Filter.scala 191:62]
  wire [3:0] _GEN_549 = 10'h17a == _T_43[9:0] ? 4'ha : _GEN_548; // @[Filter.scala 191:62]
  wire [3:0] _GEN_550 = 10'h17b == _T_43[9:0] ? 4'ha : _GEN_549; // @[Filter.scala 191:62]
  wire [3:0] _GEN_551 = 10'h17c == _T_43[9:0] ? 4'h3 : _GEN_550; // @[Filter.scala 191:62]
  wire [3:0] _GEN_552 = 10'h17d == _T_43[9:0] ? 4'h2 : _GEN_551; // @[Filter.scala 191:62]
  wire [3:0] _GEN_553 = 10'h17e == _T_43[9:0] ? 4'ha : _GEN_552; // @[Filter.scala 191:62]
  wire [3:0] _GEN_554 = 10'h17f == _T_43[9:0] ? 4'h0 : _GEN_553; // @[Filter.scala 191:62]
  wire [3:0] _GEN_555 = 10'h180 == _T_43[9:0] ? 4'h5 : _GEN_554; // @[Filter.scala 191:62]
  wire [3:0] _GEN_556 = 10'h181 == _T_43[9:0] ? 4'h5 : _GEN_555; // @[Filter.scala 191:62]
  wire [3:0] _GEN_557 = 10'h182 == _T_43[9:0] ? 4'h5 : _GEN_556; // @[Filter.scala 191:62]
  wire [3:0] _GEN_558 = 10'h183 == _T_43[9:0] ? 4'h5 : _GEN_557; // @[Filter.scala 191:62]
  wire [3:0] _GEN_559 = 10'h184 == _T_43[9:0] ? 4'h3 : _GEN_558; // @[Filter.scala 191:62]
  wire [3:0] _GEN_560 = 10'h185 == _T_43[9:0] ? 4'h1 : _GEN_559; // @[Filter.scala 191:62]
  wire [3:0] _GEN_561 = 10'h186 == _T_43[9:0] ? 4'hb : _GEN_560; // @[Filter.scala 191:62]
  wire [3:0] _GEN_562 = 10'h187 == _T_43[9:0] ? 4'h0 : _GEN_561; // @[Filter.scala 191:62]
  wire [3:0] _GEN_563 = 10'h188 == _T_43[9:0] ? 4'h5 : _GEN_562; // @[Filter.scala 191:62]
  wire [3:0] _GEN_564 = 10'h189 == _T_43[9:0] ? 4'h5 : _GEN_563; // @[Filter.scala 191:62]
  wire [3:0] _GEN_565 = 10'h18a == _T_43[9:0] ? 4'h5 : _GEN_564; // @[Filter.scala 191:62]
  wire [3:0] _GEN_566 = 10'h18b == _T_43[9:0] ? 4'h5 : _GEN_565; // @[Filter.scala 191:62]
  wire [3:0] _GEN_567 = 10'h18c == _T_43[9:0] ? 4'h5 : _GEN_566; // @[Filter.scala 191:62]
  wire [3:0] _GEN_568 = 10'h18d == _T_43[9:0] ? 4'h5 : _GEN_567; // @[Filter.scala 191:62]
  wire [3:0] _GEN_569 = 10'h18e == _T_43[9:0] ? 4'h5 : _GEN_568; // @[Filter.scala 191:62]
  wire [3:0] _GEN_570 = 10'h18f == _T_43[9:0] ? 4'h5 : _GEN_569; // @[Filter.scala 191:62]
  wire [3:0] _GEN_571 = 10'h190 == _T_43[9:0] ? 4'h5 : _GEN_570; // @[Filter.scala 191:62]
  wire [3:0] _GEN_572 = 10'h191 == _T_43[9:0] ? 4'h5 : _GEN_571; // @[Filter.scala 191:62]
  wire [3:0] _GEN_573 = 10'h192 == _T_43[9:0] ? 4'h3 : _GEN_572; // @[Filter.scala 191:62]
  wire [3:0] _GEN_574 = 10'h193 == _T_43[9:0] ? 4'h5 : _GEN_573; // @[Filter.scala 191:62]
  wire [3:0] _GEN_575 = 10'h194 == _T_43[9:0] ? 4'h5 : _GEN_574; // @[Filter.scala 191:62]
  wire [3:0] _GEN_576 = 10'h195 == _T_43[9:0] ? 4'h5 : _GEN_575; // @[Filter.scala 191:62]
  wire [3:0] _GEN_577 = 10'h196 == _T_43[9:0] ? 4'h0 : _GEN_576; // @[Filter.scala 191:62]
  wire [3:0] _GEN_578 = 10'h197 == _T_43[9:0] ? 4'ha : _GEN_577; // @[Filter.scala 191:62]
  wire [3:0] _GEN_579 = 10'h198 == _T_43[9:0] ? 4'h1 : _GEN_578; // @[Filter.scala 191:62]
  wire [3:0] _GEN_580 = 10'h199 == _T_43[9:0] ? 4'ha : _GEN_579; // @[Filter.scala 191:62]
  wire [3:0] _GEN_581 = 10'h19a == _T_43[9:0] ? 4'ha : _GEN_580; // @[Filter.scala 191:62]
  wire [3:0] _GEN_582 = 10'h19b == _T_43[9:0] ? 4'ha : _GEN_581; // @[Filter.scala 191:62]
  wire [3:0] _GEN_583 = 10'h19c == _T_43[9:0] ? 4'h3 : _GEN_582; // @[Filter.scala 191:62]
  wire [3:0] _GEN_584 = 10'h19d == _T_43[9:0] ? 4'ha : _GEN_583; // @[Filter.scala 191:62]
  wire [3:0] _GEN_585 = 10'h19e == _T_43[9:0] ? 4'ha : _GEN_584; // @[Filter.scala 191:62]
  wire [3:0] _GEN_586 = 10'h19f == _T_43[9:0] ? 4'h0 : _GEN_585; // @[Filter.scala 191:62]
  wire [3:0] _GEN_587 = 10'h1a0 == _T_43[9:0] ? 4'h5 : _GEN_586; // @[Filter.scala 191:62]
  wire [3:0] _GEN_588 = 10'h1a1 == _T_43[9:0] ? 4'h5 : _GEN_587; // @[Filter.scala 191:62]
  wire [3:0] _GEN_589 = 10'h1a2 == _T_43[9:0] ? 4'h3 : _GEN_588; // @[Filter.scala 191:62]
  wire [3:0] _GEN_590 = 10'h1a3 == _T_43[9:0] ? 4'h5 : _GEN_589; // @[Filter.scala 191:62]
  wire [3:0] _GEN_591 = 10'h1a4 == _T_43[9:0] ? 4'h3 : _GEN_590; // @[Filter.scala 191:62]
  wire [3:0] _GEN_592 = 10'h1a5 == _T_43[9:0] ? 4'h0 : _GEN_591; // @[Filter.scala 191:62]
  wire [3:0] _GEN_593 = 10'h1a6 == _T_43[9:0] ? 4'h5 : _GEN_592; // @[Filter.scala 191:62]
  wire [3:0] _GEN_594 = 10'h1a7 == _T_43[9:0] ? 4'h0 : _GEN_593; // @[Filter.scala 191:62]
  wire [3:0] _GEN_595 = 10'h1a8 == _T_43[9:0] ? 4'hb : _GEN_594; // @[Filter.scala 191:62]
  wire [3:0] _GEN_596 = 10'h1a9 == _T_43[9:0] ? 4'h5 : _GEN_595; // @[Filter.scala 191:62]
  wire [3:0] _GEN_597 = 10'h1aa == _T_43[9:0] ? 4'h5 : _GEN_596; // @[Filter.scala 191:62]
  wire [3:0] _GEN_598 = 10'h1ab == _T_43[9:0] ? 4'h3 : _GEN_597; // @[Filter.scala 191:62]
  wire [3:0] _GEN_599 = 10'h1ac == _T_43[9:0] ? 4'h5 : _GEN_598; // @[Filter.scala 191:62]
  wire [3:0] _GEN_600 = 10'h1ad == _T_43[9:0] ? 4'h5 : _GEN_599; // @[Filter.scala 191:62]
  wire [3:0] _GEN_601 = 10'h1ae == _T_43[9:0] ? 4'h5 : _GEN_600; // @[Filter.scala 191:62]
  wire [3:0] _GEN_602 = 10'h1af == _T_43[9:0] ? 4'h5 : _GEN_601; // @[Filter.scala 191:62]
  wire [3:0] _GEN_603 = 10'h1b0 == _T_43[9:0] ? 4'h5 : _GEN_602; // @[Filter.scala 191:62]
  wire [3:0] _GEN_604 = 10'h1b1 == _T_43[9:0] ? 4'h5 : _GEN_603; // @[Filter.scala 191:62]
  wire [3:0] _GEN_605 = 10'h1b2 == _T_43[9:0] ? 4'h5 : _GEN_604; // @[Filter.scala 191:62]
  wire [3:0] _GEN_606 = 10'h1b3 == _T_43[9:0] ? 4'h5 : _GEN_605; // @[Filter.scala 191:62]
  wire [3:0] _GEN_607 = 10'h1b4 == _T_43[9:0] ? 4'h5 : _GEN_606; // @[Filter.scala 191:62]
  wire [3:0] _GEN_608 = 10'h1b5 == _T_43[9:0] ? 4'h5 : _GEN_607; // @[Filter.scala 191:62]
  wire [3:0] _GEN_609 = 10'h1b6 == _T_43[9:0] ? 4'h0 : _GEN_608; // @[Filter.scala 191:62]
  wire [3:0] _GEN_610 = 10'h1b7 == _T_43[9:0] ? 4'h5 : _GEN_609; // @[Filter.scala 191:62]
  wire [3:0] _GEN_611 = 10'h1b8 == _T_43[9:0] ? 4'h0 : _GEN_610; // @[Filter.scala 191:62]
  wire [3:0] _GEN_612 = 10'h1b9 == _T_43[9:0] ? 4'h5 : _GEN_611; // @[Filter.scala 191:62]
  wire [3:0] _GEN_613 = 10'h1ba == _T_43[9:0] ? 4'h5 : _GEN_612; // @[Filter.scala 191:62]
  wire [3:0] _GEN_614 = 10'h1bb == _T_43[9:0] ? 4'h5 : _GEN_613; // @[Filter.scala 191:62]
  wire [3:0] _GEN_615 = 10'h1bc == _T_43[9:0] ? 4'h2 : _GEN_614; // @[Filter.scala 191:62]
  wire [3:0] _GEN_616 = 10'h1bd == _T_43[9:0] ? 4'h3 : _GEN_615; // @[Filter.scala 191:62]
  wire [3:0] _GEN_617 = 10'h1be == _T_43[9:0] ? 4'h5 : _GEN_616; // @[Filter.scala 191:62]
  wire [3:0] _GEN_618 = 10'h1bf == _T_43[9:0] ? 4'h0 : _GEN_617; // @[Filter.scala 191:62]
  wire [3:0] _GEN_619 = 10'h1c0 == _T_43[9:0] ? 4'h5 : _GEN_618; // @[Filter.scala 191:62]
  wire [3:0] _GEN_620 = 10'h1c1 == _T_43[9:0] ? 4'h5 : _GEN_619; // @[Filter.scala 191:62]
  wire [3:0] _GEN_621 = 10'h1c2 == _T_43[9:0] ? 4'h5 : _GEN_620; // @[Filter.scala 191:62]
  wire [3:0] _GEN_622 = 10'h1c3 == _T_43[9:0] ? 4'h2 : _GEN_621; // @[Filter.scala 191:62]
  wire [3:0] _GEN_623 = 10'h1c4 == _T_43[9:0] ? 4'h2 : _GEN_622; // @[Filter.scala 191:62]
  wire [3:0] _GEN_624 = 10'h1c5 == _T_43[9:0] ? 4'h5 : _GEN_623; // @[Filter.scala 191:62]
  wire [3:0] _GEN_625 = 10'h1c6 == _T_43[9:0] ? 4'h5 : _GEN_624; // @[Filter.scala 191:62]
  wire [3:0] _GEN_626 = 10'h1c7 == _T_43[9:0] ? 4'h5 : _GEN_625; // @[Filter.scala 191:62]
  wire [3:0] _GEN_627 = 10'h1c8 == _T_43[9:0] ? 4'h5 : _GEN_626; // @[Filter.scala 191:62]
  wire [3:0] _GEN_628 = 10'h1c9 == _T_43[9:0] ? 4'hb : _GEN_627; // @[Filter.scala 191:62]
  wire [3:0] _GEN_629 = 10'h1ca == _T_43[9:0] ? 4'hb : _GEN_628; // @[Filter.scala 191:62]
  wire [3:0] _GEN_630 = 10'h1cb == _T_43[9:0] ? 4'hb : _GEN_629; // @[Filter.scala 191:62]
  wire [3:0] _GEN_631 = 10'h1cc == _T_43[9:0] ? 4'hb : _GEN_630; // @[Filter.scala 191:62]
  wire [3:0] _GEN_632 = 10'h1cd == _T_43[9:0] ? 4'hb : _GEN_631; // @[Filter.scala 191:62]
  wire [3:0] _GEN_633 = 10'h1ce == _T_43[9:0] ? 4'hb : _GEN_632; // @[Filter.scala 191:62]
  wire [3:0] _GEN_634 = 10'h1cf == _T_43[9:0] ? 4'hb : _GEN_633; // @[Filter.scala 191:62]
  wire [3:0] _GEN_635 = 10'h1d0 == _T_43[9:0] ? 4'hb : _GEN_634; // @[Filter.scala 191:62]
  wire [3:0] _GEN_636 = 10'h1d1 == _T_43[9:0] ? 4'hb : _GEN_635; // @[Filter.scala 191:62]
  wire [3:0] _GEN_637 = 10'h1d2 == _T_43[9:0] ? 4'hb : _GEN_636; // @[Filter.scala 191:62]
  wire [3:0] _GEN_638 = 10'h1d3 == _T_43[9:0] ? 4'hb : _GEN_637; // @[Filter.scala 191:62]
  wire [3:0] _GEN_639 = 10'h1d4 == _T_43[9:0] ? 4'hb : _GEN_638; // @[Filter.scala 191:62]
  wire [3:0] _GEN_640 = 10'h1d5 == _T_43[9:0] ? 4'hb : _GEN_639; // @[Filter.scala 191:62]
  wire [3:0] _GEN_641 = 10'h1d6 == _T_43[9:0] ? 4'h5 : _GEN_640; // @[Filter.scala 191:62]
  wire [3:0] _GEN_642 = 10'h1d7 == _T_43[9:0] ? 4'h5 : _GEN_641; // @[Filter.scala 191:62]
  wire [3:0] _GEN_643 = 10'h1d8 == _T_43[9:0] ? 4'h5 : _GEN_642; // @[Filter.scala 191:62]
  wire [3:0] _GEN_644 = 10'h1d9 == _T_43[9:0] ? 4'h5 : _GEN_643; // @[Filter.scala 191:62]
  wire [3:0] _GEN_645 = 10'h1da == _T_43[9:0] ? 4'h5 : _GEN_644; // @[Filter.scala 191:62]
  wire [3:0] _GEN_646 = 10'h1db == _T_43[9:0] ? 4'h5 : _GEN_645; // @[Filter.scala 191:62]
  wire [3:0] _GEN_647 = 10'h1dc == _T_43[9:0] ? 4'h5 : _GEN_646; // @[Filter.scala 191:62]
  wire [3:0] _GEN_648 = 10'h1dd == _T_43[9:0] ? 4'h3 : _GEN_647; // @[Filter.scala 191:62]
  wire [3:0] _GEN_649 = 10'h1de == _T_43[9:0] ? 4'h5 : _GEN_648; // @[Filter.scala 191:62]
  wire [3:0] _GEN_650 = 10'h1df == _T_43[9:0] ? 4'h0 : _GEN_649; // @[Filter.scala 191:62]
  wire [3:0] _GEN_651 = 10'h1e0 == _T_43[9:0] ? 4'h3 : _GEN_650; // @[Filter.scala 191:62]
  wire [3:0] _GEN_652 = 10'h1e1 == _T_43[9:0] ? 4'h5 : _GEN_651; // @[Filter.scala 191:62]
  wire [3:0] _GEN_653 = 10'h1e2 == _T_43[9:0] ? 4'h2 : _GEN_652; // @[Filter.scala 191:62]
  wire [3:0] _GEN_654 = 10'h1e3 == _T_43[9:0] ? 4'h2 : _GEN_653; // @[Filter.scala 191:62]
  wire [3:0] _GEN_655 = 10'h1e4 == _T_43[9:0] ? 4'h5 : _GEN_654; // @[Filter.scala 191:62]
  wire [3:0] _GEN_656 = 10'h1e5 == _T_43[9:0] ? 4'h5 : _GEN_655; // @[Filter.scala 191:62]
  wire [3:0] _GEN_657 = 10'h1e6 == _T_43[9:0] ? 4'h5 : _GEN_656; // @[Filter.scala 191:62]
  wire [3:0] _GEN_658 = 10'h1e7 == _T_43[9:0] ? 4'h5 : _GEN_657; // @[Filter.scala 191:62]
  wire [3:0] _GEN_659 = 10'h1e8 == _T_43[9:0] ? 4'hb : _GEN_658; // @[Filter.scala 191:62]
  wire [3:0] _GEN_660 = 10'h1e9 == _T_43[9:0] ? 4'h5 : _GEN_659; // @[Filter.scala 191:62]
  wire [3:0] _GEN_661 = 10'h1ea == _T_43[9:0] ? 4'h5 : _GEN_660; // @[Filter.scala 191:62]
  wire [3:0] _GEN_662 = 10'h1eb == _T_43[9:0] ? 4'hb : _GEN_661; // @[Filter.scala 191:62]
  wire [3:0] _GEN_663 = 10'h1ec == _T_43[9:0] ? 4'h5 : _GEN_662; // @[Filter.scala 191:62]
  wire [3:0] _GEN_664 = 10'h1ed == _T_43[9:0] ? 4'hb : _GEN_663; // @[Filter.scala 191:62]
  wire [3:0] _GEN_665 = 10'h1ee == _T_43[9:0] ? 4'h5 : _GEN_664; // @[Filter.scala 191:62]
  wire [3:0] _GEN_666 = 10'h1ef == _T_43[9:0] ? 4'hb : _GEN_665; // @[Filter.scala 191:62]
  wire [3:0] _GEN_667 = 10'h1f0 == _T_43[9:0] ? 4'h5 : _GEN_666; // @[Filter.scala 191:62]
  wire [3:0] _GEN_668 = 10'h1f1 == _T_43[9:0] ? 4'hb : _GEN_667; // @[Filter.scala 191:62]
  wire [3:0] _GEN_669 = 10'h1f2 == _T_43[9:0] ? 4'hb : _GEN_668; // @[Filter.scala 191:62]
  wire [3:0] _GEN_670 = 10'h1f3 == _T_43[9:0] ? 4'h5 : _GEN_669; // @[Filter.scala 191:62]
  wire [3:0] _GEN_671 = 10'h1f4 == _T_43[9:0] ? 4'hb : _GEN_670; // @[Filter.scala 191:62]
  wire [3:0] _GEN_672 = 10'h1f5 == _T_43[9:0] ? 4'hb : _GEN_671; // @[Filter.scala 191:62]
  wire [3:0] _GEN_673 = 10'h1f6 == _T_43[9:0] ? 4'h5 : _GEN_672; // @[Filter.scala 191:62]
  wire [3:0] _GEN_674 = 10'h1f7 == _T_43[9:0] ? 4'h5 : _GEN_673; // @[Filter.scala 191:62]
  wire [3:0] _GEN_675 = 10'h1f8 == _T_43[9:0] ? 4'h5 : _GEN_674; // @[Filter.scala 191:62]
  wire [3:0] _GEN_676 = 10'h1f9 == _T_43[9:0] ? 4'h5 : _GEN_675; // @[Filter.scala 191:62]
  wire [3:0] _GEN_677 = 10'h1fa == _T_43[9:0] ? 4'h3 : _GEN_676; // @[Filter.scala 191:62]
  wire [3:0] _GEN_678 = 10'h1fb == _T_43[9:0] ? 4'h5 : _GEN_677; // @[Filter.scala 191:62]
  wire [3:0] _GEN_679 = 10'h1fc == _T_43[9:0] ? 4'h5 : _GEN_678; // @[Filter.scala 191:62]
  wire [3:0] _GEN_680 = 10'h1fd == _T_43[9:0] ? 4'h2 : _GEN_679; // @[Filter.scala 191:62]
  wire [3:0] _GEN_681 = 10'h1fe == _T_43[9:0] ? 4'h5 : _GEN_680; // @[Filter.scala 191:62]
  wire [3:0] _GEN_682 = 10'h1ff == _T_43[9:0] ? 4'h0 : _GEN_681; // @[Filter.scala 191:62]
  wire [3:0] _GEN_683 = 10'h200 == _T_43[9:0] ? 4'h5 : _GEN_682; // @[Filter.scala 191:62]
  wire [3:0] _GEN_684 = 10'h201 == _T_43[9:0] ? 4'h5 : _GEN_683; // @[Filter.scala 191:62]
  wire [3:0] _GEN_685 = 10'h202 == _T_43[9:0] ? 4'h3 : _GEN_684; // @[Filter.scala 191:62]
  wire [3:0] _GEN_686 = 10'h203 == _T_43[9:0] ? 4'h5 : _GEN_685; // @[Filter.scala 191:62]
  wire [3:0] _GEN_687 = 10'h204 == _T_43[9:0] ? 4'h5 : _GEN_686; // @[Filter.scala 191:62]
  wire [3:0] _GEN_688 = 10'h205 == _T_43[9:0] ? 4'h5 : _GEN_687; // @[Filter.scala 191:62]
  wire [3:0] _GEN_689 = 10'h206 == _T_43[9:0] ? 4'hb : _GEN_688; // @[Filter.scala 191:62]
  wire [3:0] _GEN_690 = 10'h207 == _T_43[9:0] ? 4'hb : _GEN_689; // @[Filter.scala 191:62]
  wire [3:0] _GEN_691 = 10'h208 == _T_43[9:0] ? 4'h5 : _GEN_690; // @[Filter.scala 191:62]
  wire [3:0] _GEN_692 = 10'h209 == _T_43[9:0] ? 4'h5 : _GEN_691; // @[Filter.scala 191:62]
  wire [3:0] _GEN_693 = 10'h20a == _T_43[9:0] ? 4'h5 : _GEN_692; // @[Filter.scala 191:62]
  wire [3:0] _GEN_694 = 10'h20b == _T_43[9:0] ? 4'hb : _GEN_693; // @[Filter.scala 191:62]
  wire [3:0] _GEN_695 = 10'h20c == _T_43[9:0] ? 4'h5 : _GEN_694; // @[Filter.scala 191:62]
  wire [3:0] _GEN_696 = 10'h20d == _T_43[9:0] ? 4'hb : _GEN_695; // @[Filter.scala 191:62]
  wire [3:0] _GEN_697 = 10'h20e == _T_43[9:0] ? 4'h5 : _GEN_696; // @[Filter.scala 191:62]
  wire [3:0] _GEN_698 = 10'h20f == _T_43[9:0] ? 4'hb : _GEN_697; // @[Filter.scala 191:62]
  wire [3:0] _GEN_699 = 10'h210 == _T_43[9:0] ? 4'h5 : _GEN_698; // @[Filter.scala 191:62]
  wire [3:0] _GEN_700 = 10'h211 == _T_43[9:0] ? 4'h5 : _GEN_699; // @[Filter.scala 191:62]
  wire [3:0] _GEN_701 = 10'h212 == _T_43[9:0] ? 4'hb : _GEN_700; // @[Filter.scala 191:62]
  wire [3:0] _GEN_702 = 10'h213 == _T_43[9:0] ? 4'hb : _GEN_701; // @[Filter.scala 191:62]
  wire [3:0] _GEN_703 = 10'h214 == _T_43[9:0] ? 4'hb : _GEN_702; // @[Filter.scala 191:62]
  wire [3:0] _GEN_704 = 10'h215 == _T_43[9:0] ? 4'h5 : _GEN_703; // @[Filter.scala 191:62]
  wire [3:0] _GEN_705 = 10'h216 == _T_43[9:0] ? 4'h5 : _GEN_704; // @[Filter.scala 191:62]
  wire [3:0] _GEN_706 = 10'h217 == _T_43[9:0] ? 4'h5 : _GEN_705; // @[Filter.scala 191:62]
  wire [3:0] _GEN_707 = 10'h218 == _T_43[9:0] ? 4'h5 : _GEN_706; // @[Filter.scala 191:62]
  wire [3:0] _GEN_708 = 10'h219 == _T_43[9:0] ? 4'h5 : _GEN_707; // @[Filter.scala 191:62]
  wire [3:0] _GEN_709 = 10'h21a == _T_43[9:0] ? 4'h5 : _GEN_708; // @[Filter.scala 191:62]
  wire [3:0] _GEN_710 = 10'h21b == _T_43[9:0] ? 4'h5 : _GEN_709; // @[Filter.scala 191:62]
  wire [3:0] _GEN_711 = 10'h21c == _T_43[9:0] ? 4'h3 : _GEN_710; // @[Filter.scala 191:62]
  wire [3:0] _GEN_712 = 10'h21d == _T_43[9:0] ? 4'h2 : _GEN_711; // @[Filter.scala 191:62]
  wire [3:0] _GEN_713 = 10'h21e == _T_43[9:0] ? 4'h5 : _GEN_712; // @[Filter.scala 191:62]
  wire [3:0] _GEN_714 = 10'h21f == _T_43[9:0] ? 4'h0 : _GEN_713; // @[Filter.scala 191:62]
  wire [3:0] _GEN_715 = 10'h220 == _T_43[9:0] ? 4'h0 : _GEN_714; // @[Filter.scala 191:62]
  wire [3:0] _GEN_716 = 10'h221 == _T_43[9:0] ? 4'h0 : _GEN_715; // @[Filter.scala 191:62]
  wire [3:0] _GEN_717 = 10'h222 == _T_43[9:0] ? 4'h0 : _GEN_716; // @[Filter.scala 191:62]
  wire [3:0] _GEN_718 = 10'h223 == _T_43[9:0] ? 4'h0 : _GEN_717; // @[Filter.scala 191:62]
  wire [3:0] _GEN_719 = 10'h224 == _T_43[9:0] ? 4'h0 : _GEN_718; // @[Filter.scala 191:62]
  wire [3:0] _GEN_720 = 10'h225 == _T_43[9:0] ? 4'h0 : _GEN_719; // @[Filter.scala 191:62]
  wire [3:0] _GEN_721 = 10'h226 == _T_43[9:0] ? 4'h0 : _GEN_720; // @[Filter.scala 191:62]
  wire [3:0] _GEN_722 = 10'h227 == _T_43[9:0] ? 4'h0 : _GEN_721; // @[Filter.scala 191:62]
  wire [3:0] _GEN_723 = 10'h228 == _T_43[9:0] ? 4'h0 : _GEN_722; // @[Filter.scala 191:62]
  wire [3:0] _GEN_724 = 10'h229 == _T_43[9:0] ? 4'h0 : _GEN_723; // @[Filter.scala 191:62]
  wire [3:0] _GEN_725 = 10'h22a == _T_43[9:0] ? 4'h0 : _GEN_724; // @[Filter.scala 191:62]
  wire [3:0] _GEN_726 = 10'h22b == _T_43[9:0] ? 4'h0 : _GEN_725; // @[Filter.scala 191:62]
  wire [3:0] _GEN_727 = 10'h22c == _T_43[9:0] ? 4'h0 : _GEN_726; // @[Filter.scala 191:62]
  wire [3:0] _GEN_728 = 10'h22d == _T_43[9:0] ? 4'h0 : _GEN_727; // @[Filter.scala 191:62]
  wire [3:0] _GEN_729 = 10'h22e == _T_43[9:0] ? 4'h0 : _GEN_728; // @[Filter.scala 191:62]
  wire [3:0] _GEN_730 = 10'h22f == _T_43[9:0] ? 4'h0 : _GEN_729; // @[Filter.scala 191:62]
  wire [3:0] _GEN_731 = 10'h230 == _T_43[9:0] ? 4'h0 : _GEN_730; // @[Filter.scala 191:62]
  wire [3:0] _GEN_732 = 10'h231 == _T_43[9:0] ? 4'h0 : _GEN_731; // @[Filter.scala 191:62]
  wire [3:0] _GEN_733 = 10'h232 == _T_43[9:0] ? 4'h0 : _GEN_732; // @[Filter.scala 191:62]
  wire [3:0] _GEN_734 = 10'h233 == _T_43[9:0] ? 4'h0 : _GEN_733; // @[Filter.scala 191:62]
  wire [3:0] _GEN_735 = 10'h234 == _T_43[9:0] ? 4'h0 : _GEN_734; // @[Filter.scala 191:62]
  wire [3:0] _GEN_736 = 10'h235 == _T_43[9:0] ? 4'h0 : _GEN_735; // @[Filter.scala 191:62]
  wire [3:0] _GEN_737 = 10'h236 == _T_43[9:0] ? 4'h0 : _GEN_736; // @[Filter.scala 191:62]
  wire [3:0] _GEN_738 = 10'h237 == _T_43[9:0] ? 4'h0 : _GEN_737; // @[Filter.scala 191:62]
  wire [3:0] _GEN_739 = 10'h238 == _T_43[9:0] ? 4'h0 : _GEN_738; // @[Filter.scala 191:62]
  wire [3:0] _GEN_740 = 10'h239 == _T_43[9:0] ? 4'h0 : _GEN_739; // @[Filter.scala 191:62]
  wire [3:0] _GEN_741 = 10'h23a == _T_43[9:0] ? 4'h0 : _GEN_740; // @[Filter.scala 191:62]
  wire [3:0] _GEN_742 = 10'h23b == _T_43[9:0] ? 4'h0 : _GEN_741; // @[Filter.scala 191:62]
  wire [3:0] _GEN_743 = 10'h23c == _T_43[9:0] ? 4'h0 : _GEN_742; // @[Filter.scala 191:62]
  wire [3:0] _GEN_744 = 10'h23d == _T_43[9:0] ? 4'h0 : _GEN_743; // @[Filter.scala 191:62]
  wire [3:0] _GEN_745 = 10'h23e == _T_43[9:0] ? 4'h0 : _GEN_744; // @[Filter.scala 191:62]
  wire [3:0] _GEN_746 = 10'h23f == _T_43[9:0] ? 4'h0 : _GEN_745; // @[Filter.scala 191:62]
  wire [4:0] _GEN_28298 = {{1'd0}, _GEN_746}; // @[Filter.scala 191:62]
  wire [8:0] _T_45 = _GEN_28298 * 5'h14; // @[Filter.scala 191:62]
  wire [3:0] _GEN_750 = 10'h3 == _T_43[9:0] ? 4'ha : 4'h3; // @[Filter.scala 191:102]
  wire [3:0] _GEN_751 = 10'h4 == _T_43[9:0] ? 4'h3 : _GEN_750; // @[Filter.scala 191:102]
  wire [3:0] _GEN_752 = 10'h5 == _T_43[9:0] ? 4'h3 : _GEN_751; // @[Filter.scala 191:102]
  wire [3:0] _GEN_753 = 10'h6 == _T_43[9:0] ? 4'h3 : _GEN_752; // @[Filter.scala 191:102]
  wire [3:0] _GEN_754 = 10'h7 == _T_43[9:0] ? 4'h3 : _GEN_753; // @[Filter.scala 191:102]
  wire [3:0] _GEN_755 = 10'h8 == _T_43[9:0] ? 4'h3 : _GEN_754; // @[Filter.scala 191:102]
  wire [3:0] _GEN_756 = 10'h9 == _T_43[9:0] ? 4'h3 : _GEN_755; // @[Filter.scala 191:102]
  wire [3:0] _GEN_757 = 10'ha == _T_43[9:0] ? 4'h3 : _GEN_756; // @[Filter.scala 191:102]
  wire [3:0] _GEN_758 = 10'hb == _T_43[9:0] ? 4'h3 : _GEN_757; // @[Filter.scala 191:102]
  wire [3:0] _GEN_759 = 10'hc == _T_43[9:0] ? 4'h5 : _GEN_758; // @[Filter.scala 191:102]
  wire [3:0] _GEN_760 = 10'hd == _T_43[9:0] ? 4'h3 : _GEN_759; // @[Filter.scala 191:102]
  wire [3:0] _GEN_761 = 10'he == _T_43[9:0] ? 4'h3 : _GEN_760; // @[Filter.scala 191:102]
  wire [3:0] _GEN_762 = 10'hf == _T_43[9:0] ? 4'h3 : _GEN_761; // @[Filter.scala 191:102]
  wire [3:0] _GEN_763 = 10'h10 == _T_43[9:0] ? 4'h3 : _GEN_762; // @[Filter.scala 191:102]
  wire [3:0] _GEN_764 = 10'h11 == _T_43[9:0] ? 4'h3 : _GEN_763; // @[Filter.scala 191:102]
  wire [3:0] _GEN_765 = 10'h12 == _T_43[9:0] ? 4'h3 : _GEN_764; // @[Filter.scala 191:102]
  wire [3:0] _GEN_766 = 10'h13 == _T_43[9:0] ? 4'h3 : _GEN_765; // @[Filter.scala 191:102]
  wire [3:0] _GEN_767 = 10'h14 == _T_43[9:0] ? 4'h3 : _GEN_766; // @[Filter.scala 191:102]
  wire [3:0] _GEN_768 = 10'h15 == _T_43[9:0] ? 4'h3 : _GEN_767; // @[Filter.scala 191:102]
  wire [3:0] _GEN_769 = 10'h16 == _T_43[9:0] ? 4'h3 : _GEN_768; // @[Filter.scala 191:102]
  wire [3:0] _GEN_770 = 10'h17 == _T_43[9:0] ? 4'h3 : _GEN_769; // @[Filter.scala 191:102]
  wire [3:0] _GEN_771 = 10'h18 == _T_43[9:0] ? 4'h3 : _GEN_770; // @[Filter.scala 191:102]
  wire [3:0] _GEN_772 = 10'h19 == _T_43[9:0] ? 4'h3 : _GEN_771; // @[Filter.scala 191:102]
  wire [3:0] _GEN_773 = 10'h1a == _T_43[9:0] ? 4'h3 : _GEN_772; // @[Filter.scala 191:102]
  wire [3:0] _GEN_774 = 10'h1b == _T_43[9:0] ? 4'h3 : _GEN_773; // @[Filter.scala 191:102]
  wire [3:0] _GEN_775 = 10'h1c == _T_43[9:0] ? 4'h3 : _GEN_774; // @[Filter.scala 191:102]
  wire [3:0] _GEN_776 = 10'h1d == _T_43[9:0] ? 4'h3 : _GEN_775; // @[Filter.scala 191:102]
  wire [3:0] _GEN_777 = 10'h1e == _T_43[9:0] ? 4'h3 : _GEN_776; // @[Filter.scala 191:102]
  wire [3:0] _GEN_778 = 10'h1f == _T_43[9:0] ? 4'h0 : _GEN_777; // @[Filter.scala 191:102]
  wire [3:0] _GEN_779 = 10'h20 == _T_43[9:0] ? 4'h3 : _GEN_778; // @[Filter.scala 191:102]
  wire [3:0] _GEN_780 = 10'h21 == _T_43[9:0] ? 4'h5 : _GEN_779; // @[Filter.scala 191:102]
  wire [3:0] _GEN_781 = 10'h22 == _T_43[9:0] ? 4'h3 : _GEN_780; // @[Filter.scala 191:102]
  wire [3:0] _GEN_782 = 10'h23 == _T_43[9:0] ? 4'ha : _GEN_781; // @[Filter.scala 191:102]
  wire [3:0] _GEN_783 = 10'h24 == _T_43[9:0] ? 4'h3 : _GEN_782; // @[Filter.scala 191:102]
  wire [3:0] _GEN_784 = 10'h25 == _T_43[9:0] ? 4'h3 : _GEN_783; // @[Filter.scala 191:102]
  wire [3:0] _GEN_785 = 10'h26 == _T_43[9:0] ? 4'h3 : _GEN_784; // @[Filter.scala 191:102]
  wire [3:0] _GEN_786 = 10'h27 == _T_43[9:0] ? 4'h1 : _GEN_785; // @[Filter.scala 191:102]
  wire [3:0] _GEN_787 = 10'h28 == _T_43[9:0] ? 4'h1 : _GEN_786; // @[Filter.scala 191:102]
  wire [3:0] _GEN_788 = 10'h29 == _T_43[9:0] ? 4'h3 : _GEN_787; // @[Filter.scala 191:102]
  wire [3:0] _GEN_789 = 10'h2a == _T_43[9:0] ? 4'h3 : _GEN_788; // @[Filter.scala 191:102]
  wire [3:0] _GEN_790 = 10'h2b == _T_43[9:0] ? 4'h3 : _GEN_789; // @[Filter.scala 191:102]
  wire [3:0] _GEN_791 = 10'h2c == _T_43[9:0] ? 4'h3 : _GEN_790; // @[Filter.scala 191:102]
  wire [3:0] _GEN_792 = 10'h2d == _T_43[9:0] ? 4'h3 : _GEN_791; // @[Filter.scala 191:102]
  wire [3:0] _GEN_793 = 10'h2e == _T_43[9:0] ? 4'h3 : _GEN_792; // @[Filter.scala 191:102]
  wire [3:0] _GEN_794 = 10'h2f == _T_43[9:0] ? 4'h3 : _GEN_793; // @[Filter.scala 191:102]
  wire [3:0] _GEN_795 = 10'h30 == _T_43[9:0] ? 4'h3 : _GEN_794; // @[Filter.scala 191:102]
  wire [3:0] _GEN_796 = 10'h31 == _T_43[9:0] ? 4'h5 : _GEN_795; // @[Filter.scala 191:102]
  wire [3:0] _GEN_797 = 10'h32 == _T_43[9:0] ? 4'h3 : _GEN_796; // @[Filter.scala 191:102]
  wire [3:0] _GEN_798 = 10'h33 == _T_43[9:0] ? 4'h3 : _GEN_797; // @[Filter.scala 191:102]
  wire [3:0] _GEN_799 = 10'h34 == _T_43[9:0] ? 4'h3 : _GEN_798; // @[Filter.scala 191:102]
  wire [3:0] _GEN_800 = 10'h35 == _T_43[9:0] ? 4'h3 : _GEN_799; // @[Filter.scala 191:102]
  wire [3:0] _GEN_801 = 10'h36 == _T_43[9:0] ? 4'h3 : _GEN_800; // @[Filter.scala 191:102]
  wire [3:0] _GEN_802 = 10'h37 == _T_43[9:0] ? 4'h1 : _GEN_801; // @[Filter.scala 191:102]
  wire [3:0] _GEN_803 = 10'h38 == _T_43[9:0] ? 4'h1 : _GEN_802; // @[Filter.scala 191:102]
  wire [3:0] _GEN_804 = 10'h39 == _T_43[9:0] ? 4'h3 : _GEN_803; // @[Filter.scala 191:102]
  wire [3:0] _GEN_805 = 10'h3a == _T_43[9:0] ? 4'h3 : _GEN_804; // @[Filter.scala 191:102]
  wire [3:0] _GEN_806 = 10'h3b == _T_43[9:0] ? 4'h5 : _GEN_805; // @[Filter.scala 191:102]
  wire [3:0] _GEN_807 = 10'h3c == _T_43[9:0] ? 4'h3 : _GEN_806; // @[Filter.scala 191:102]
  wire [3:0] _GEN_808 = 10'h3d == _T_43[9:0] ? 4'ha : _GEN_807; // @[Filter.scala 191:102]
  wire [3:0] _GEN_809 = 10'h3e == _T_43[9:0] ? 4'h3 : _GEN_808; // @[Filter.scala 191:102]
  wire [3:0] _GEN_810 = 10'h3f == _T_43[9:0] ? 4'h0 : _GEN_809; // @[Filter.scala 191:102]
  wire [3:0] _GEN_811 = 10'h40 == _T_43[9:0] ? 4'h3 : _GEN_810; // @[Filter.scala 191:102]
  wire [3:0] _GEN_812 = 10'h41 == _T_43[9:0] ? 4'h3 : _GEN_811; // @[Filter.scala 191:102]
  wire [3:0] _GEN_813 = 10'h42 == _T_43[9:0] ? 4'h3 : _GEN_812; // @[Filter.scala 191:102]
  wire [3:0] _GEN_814 = 10'h43 == _T_43[9:0] ? 4'h7 : _GEN_813; // @[Filter.scala 191:102]
  wire [3:0] _GEN_815 = 10'h44 == _T_43[9:0] ? 4'ha : _GEN_814; // @[Filter.scala 191:102]
  wire [3:0] _GEN_816 = 10'h45 == _T_43[9:0] ? 4'h0 : _GEN_815; // @[Filter.scala 191:102]
  wire [3:0] _GEN_817 = 10'h46 == _T_43[9:0] ? 4'h0 : _GEN_816; // @[Filter.scala 191:102]
  wire [3:0] _GEN_818 = 10'h47 == _T_43[9:0] ? 4'h0 : _GEN_817; // @[Filter.scala 191:102]
  wire [3:0] _GEN_819 = 10'h48 == _T_43[9:0] ? 4'h0 : _GEN_818; // @[Filter.scala 191:102]
  wire [3:0] _GEN_820 = 10'h49 == _T_43[9:0] ? 4'h3 : _GEN_819; // @[Filter.scala 191:102]
  wire [3:0] _GEN_821 = 10'h4a == _T_43[9:0] ? 4'h3 : _GEN_820; // @[Filter.scala 191:102]
  wire [3:0] _GEN_822 = 10'h4b == _T_43[9:0] ? 4'h3 : _GEN_821; // @[Filter.scala 191:102]
  wire [3:0] _GEN_823 = 10'h4c == _T_43[9:0] ? 4'h3 : _GEN_822; // @[Filter.scala 191:102]
  wire [3:0] _GEN_824 = 10'h4d == _T_43[9:0] ? 4'h5 : _GEN_823; // @[Filter.scala 191:102]
  wire [3:0] _GEN_825 = 10'h4e == _T_43[9:0] ? 4'h3 : _GEN_824; // @[Filter.scala 191:102]
  wire [3:0] _GEN_826 = 10'h4f == _T_43[9:0] ? 4'h3 : _GEN_825; // @[Filter.scala 191:102]
  wire [3:0] _GEN_827 = 10'h50 == _T_43[9:0] ? 4'h3 : _GEN_826; // @[Filter.scala 191:102]
  wire [3:0] _GEN_828 = 10'h51 == _T_43[9:0] ? 4'h3 : _GEN_827; // @[Filter.scala 191:102]
  wire [3:0] _GEN_829 = 10'h52 == _T_43[9:0] ? 4'h3 : _GEN_828; // @[Filter.scala 191:102]
  wire [3:0] _GEN_830 = 10'h53 == _T_43[9:0] ? 4'h3 : _GEN_829; // @[Filter.scala 191:102]
  wire [3:0] _GEN_831 = 10'h54 == _T_43[9:0] ? 4'h1 : _GEN_830; // @[Filter.scala 191:102]
  wire [3:0] _GEN_832 = 10'h55 == _T_43[9:0] ? 4'h1 : _GEN_831; // @[Filter.scala 191:102]
  wire [3:0] _GEN_833 = 10'h56 == _T_43[9:0] ? 4'h1 : _GEN_832; // @[Filter.scala 191:102]
  wire [3:0] _GEN_834 = 10'h57 == _T_43[9:0] ? 4'h0 : _GEN_833; // @[Filter.scala 191:102]
  wire [3:0] _GEN_835 = 10'h58 == _T_43[9:0] ? 4'h3 : _GEN_834; // @[Filter.scala 191:102]
  wire [3:0] _GEN_836 = 10'h59 == _T_43[9:0] ? 4'h0 : _GEN_835; // @[Filter.scala 191:102]
  wire [3:0] _GEN_837 = 10'h5a == _T_43[9:0] ? 4'h3 : _GEN_836; // @[Filter.scala 191:102]
  wire [3:0] _GEN_838 = 10'h5b == _T_43[9:0] ? 4'h3 : _GEN_837; // @[Filter.scala 191:102]
  wire [3:0] _GEN_839 = 10'h5c == _T_43[9:0] ? 4'h3 : _GEN_838; // @[Filter.scala 191:102]
  wire [3:0] _GEN_840 = 10'h5d == _T_43[9:0] ? 4'ha : _GEN_839; // @[Filter.scala 191:102]
  wire [3:0] _GEN_841 = 10'h5e == _T_43[9:0] ? 4'h3 : _GEN_840; // @[Filter.scala 191:102]
  wire [3:0] _GEN_842 = 10'h5f == _T_43[9:0] ? 4'h0 : _GEN_841; // @[Filter.scala 191:102]
  wire [3:0] _GEN_843 = 10'h60 == _T_43[9:0] ? 4'h3 : _GEN_842; // @[Filter.scala 191:102]
  wire [3:0] _GEN_844 = 10'h61 == _T_43[9:0] ? 4'h3 : _GEN_843; // @[Filter.scala 191:102]
  wire [3:0] _GEN_845 = 10'h62 == _T_43[9:0] ? 4'h3 : _GEN_844; // @[Filter.scala 191:102]
  wire [3:0] _GEN_846 = 10'h63 == _T_43[9:0] ? 4'h3 : _GEN_845; // @[Filter.scala 191:102]
  wire [3:0] _GEN_847 = 10'h64 == _T_43[9:0] ? 4'ha : _GEN_846; // @[Filter.scala 191:102]
  wire [3:0] _GEN_848 = 10'h65 == _T_43[9:0] ? 4'h0 : _GEN_847; // @[Filter.scala 191:102]
  wire [3:0] _GEN_849 = 10'h66 == _T_43[9:0] ? 4'h3 : _GEN_848; // @[Filter.scala 191:102]
  wire [3:0] _GEN_850 = 10'h67 == _T_43[9:0] ? 4'h3 : _GEN_849; // @[Filter.scala 191:102]
  wire [3:0] _GEN_851 = 10'h68 == _T_43[9:0] ? 4'h3 : _GEN_850; // @[Filter.scala 191:102]
  wire [3:0] _GEN_852 = 10'h69 == _T_43[9:0] ? 4'h0 : _GEN_851; // @[Filter.scala 191:102]
  wire [3:0] _GEN_853 = 10'h6a == _T_43[9:0] ? 4'h1 : _GEN_852; // @[Filter.scala 191:102]
  wire [3:0] _GEN_854 = 10'h6b == _T_43[9:0] ? 4'h1 : _GEN_853; // @[Filter.scala 191:102]
  wire [3:0] _GEN_855 = 10'h6c == _T_43[9:0] ? 4'h3 : _GEN_854; // @[Filter.scala 191:102]
  wire [3:0] _GEN_856 = 10'h6d == _T_43[9:0] ? 4'h3 : _GEN_855; // @[Filter.scala 191:102]
  wire [3:0] _GEN_857 = 10'h6e == _T_43[9:0] ? 4'h3 : _GEN_856; // @[Filter.scala 191:102]
  wire [3:0] _GEN_858 = 10'h6f == _T_43[9:0] ? 4'h3 : _GEN_857; // @[Filter.scala 191:102]
  wire [3:0] _GEN_859 = 10'h70 == _T_43[9:0] ? 4'h3 : _GEN_858; // @[Filter.scala 191:102]
  wire [3:0] _GEN_860 = 10'h71 == _T_43[9:0] ? 4'h3 : _GEN_859; // @[Filter.scala 191:102]
  wire [3:0] _GEN_861 = 10'h72 == _T_43[9:0] ? 4'h3 : _GEN_860; // @[Filter.scala 191:102]
  wire [3:0] _GEN_862 = 10'h73 == _T_43[9:0] ? 4'h1 : _GEN_861; // @[Filter.scala 191:102]
  wire [3:0] _GEN_863 = 10'h74 == _T_43[9:0] ? 4'h0 : _GEN_862; // @[Filter.scala 191:102]
  wire [3:0] _GEN_864 = 10'h75 == _T_43[9:0] ? 4'h0 : _GEN_863; // @[Filter.scala 191:102]
  wire [3:0] _GEN_865 = 10'h76 == _T_43[9:0] ? 4'h0 : _GEN_864; // @[Filter.scala 191:102]
  wire [3:0] _GEN_866 = 10'h77 == _T_43[9:0] ? 4'h3 : _GEN_865; // @[Filter.scala 191:102]
  wire [3:0] _GEN_867 = 10'h78 == _T_43[9:0] ? 4'h3 : _GEN_866; // @[Filter.scala 191:102]
  wire [3:0] _GEN_868 = 10'h79 == _T_43[9:0] ? 4'h3 : _GEN_867; // @[Filter.scala 191:102]
  wire [3:0] _GEN_869 = 10'h7a == _T_43[9:0] ? 4'h0 : _GEN_868; // @[Filter.scala 191:102]
  wire [3:0] _GEN_870 = 10'h7b == _T_43[9:0] ? 4'h3 : _GEN_869; // @[Filter.scala 191:102]
  wire [3:0] _GEN_871 = 10'h7c == _T_43[9:0] ? 4'h3 : _GEN_870; // @[Filter.scala 191:102]
  wire [3:0] _GEN_872 = 10'h7d == _T_43[9:0] ? 4'h7 : _GEN_871; // @[Filter.scala 191:102]
  wire [3:0] _GEN_873 = 10'h7e == _T_43[9:0] ? 4'ha : _GEN_872; // @[Filter.scala 191:102]
  wire [3:0] _GEN_874 = 10'h7f == _T_43[9:0] ? 4'h0 : _GEN_873; // @[Filter.scala 191:102]
  wire [3:0] _GEN_875 = 10'h80 == _T_43[9:0] ? 4'h3 : _GEN_874; // @[Filter.scala 191:102]
  wire [3:0] _GEN_876 = 10'h81 == _T_43[9:0] ? 4'h3 : _GEN_875; // @[Filter.scala 191:102]
  wire [3:0] _GEN_877 = 10'h82 == _T_43[9:0] ? 4'h1 : _GEN_876; // @[Filter.scala 191:102]
  wire [3:0] _GEN_878 = 10'h83 == _T_43[9:0] ? 4'h0 : _GEN_877; // @[Filter.scala 191:102]
  wire [3:0] _GEN_879 = 10'h84 == _T_43[9:0] ? 4'h7 : _GEN_878; // @[Filter.scala 191:102]
  wire [3:0] _GEN_880 = 10'h85 == _T_43[9:0] ? 4'h1 : _GEN_879; // @[Filter.scala 191:102]
  wire [3:0] _GEN_881 = 10'h86 == _T_43[9:0] ? 4'h1 : _GEN_880; // @[Filter.scala 191:102]
  wire [3:0] _GEN_882 = 10'h87 == _T_43[9:0] ? 4'h3 : _GEN_881; // @[Filter.scala 191:102]
  wire [3:0] _GEN_883 = 10'h88 == _T_43[9:0] ? 4'h3 : _GEN_882; // @[Filter.scala 191:102]
  wire [3:0] _GEN_884 = 10'h89 == _T_43[9:0] ? 4'h0 : _GEN_883; // @[Filter.scala 191:102]
  wire [3:0] _GEN_885 = 10'h8a == _T_43[9:0] ? 4'h0 : _GEN_884; // @[Filter.scala 191:102]
  wire [3:0] _GEN_886 = 10'h8b == _T_43[9:0] ? 4'h1 : _GEN_885; // @[Filter.scala 191:102]
  wire [3:0] _GEN_887 = 10'h8c == _T_43[9:0] ? 4'h1 : _GEN_886; // @[Filter.scala 191:102]
  wire [3:0] _GEN_888 = 10'h8d == _T_43[9:0] ? 4'h1 : _GEN_887; // @[Filter.scala 191:102]
  wire [3:0] _GEN_889 = 10'h8e == _T_43[9:0] ? 4'h1 : _GEN_888; // @[Filter.scala 191:102]
  wire [3:0] _GEN_890 = 10'h8f == _T_43[9:0] ? 4'h1 : _GEN_889; // @[Filter.scala 191:102]
  wire [3:0] _GEN_891 = 10'h90 == _T_43[9:0] ? 4'h1 : _GEN_890; // @[Filter.scala 191:102]
  wire [3:0] _GEN_892 = 10'h91 == _T_43[9:0] ? 4'h1 : _GEN_891; // @[Filter.scala 191:102]
  wire [3:0] _GEN_893 = 10'h92 == _T_43[9:0] ? 4'h1 : _GEN_892; // @[Filter.scala 191:102]
  wire [3:0] _GEN_894 = 10'h93 == _T_43[9:0] ? 4'h0 : _GEN_893; // @[Filter.scala 191:102]
  wire [3:0] _GEN_895 = 10'h94 == _T_43[9:0] ? 4'h0 : _GEN_894; // @[Filter.scala 191:102]
  wire [3:0] _GEN_896 = 10'h95 == _T_43[9:0] ? 4'h3 : _GEN_895; // @[Filter.scala 191:102]
  wire [3:0] _GEN_897 = 10'h96 == _T_43[9:0] ? 4'h3 : _GEN_896; // @[Filter.scala 191:102]
  wire [3:0] _GEN_898 = 10'h97 == _T_43[9:0] ? 4'h3 : _GEN_897; // @[Filter.scala 191:102]
  wire [3:0] _GEN_899 = 10'h98 == _T_43[9:0] ? 4'h1 : _GEN_898; // @[Filter.scala 191:102]
  wire [3:0] _GEN_900 = 10'h99 == _T_43[9:0] ? 4'h0 : _GEN_899; // @[Filter.scala 191:102]
  wire [3:0] _GEN_901 = 10'h9a == _T_43[9:0] ? 4'h1 : _GEN_900; // @[Filter.scala 191:102]
  wire [3:0] _GEN_902 = 10'h9b == _T_43[9:0] ? 4'h1 : _GEN_901; // @[Filter.scala 191:102]
  wire [3:0] _GEN_903 = 10'h9c == _T_43[9:0] ? 4'h3 : _GEN_902; // @[Filter.scala 191:102]
  wire [3:0] _GEN_904 = 10'h9d == _T_43[9:0] ? 4'h3 : _GEN_903; // @[Filter.scala 191:102]
  wire [3:0] _GEN_905 = 10'h9e == _T_43[9:0] ? 4'ha : _GEN_904; // @[Filter.scala 191:102]
  wire [3:0] _GEN_906 = 10'h9f == _T_43[9:0] ? 4'h0 : _GEN_905; // @[Filter.scala 191:102]
  wire [3:0] _GEN_907 = 10'ha0 == _T_43[9:0] ? 4'h3 : _GEN_906; // @[Filter.scala 191:102]
  wire [3:0] _GEN_908 = 10'ha1 == _T_43[9:0] ? 4'h1 : _GEN_907; // @[Filter.scala 191:102]
  wire [3:0] _GEN_909 = 10'ha2 == _T_43[9:0] ? 4'h0 : _GEN_908; // @[Filter.scala 191:102]
  wire [3:0] _GEN_910 = 10'ha3 == _T_43[9:0] ? 4'ha : _GEN_909; // @[Filter.scala 191:102]
  wire [3:0] _GEN_911 = 10'ha4 == _T_43[9:0] ? 4'h3 : _GEN_910; // @[Filter.scala 191:102]
  wire [3:0] _GEN_912 = 10'ha5 == _T_43[9:0] ? 4'h3 : _GEN_911; // @[Filter.scala 191:102]
  wire [3:0] _GEN_913 = 10'ha6 == _T_43[9:0] ? 4'h3 : _GEN_912; // @[Filter.scala 191:102]
  wire [3:0] _GEN_914 = 10'ha7 == _T_43[9:0] ? 4'h0 : _GEN_913; // @[Filter.scala 191:102]
  wire [3:0] _GEN_915 = 10'ha8 == _T_43[9:0] ? 4'h3 : _GEN_914; // @[Filter.scala 191:102]
  wire [3:0] _GEN_916 = 10'ha9 == _T_43[9:0] ? 4'h1 : _GEN_915; // @[Filter.scala 191:102]
  wire [3:0] _GEN_917 = 10'haa == _T_43[9:0] ? 4'h0 : _GEN_916; // @[Filter.scala 191:102]
  wire [3:0] _GEN_918 = 10'hab == _T_43[9:0] ? 4'h0 : _GEN_917; // @[Filter.scala 191:102]
  wire [3:0] _GEN_919 = 10'hac == _T_43[9:0] ? 4'h0 : _GEN_918; // @[Filter.scala 191:102]
  wire [3:0] _GEN_920 = 10'had == _T_43[9:0] ? 4'h0 : _GEN_919; // @[Filter.scala 191:102]
  wire [3:0] _GEN_921 = 10'hae == _T_43[9:0] ? 4'h0 : _GEN_920; // @[Filter.scala 191:102]
  wire [3:0] _GEN_922 = 10'haf == _T_43[9:0] ? 4'h0 : _GEN_921; // @[Filter.scala 191:102]
  wire [3:0] _GEN_923 = 10'hb0 == _T_43[9:0] ? 4'h0 : _GEN_922; // @[Filter.scala 191:102]
  wire [3:0] _GEN_924 = 10'hb1 == _T_43[9:0] ? 4'h0 : _GEN_923; // @[Filter.scala 191:102]
  wire [3:0] _GEN_925 = 10'hb2 == _T_43[9:0] ? 4'h0 : _GEN_924; // @[Filter.scala 191:102]
  wire [3:0] _GEN_926 = 10'hb3 == _T_43[9:0] ? 4'h0 : _GEN_925; // @[Filter.scala 191:102]
  wire [3:0] _GEN_927 = 10'hb4 == _T_43[9:0] ? 4'h1 : _GEN_926; // @[Filter.scala 191:102]
  wire [3:0] _GEN_928 = 10'hb5 == _T_43[9:0] ? 4'h1 : _GEN_927; // @[Filter.scala 191:102]
  wire [3:0] _GEN_929 = 10'hb6 == _T_43[9:0] ? 4'h3 : _GEN_928; // @[Filter.scala 191:102]
  wire [3:0] _GEN_930 = 10'hb7 == _T_43[9:0] ? 4'h0 : _GEN_929; // @[Filter.scala 191:102]
  wire [3:0] _GEN_931 = 10'hb8 == _T_43[9:0] ? 4'h3 : _GEN_930; // @[Filter.scala 191:102]
  wire [3:0] _GEN_932 = 10'hb9 == _T_43[9:0] ? 4'h3 : _GEN_931; // @[Filter.scala 191:102]
  wire [3:0] _GEN_933 = 10'hba == _T_43[9:0] ? 4'h3 : _GEN_932; // @[Filter.scala 191:102]
  wire [3:0] _GEN_934 = 10'hbb == _T_43[9:0] ? 4'h0 : _GEN_933; // @[Filter.scala 191:102]
  wire [3:0] _GEN_935 = 10'hbc == _T_43[9:0] ? 4'h3 : _GEN_934; // @[Filter.scala 191:102]
  wire [3:0] _GEN_936 = 10'hbd == _T_43[9:0] ? 4'h3 : _GEN_935; // @[Filter.scala 191:102]
  wire [3:0] _GEN_937 = 10'hbe == _T_43[9:0] ? 4'ha : _GEN_936; // @[Filter.scala 191:102]
  wire [3:0] _GEN_938 = 10'hbf == _T_43[9:0] ? 4'h0 : _GEN_937; // @[Filter.scala 191:102]
  wire [3:0] _GEN_939 = 10'hc0 == _T_43[9:0] ? 4'h3 : _GEN_938; // @[Filter.scala 191:102]
  wire [3:0] _GEN_940 = 10'hc1 == _T_43[9:0] ? 4'h3 : _GEN_939; // @[Filter.scala 191:102]
  wire [3:0] _GEN_941 = 10'hc2 == _T_43[9:0] ? 4'ha : _GEN_940; // @[Filter.scala 191:102]
  wire [3:0] _GEN_942 = 10'hc3 == _T_43[9:0] ? 4'h7 : _GEN_941; // @[Filter.scala 191:102]
  wire [3:0] _GEN_943 = 10'hc4 == _T_43[9:0] ? 4'h0 : _GEN_942; // @[Filter.scala 191:102]
  wire [3:0] _GEN_944 = 10'hc5 == _T_43[9:0] ? 4'h0 : _GEN_943; // @[Filter.scala 191:102]
  wire [3:0] _GEN_945 = 10'hc6 == _T_43[9:0] ? 4'h0 : _GEN_944; // @[Filter.scala 191:102]
  wire [3:0] _GEN_946 = 10'hc7 == _T_43[9:0] ? 4'h3 : _GEN_945; // @[Filter.scala 191:102]
  wire [3:0] _GEN_947 = 10'hc8 == _T_43[9:0] ? 4'h1 : _GEN_946; // @[Filter.scala 191:102]
  wire [3:0] _GEN_948 = 10'hc9 == _T_43[9:0] ? 4'h0 : _GEN_947; // @[Filter.scala 191:102]
  wire [3:0] _GEN_949 = 10'hca == _T_43[9:0] ? 4'h0 : _GEN_948; // @[Filter.scala 191:102]
  wire [3:0] _GEN_950 = 10'hcb == _T_43[9:0] ? 4'h0 : _GEN_949; // @[Filter.scala 191:102]
  wire [3:0] _GEN_951 = 10'hcc == _T_43[9:0] ? 4'h0 : _GEN_950; // @[Filter.scala 191:102]
  wire [3:0] _GEN_952 = 10'hcd == _T_43[9:0] ? 4'h0 : _GEN_951; // @[Filter.scala 191:102]
  wire [3:0] _GEN_953 = 10'hce == _T_43[9:0] ? 4'h0 : _GEN_952; // @[Filter.scala 191:102]
  wire [3:0] _GEN_954 = 10'hcf == _T_43[9:0] ? 4'h0 : _GEN_953; // @[Filter.scala 191:102]
  wire [3:0] _GEN_955 = 10'hd0 == _T_43[9:0] ? 4'h0 : _GEN_954; // @[Filter.scala 191:102]
  wire [3:0] _GEN_956 = 10'hd1 == _T_43[9:0] ? 4'h0 : _GEN_955; // @[Filter.scala 191:102]
  wire [3:0] _GEN_957 = 10'hd2 == _T_43[9:0] ? 4'h0 : _GEN_956; // @[Filter.scala 191:102]
  wire [3:0] _GEN_958 = 10'hd3 == _T_43[9:0] ? 4'h0 : _GEN_957; // @[Filter.scala 191:102]
  wire [3:0] _GEN_959 = 10'hd4 == _T_43[9:0] ? 4'h0 : _GEN_958; // @[Filter.scala 191:102]
  wire [3:0] _GEN_960 = 10'hd5 == _T_43[9:0] ? 4'h0 : _GEN_959; // @[Filter.scala 191:102]
  wire [3:0] _GEN_961 = 10'hd6 == _T_43[9:0] ? 4'h1 : _GEN_960; // @[Filter.scala 191:102]
  wire [3:0] _GEN_962 = 10'hd7 == _T_43[9:0] ? 4'h3 : _GEN_961; // @[Filter.scala 191:102]
  wire [3:0] _GEN_963 = 10'hd8 == _T_43[9:0] ? 4'h0 : _GEN_962; // @[Filter.scala 191:102]
  wire [3:0] _GEN_964 = 10'hd9 == _T_43[9:0] ? 4'h3 : _GEN_963; // @[Filter.scala 191:102]
  wire [3:0] _GEN_965 = 10'hda == _T_43[9:0] ? 4'h3 : _GEN_964; // @[Filter.scala 191:102]
  wire [3:0] _GEN_966 = 10'hdb == _T_43[9:0] ? 4'h3 : _GEN_965; // @[Filter.scala 191:102]
  wire [3:0] _GEN_967 = 10'hdc == _T_43[9:0] ? 4'h3 : _GEN_966; // @[Filter.scala 191:102]
  wire [3:0] _GEN_968 = 10'hdd == _T_43[9:0] ? 4'ha : _GEN_967; // @[Filter.scala 191:102]
  wire [3:0] _GEN_969 = 10'hde == _T_43[9:0] ? 4'h7 : _GEN_968; // @[Filter.scala 191:102]
  wire [3:0] _GEN_970 = 10'hdf == _T_43[9:0] ? 4'h0 : _GEN_969; // @[Filter.scala 191:102]
  wire [3:0] _GEN_971 = 10'he0 == _T_43[9:0] ? 4'h3 : _GEN_970; // @[Filter.scala 191:102]
  wire [3:0] _GEN_972 = 10'he1 == _T_43[9:0] ? 4'h3 : _GEN_971; // @[Filter.scala 191:102]
  wire [3:0] _GEN_973 = 10'he2 == _T_43[9:0] ? 4'ha : _GEN_972; // @[Filter.scala 191:102]
  wire [3:0] _GEN_974 = 10'he3 == _T_43[9:0] ? 4'h3 : _GEN_973; // @[Filter.scala 191:102]
  wire [3:0] _GEN_975 = 10'he4 == _T_43[9:0] ? 4'h3 : _GEN_974; // @[Filter.scala 191:102]
  wire [3:0] _GEN_976 = 10'he5 == _T_43[9:0] ? 4'h3 : _GEN_975; // @[Filter.scala 191:102]
  wire [3:0] _GEN_977 = 10'he6 == _T_43[9:0] ? 4'h3 : _GEN_976; // @[Filter.scala 191:102]
  wire [3:0] _GEN_978 = 10'he7 == _T_43[9:0] ? 4'h1 : _GEN_977; // @[Filter.scala 191:102]
  wire [3:0] _GEN_979 = 10'he8 == _T_43[9:0] ? 4'h1 : _GEN_978; // @[Filter.scala 191:102]
  wire [3:0] _GEN_980 = 10'he9 == _T_43[9:0] ? 4'h1 : _GEN_979; // @[Filter.scala 191:102]
  wire [3:0] _GEN_981 = 10'hea == _T_43[9:0] ? 4'h0 : _GEN_980; // @[Filter.scala 191:102]
  wire [3:0] _GEN_982 = 10'heb == _T_43[9:0] ? 4'h0 : _GEN_981; // @[Filter.scala 191:102]
  wire [3:0] _GEN_983 = 10'hec == _T_43[9:0] ? 4'h0 : _GEN_982; // @[Filter.scala 191:102]
  wire [3:0] _GEN_984 = 10'hed == _T_43[9:0] ? 4'h0 : _GEN_983; // @[Filter.scala 191:102]
  wire [3:0] _GEN_985 = 10'hee == _T_43[9:0] ? 4'h0 : _GEN_984; // @[Filter.scala 191:102]
  wire [3:0] _GEN_986 = 10'hef == _T_43[9:0] ? 4'h0 : _GEN_985; // @[Filter.scala 191:102]
  wire [3:0] _GEN_987 = 10'hf0 == _T_43[9:0] ? 4'h0 : _GEN_986; // @[Filter.scala 191:102]
  wire [3:0] _GEN_988 = 10'hf1 == _T_43[9:0] ? 4'h0 : _GEN_987; // @[Filter.scala 191:102]
  wire [3:0] _GEN_989 = 10'hf2 == _T_43[9:0] ? 4'h0 : _GEN_988; // @[Filter.scala 191:102]
  wire [3:0] _GEN_990 = 10'hf3 == _T_43[9:0] ? 4'h0 : _GEN_989; // @[Filter.scala 191:102]
  wire [3:0] _GEN_991 = 10'hf4 == _T_43[9:0] ? 4'h0 : _GEN_990; // @[Filter.scala 191:102]
  wire [3:0] _GEN_992 = 10'hf5 == _T_43[9:0] ? 4'h1 : _GEN_991; // @[Filter.scala 191:102]
  wire [3:0] _GEN_993 = 10'hf6 == _T_43[9:0] ? 4'h0 : _GEN_992; // @[Filter.scala 191:102]
  wire [3:0] _GEN_994 = 10'hf7 == _T_43[9:0] ? 4'h0 : _GEN_993; // @[Filter.scala 191:102]
  wire [3:0] _GEN_995 = 10'hf8 == _T_43[9:0] ? 4'h1 : _GEN_994; // @[Filter.scala 191:102]
  wire [3:0] _GEN_996 = 10'hf9 == _T_43[9:0] ? 4'h0 : _GEN_995; // @[Filter.scala 191:102]
  wire [3:0] _GEN_997 = 10'hfa == _T_43[9:0] ? 4'h3 : _GEN_996; // @[Filter.scala 191:102]
  wire [3:0] _GEN_998 = 10'hfb == _T_43[9:0] ? 4'h3 : _GEN_997; // @[Filter.scala 191:102]
  wire [3:0] _GEN_999 = 10'hfc == _T_43[9:0] ? 4'h3 : _GEN_998; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1000 = 10'hfd == _T_43[9:0] ? 4'ha : _GEN_999; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1001 = 10'hfe == _T_43[9:0] ? 4'h3 : _GEN_1000; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1002 = 10'hff == _T_43[9:0] ? 4'h0 : _GEN_1001; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1003 = 10'h100 == _T_43[9:0] ? 4'h3 : _GEN_1002; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1004 = 10'h101 == _T_43[9:0] ? 4'h0 : _GEN_1003; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1005 = 10'h102 == _T_43[9:0] ? 4'ha : _GEN_1004; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1006 = 10'h103 == _T_43[9:0] ? 4'h3 : _GEN_1005; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1007 = 10'h104 == _T_43[9:0] ? 4'h3 : _GEN_1006; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1008 = 10'h105 == _T_43[9:0] ? 4'h3 : _GEN_1007; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1009 = 10'h106 == _T_43[9:0] ? 4'h3 : _GEN_1008; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1010 = 10'h107 == _T_43[9:0] ? 4'h3 : _GEN_1009; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1011 = 10'h108 == _T_43[9:0] ? 4'h1 : _GEN_1010; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1012 = 10'h109 == _T_43[9:0] ? 4'h0 : _GEN_1011; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1013 = 10'h10a == _T_43[9:0] ? 4'h0 : _GEN_1012; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1014 = 10'h10b == _T_43[9:0] ? 4'h0 : _GEN_1013; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1015 = 10'h10c == _T_43[9:0] ? 4'h0 : _GEN_1014; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1016 = 10'h10d == _T_43[9:0] ? 4'h0 : _GEN_1015; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1017 = 10'h10e == _T_43[9:0] ? 4'h0 : _GEN_1016; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1018 = 10'h10f == _T_43[9:0] ? 4'h0 : _GEN_1017; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1019 = 10'h110 == _T_43[9:0] ? 4'h0 : _GEN_1018; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1020 = 10'h111 == _T_43[9:0] ? 4'h0 : _GEN_1019; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1021 = 10'h112 == _T_43[9:0] ? 4'h0 : _GEN_1020; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1022 = 10'h113 == _T_43[9:0] ? 4'h0 : _GEN_1021; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1023 = 10'h114 == _T_43[9:0] ? 4'h0 : _GEN_1022; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1024 = 10'h115 == _T_43[9:0] ? 4'h0 : _GEN_1023; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1025 = 10'h116 == _T_43[9:0] ? 4'h1 : _GEN_1024; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1026 = 10'h117 == _T_43[9:0] ? 4'h3 : _GEN_1025; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1027 = 10'h118 == _T_43[9:0] ? 4'h3 : _GEN_1026; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1028 = 10'h119 == _T_43[9:0] ? 4'h3 : _GEN_1027; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1029 = 10'h11a == _T_43[9:0] ? 4'h0 : _GEN_1028; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1030 = 10'h11b == _T_43[9:0] ? 4'h3 : _GEN_1029; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1031 = 10'h11c == _T_43[9:0] ? 4'h3 : _GEN_1030; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1032 = 10'h11d == _T_43[9:0] ? 4'h7 : _GEN_1031; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1033 = 10'h11e == _T_43[9:0] ? 4'ha : _GEN_1032; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1034 = 10'h11f == _T_43[9:0] ? 4'h0 : _GEN_1033; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1035 = 10'h120 == _T_43[9:0] ? 4'h3 : _GEN_1034; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1036 = 10'h121 == _T_43[9:0] ? 4'h3 : _GEN_1035; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1037 = 10'h122 == _T_43[9:0] ? 4'ha : _GEN_1036; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1038 = 10'h123 == _T_43[9:0] ? 4'h3 : _GEN_1037; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1039 = 10'h124 == _T_43[9:0] ? 4'h3 : _GEN_1038; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1040 = 10'h125 == _T_43[9:0] ? 4'h3 : _GEN_1039; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1041 = 10'h126 == _T_43[9:0] ? 4'h3 : _GEN_1040; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1042 = 10'h127 == _T_43[9:0] ? 4'h1 : _GEN_1041; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1043 = 10'h128 == _T_43[9:0] ? 4'h0 : _GEN_1042; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1044 = 10'h129 == _T_43[9:0] ? 4'h3 : _GEN_1043; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1045 = 10'h12a == _T_43[9:0] ? 4'h3 : _GEN_1044; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1046 = 10'h12b == _T_43[9:0] ? 4'h0 : _GEN_1045; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1047 = 10'h12c == _T_43[9:0] ? 4'h0 : _GEN_1046; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1048 = 10'h12d == _T_43[9:0] ? 4'h0 : _GEN_1047; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1049 = 10'h12e == _T_43[9:0] ? 4'h0 : _GEN_1048; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1050 = 10'h12f == _T_43[9:0] ? 4'h0 : _GEN_1049; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1051 = 10'h130 == _T_43[9:0] ? 4'h0 : _GEN_1050; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1052 = 10'h131 == _T_43[9:0] ? 4'h0 : _GEN_1051; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1053 = 10'h132 == _T_43[9:0] ? 4'h0 : _GEN_1052; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1054 = 10'h133 == _T_43[9:0] ? 4'h0 : _GEN_1053; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1055 = 10'h134 == _T_43[9:0] ? 4'h3 : _GEN_1054; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1056 = 10'h135 == _T_43[9:0] ? 4'h3 : _GEN_1055; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1057 = 10'h136 == _T_43[9:0] ? 4'h0 : _GEN_1056; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1058 = 10'h137 == _T_43[9:0] ? 4'h1 : _GEN_1057; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1059 = 10'h138 == _T_43[9:0] ? 4'h3 : _GEN_1058; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1060 = 10'h139 == _T_43[9:0] ? 4'h3 : _GEN_1059; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1061 = 10'h13a == _T_43[9:0] ? 4'h3 : _GEN_1060; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1062 = 10'h13b == _T_43[9:0] ? 4'h3 : _GEN_1061; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1063 = 10'h13c == _T_43[9:0] ? 4'h3 : _GEN_1062; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1064 = 10'h13d == _T_43[9:0] ? 4'h3 : _GEN_1063; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1065 = 10'h13e == _T_43[9:0] ? 4'ha : _GEN_1064; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1066 = 10'h13f == _T_43[9:0] ? 4'h0 : _GEN_1065; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1067 = 10'h140 == _T_43[9:0] ? 4'h5 : _GEN_1066; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1068 = 10'h141 == _T_43[9:0] ? 4'h3 : _GEN_1067; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1069 = 10'h142 == _T_43[9:0] ? 4'h7 : _GEN_1068; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1070 = 10'h143 == _T_43[9:0] ? 4'ha : _GEN_1069; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1071 = 10'h144 == _T_43[9:0] ? 4'h3 : _GEN_1070; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1072 = 10'h145 == _T_43[9:0] ? 4'h3 : _GEN_1071; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1073 = 10'h146 == _T_43[9:0] ? 4'h1 : _GEN_1072; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1074 = 10'h147 == _T_43[9:0] ? 4'h0 : _GEN_1073; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1075 = 10'h148 == _T_43[9:0] ? 4'h3 : _GEN_1074; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1076 = 10'h149 == _T_43[9:0] ? 4'h3 : _GEN_1075; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1077 = 10'h14a == _T_43[9:0] ? 4'h3 : _GEN_1076; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1078 = 10'h14b == _T_43[9:0] ? 4'h3 : _GEN_1077; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1079 = 10'h14c == _T_43[9:0] ? 4'h3 : _GEN_1078; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1080 = 10'h14d == _T_43[9:0] ? 4'h3 : _GEN_1079; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1081 = 10'h14e == _T_43[9:0] ? 4'h3 : _GEN_1080; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1082 = 10'h14f == _T_43[9:0] ? 4'h3 : _GEN_1081; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1083 = 10'h150 == _T_43[9:0] ? 4'h3 : _GEN_1082; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1084 = 10'h151 == _T_43[9:0] ? 4'h3 : _GEN_1083; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1085 = 10'h152 == _T_43[9:0] ? 4'h3 : _GEN_1084; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1086 = 10'h153 == _T_43[9:0] ? 4'h3 : _GEN_1085; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1087 = 10'h154 == _T_43[9:0] ? 4'h3 : _GEN_1086; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1088 = 10'h155 == _T_43[9:0] ? 4'h3 : _GEN_1087; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1089 = 10'h156 == _T_43[9:0] ? 4'h3 : _GEN_1088; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1090 = 10'h157 == _T_43[9:0] ? 4'h0 : _GEN_1089; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1091 = 10'h158 == _T_43[9:0] ? 4'h3 : _GEN_1090; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1092 = 10'h159 == _T_43[9:0] ? 4'h3 : _GEN_1091; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1093 = 10'h15a == _T_43[9:0] ? 4'h3 : _GEN_1092; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1094 = 10'h15b == _T_43[9:0] ? 4'h3 : _GEN_1093; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1095 = 10'h15c == _T_43[9:0] ? 4'h3 : _GEN_1094; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1096 = 10'h15d == _T_43[9:0] ? 4'ha : _GEN_1095; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1097 = 10'h15e == _T_43[9:0] ? 4'h7 : _GEN_1096; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1098 = 10'h15f == _T_43[9:0] ? 4'h0 : _GEN_1097; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1099 = 10'h160 == _T_43[9:0] ? 4'h3 : _GEN_1098; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1100 = 10'h161 == _T_43[9:0] ? 4'h3 : _GEN_1099; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1101 = 10'h162 == _T_43[9:0] ? 4'h3 : _GEN_1100; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1102 = 10'h163 == _T_43[9:0] ? 4'h7 : _GEN_1101; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1103 = 10'h164 == _T_43[9:0] ? 4'ha : _GEN_1102; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1104 = 10'h165 == _T_43[9:0] ? 4'h1 : _GEN_1103; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1105 = 10'h166 == _T_43[9:0] ? 4'h0 : _GEN_1104; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1106 = 10'h167 == _T_43[9:0] ? 4'h0 : _GEN_1105; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1107 = 10'h168 == _T_43[9:0] ? 4'hc : _GEN_1106; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1108 = 10'h169 == _T_43[9:0] ? 4'h9 : _GEN_1107; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1109 = 10'h16a == _T_43[9:0] ? 4'hc : _GEN_1108; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1110 = 10'h16b == _T_43[9:0] ? 4'hc : _GEN_1109; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1111 = 10'h16c == _T_43[9:0] ? 4'h3 : _GEN_1110; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1112 = 10'h16d == _T_43[9:0] ? 4'h3 : _GEN_1111; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1113 = 10'h16e == _T_43[9:0] ? 4'h3 : _GEN_1112; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1114 = 10'h16f == _T_43[9:0] ? 4'h3 : _GEN_1113; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1115 = 10'h170 == _T_43[9:0] ? 4'h5 : _GEN_1114; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1116 = 10'h171 == _T_43[9:0] ? 4'h3 : _GEN_1115; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1117 = 10'h172 == _T_43[9:0] ? 4'h3 : _GEN_1116; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1118 = 10'h173 == _T_43[9:0] ? 4'h3 : _GEN_1117; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1119 = 10'h174 == _T_43[9:0] ? 4'h3 : _GEN_1118; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1120 = 10'h175 == _T_43[9:0] ? 4'h3 : _GEN_1119; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1121 = 10'h176 == _T_43[9:0] ? 4'h0 : _GEN_1120; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1122 = 10'h177 == _T_43[9:0] ? 4'h0 : _GEN_1121; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1123 = 10'h178 == _T_43[9:0] ? 4'h1 : _GEN_1122; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1124 = 10'h179 == _T_43[9:0] ? 4'h3 : _GEN_1123; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1125 = 10'h17a == _T_43[9:0] ? 4'h5 : _GEN_1124; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1126 = 10'h17b == _T_43[9:0] ? 4'h3 : _GEN_1125; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1127 = 10'h17c == _T_43[9:0] ? 4'ha : _GEN_1126; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1128 = 10'h17d == _T_43[9:0] ? 4'h7 : _GEN_1127; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1129 = 10'h17e == _T_43[9:0] ? 4'h3 : _GEN_1128; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1130 = 10'h17f == _T_43[9:0] ? 4'h0 : _GEN_1129; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1131 = 10'h180 == _T_43[9:0] ? 4'hc : _GEN_1130; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1132 = 10'h181 == _T_43[9:0] ? 4'hc : _GEN_1131; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1133 = 10'h182 == _T_43[9:0] ? 4'hc : _GEN_1132; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1134 = 10'h183 == _T_43[9:0] ? 4'hc : _GEN_1133; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1135 = 10'h184 == _T_43[9:0] ? 4'ha : _GEN_1134; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1136 = 10'h185 == _T_43[9:0] ? 4'h1 : _GEN_1135; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1137 = 10'h186 == _T_43[9:0] ? 4'hc : _GEN_1136; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1138 = 10'h187 == _T_43[9:0] ? 4'h0 : _GEN_1137; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1139 = 10'h188 == _T_43[9:0] ? 4'hc : _GEN_1138; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1140 = 10'h189 == _T_43[9:0] ? 4'hc : _GEN_1139; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1141 = 10'h18a == _T_43[9:0] ? 4'hc : _GEN_1140; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1142 = 10'h18b == _T_43[9:0] ? 4'hc : _GEN_1141; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1143 = 10'h18c == _T_43[9:0] ? 4'hc : _GEN_1142; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1144 = 10'h18d == _T_43[9:0] ? 4'hc : _GEN_1143; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1145 = 10'h18e == _T_43[9:0] ? 4'hc : _GEN_1144; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1146 = 10'h18f == _T_43[9:0] ? 4'hc : _GEN_1145; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1147 = 10'h190 == _T_43[9:0] ? 4'hc : _GEN_1146; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1148 = 10'h191 == _T_43[9:0] ? 4'hc : _GEN_1147; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1149 = 10'h192 == _T_43[9:0] ? 4'h9 : _GEN_1148; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1150 = 10'h193 == _T_43[9:0] ? 4'hc : _GEN_1149; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1151 = 10'h194 == _T_43[9:0] ? 4'hc : _GEN_1150; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1152 = 10'h195 == _T_43[9:0] ? 4'hc : _GEN_1151; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1153 = 10'h196 == _T_43[9:0] ? 4'h0 : _GEN_1152; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1154 = 10'h197 == _T_43[9:0] ? 4'h3 : _GEN_1153; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1155 = 10'h198 == _T_43[9:0] ? 4'h1 : _GEN_1154; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1156 = 10'h199 == _T_43[9:0] ? 4'h3 : _GEN_1155; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1157 = 10'h19a == _T_43[9:0] ? 4'h3 : _GEN_1156; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1158 = 10'h19b == _T_43[9:0] ? 4'h3 : _GEN_1157; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1159 = 10'h19c == _T_43[9:0] ? 4'ha : _GEN_1158; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1160 = 10'h19d == _T_43[9:0] ? 4'h3 : _GEN_1159; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1161 = 10'h19e == _T_43[9:0] ? 4'h3 : _GEN_1160; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1162 = 10'h19f == _T_43[9:0] ? 4'h0 : _GEN_1161; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1163 = 10'h1a0 == _T_43[9:0] ? 4'hc : _GEN_1162; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1164 = 10'h1a1 == _T_43[9:0] ? 4'hc : _GEN_1163; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1165 = 10'h1a2 == _T_43[9:0] ? 4'h9 : _GEN_1164; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1166 = 10'h1a3 == _T_43[9:0] ? 4'hc : _GEN_1165; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1167 = 10'h1a4 == _T_43[9:0] ? 4'ha : _GEN_1166; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1168 = 10'h1a5 == _T_43[9:0] ? 4'h0 : _GEN_1167; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1169 = 10'h1a6 == _T_43[9:0] ? 4'hc : _GEN_1168; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1170 = 10'h1a7 == _T_43[9:0] ? 4'h0 : _GEN_1169; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1171 = 10'h1a8 == _T_43[9:0] ? 4'hc : _GEN_1170; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1172 = 10'h1a9 == _T_43[9:0] ? 4'hc : _GEN_1171; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1173 = 10'h1aa == _T_43[9:0] ? 4'hc : _GEN_1172; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1174 = 10'h1ab == _T_43[9:0] ? 4'h9 : _GEN_1173; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1175 = 10'h1ac == _T_43[9:0] ? 4'hc : _GEN_1174; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1176 = 10'h1ad == _T_43[9:0] ? 4'hc : _GEN_1175; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1177 = 10'h1ae == _T_43[9:0] ? 4'hc : _GEN_1176; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1178 = 10'h1af == _T_43[9:0] ? 4'hc : _GEN_1177; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1179 = 10'h1b0 == _T_43[9:0] ? 4'hc : _GEN_1178; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1180 = 10'h1b1 == _T_43[9:0] ? 4'hc : _GEN_1179; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1181 = 10'h1b2 == _T_43[9:0] ? 4'hc : _GEN_1180; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1182 = 10'h1b3 == _T_43[9:0] ? 4'hc : _GEN_1181; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1183 = 10'h1b4 == _T_43[9:0] ? 4'hc : _GEN_1182; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1184 = 10'h1b5 == _T_43[9:0] ? 4'hc : _GEN_1183; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1185 = 10'h1b6 == _T_43[9:0] ? 4'h0 : _GEN_1184; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1186 = 10'h1b7 == _T_43[9:0] ? 4'hc : _GEN_1185; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1187 = 10'h1b8 == _T_43[9:0] ? 4'h0 : _GEN_1186; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1188 = 10'h1b9 == _T_43[9:0] ? 4'hc : _GEN_1187; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1189 = 10'h1ba == _T_43[9:0] ? 4'hc : _GEN_1188; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1190 = 10'h1bb == _T_43[9:0] ? 4'hc : _GEN_1189; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1191 = 10'h1bc == _T_43[9:0] ? 4'h7 : _GEN_1190; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1192 = 10'h1bd == _T_43[9:0] ? 4'ha : _GEN_1191; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1193 = 10'h1be == _T_43[9:0] ? 4'hc : _GEN_1192; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1194 = 10'h1bf == _T_43[9:0] ? 4'h0 : _GEN_1193; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1195 = 10'h1c0 == _T_43[9:0] ? 4'hc : _GEN_1194; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1196 = 10'h1c1 == _T_43[9:0] ? 4'hc : _GEN_1195; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1197 = 10'h1c2 == _T_43[9:0] ? 4'hc : _GEN_1196; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1198 = 10'h1c3 == _T_43[9:0] ? 4'h7 : _GEN_1197; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1199 = 10'h1c4 == _T_43[9:0] ? 4'h7 : _GEN_1198; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1200 = 10'h1c5 == _T_43[9:0] ? 4'hc : _GEN_1199; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1201 = 10'h1c6 == _T_43[9:0] ? 4'hc : _GEN_1200; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1202 = 10'h1c7 == _T_43[9:0] ? 4'hc : _GEN_1201; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1203 = 10'h1c8 == _T_43[9:0] ? 4'hc : _GEN_1202; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1204 = 10'h1c9 == _T_43[9:0] ? 4'hc : _GEN_1203; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1205 = 10'h1ca == _T_43[9:0] ? 4'hc : _GEN_1204; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1206 = 10'h1cb == _T_43[9:0] ? 4'hc : _GEN_1205; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1207 = 10'h1cc == _T_43[9:0] ? 4'hc : _GEN_1206; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1208 = 10'h1cd == _T_43[9:0] ? 4'hc : _GEN_1207; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1209 = 10'h1ce == _T_43[9:0] ? 4'hc : _GEN_1208; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1210 = 10'h1cf == _T_43[9:0] ? 4'hc : _GEN_1209; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1211 = 10'h1d0 == _T_43[9:0] ? 4'hc : _GEN_1210; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1212 = 10'h1d1 == _T_43[9:0] ? 4'hc : _GEN_1211; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1213 = 10'h1d2 == _T_43[9:0] ? 4'hc : _GEN_1212; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1214 = 10'h1d3 == _T_43[9:0] ? 4'hc : _GEN_1213; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1215 = 10'h1d4 == _T_43[9:0] ? 4'hc : _GEN_1214; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1216 = 10'h1d5 == _T_43[9:0] ? 4'hc : _GEN_1215; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1217 = 10'h1d6 == _T_43[9:0] ? 4'hc : _GEN_1216; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1218 = 10'h1d7 == _T_43[9:0] ? 4'hc : _GEN_1217; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1219 = 10'h1d8 == _T_43[9:0] ? 4'hc : _GEN_1218; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1220 = 10'h1d9 == _T_43[9:0] ? 4'hc : _GEN_1219; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1221 = 10'h1da == _T_43[9:0] ? 4'hc : _GEN_1220; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1222 = 10'h1db == _T_43[9:0] ? 4'hc : _GEN_1221; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1223 = 10'h1dc == _T_43[9:0] ? 4'hc : _GEN_1222; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1224 = 10'h1dd == _T_43[9:0] ? 4'ha : _GEN_1223; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1225 = 10'h1de == _T_43[9:0] ? 4'hc : _GEN_1224; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1226 = 10'h1df == _T_43[9:0] ? 4'h0 : _GEN_1225; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1227 = 10'h1e0 == _T_43[9:0] ? 4'h9 : _GEN_1226; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1228 = 10'h1e1 == _T_43[9:0] ? 4'hc : _GEN_1227; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1229 = 10'h1e2 == _T_43[9:0] ? 4'h7 : _GEN_1228; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1230 = 10'h1e3 == _T_43[9:0] ? 4'h7 : _GEN_1229; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1231 = 10'h1e4 == _T_43[9:0] ? 4'hc : _GEN_1230; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1232 = 10'h1e5 == _T_43[9:0] ? 4'hc : _GEN_1231; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1233 = 10'h1e6 == _T_43[9:0] ? 4'hc : _GEN_1232; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1234 = 10'h1e7 == _T_43[9:0] ? 4'hc : _GEN_1233; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1235 = 10'h1e8 == _T_43[9:0] ? 4'hc : _GEN_1234; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1236 = 10'h1e9 == _T_43[9:0] ? 4'hc : _GEN_1235; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1237 = 10'h1ea == _T_43[9:0] ? 4'hc : _GEN_1236; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1238 = 10'h1eb == _T_43[9:0] ? 4'hc : _GEN_1237; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1239 = 10'h1ec == _T_43[9:0] ? 4'hc : _GEN_1238; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1240 = 10'h1ed == _T_43[9:0] ? 4'hc : _GEN_1239; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1241 = 10'h1ee == _T_43[9:0] ? 4'hc : _GEN_1240; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1242 = 10'h1ef == _T_43[9:0] ? 4'hc : _GEN_1241; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1243 = 10'h1f0 == _T_43[9:0] ? 4'hc : _GEN_1242; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1244 = 10'h1f1 == _T_43[9:0] ? 4'hc : _GEN_1243; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1245 = 10'h1f2 == _T_43[9:0] ? 4'hc : _GEN_1244; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1246 = 10'h1f3 == _T_43[9:0] ? 4'hc : _GEN_1245; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1247 = 10'h1f4 == _T_43[9:0] ? 4'hc : _GEN_1246; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1248 = 10'h1f5 == _T_43[9:0] ? 4'hc : _GEN_1247; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1249 = 10'h1f6 == _T_43[9:0] ? 4'hc : _GEN_1248; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1250 = 10'h1f7 == _T_43[9:0] ? 4'hc : _GEN_1249; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1251 = 10'h1f8 == _T_43[9:0] ? 4'hc : _GEN_1250; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1252 = 10'h1f9 == _T_43[9:0] ? 4'hc : _GEN_1251; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1253 = 10'h1fa == _T_43[9:0] ? 4'h9 : _GEN_1252; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1254 = 10'h1fb == _T_43[9:0] ? 4'hc : _GEN_1253; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1255 = 10'h1fc == _T_43[9:0] ? 4'hc : _GEN_1254; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1256 = 10'h1fd == _T_43[9:0] ? 4'h7 : _GEN_1255; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1257 = 10'h1fe == _T_43[9:0] ? 4'hc : _GEN_1256; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1258 = 10'h1ff == _T_43[9:0] ? 4'h0 : _GEN_1257; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1259 = 10'h200 == _T_43[9:0] ? 4'hc : _GEN_1258; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1260 = 10'h201 == _T_43[9:0] ? 4'hc : _GEN_1259; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1261 = 10'h202 == _T_43[9:0] ? 4'ha : _GEN_1260; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1262 = 10'h203 == _T_43[9:0] ? 4'hc : _GEN_1261; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1263 = 10'h204 == _T_43[9:0] ? 4'hc : _GEN_1262; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1264 = 10'h205 == _T_43[9:0] ? 4'hc : _GEN_1263; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1265 = 10'h206 == _T_43[9:0] ? 4'hc : _GEN_1264; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1266 = 10'h207 == _T_43[9:0] ? 4'hc : _GEN_1265; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1267 = 10'h208 == _T_43[9:0] ? 4'hc : _GEN_1266; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1268 = 10'h209 == _T_43[9:0] ? 4'hc : _GEN_1267; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1269 = 10'h20a == _T_43[9:0] ? 4'hc : _GEN_1268; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1270 = 10'h20b == _T_43[9:0] ? 4'hc : _GEN_1269; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1271 = 10'h20c == _T_43[9:0] ? 4'hc : _GEN_1270; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1272 = 10'h20d == _T_43[9:0] ? 4'hc : _GEN_1271; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1273 = 10'h20e == _T_43[9:0] ? 4'hc : _GEN_1272; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1274 = 10'h20f == _T_43[9:0] ? 4'hc : _GEN_1273; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1275 = 10'h210 == _T_43[9:0] ? 4'hc : _GEN_1274; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1276 = 10'h211 == _T_43[9:0] ? 4'hc : _GEN_1275; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1277 = 10'h212 == _T_43[9:0] ? 4'hc : _GEN_1276; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1278 = 10'h213 == _T_43[9:0] ? 4'hc : _GEN_1277; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1279 = 10'h214 == _T_43[9:0] ? 4'hc : _GEN_1278; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1280 = 10'h215 == _T_43[9:0] ? 4'hc : _GEN_1279; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1281 = 10'h216 == _T_43[9:0] ? 4'hc : _GEN_1280; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1282 = 10'h217 == _T_43[9:0] ? 4'hc : _GEN_1281; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1283 = 10'h218 == _T_43[9:0] ? 4'hc : _GEN_1282; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1284 = 10'h219 == _T_43[9:0] ? 4'hc : _GEN_1283; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1285 = 10'h21a == _T_43[9:0] ? 4'hc : _GEN_1284; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1286 = 10'h21b == _T_43[9:0] ? 4'hc : _GEN_1285; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1287 = 10'h21c == _T_43[9:0] ? 4'ha : _GEN_1286; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1288 = 10'h21d == _T_43[9:0] ? 4'h7 : _GEN_1287; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1289 = 10'h21e == _T_43[9:0] ? 4'hc : _GEN_1288; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1290 = 10'h21f == _T_43[9:0] ? 4'h0 : _GEN_1289; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1291 = 10'h220 == _T_43[9:0] ? 4'h0 : _GEN_1290; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1292 = 10'h221 == _T_43[9:0] ? 4'h0 : _GEN_1291; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1293 = 10'h222 == _T_43[9:0] ? 4'h0 : _GEN_1292; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1294 = 10'h223 == _T_43[9:0] ? 4'h0 : _GEN_1293; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1295 = 10'h224 == _T_43[9:0] ? 4'h0 : _GEN_1294; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1296 = 10'h225 == _T_43[9:0] ? 4'h0 : _GEN_1295; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1297 = 10'h226 == _T_43[9:0] ? 4'h0 : _GEN_1296; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1298 = 10'h227 == _T_43[9:0] ? 4'h0 : _GEN_1297; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1299 = 10'h228 == _T_43[9:0] ? 4'h0 : _GEN_1298; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1300 = 10'h229 == _T_43[9:0] ? 4'h0 : _GEN_1299; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1301 = 10'h22a == _T_43[9:0] ? 4'h0 : _GEN_1300; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1302 = 10'h22b == _T_43[9:0] ? 4'h0 : _GEN_1301; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1303 = 10'h22c == _T_43[9:0] ? 4'h0 : _GEN_1302; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1304 = 10'h22d == _T_43[9:0] ? 4'h0 : _GEN_1303; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1305 = 10'h22e == _T_43[9:0] ? 4'h0 : _GEN_1304; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1306 = 10'h22f == _T_43[9:0] ? 4'h0 : _GEN_1305; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1307 = 10'h230 == _T_43[9:0] ? 4'h0 : _GEN_1306; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1308 = 10'h231 == _T_43[9:0] ? 4'h0 : _GEN_1307; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1309 = 10'h232 == _T_43[9:0] ? 4'h0 : _GEN_1308; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1310 = 10'h233 == _T_43[9:0] ? 4'h0 : _GEN_1309; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1311 = 10'h234 == _T_43[9:0] ? 4'h0 : _GEN_1310; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1312 = 10'h235 == _T_43[9:0] ? 4'h0 : _GEN_1311; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1313 = 10'h236 == _T_43[9:0] ? 4'h0 : _GEN_1312; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1314 = 10'h237 == _T_43[9:0] ? 4'h0 : _GEN_1313; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1315 = 10'h238 == _T_43[9:0] ? 4'h0 : _GEN_1314; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1316 = 10'h239 == _T_43[9:0] ? 4'h0 : _GEN_1315; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1317 = 10'h23a == _T_43[9:0] ? 4'h0 : _GEN_1316; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1318 = 10'h23b == _T_43[9:0] ? 4'h0 : _GEN_1317; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1319 = 10'h23c == _T_43[9:0] ? 4'h0 : _GEN_1318; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1320 = 10'h23d == _T_43[9:0] ? 4'h0 : _GEN_1319; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1321 = 10'h23e == _T_43[9:0] ? 4'h0 : _GEN_1320; // @[Filter.scala 191:102]
  wire [3:0] _GEN_1322 = 10'h23f == _T_43[9:0] ? 4'h0 : _GEN_1321; // @[Filter.scala 191:102]
  wire [6:0] _GEN_28300 = {{3'd0}, _GEN_1322}; // @[Filter.scala 191:102]
  wire [10:0] _T_50 = _GEN_28300 * 7'h46; // @[Filter.scala 191:102]
  wire [10:0] _GEN_28301 = {{2'd0}, _T_45}; // @[Filter.scala 191:69]
  wire [10:0] _T_52 = _GEN_28301 + _T_50; // @[Filter.scala 191:69]
  wire [3:0] _GEN_1354 = 10'h1f == _T_43[9:0] ? 4'h0 : 4'h3; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1355 = 10'h20 == _T_43[9:0] ? 4'h3 : _GEN_1354; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1356 = 10'h21 == _T_43[9:0] ? 4'h3 : _GEN_1355; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1357 = 10'h22 == _T_43[9:0] ? 4'h3 : _GEN_1356; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1358 = 10'h23 == _T_43[9:0] ? 4'h3 : _GEN_1357; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1359 = 10'h24 == _T_43[9:0] ? 4'h3 : _GEN_1358; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1360 = 10'h25 == _T_43[9:0] ? 4'h3 : _GEN_1359; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1361 = 10'h26 == _T_43[9:0] ? 4'h3 : _GEN_1360; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1362 = 10'h27 == _T_43[9:0] ? 4'h9 : _GEN_1361; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1363 = 10'h28 == _T_43[9:0] ? 4'h9 : _GEN_1362; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1364 = 10'h29 == _T_43[9:0] ? 4'h3 : _GEN_1363; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1365 = 10'h2a == _T_43[9:0] ? 4'h3 : _GEN_1364; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1366 = 10'h2b == _T_43[9:0] ? 4'h3 : _GEN_1365; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1367 = 10'h2c == _T_43[9:0] ? 4'h3 : _GEN_1366; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1368 = 10'h2d == _T_43[9:0] ? 4'h3 : _GEN_1367; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1369 = 10'h2e == _T_43[9:0] ? 4'h3 : _GEN_1368; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1370 = 10'h2f == _T_43[9:0] ? 4'h3 : _GEN_1369; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1371 = 10'h30 == _T_43[9:0] ? 4'h3 : _GEN_1370; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1372 = 10'h31 == _T_43[9:0] ? 4'h3 : _GEN_1371; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1373 = 10'h32 == _T_43[9:0] ? 4'h3 : _GEN_1372; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1374 = 10'h33 == _T_43[9:0] ? 4'h3 : _GEN_1373; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1375 = 10'h34 == _T_43[9:0] ? 4'h3 : _GEN_1374; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1376 = 10'h35 == _T_43[9:0] ? 4'h3 : _GEN_1375; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1377 = 10'h36 == _T_43[9:0] ? 4'h3 : _GEN_1376; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1378 = 10'h37 == _T_43[9:0] ? 4'h9 : _GEN_1377; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1379 = 10'h38 == _T_43[9:0] ? 4'h9 : _GEN_1378; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1380 = 10'h39 == _T_43[9:0] ? 4'h3 : _GEN_1379; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1381 = 10'h3a == _T_43[9:0] ? 4'h3 : _GEN_1380; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1382 = 10'h3b == _T_43[9:0] ? 4'h3 : _GEN_1381; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1383 = 10'h3c == _T_43[9:0] ? 4'h3 : _GEN_1382; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1384 = 10'h3d == _T_43[9:0] ? 4'h3 : _GEN_1383; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1385 = 10'h3e == _T_43[9:0] ? 4'h3 : _GEN_1384; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1386 = 10'h3f == _T_43[9:0] ? 4'h0 : _GEN_1385; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1387 = 10'h40 == _T_43[9:0] ? 4'h3 : _GEN_1386; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1388 = 10'h41 == _T_43[9:0] ? 4'h3 : _GEN_1387; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1389 = 10'h42 == _T_43[9:0] ? 4'h3 : _GEN_1388; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1390 = 10'h43 == _T_43[9:0] ? 4'h2 : _GEN_1389; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1391 = 10'h44 == _T_43[9:0] ? 4'h3 : _GEN_1390; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1392 = 10'h45 == _T_43[9:0] ? 4'hf : _GEN_1391; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1393 = 10'h46 == _T_43[9:0] ? 4'hf : _GEN_1392; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1394 = 10'h47 == _T_43[9:0] ? 4'hf : _GEN_1393; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1395 = 10'h48 == _T_43[9:0] ? 4'hf : _GEN_1394; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1396 = 10'h49 == _T_43[9:0] ? 4'h3 : _GEN_1395; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1397 = 10'h4a == _T_43[9:0] ? 4'h3 : _GEN_1396; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1398 = 10'h4b == _T_43[9:0] ? 4'h3 : _GEN_1397; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1399 = 10'h4c == _T_43[9:0] ? 4'h3 : _GEN_1398; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1400 = 10'h4d == _T_43[9:0] ? 4'h3 : _GEN_1399; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1401 = 10'h4e == _T_43[9:0] ? 4'h3 : _GEN_1400; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1402 = 10'h4f == _T_43[9:0] ? 4'h3 : _GEN_1401; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1403 = 10'h50 == _T_43[9:0] ? 4'h3 : _GEN_1402; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1404 = 10'h51 == _T_43[9:0] ? 4'h3 : _GEN_1403; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1405 = 10'h52 == _T_43[9:0] ? 4'h3 : _GEN_1404; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1406 = 10'h53 == _T_43[9:0] ? 4'h3 : _GEN_1405; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1407 = 10'h54 == _T_43[9:0] ? 4'h9 : _GEN_1406; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1408 = 10'h55 == _T_43[9:0] ? 4'h9 : _GEN_1407; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1409 = 10'h56 == _T_43[9:0] ? 4'h9 : _GEN_1408; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1410 = 10'h57 == _T_43[9:0] ? 4'hf : _GEN_1409; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1411 = 10'h58 == _T_43[9:0] ? 4'h3 : _GEN_1410; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1412 = 10'h59 == _T_43[9:0] ? 4'hf : _GEN_1411; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1413 = 10'h5a == _T_43[9:0] ? 4'h3 : _GEN_1412; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1414 = 10'h5b == _T_43[9:0] ? 4'h3 : _GEN_1413; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1415 = 10'h5c == _T_43[9:0] ? 4'h3 : _GEN_1414; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1416 = 10'h5d == _T_43[9:0] ? 4'h3 : _GEN_1415; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1417 = 10'h5e == _T_43[9:0] ? 4'h3 : _GEN_1416; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1418 = 10'h5f == _T_43[9:0] ? 4'h0 : _GEN_1417; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1419 = 10'h60 == _T_43[9:0] ? 4'h3 : _GEN_1418; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1420 = 10'h61 == _T_43[9:0] ? 4'h3 : _GEN_1419; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1421 = 10'h62 == _T_43[9:0] ? 4'h3 : _GEN_1420; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1422 = 10'h63 == _T_43[9:0] ? 4'h3 : _GEN_1421; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1423 = 10'h64 == _T_43[9:0] ? 4'h3 : _GEN_1422; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1424 = 10'h65 == _T_43[9:0] ? 4'hf : _GEN_1423; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1425 = 10'h66 == _T_43[9:0] ? 4'h3 : _GEN_1424; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1426 = 10'h67 == _T_43[9:0] ? 4'h3 : _GEN_1425; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1427 = 10'h68 == _T_43[9:0] ? 4'h3 : _GEN_1426; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1428 = 10'h69 == _T_43[9:0] ? 4'hf : _GEN_1427; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1429 = 10'h6a == _T_43[9:0] ? 4'h9 : _GEN_1428; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1430 = 10'h6b == _T_43[9:0] ? 4'h9 : _GEN_1429; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1431 = 10'h6c == _T_43[9:0] ? 4'h3 : _GEN_1430; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1432 = 10'h6d == _T_43[9:0] ? 4'h3 : _GEN_1431; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1433 = 10'h6e == _T_43[9:0] ? 4'h3 : _GEN_1432; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1434 = 10'h6f == _T_43[9:0] ? 4'h3 : _GEN_1433; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1435 = 10'h70 == _T_43[9:0] ? 4'h3 : _GEN_1434; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1436 = 10'h71 == _T_43[9:0] ? 4'h3 : _GEN_1435; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1437 = 10'h72 == _T_43[9:0] ? 4'h3 : _GEN_1436; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1438 = 10'h73 == _T_43[9:0] ? 4'h9 : _GEN_1437; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1439 = 10'h74 == _T_43[9:0] ? 4'hf : _GEN_1438; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1440 = 10'h75 == _T_43[9:0] ? 4'hf : _GEN_1439; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1441 = 10'h76 == _T_43[9:0] ? 4'hf : _GEN_1440; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1442 = 10'h77 == _T_43[9:0] ? 4'h3 : _GEN_1441; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1443 = 10'h78 == _T_43[9:0] ? 4'h3 : _GEN_1442; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1444 = 10'h79 == _T_43[9:0] ? 4'h3 : _GEN_1443; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1445 = 10'h7a == _T_43[9:0] ? 4'hf : _GEN_1444; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1446 = 10'h7b == _T_43[9:0] ? 4'h3 : _GEN_1445; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1447 = 10'h7c == _T_43[9:0] ? 4'h3 : _GEN_1446; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1448 = 10'h7d == _T_43[9:0] ? 4'h2 : _GEN_1447; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1449 = 10'h7e == _T_43[9:0] ? 4'h3 : _GEN_1448; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1450 = 10'h7f == _T_43[9:0] ? 4'h0 : _GEN_1449; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1451 = 10'h80 == _T_43[9:0] ? 4'h3 : _GEN_1450; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1452 = 10'h81 == _T_43[9:0] ? 4'h3 : _GEN_1451; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1453 = 10'h82 == _T_43[9:0] ? 4'h9 : _GEN_1452; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1454 = 10'h83 == _T_43[9:0] ? 4'hf : _GEN_1453; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1455 = 10'h84 == _T_43[9:0] ? 4'h2 : _GEN_1454; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1456 = 10'h85 == _T_43[9:0] ? 4'h9 : _GEN_1455; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1457 = 10'h86 == _T_43[9:0] ? 4'h9 : _GEN_1456; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1458 = 10'h87 == _T_43[9:0] ? 4'h3 : _GEN_1457; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1459 = 10'h88 == _T_43[9:0] ? 4'h3 : _GEN_1458; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1460 = 10'h89 == _T_43[9:0] ? 4'hf : _GEN_1459; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1461 = 10'h8a == _T_43[9:0] ? 4'hf : _GEN_1460; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1462 = 10'h8b == _T_43[9:0] ? 4'h9 : _GEN_1461; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1463 = 10'h8c == _T_43[9:0] ? 4'h9 : _GEN_1462; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1464 = 10'h8d == _T_43[9:0] ? 4'h9 : _GEN_1463; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1465 = 10'h8e == _T_43[9:0] ? 4'h9 : _GEN_1464; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1466 = 10'h8f == _T_43[9:0] ? 4'h9 : _GEN_1465; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1467 = 10'h90 == _T_43[9:0] ? 4'h9 : _GEN_1466; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1468 = 10'h91 == _T_43[9:0] ? 4'h9 : _GEN_1467; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1469 = 10'h92 == _T_43[9:0] ? 4'h9 : _GEN_1468; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1470 = 10'h93 == _T_43[9:0] ? 4'hf : _GEN_1469; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1471 = 10'h94 == _T_43[9:0] ? 4'hf : _GEN_1470; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1472 = 10'h95 == _T_43[9:0] ? 4'h3 : _GEN_1471; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1473 = 10'h96 == _T_43[9:0] ? 4'h3 : _GEN_1472; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1474 = 10'h97 == _T_43[9:0] ? 4'h3 : _GEN_1473; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1475 = 10'h98 == _T_43[9:0] ? 4'h9 : _GEN_1474; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1476 = 10'h99 == _T_43[9:0] ? 4'hf : _GEN_1475; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1477 = 10'h9a == _T_43[9:0] ? 4'h9 : _GEN_1476; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1478 = 10'h9b == _T_43[9:0] ? 4'h9 : _GEN_1477; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1479 = 10'h9c == _T_43[9:0] ? 4'h3 : _GEN_1478; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1480 = 10'h9d == _T_43[9:0] ? 4'h3 : _GEN_1479; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1481 = 10'h9e == _T_43[9:0] ? 4'h3 : _GEN_1480; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1482 = 10'h9f == _T_43[9:0] ? 4'h0 : _GEN_1481; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1483 = 10'ha0 == _T_43[9:0] ? 4'h3 : _GEN_1482; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1484 = 10'ha1 == _T_43[9:0] ? 4'h9 : _GEN_1483; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1485 = 10'ha2 == _T_43[9:0] ? 4'hf : _GEN_1484; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1486 = 10'ha3 == _T_43[9:0] ? 4'h3 : _GEN_1485; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1487 = 10'ha4 == _T_43[9:0] ? 4'h3 : _GEN_1486; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1488 = 10'ha5 == _T_43[9:0] ? 4'h3 : _GEN_1487; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1489 = 10'ha6 == _T_43[9:0] ? 4'h3 : _GEN_1488; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1490 = 10'ha7 == _T_43[9:0] ? 4'hf : _GEN_1489; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1491 = 10'ha8 == _T_43[9:0] ? 4'h3 : _GEN_1490; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1492 = 10'ha9 == _T_43[9:0] ? 4'h9 : _GEN_1491; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1493 = 10'haa == _T_43[9:0] ? 4'hf : _GEN_1492; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1494 = 10'hab == _T_43[9:0] ? 4'hf : _GEN_1493; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1495 = 10'hac == _T_43[9:0] ? 4'hf : _GEN_1494; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1496 = 10'had == _T_43[9:0] ? 4'hf : _GEN_1495; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1497 = 10'hae == _T_43[9:0] ? 4'hf : _GEN_1496; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1498 = 10'haf == _T_43[9:0] ? 4'hf : _GEN_1497; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1499 = 10'hb0 == _T_43[9:0] ? 4'hf : _GEN_1498; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1500 = 10'hb1 == _T_43[9:0] ? 4'hf : _GEN_1499; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1501 = 10'hb2 == _T_43[9:0] ? 4'hf : _GEN_1500; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1502 = 10'hb3 == _T_43[9:0] ? 4'hf : _GEN_1501; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1503 = 10'hb4 == _T_43[9:0] ? 4'h9 : _GEN_1502; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1504 = 10'hb5 == _T_43[9:0] ? 4'h9 : _GEN_1503; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1505 = 10'hb6 == _T_43[9:0] ? 4'h3 : _GEN_1504; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1506 = 10'hb7 == _T_43[9:0] ? 4'hf : _GEN_1505; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1507 = 10'hb8 == _T_43[9:0] ? 4'h3 : _GEN_1506; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1508 = 10'hb9 == _T_43[9:0] ? 4'h3 : _GEN_1507; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1509 = 10'hba == _T_43[9:0] ? 4'h3 : _GEN_1508; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1510 = 10'hbb == _T_43[9:0] ? 4'hf : _GEN_1509; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1511 = 10'hbc == _T_43[9:0] ? 4'h3 : _GEN_1510; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1512 = 10'hbd == _T_43[9:0] ? 4'h3 : _GEN_1511; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1513 = 10'hbe == _T_43[9:0] ? 4'h3 : _GEN_1512; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1514 = 10'hbf == _T_43[9:0] ? 4'h0 : _GEN_1513; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1515 = 10'hc0 == _T_43[9:0] ? 4'h3 : _GEN_1514; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1516 = 10'hc1 == _T_43[9:0] ? 4'h3 : _GEN_1515; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1517 = 10'hc2 == _T_43[9:0] ? 4'h3 : _GEN_1516; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1518 = 10'hc3 == _T_43[9:0] ? 4'h2 : _GEN_1517; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1519 = 10'hc4 == _T_43[9:0] ? 4'hf : _GEN_1518; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1520 = 10'hc5 == _T_43[9:0] ? 4'hf : _GEN_1519; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1521 = 10'hc6 == _T_43[9:0] ? 4'hf : _GEN_1520; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1522 = 10'hc7 == _T_43[9:0] ? 4'h3 : _GEN_1521; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1523 = 10'hc8 == _T_43[9:0] ? 4'h9 : _GEN_1522; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1524 = 10'hc9 == _T_43[9:0] ? 4'hf : _GEN_1523; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1525 = 10'hca == _T_43[9:0] ? 4'hf : _GEN_1524; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1526 = 10'hcb == _T_43[9:0] ? 4'hf : _GEN_1525; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1527 = 10'hcc == _T_43[9:0] ? 4'hf : _GEN_1526; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1528 = 10'hcd == _T_43[9:0] ? 4'hf : _GEN_1527; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1529 = 10'hce == _T_43[9:0] ? 4'hf : _GEN_1528; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1530 = 10'hcf == _T_43[9:0] ? 4'hf : _GEN_1529; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1531 = 10'hd0 == _T_43[9:0] ? 4'hf : _GEN_1530; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1532 = 10'hd1 == _T_43[9:0] ? 4'hf : _GEN_1531; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1533 = 10'hd2 == _T_43[9:0] ? 4'hf : _GEN_1532; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1534 = 10'hd3 == _T_43[9:0] ? 4'hf : _GEN_1533; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1535 = 10'hd4 == _T_43[9:0] ? 4'hf : _GEN_1534; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1536 = 10'hd5 == _T_43[9:0] ? 4'hf : _GEN_1535; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1537 = 10'hd6 == _T_43[9:0] ? 4'h9 : _GEN_1536; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1538 = 10'hd7 == _T_43[9:0] ? 4'h3 : _GEN_1537; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1539 = 10'hd8 == _T_43[9:0] ? 4'hf : _GEN_1538; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1540 = 10'hd9 == _T_43[9:0] ? 4'h3 : _GEN_1539; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1541 = 10'hda == _T_43[9:0] ? 4'h3 : _GEN_1540; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1542 = 10'hdb == _T_43[9:0] ? 4'h3 : _GEN_1541; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1543 = 10'hdc == _T_43[9:0] ? 4'h3 : _GEN_1542; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1544 = 10'hdd == _T_43[9:0] ? 4'h3 : _GEN_1543; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1545 = 10'hde == _T_43[9:0] ? 4'h2 : _GEN_1544; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1546 = 10'hdf == _T_43[9:0] ? 4'h0 : _GEN_1545; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1547 = 10'he0 == _T_43[9:0] ? 4'h3 : _GEN_1546; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1548 = 10'he1 == _T_43[9:0] ? 4'h3 : _GEN_1547; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1549 = 10'he2 == _T_43[9:0] ? 4'h3 : _GEN_1548; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1550 = 10'he3 == _T_43[9:0] ? 4'h3 : _GEN_1549; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1551 = 10'he4 == _T_43[9:0] ? 4'h3 : _GEN_1550; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1552 = 10'he5 == _T_43[9:0] ? 4'h3 : _GEN_1551; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1553 = 10'he6 == _T_43[9:0] ? 4'h3 : _GEN_1552; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1554 = 10'he7 == _T_43[9:0] ? 4'h9 : _GEN_1553; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1555 = 10'he8 == _T_43[9:0] ? 4'h9 : _GEN_1554; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1556 = 10'he9 == _T_43[9:0] ? 4'h9 : _GEN_1555; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1557 = 10'hea == _T_43[9:0] ? 4'hf : _GEN_1556; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1558 = 10'heb == _T_43[9:0] ? 4'hf : _GEN_1557; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1559 = 10'hec == _T_43[9:0] ? 4'hf : _GEN_1558; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1560 = 10'hed == _T_43[9:0] ? 4'hf : _GEN_1559; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1561 = 10'hee == _T_43[9:0] ? 4'hf : _GEN_1560; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1562 = 10'hef == _T_43[9:0] ? 4'hf : _GEN_1561; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1563 = 10'hf0 == _T_43[9:0] ? 4'hf : _GEN_1562; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1564 = 10'hf1 == _T_43[9:0] ? 4'hf : _GEN_1563; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1565 = 10'hf2 == _T_43[9:0] ? 4'hf : _GEN_1564; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1566 = 10'hf3 == _T_43[9:0] ? 4'hf : _GEN_1565; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1567 = 10'hf4 == _T_43[9:0] ? 4'hf : _GEN_1566; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1568 = 10'hf5 == _T_43[9:0] ? 4'h9 : _GEN_1567; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1569 = 10'hf6 == _T_43[9:0] ? 4'hf : _GEN_1568; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1570 = 10'hf7 == _T_43[9:0] ? 4'hf : _GEN_1569; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1571 = 10'hf8 == _T_43[9:0] ? 4'h9 : _GEN_1570; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1572 = 10'hf9 == _T_43[9:0] ? 4'hf : _GEN_1571; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1573 = 10'hfa == _T_43[9:0] ? 4'h3 : _GEN_1572; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1574 = 10'hfb == _T_43[9:0] ? 4'h3 : _GEN_1573; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1575 = 10'hfc == _T_43[9:0] ? 4'h3 : _GEN_1574; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1576 = 10'hfd == _T_43[9:0] ? 4'h3 : _GEN_1575; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1577 = 10'hfe == _T_43[9:0] ? 4'h3 : _GEN_1576; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1578 = 10'hff == _T_43[9:0] ? 4'h0 : _GEN_1577; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1579 = 10'h100 == _T_43[9:0] ? 4'h3 : _GEN_1578; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1580 = 10'h101 == _T_43[9:0] ? 4'hf : _GEN_1579; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1581 = 10'h102 == _T_43[9:0] ? 4'h3 : _GEN_1580; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1582 = 10'h103 == _T_43[9:0] ? 4'h3 : _GEN_1581; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1583 = 10'h104 == _T_43[9:0] ? 4'h3 : _GEN_1582; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1584 = 10'h105 == _T_43[9:0] ? 4'h3 : _GEN_1583; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1585 = 10'h106 == _T_43[9:0] ? 4'h3 : _GEN_1584; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1586 = 10'h107 == _T_43[9:0] ? 4'h3 : _GEN_1585; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1587 = 10'h108 == _T_43[9:0] ? 4'h9 : _GEN_1586; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1588 = 10'h109 == _T_43[9:0] ? 4'hf : _GEN_1587; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1589 = 10'h10a == _T_43[9:0] ? 4'hf : _GEN_1588; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1590 = 10'h10b == _T_43[9:0] ? 4'hf : _GEN_1589; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1591 = 10'h10c == _T_43[9:0] ? 4'hf : _GEN_1590; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1592 = 10'h10d == _T_43[9:0] ? 4'h0 : _GEN_1591; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1593 = 10'h10e == _T_43[9:0] ? 4'hf : _GEN_1592; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1594 = 10'h10f == _T_43[9:0] ? 4'hf : _GEN_1593; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1595 = 10'h110 == _T_43[9:0] ? 4'hf : _GEN_1594; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1596 = 10'h111 == _T_43[9:0] ? 4'h0 : _GEN_1595; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1597 = 10'h112 == _T_43[9:0] ? 4'hf : _GEN_1596; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1598 = 10'h113 == _T_43[9:0] ? 4'hf : _GEN_1597; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1599 = 10'h114 == _T_43[9:0] ? 4'hf : _GEN_1598; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1600 = 10'h115 == _T_43[9:0] ? 4'hf : _GEN_1599; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1601 = 10'h116 == _T_43[9:0] ? 4'h9 : _GEN_1600; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1602 = 10'h117 == _T_43[9:0] ? 4'h3 : _GEN_1601; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1603 = 10'h118 == _T_43[9:0] ? 4'h3 : _GEN_1602; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1604 = 10'h119 == _T_43[9:0] ? 4'h3 : _GEN_1603; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1605 = 10'h11a == _T_43[9:0] ? 4'hf : _GEN_1604; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1606 = 10'h11b == _T_43[9:0] ? 4'h3 : _GEN_1605; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1607 = 10'h11c == _T_43[9:0] ? 4'h3 : _GEN_1606; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1608 = 10'h11d == _T_43[9:0] ? 4'h2 : _GEN_1607; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1609 = 10'h11e == _T_43[9:0] ? 4'h3 : _GEN_1608; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1610 = 10'h11f == _T_43[9:0] ? 4'h0 : _GEN_1609; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1611 = 10'h120 == _T_43[9:0] ? 4'h3 : _GEN_1610; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1612 = 10'h121 == _T_43[9:0] ? 4'h3 : _GEN_1611; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1613 = 10'h122 == _T_43[9:0] ? 4'h3 : _GEN_1612; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1614 = 10'h123 == _T_43[9:0] ? 4'h3 : _GEN_1613; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1615 = 10'h124 == _T_43[9:0] ? 4'h3 : _GEN_1614; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1616 = 10'h125 == _T_43[9:0] ? 4'h3 : _GEN_1615; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1617 = 10'h126 == _T_43[9:0] ? 4'h3 : _GEN_1616; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1618 = 10'h127 == _T_43[9:0] ? 4'h9 : _GEN_1617; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1619 = 10'h128 == _T_43[9:0] ? 4'hf : _GEN_1618; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1620 = 10'h129 == _T_43[9:0] ? 4'h3 : _GEN_1619; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1621 = 10'h12a == _T_43[9:0] ? 4'h3 : _GEN_1620; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1622 = 10'h12b == _T_43[9:0] ? 4'hf : _GEN_1621; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1623 = 10'h12c == _T_43[9:0] ? 4'hf : _GEN_1622; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1624 = 10'h12d == _T_43[9:0] ? 4'hf : _GEN_1623; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1625 = 10'h12e == _T_43[9:0] ? 4'hf : _GEN_1624; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1626 = 10'h12f == _T_43[9:0] ? 4'hf : _GEN_1625; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1627 = 10'h130 == _T_43[9:0] ? 4'hf : _GEN_1626; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1628 = 10'h131 == _T_43[9:0] ? 4'hf : _GEN_1627; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1629 = 10'h132 == _T_43[9:0] ? 4'hf : _GEN_1628; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1630 = 10'h133 == _T_43[9:0] ? 4'hf : _GEN_1629; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1631 = 10'h134 == _T_43[9:0] ? 4'h3 : _GEN_1630; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1632 = 10'h135 == _T_43[9:0] ? 4'h3 : _GEN_1631; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1633 = 10'h136 == _T_43[9:0] ? 4'hf : _GEN_1632; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1634 = 10'h137 == _T_43[9:0] ? 4'h9 : _GEN_1633; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1635 = 10'h138 == _T_43[9:0] ? 4'h3 : _GEN_1634; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1636 = 10'h139 == _T_43[9:0] ? 4'h3 : _GEN_1635; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1637 = 10'h13a == _T_43[9:0] ? 4'h3 : _GEN_1636; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1638 = 10'h13b == _T_43[9:0] ? 4'h3 : _GEN_1637; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1639 = 10'h13c == _T_43[9:0] ? 4'h3 : _GEN_1638; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1640 = 10'h13d == _T_43[9:0] ? 4'h3 : _GEN_1639; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1641 = 10'h13e == _T_43[9:0] ? 4'h3 : _GEN_1640; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1642 = 10'h13f == _T_43[9:0] ? 4'h0 : _GEN_1641; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1643 = 10'h140 == _T_43[9:0] ? 4'h3 : _GEN_1642; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1644 = 10'h141 == _T_43[9:0] ? 4'h3 : _GEN_1643; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1645 = 10'h142 == _T_43[9:0] ? 4'h2 : _GEN_1644; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1646 = 10'h143 == _T_43[9:0] ? 4'h3 : _GEN_1645; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1647 = 10'h144 == _T_43[9:0] ? 4'h3 : _GEN_1646; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1648 = 10'h145 == _T_43[9:0] ? 4'h3 : _GEN_1647; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1649 = 10'h146 == _T_43[9:0] ? 4'h9 : _GEN_1648; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1650 = 10'h147 == _T_43[9:0] ? 4'hf : _GEN_1649; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1651 = 10'h148 == _T_43[9:0] ? 4'h3 : _GEN_1650; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1652 = 10'h149 == _T_43[9:0] ? 4'h3 : _GEN_1651; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1653 = 10'h14a == _T_43[9:0] ? 4'h3 : _GEN_1652; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1654 = 10'h14b == _T_43[9:0] ? 4'h3 : _GEN_1653; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1655 = 10'h14c == _T_43[9:0] ? 4'h3 : _GEN_1654; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1656 = 10'h14d == _T_43[9:0] ? 4'h3 : _GEN_1655; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1657 = 10'h14e == _T_43[9:0] ? 4'h3 : _GEN_1656; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1658 = 10'h14f == _T_43[9:0] ? 4'h3 : _GEN_1657; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1659 = 10'h150 == _T_43[9:0] ? 4'h3 : _GEN_1658; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1660 = 10'h151 == _T_43[9:0] ? 4'h3 : _GEN_1659; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1661 = 10'h152 == _T_43[9:0] ? 4'h3 : _GEN_1660; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1662 = 10'h153 == _T_43[9:0] ? 4'h3 : _GEN_1661; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1663 = 10'h154 == _T_43[9:0] ? 4'h3 : _GEN_1662; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1664 = 10'h155 == _T_43[9:0] ? 4'h3 : _GEN_1663; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1665 = 10'h156 == _T_43[9:0] ? 4'h3 : _GEN_1664; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1666 = 10'h157 == _T_43[9:0] ? 4'hf : _GEN_1665; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1667 = 10'h158 == _T_43[9:0] ? 4'h3 : _GEN_1666; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1668 = 10'h159 == _T_43[9:0] ? 4'h3 : _GEN_1667; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1669 = 10'h15a == _T_43[9:0] ? 4'h3 : _GEN_1668; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1670 = 10'h15b == _T_43[9:0] ? 4'h3 : _GEN_1669; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1671 = 10'h15c == _T_43[9:0] ? 4'h3 : _GEN_1670; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1672 = 10'h15d == _T_43[9:0] ? 4'h3 : _GEN_1671; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1673 = 10'h15e == _T_43[9:0] ? 4'h2 : _GEN_1672; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1674 = 10'h15f == _T_43[9:0] ? 4'h0 : _GEN_1673; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1675 = 10'h160 == _T_43[9:0] ? 4'h3 : _GEN_1674; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1676 = 10'h161 == _T_43[9:0] ? 4'h3 : _GEN_1675; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1677 = 10'h162 == _T_43[9:0] ? 4'h3 : _GEN_1676; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1678 = 10'h163 == _T_43[9:0] ? 4'h2 : _GEN_1677; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1679 = 10'h164 == _T_43[9:0] ? 4'h3 : _GEN_1678; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1680 = 10'h165 == _T_43[9:0] ? 4'h9 : _GEN_1679; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1681 = 10'h166 == _T_43[9:0] ? 4'hf : _GEN_1680; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1682 = 10'h167 == _T_43[9:0] ? 4'hf : _GEN_1681; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1683 = 10'h168 == _T_43[9:0] ? 4'hd : _GEN_1682; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1684 = 10'h169 == _T_43[9:0] ? 4'h9 : _GEN_1683; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1685 = 10'h16a == _T_43[9:0] ? 4'hd : _GEN_1684; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1686 = 10'h16b == _T_43[9:0] ? 4'hd : _GEN_1685; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1687 = 10'h16c == _T_43[9:0] ? 4'h3 : _GEN_1686; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1688 = 10'h16d == _T_43[9:0] ? 4'h3 : _GEN_1687; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1689 = 10'h16e == _T_43[9:0] ? 4'h3 : _GEN_1688; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1690 = 10'h16f == _T_43[9:0] ? 4'h3 : _GEN_1689; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1691 = 10'h170 == _T_43[9:0] ? 4'h3 : _GEN_1690; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1692 = 10'h171 == _T_43[9:0] ? 4'h3 : _GEN_1691; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1693 = 10'h172 == _T_43[9:0] ? 4'h3 : _GEN_1692; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1694 = 10'h173 == _T_43[9:0] ? 4'h3 : _GEN_1693; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1695 = 10'h174 == _T_43[9:0] ? 4'h3 : _GEN_1694; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1696 = 10'h175 == _T_43[9:0] ? 4'h3 : _GEN_1695; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1697 = 10'h176 == _T_43[9:0] ? 4'hf : _GEN_1696; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1698 = 10'h177 == _T_43[9:0] ? 4'hf : _GEN_1697; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1699 = 10'h178 == _T_43[9:0] ? 4'h9 : _GEN_1698; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1700 = 10'h179 == _T_43[9:0] ? 4'h3 : _GEN_1699; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1701 = 10'h17a == _T_43[9:0] ? 4'h3 : _GEN_1700; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1702 = 10'h17b == _T_43[9:0] ? 4'h3 : _GEN_1701; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1703 = 10'h17c == _T_43[9:0] ? 4'h3 : _GEN_1702; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1704 = 10'h17d == _T_43[9:0] ? 4'h2 : _GEN_1703; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1705 = 10'h17e == _T_43[9:0] ? 4'h3 : _GEN_1704; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1706 = 10'h17f == _T_43[9:0] ? 4'h0 : _GEN_1705; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1707 = 10'h180 == _T_43[9:0] ? 4'hd : _GEN_1706; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1708 = 10'h181 == _T_43[9:0] ? 4'hd : _GEN_1707; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1709 = 10'h182 == _T_43[9:0] ? 4'hd : _GEN_1708; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1710 = 10'h183 == _T_43[9:0] ? 4'hd : _GEN_1709; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1711 = 10'h184 == _T_43[9:0] ? 4'h3 : _GEN_1710; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1712 = 10'h185 == _T_43[9:0] ? 4'h9 : _GEN_1711; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1713 = 10'h186 == _T_43[9:0] ? 4'hb : _GEN_1712; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1714 = 10'h187 == _T_43[9:0] ? 4'hf : _GEN_1713; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1715 = 10'h188 == _T_43[9:0] ? 4'hd : _GEN_1714; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1716 = 10'h189 == _T_43[9:0] ? 4'hd : _GEN_1715; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1717 = 10'h18a == _T_43[9:0] ? 4'hd : _GEN_1716; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1718 = 10'h18b == _T_43[9:0] ? 4'hd : _GEN_1717; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1719 = 10'h18c == _T_43[9:0] ? 4'hd : _GEN_1718; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1720 = 10'h18d == _T_43[9:0] ? 4'hd : _GEN_1719; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1721 = 10'h18e == _T_43[9:0] ? 4'hd : _GEN_1720; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1722 = 10'h18f == _T_43[9:0] ? 4'hd : _GEN_1721; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1723 = 10'h190 == _T_43[9:0] ? 4'hd : _GEN_1722; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1724 = 10'h191 == _T_43[9:0] ? 4'hd : _GEN_1723; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1725 = 10'h192 == _T_43[9:0] ? 4'h9 : _GEN_1724; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1726 = 10'h193 == _T_43[9:0] ? 4'hd : _GEN_1725; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1727 = 10'h194 == _T_43[9:0] ? 4'hd : _GEN_1726; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1728 = 10'h195 == _T_43[9:0] ? 4'hd : _GEN_1727; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1729 = 10'h196 == _T_43[9:0] ? 4'hf : _GEN_1728; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1730 = 10'h197 == _T_43[9:0] ? 4'h3 : _GEN_1729; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1731 = 10'h198 == _T_43[9:0] ? 4'h9 : _GEN_1730; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1732 = 10'h199 == _T_43[9:0] ? 4'h3 : _GEN_1731; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1733 = 10'h19a == _T_43[9:0] ? 4'h3 : _GEN_1732; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1734 = 10'h19b == _T_43[9:0] ? 4'h3 : _GEN_1733; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1735 = 10'h19c == _T_43[9:0] ? 4'h3 : _GEN_1734; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1736 = 10'h19d == _T_43[9:0] ? 4'h3 : _GEN_1735; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1737 = 10'h19e == _T_43[9:0] ? 4'h3 : _GEN_1736; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1738 = 10'h19f == _T_43[9:0] ? 4'h0 : _GEN_1737; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1739 = 10'h1a0 == _T_43[9:0] ? 4'hd : _GEN_1738; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1740 = 10'h1a1 == _T_43[9:0] ? 4'hd : _GEN_1739; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1741 = 10'h1a2 == _T_43[9:0] ? 4'h9 : _GEN_1740; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1742 = 10'h1a3 == _T_43[9:0] ? 4'hd : _GEN_1741; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1743 = 10'h1a4 == _T_43[9:0] ? 4'h3 : _GEN_1742; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1744 = 10'h1a5 == _T_43[9:0] ? 4'hf : _GEN_1743; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1745 = 10'h1a6 == _T_43[9:0] ? 4'hd : _GEN_1744; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1746 = 10'h1a7 == _T_43[9:0] ? 4'hf : _GEN_1745; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1747 = 10'h1a8 == _T_43[9:0] ? 4'hb : _GEN_1746; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1748 = 10'h1a9 == _T_43[9:0] ? 4'hd : _GEN_1747; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1749 = 10'h1aa == _T_43[9:0] ? 4'hd : _GEN_1748; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1750 = 10'h1ab == _T_43[9:0] ? 4'h9 : _GEN_1749; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1751 = 10'h1ac == _T_43[9:0] ? 4'hd : _GEN_1750; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1752 = 10'h1ad == _T_43[9:0] ? 4'hd : _GEN_1751; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1753 = 10'h1ae == _T_43[9:0] ? 4'hd : _GEN_1752; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1754 = 10'h1af == _T_43[9:0] ? 4'hd : _GEN_1753; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1755 = 10'h1b0 == _T_43[9:0] ? 4'hd : _GEN_1754; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1756 = 10'h1b1 == _T_43[9:0] ? 4'hd : _GEN_1755; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1757 = 10'h1b2 == _T_43[9:0] ? 4'hd : _GEN_1756; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1758 = 10'h1b3 == _T_43[9:0] ? 4'hd : _GEN_1757; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1759 = 10'h1b4 == _T_43[9:0] ? 4'hd : _GEN_1758; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1760 = 10'h1b5 == _T_43[9:0] ? 4'hd : _GEN_1759; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1761 = 10'h1b6 == _T_43[9:0] ? 4'hf : _GEN_1760; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1762 = 10'h1b7 == _T_43[9:0] ? 4'hd : _GEN_1761; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1763 = 10'h1b8 == _T_43[9:0] ? 4'hf : _GEN_1762; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1764 = 10'h1b9 == _T_43[9:0] ? 4'hd : _GEN_1763; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1765 = 10'h1ba == _T_43[9:0] ? 4'hd : _GEN_1764; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1766 = 10'h1bb == _T_43[9:0] ? 4'hd : _GEN_1765; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1767 = 10'h1bc == _T_43[9:0] ? 4'h2 : _GEN_1766; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1768 = 10'h1bd == _T_43[9:0] ? 4'h3 : _GEN_1767; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1769 = 10'h1be == _T_43[9:0] ? 4'hd : _GEN_1768; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1770 = 10'h1bf == _T_43[9:0] ? 4'h0 : _GEN_1769; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1771 = 10'h1c0 == _T_43[9:0] ? 4'hd : _GEN_1770; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1772 = 10'h1c1 == _T_43[9:0] ? 4'hd : _GEN_1771; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1773 = 10'h1c2 == _T_43[9:0] ? 4'hd : _GEN_1772; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1774 = 10'h1c3 == _T_43[9:0] ? 4'h2 : _GEN_1773; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1775 = 10'h1c4 == _T_43[9:0] ? 4'h2 : _GEN_1774; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1776 = 10'h1c5 == _T_43[9:0] ? 4'hd : _GEN_1775; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1777 = 10'h1c6 == _T_43[9:0] ? 4'hd : _GEN_1776; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1778 = 10'h1c7 == _T_43[9:0] ? 4'hd : _GEN_1777; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1779 = 10'h1c8 == _T_43[9:0] ? 4'hd : _GEN_1778; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1780 = 10'h1c9 == _T_43[9:0] ? 4'hb : _GEN_1779; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1781 = 10'h1ca == _T_43[9:0] ? 4'hb : _GEN_1780; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1782 = 10'h1cb == _T_43[9:0] ? 4'hb : _GEN_1781; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1783 = 10'h1cc == _T_43[9:0] ? 4'hb : _GEN_1782; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1784 = 10'h1cd == _T_43[9:0] ? 4'hb : _GEN_1783; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1785 = 10'h1ce == _T_43[9:0] ? 4'hb : _GEN_1784; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1786 = 10'h1cf == _T_43[9:0] ? 4'hb : _GEN_1785; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1787 = 10'h1d0 == _T_43[9:0] ? 4'hb : _GEN_1786; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1788 = 10'h1d1 == _T_43[9:0] ? 4'hb : _GEN_1787; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1789 = 10'h1d2 == _T_43[9:0] ? 4'hb : _GEN_1788; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1790 = 10'h1d3 == _T_43[9:0] ? 4'hb : _GEN_1789; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1791 = 10'h1d4 == _T_43[9:0] ? 4'hb : _GEN_1790; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1792 = 10'h1d5 == _T_43[9:0] ? 4'hb : _GEN_1791; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1793 = 10'h1d6 == _T_43[9:0] ? 4'hd : _GEN_1792; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1794 = 10'h1d7 == _T_43[9:0] ? 4'hd : _GEN_1793; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1795 = 10'h1d8 == _T_43[9:0] ? 4'hd : _GEN_1794; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1796 = 10'h1d9 == _T_43[9:0] ? 4'hd : _GEN_1795; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1797 = 10'h1da == _T_43[9:0] ? 4'hd : _GEN_1796; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1798 = 10'h1db == _T_43[9:0] ? 4'hd : _GEN_1797; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1799 = 10'h1dc == _T_43[9:0] ? 4'hd : _GEN_1798; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1800 = 10'h1dd == _T_43[9:0] ? 4'h3 : _GEN_1799; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1801 = 10'h1de == _T_43[9:0] ? 4'hd : _GEN_1800; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1802 = 10'h1df == _T_43[9:0] ? 4'h0 : _GEN_1801; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1803 = 10'h1e0 == _T_43[9:0] ? 4'h9 : _GEN_1802; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1804 = 10'h1e1 == _T_43[9:0] ? 4'hd : _GEN_1803; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1805 = 10'h1e2 == _T_43[9:0] ? 4'h2 : _GEN_1804; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1806 = 10'h1e3 == _T_43[9:0] ? 4'h2 : _GEN_1805; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1807 = 10'h1e4 == _T_43[9:0] ? 4'hd : _GEN_1806; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1808 = 10'h1e5 == _T_43[9:0] ? 4'hd : _GEN_1807; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1809 = 10'h1e6 == _T_43[9:0] ? 4'hd : _GEN_1808; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1810 = 10'h1e7 == _T_43[9:0] ? 4'hd : _GEN_1809; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1811 = 10'h1e8 == _T_43[9:0] ? 4'hb : _GEN_1810; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1812 = 10'h1e9 == _T_43[9:0] ? 4'hd : _GEN_1811; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1813 = 10'h1ea == _T_43[9:0] ? 4'hd : _GEN_1812; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1814 = 10'h1eb == _T_43[9:0] ? 4'hb : _GEN_1813; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1815 = 10'h1ec == _T_43[9:0] ? 4'hd : _GEN_1814; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1816 = 10'h1ed == _T_43[9:0] ? 4'hb : _GEN_1815; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1817 = 10'h1ee == _T_43[9:0] ? 4'hd : _GEN_1816; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1818 = 10'h1ef == _T_43[9:0] ? 4'hb : _GEN_1817; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1819 = 10'h1f0 == _T_43[9:0] ? 4'hd : _GEN_1818; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1820 = 10'h1f1 == _T_43[9:0] ? 4'hb : _GEN_1819; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1821 = 10'h1f2 == _T_43[9:0] ? 4'hb : _GEN_1820; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1822 = 10'h1f3 == _T_43[9:0] ? 4'hd : _GEN_1821; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1823 = 10'h1f4 == _T_43[9:0] ? 4'hb : _GEN_1822; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1824 = 10'h1f5 == _T_43[9:0] ? 4'hb : _GEN_1823; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1825 = 10'h1f6 == _T_43[9:0] ? 4'hd : _GEN_1824; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1826 = 10'h1f7 == _T_43[9:0] ? 4'hd : _GEN_1825; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1827 = 10'h1f8 == _T_43[9:0] ? 4'hd : _GEN_1826; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1828 = 10'h1f9 == _T_43[9:0] ? 4'hd : _GEN_1827; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1829 = 10'h1fa == _T_43[9:0] ? 4'h9 : _GEN_1828; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1830 = 10'h1fb == _T_43[9:0] ? 4'hd : _GEN_1829; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1831 = 10'h1fc == _T_43[9:0] ? 4'hd : _GEN_1830; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1832 = 10'h1fd == _T_43[9:0] ? 4'h2 : _GEN_1831; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1833 = 10'h1fe == _T_43[9:0] ? 4'hd : _GEN_1832; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1834 = 10'h1ff == _T_43[9:0] ? 4'h0 : _GEN_1833; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1835 = 10'h200 == _T_43[9:0] ? 4'hd : _GEN_1834; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1836 = 10'h201 == _T_43[9:0] ? 4'hd : _GEN_1835; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1837 = 10'h202 == _T_43[9:0] ? 4'h3 : _GEN_1836; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1838 = 10'h203 == _T_43[9:0] ? 4'hd : _GEN_1837; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1839 = 10'h204 == _T_43[9:0] ? 4'hd : _GEN_1838; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1840 = 10'h205 == _T_43[9:0] ? 4'hd : _GEN_1839; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1841 = 10'h206 == _T_43[9:0] ? 4'hb : _GEN_1840; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1842 = 10'h207 == _T_43[9:0] ? 4'hb : _GEN_1841; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1843 = 10'h208 == _T_43[9:0] ? 4'hd : _GEN_1842; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1844 = 10'h209 == _T_43[9:0] ? 4'hd : _GEN_1843; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1845 = 10'h20a == _T_43[9:0] ? 4'hd : _GEN_1844; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1846 = 10'h20b == _T_43[9:0] ? 4'hb : _GEN_1845; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1847 = 10'h20c == _T_43[9:0] ? 4'hd : _GEN_1846; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1848 = 10'h20d == _T_43[9:0] ? 4'hb : _GEN_1847; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1849 = 10'h20e == _T_43[9:0] ? 4'hd : _GEN_1848; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1850 = 10'h20f == _T_43[9:0] ? 4'hb : _GEN_1849; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1851 = 10'h210 == _T_43[9:0] ? 4'hd : _GEN_1850; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1852 = 10'h211 == _T_43[9:0] ? 4'hd : _GEN_1851; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1853 = 10'h212 == _T_43[9:0] ? 4'hb : _GEN_1852; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1854 = 10'h213 == _T_43[9:0] ? 4'hb : _GEN_1853; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1855 = 10'h214 == _T_43[9:0] ? 4'hb : _GEN_1854; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1856 = 10'h215 == _T_43[9:0] ? 4'hd : _GEN_1855; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1857 = 10'h216 == _T_43[9:0] ? 4'hd : _GEN_1856; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1858 = 10'h217 == _T_43[9:0] ? 4'hd : _GEN_1857; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1859 = 10'h218 == _T_43[9:0] ? 4'hd : _GEN_1858; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1860 = 10'h219 == _T_43[9:0] ? 4'hd : _GEN_1859; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1861 = 10'h21a == _T_43[9:0] ? 4'hd : _GEN_1860; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1862 = 10'h21b == _T_43[9:0] ? 4'hd : _GEN_1861; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1863 = 10'h21c == _T_43[9:0] ? 4'h3 : _GEN_1862; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1864 = 10'h21d == _T_43[9:0] ? 4'h2 : _GEN_1863; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1865 = 10'h21e == _T_43[9:0] ? 4'hd : _GEN_1864; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1866 = 10'h21f == _T_43[9:0] ? 4'h0 : _GEN_1865; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1867 = 10'h220 == _T_43[9:0] ? 4'h0 : _GEN_1866; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1868 = 10'h221 == _T_43[9:0] ? 4'h0 : _GEN_1867; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1869 = 10'h222 == _T_43[9:0] ? 4'h0 : _GEN_1868; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1870 = 10'h223 == _T_43[9:0] ? 4'h0 : _GEN_1869; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1871 = 10'h224 == _T_43[9:0] ? 4'h0 : _GEN_1870; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1872 = 10'h225 == _T_43[9:0] ? 4'h0 : _GEN_1871; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1873 = 10'h226 == _T_43[9:0] ? 4'h0 : _GEN_1872; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1874 = 10'h227 == _T_43[9:0] ? 4'h0 : _GEN_1873; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1875 = 10'h228 == _T_43[9:0] ? 4'h0 : _GEN_1874; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1876 = 10'h229 == _T_43[9:0] ? 4'h0 : _GEN_1875; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1877 = 10'h22a == _T_43[9:0] ? 4'h0 : _GEN_1876; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1878 = 10'h22b == _T_43[9:0] ? 4'h0 : _GEN_1877; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1879 = 10'h22c == _T_43[9:0] ? 4'h0 : _GEN_1878; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1880 = 10'h22d == _T_43[9:0] ? 4'h0 : _GEN_1879; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1881 = 10'h22e == _T_43[9:0] ? 4'h0 : _GEN_1880; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1882 = 10'h22f == _T_43[9:0] ? 4'h0 : _GEN_1881; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1883 = 10'h230 == _T_43[9:0] ? 4'h0 : _GEN_1882; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1884 = 10'h231 == _T_43[9:0] ? 4'h0 : _GEN_1883; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1885 = 10'h232 == _T_43[9:0] ? 4'h0 : _GEN_1884; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1886 = 10'h233 == _T_43[9:0] ? 4'h0 : _GEN_1885; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1887 = 10'h234 == _T_43[9:0] ? 4'h0 : _GEN_1886; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1888 = 10'h235 == _T_43[9:0] ? 4'h0 : _GEN_1887; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1889 = 10'h236 == _T_43[9:0] ? 4'h0 : _GEN_1888; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1890 = 10'h237 == _T_43[9:0] ? 4'h0 : _GEN_1889; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1891 = 10'h238 == _T_43[9:0] ? 4'h0 : _GEN_1890; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1892 = 10'h239 == _T_43[9:0] ? 4'h0 : _GEN_1891; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1893 = 10'h23a == _T_43[9:0] ? 4'h0 : _GEN_1892; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1894 = 10'h23b == _T_43[9:0] ? 4'h0 : _GEN_1893; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1895 = 10'h23c == _T_43[9:0] ? 4'h0 : _GEN_1894; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1896 = 10'h23d == _T_43[9:0] ? 4'h0 : _GEN_1895; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1897 = 10'h23e == _T_43[9:0] ? 4'h0 : _GEN_1896; // @[Filter.scala 191:142]
  wire [3:0] _GEN_1898 = 10'h23f == _T_43[9:0] ? 4'h0 : _GEN_1897; // @[Filter.scala 191:142]
  wire [7:0] _T_57 = _GEN_1898 * 4'ha; // @[Filter.scala 191:142]
  wire [10:0] _GEN_28303 = {{3'd0}, _T_57}; // @[Filter.scala 191:109]
  wire [10:0] _T_59 = _T_52 + _GEN_28303; // @[Filter.scala 191:109]
  wire [10:0] _T_60 = _T_59 / 11'h64; // @[Filter.scala 191:150]
  wire  _T_62 = _T_33 >= 6'h20; // @[Filter.scala 194:31]
  wire  _T_66 = _T_40 >= 32'h12; // @[Filter.scala 194:63]
  wire  _T_67 = _T_62 | _T_66; // @[Filter.scala 194:58]
  wire [10:0] _GEN_2475 = io_SPI_distort ? _T_60 : {{7'd0}, _GEN_746}; // @[Filter.scala 196:35]
  wire [10:0] _GEN_2476 = _T_67 ? 11'h0 : _GEN_2475; // @[Filter.scala 194:80]
  wire [10:0] _GEN_3053 = io_SPI_distort ? _T_60 : {{7'd0}, _GEN_1322}; // @[Filter.scala 196:35]
  wire [10:0] _GEN_3054 = _T_67 ? 11'h0 : _GEN_3053; // @[Filter.scala 194:80]
  wire [10:0] _GEN_3631 = io_SPI_distort ? _T_60 : {{7'd0}, _GEN_1898}; // @[Filter.scala 196:35]
  wire [10:0] _GEN_3632 = _T_67 ? 11'h0 : _GEN_3631; // @[Filter.scala 194:80]
  wire [31:0] _T_95 = pixelIndex + 32'h1; // @[Filter.scala 189:31]
  wire [31:0] _GEN_1 = _T_95 % 32'h20; // @[Filter.scala 189:38]
  wire [5:0] _T_96 = _GEN_1[5:0]; // @[Filter.scala 189:38]
  wire [5:0] _T_98 = _T_96 + _GEN_28295; // @[Filter.scala 189:53]
  wire [5:0] _T_100 = _T_98 - 6'h1; // @[Filter.scala 189:69]
  wire [31:0] _T_103 = _T_95 / 32'h20; // @[Filter.scala 190:38]
  wire [31:0] _T_105 = _T_103 + _GEN_28296; // @[Filter.scala 190:53]
  wire [31:0] _T_107 = _T_105 - 32'h1; // @[Filter.scala 190:69]
  wire [37:0] _T_108 = _T_107 * 32'h20; // @[Filter.scala 191:42]
  wire [37:0] _GEN_28309 = {{32'd0}, _T_100}; // @[Filter.scala 191:57]
  wire [37:0] _T_110 = _T_108 + _GEN_28309; // @[Filter.scala 191:57]
  wire [3:0] _GEN_3636 = 10'h3 == _T_110[9:0] ? 4'h3 : 4'ha; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3637 = 10'h4 == _T_110[9:0] ? 4'ha : _GEN_3636; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3638 = 10'h5 == _T_110[9:0] ? 4'ha : _GEN_3637; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3639 = 10'h6 == _T_110[9:0] ? 4'ha : _GEN_3638; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3640 = 10'h7 == _T_110[9:0] ? 4'ha : _GEN_3639; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3641 = 10'h8 == _T_110[9:0] ? 4'ha : _GEN_3640; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3642 = 10'h9 == _T_110[9:0] ? 4'ha : _GEN_3641; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3643 = 10'ha == _T_110[9:0] ? 4'ha : _GEN_3642; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3644 = 10'hb == _T_110[9:0] ? 4'ha : _GEN_3643; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3645 = 10'hc == _T_110[9:0] ? 4'ha : _GEN_3644; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3646 = 10'hd == _T_110[9:0] ? 4'ha : _GEN_3645; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3647 = 10'he == _T_110[9:0] ? 4'ha : _GEN_3646; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3648 = 10'hf == _T_110[9:0] ? 4'ha : _GEN_3647; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3649 = 10'h10 == _T_110[9:0] ? 4'ha : _GEN_3648; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3650 = 10'h11 == _T_110[9:0] ? 4'ha : _GEN_3649; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3651 = 10'h12 == _T_110[9:0] ? 4'ha : _GEN_3650; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3652 = 10'h13 == _T_110[9:0] ? 4'ha : _GEN_3651; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3653 = 10'h14 == _T_110[9:0] ? 4'ha : _GEN_3652; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3654 = 10'h15 == _T_110[9:0] ? 4'ha : _GEN_3653; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3655 = 10'h16 == _T_110[9:0] ? 4'ha : _GEN_3654; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3656 = 10'h17 == _T_110[9:0] ? 4'ha : _GEN_3655; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3657 = 10'h18 == _T_110[9:0] ? 4'ha : _GEN_3656; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3658 = 10'h19 == _T_110[9:0] ? 4'ha : _GEN_3657; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3659 = 10'h1a == _T_110[9:0] ? 4'ha : _GEN_3658; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3660 = 10'h1b == _T_110[9:0] ? 4'ha : _GEN_3659; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3661 = 10'h1c == _T_110[9:0] ? 4'ha : _GEN_3660; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3662 = 10'h1d == _T_110[9:0] ? 4'ha : _GEN_3661; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3663 = 10'h1e == _T_110[9:0] ? 4'ha : _GEN_3662; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3664 = 10'h1f == _T_110[9:0] ? 4'h0 : _GEN_3663; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3665 = 10'h20 == _T_110[9:0] ? 4'ha : _GEN_3664; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3666 = 10'h21 == _T_110[9:0] ? 4'ha : _GEN_3665; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3667 = 10'h22 == _T_110[9:0] ? 4'ha : _GEN_3666; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3668 = 10'h23 == _T_110[9:0] ? 4'h3 : _GEN_3667; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3669 = 10'h24 == _T_110[9:0] ? 4'ha : _GEN_3668; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3670 = 10'h25 == _T_110[9:0] ? 4'ha : _GEN_3669; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3671 = 10'h26 == _T_110[9:0] ? 4'ha : _GEN_3670; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3672 = 10'h27 == _T_110[9:0] ? 4'h1 : _GEN_3671; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3673 = 10'h28 == _T_110[9:0] ? 4'h1 : _GEN_3672; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3674 = 10'h29 == _T_110[9:0] ? 4'ha : _GEN_3673; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3675 = 10'h2a == _T_110[9:0] ? 4'ha : _GEN_3674; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3676 = 10'h2b == _T_110[9:0] ? 4'ha : _GEN_3675; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3677 = 10'h2c == _T_110[9:0] ? 4'ha : _GEN_3676; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3678 = 10'h2d == _T_110[9:0] ? 4'ha : _GEN_3677; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3679 = 10'h2e == _T_110[9:0] ? 4'ha : _GEN_3678; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3680 = 10'h2f == _T_110[9:0] ? 4'ha : _GEN_3679; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3681 = 10'h30 == _T_110[9:0] ? 4'ha : _GEN_3680; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3682 = 10'h31 == _T_110[9:0] ? 4'ha : _GEN_3681; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3683 = 10'h32 == _T_110[9:0] ? 4'ha : _GEN_3682; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3684 = 10'h33 == _T_110[9:0] ? 4'ha : _GEN_3683; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3685 = 10'h34 == _T_110[9:0] ? 4'ha : _GEN_3684; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3686 = 10'h35 == _T_110[9:0] ? 4'ha : _GEN_3685; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3687 = 10'h36 == _T_110[9:0] ? 4'ha : _GEN_3686; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3688 = 10'h37 == _T_110[9:0] ? 4'h1 : _GEN_3687; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3689 = 10'h38 == _T_110[9:0] ? 4'h1 : _GEN_3688; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3690 = 10'h39 == _T_110[9:0] ? 4'ha : _GEN_3689; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3691 = 10'h3a == _T_110[9:0] ? 4'ha : _GEN_3690; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3692 = 10'h3b == _T_110[9:0] ? 4'ha : _GEN_3691; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3693 = 10'h3c == _T_110[9:0] ? 4'ha : _GEN_3692; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3694 = 10'h3d == _T_110[9:0] ? 4'h3 : _GEN_3693; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3695 = 10'h3e == _T_110[9:0] ? 4'ha : _GEN_3694; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3696 = 10'h3f == _T_110[9:0] ? 4'h0 : _GEN_3695; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3697 = 10'h40 == _T_110[9:0] ? 4'ha : _GEN_3696; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3698 = 10'h41 == _T_110[9:0] ? 4'ha : _GEN_3697; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3699 = 10'h42 == _T_110[9:0] ? 4'ha : _GEN_3698; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3700 = 10'h43 == _T_110[9:0] ? 4'h2 : _GEN_3699; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3701 = 10'h44 == _T_110[9:0] ? 4'h3 : _GEN_3700; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3702 = 10'h45 == _T_110[9:0] ? 4'h0 : _GEN_3701; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3703 = 10'h46 == _T_110[9:0] ? 4'h0 : _GEN_3702; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3704 = 10'h47 == _T_110[9:0] ? 4'h0 : _GEN_3703; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3705 = 10'h48 == _T_110[9:0] ? 4'h0 : _GEN_3704; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3706 = 10'h49 == _T_110[9:0] ? 4'ha : _GEN_3705; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3707 = 10'h4a == _T_110[9:0] ? 4'ha : _GEN_3706; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3708 = 10'h4b == _T_110[9:0] ? 4'ha : _GEN_3707; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3709 = 10'h4c == _T_110[9:0] ? 4'ha : _GEN_3708; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3710 = 10'h4d == _T_110[9:0] ? 4'ha : _GEN_3709; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3711 = 10'h4e == _T_110[9:0] ? 4'ha : _GEN_3710; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3712 = 10'h4f == _T_110[9:0] ? 4'ha : _GEN_3711; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3713 = 10'h50 == _T_110[9:0] ? 4'ha : _GEN_3712; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3714 = 10'h51 == _T_110[9:0] ? 4'ha : _GEN_3713; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3715 = 10'h52 == _T_110[9:0] ? 4'ha : _GEN_3714; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3716 = 10'h53 == _T_110[9:0] ? 4'ha : _GEN_3715; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3717 = 10'h54 == _T_110[9:0] ? 4'h1 : _GEN_3716; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3718 = 10'h55 == _T_110[9:0] ? 4'h1 : _GEN_3717; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3719 = 10'h56 == _T_110[9:0] ? 4'h1 : _GEN_3718; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3720 = 10'h57 == _T_110[9:0] ? 4'h0 : _GEN_3719; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3721 = 10'h58 == _T_110[9:0] ? 4'ha : _GEN_3720; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3722 = 10'h59 == _T_110[9:0] ? 4'h0 : _GEN_3721; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3723 = 10'h5a == _T_110[9:0] ? 4'ha : _GEN_3722; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3724 = 10'h5b == _T_110[9:0] ? 4'ha : _GEN_3723; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3725 = 10'h5c == _T_110[9:0] ? 4'ha : _GEN_3724; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3726 = 10'h5d == _T_110[9:0] ? 4'h3 : _GEN_3725; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3727 = 10'h5e == _T_110[9:0] ? 4'ha : _GEN_3726; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3728 = 10'h5f == _T_110[9:0] ? 4'h0 : _GEN_3727; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3729 = 10'h60 == _T_110[9:0] ? 4'ha : _GEN_3728; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3730 = 10'h61 == _T_110[9:0] ? 4'ha : _GEN_3729; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3731 = 10'h62 == _T_110[9:0] ? 4'ha : _GEN_3730; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3732 = 10'h63 == _T_110[9:0] ? 4'ha : _GEN_3731; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3733 = 10'h64 == _T_110[9:0] ? 4'h3 : _GEN_3732; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3734 = 10'h65 == _T_110[9:0] ? 4'h0 : _GEN_3733; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3735 = 10'h66 == _T_110[9:0] ? 4'ha : _GEN_3734; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3736 = 10'h67 == _T_110[9:0] ? 4'ha : _GEN_3735; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3737 = 10'h68 == _T_110[9:0] ? 4'ha : _GEN_3736; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3738 = 10'h69 == _T_110[9:0] ? 4'h0 : _GEN_3737; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3739 = 10'h6a == _T_110[9:0] ? 4'h1 : _GEN_3738; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3740 = 10'h6b == _T_110[9:0] ? 4'h1 : _GEN_3739; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3741 = 10'h6c == _T_110[9:0] ? 4'ha : _GEN_3740; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3742 = 10'h6d == _T_110[9:0] ? 4'ha : _GEN_3741; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3743 = 10'h6e == _T_110[9:0] ? 4'ha : _GEN_3742; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3744 = 10'h6f == _T_110[9:0] ? 4'ha : _GEN_3743; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3745 = 10'h70 == _T_110[9:0] ? 4'ha : _GEN_3744; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3746 = 10'h71 == _T_110[9:0] ? 4'ha : _GEN_3745; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3747 = 10'h72 == _T_110[9:0] ? 4'ha : _GEN_3746; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3748 = 10'h73 == _T_110[9:0] ? 4'h1 : _GEN_3747; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3749 = 10'h74 == _T_110[9:0] ? 4'h0 : _GEN_3748; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3750 = 10'h75 == _T_110[9:0] ? 4'h0 : _GEN_3749; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3751 = 10'h76 == _T_110[9:0] ? 4'h0 : _GEN_3750; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3752 = 10'h77 == _T_110[9:0] ? 4'ha : _GEN_3751; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3753 = 10'h78 == _T_110[9:0] ? 4'ha : _GEN_3752; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3754 = 10'h79 == _T_110[9:0] ? 4'ha : _GEN_3753; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3755 = 10'h7a == _T_110[9:0] ? 4'h0 : _GEN_3754; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3756 = 10'h7b == _T_110[9:0] ? 4'ha : _GEN_3755; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3757 = 10'h7c == _T_110[9:0] ? 4'ha : _GEN_3756; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3758 = 10'h7d == _T_110[9:0] ? 4'h2 : _GEN_3757; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3759 = 10'h7e == _T_110[9:0] ? 4'h3 : _GEN_3758; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3760 = 10'h7f == _T_110[9:0] ? 4'h0 : _GEN_3759; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3761 = 10'h80 == _T_110[9:0] ? 4'ha : _GEN_3760; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3762 = 10'h81 == _T_110[9:0] ? 4'ha : _GEN_3761; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3763 = 10'h82 == _T_110[9:0] ? 4'h1 : _GEN_3762; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3764 = 10'h83 == _T_110[9:0] ? 4'h0 : _GEN_3763; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3765 = 10'h84 == _T_110[9:0] ? 4'h2 : _GEN_3764; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3766 = 10'h85 == _T_110[9:0] ? 4'h1 : _GEN_3765; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3767 = 10'h86 == _T_110[9:0] ? 4'h1 : _GEN_3766; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3768 = 10'h87 == _T_110[9:0] ? 4'ha : _GEN_3767; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3769 = 10'h88 == _T_110[9:0] ? 4'ha : _GEN_3768; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3770 = 10'h89 == _T_110[9:0] ? 4'h0 : _GEN_3769; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3771 = 10'h8a == _T_110[9:0] ? 4'h0 : _GEN_3770; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3772 = 10'h8b == _T_110[9:0] ? 4'h1 : _GEN_3771; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3773 = 10'h8c == _T_110[9:0] ? 4'h1 : _GEN_3772; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3774 = 10'h8d == _T_110[9:0] ? 4'h1 : _GEN_3773; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3775 = 10'h8e == _T_110[9:0] ? 4'h1 : _GEN_3774; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3776 = 10'h8f == _T_110[9:0] ? 4'h1 : _GEN_3775; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3777 = 10'h90 == _T_110[9:0] ? 4'h1 : _GEN_3776; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3778 = 10'h91 == _T_110[9:0] ? 4'h1 : _GEN_3777; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3779 = 10'h92 == _T_110[9:0] ? 4'h1 : _GEN_3778; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3780 = 10'h93 == _T_110[9:0] ? 4'h0 : _GEN_3779; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3781 = 10'h94 == _T_110[9:0] ? 4'h0 : _GEN_3780; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3782 = 10'h95 == _T_110[9:0] ? 4'ha : _GEN_3781; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3783 = 10'h96 == _T_110[9:0] ? 4'ha : _GEN_3782; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3784 = 10'h97 == _T_110[9:0] ? 4'ha : _GEN_3783; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3785 = 10'h98 == _T_110[9:0] ? 4'h1 : _GEN_3784; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3786 = 10'h99 == _T_110[9:0] ? 4'h0 : _GEN_3785; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3787 = 10'h9a == _T_110[9:0] ? 4'h1 : _GEN_3786; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3788 = 10'h9b == _T_110[9:0] ? 4'h1 : _GEN_3787; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3789 = 10'h9c == _T_110[9:0] ? 4'ha : _GEN_3788; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3790 = 10'h9d == _T_110[9:0] ? 4'ha : _GEN_3789; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3791 = 10'h9e == _T_110[9:0] ? 4'h3 : _GEN_3790; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3792 = 10'h9f == _T_110[9:0] ? 4'h0 : _GEN_3791; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3793 = 10'ha0 == _T_110[9:0] ? 4'ha : _GEN_3792; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3794 = 10'ha1 == _T_110[9:0] ? 4'h1 : _GEN_3793; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3795 = 10'ha2 == _T_110[9:0] ? 4'h0 : _GEN_3794; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3796 = 10'ha3 == _T_110[9:0] ? 4'h3 : _GEN_3795; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3797 = 10'ha4 == _T_110[9:0] ? 4'ha : _GEN_3796; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3798 = 10'ha5 == _T_110[9:0] ? 4'ha : _GEN_3797; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3799 = 10'ha6 == _T_110[9:0] ? 4'ha : _GEN_3798; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3800 = 10'ha7 == _T_110[9:0] ? 4'h0 : _GEN_3799; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3801 = 10'ha8 == _T_110[9:0] ? 4'ha : _GEN_3800; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3802 = 10'ha9 == _T_110[9:0] ? 4'h1 : _GEN_3801; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3803 = 10'haa == _T_110[9:0] ? 4'h0 : _GEN_3802; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3804 = 10'hab == _T_110[9:0] ? 4'h0 : _GEN_3803; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3805 = 10'hac == _T_110[9:0] ? 4'h0 : _GEN_3804; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3806 = 10'had == _T_110[9:0] ? 4'h0 : _GEN_3805; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3807 = 10'hae == _T_110[9:0] ? 4'h0 : _GEN_3806; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3808 = 10'haf == _T_110[9:0] ? 4'h0 : _GEN_3807; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3809 = 10'hb0 == _T_110[9:0] ? 4'h0 : _GEN_3808; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3810 = 10'hb1 == _T_110[9:0] ? 4'h0 : _GEN_3809; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3811 = 10'hb2 == _T_110[9:0] ? 4'h0 : _GEN_3810; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3812 = 10'hb3 == _T_110[9:0] ? 4'h0 : _GEN_3811; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3813 = 10'hb4 == _T_110[9:0] ? 4'h1 : _GEN_3812; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3814 = 10'hb5 == _T_110[9:0] ? 4'h1 : _GEN_3813; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3815 = 10'hb6 == _T_110[9:0] ? 4'ha : _GEN_3814; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3816 = 10'hb7 == _T_110[9:0] ? 4'h0 : _GEN_3815; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3817 = 10'hb8 == _T_110[9:0] ? 4'ha : _GEN_3816; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3818 = 10'hb9 == _T_110[9:0] ? 4'ha : _GEN_3817; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3819 = 10'hba == _T_110[9:0] ? 4'ha : _GEN_3818; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3820 = 10'hbb == _T_110[9:0] ? 4'h0 : _GEN_3819; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3821 = 10'hbc == _T_110[9:0] ? 4'ha : _GEN_3820; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3822 = 10'hbd == _T_110[9:0] ? 4'ha : _GEN_3821; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3823 = 10'hbe == _T_110[9:0] ? 4'h3 : _GEN_3822; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3824 = 10'hbf == _T_110[9:0] ? 4'h0 : _GEN_3823; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3825 = 10'hc0 == _T_110[9:0] ? 4'ha : _GEN_3824; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3826 = 10'hc1 == _T_110[9:0] ? 4'ha : _GEN_3825; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3827 = 10'hc2 == _T_110[9:0] ? 4'h3 : _GEN_3826; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3828 = 10'hc3 == _T_110[9:0] ? 4'h2 : _GEN_3827; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3829 = 10'hc4 == _T_110[9:0] ? 4'h0 : _GEN_3828; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3830 = 10'hc5 == _T_110[9:0] ? 4'h0 : _GEN_3829; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3831 = 10'hc6 == _T_110[9:0] ? 4'h0 : _GEN_3830; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3832 = 10'hc7 == _T_110[9:0] ? 4'ha : _GEN_3831; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3833 = 10'hc8 == _T_110[9:0] ? 4'h1 : _GEN_3832; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3834 = 10'hc9 == _T_110[9:0] ? 4'h0 : _GEN_3833; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3835 = 10'hca == _T_110[9:0] ? 4'h0 : _GEN_3834; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3836 = 10'hcb == _T_110[9:0] ? 4'h0 : _GEN_3835; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3837 = 10'hcc == _T_110[9:0] ? 4'h0 : _GEN_3836; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3838 = 10'hcd == _T_110[9:0] ? 4'h0 : _GEN_3837; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3839 = 10'hce == _T_110[9:0] ? 4'h0 : _GEN_3838; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3840 = 10'hcf == _T_110[9:0] ? 4'h0 : _GEN_3839; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3841 = 10'hd0 == _T_110[9:0] ? 4'h0 : _GEN_3840; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3842 = 10'hd1 == _T_110[9:0] ? 4'h0 : _GEN_3841; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3843 = 10'hd2 == _T_110[9:0] ? 4'h0 : _GEN_3842; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3844 = 10'hd3 == _T_110[9:0] ? 4'h0 : _GEN_3843; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3845 = 10'hd4 == _T_110[9:0] ? 4'h0 : _GEN_3844; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3846 = 10'hd5 == _T_110[9:0] ? 4'h0 : _GEN_3845; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3847 = 10'hd6 == _T_110[9:0] ? 4'h1 : _GEN_3846; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3848 = 10'hd7 == _T_110[9:0] ? 4'ha : _GEN_3847; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3849 = 10'hd8 == _T_110[9:0] ? 4'h0 : _GEN_3848; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3850 = 10'hd9 == _T_110[9:0] ? 4'ha : _GEN_3849; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3851 = 10'hda == _T_110[9:0] ? 4'ha : _GEN_3850; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3852 = 10'hdb == _T_110[9:0] ? 4'ha : _GEN_3851; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3853 = 10'hdc == _T_110[9:0] ? 4'ha : _GEN_3852; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3854 = 10'hdd == _T_110[9:0] ? 4'h3 : _GEN_3853; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3855 = 10'hde == _T_110[9:0] ? 4'h2 : _GEN_3854; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3856 = 10'hdf == _T_110[9:0] ? 4'h0 : _GEN_3855; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3857 = 10'he0 == _T_110[9:0] ? 4'ha : _GEN_3856; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3858 = 10'he1 == _T_110[9:0] ? 4'ha : _GEN_3857; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3859 = 10'he2 == _T_110[9:0] ? 4'h3 : _GEN_3858; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3860 = 10'he3 == _T_110[9:0] ? 4'ha : _GEN_3859; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3861 = 10'he4 == _T_110[9:0] ? 4'ha : _GEN_3860; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3862 = 10'he5 == _T_110[9:0] ? 4'ha : _GEN_3861; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3863 = 10'he6 == _T_110[9:0] ? 4'ha : _GEN_3862; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3864 = 10'he7 == _T_110[9:0] ? 4'h1 : _GEN_3863; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3865 = 10'he8 == _T_110[9:0] ? 4'h1 : _GEN_3864; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3866 = 10'he9 == _T_110[9:0] ? 4'h1 : _GEN_3865; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3867 = 10'hea == _T_110[9:0] ? 4'h0 : _GEN_3866; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3868 = 10'heb == _T_110[9:0] ? 4'h0 : _GEN_3867; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3869 = 10'hec == _T_110[9:0] ? 4'h0 : _GEN_3868; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3870 = 10'hed == _T_110[9:0] ? 4'h0 : _GEN_3869; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3871 = 10'hee == _T_110[9:0] ? 4'h0 : _GEN_3870; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3872 = 10'hef == _T_110[9:0] ? 4'h0 : _GEN_3871; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3873 = 10'hf0 == _T_110[9:0] ? 4'h0 : _GEN_3872; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3874 = 10'hf1 == _T_110[9:0] ? 4'h0 : _GEN_3873; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3875 = 10'hf2 == _T_110[9:0] ? 4'h0 : _GEN_3874; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3876 = 10'hf3 == _T_110[9:0] ? 4'h0 : _GEN_3875; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3877 = 10'hf4 == _T_110[9:0] ? 4'h0 : _GEN_3876; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3878 = 10'hf5 == _T_110[9:0] ? 4'h1 : _GEN_3877; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3879 = 10'hf6 == _T_110[9:0] ? 4'h0 : _GEN_3878; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3880 = 10'hf7 == _T_110[9:0] ? 4'h0 : _GEN_3879; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3881 = 10'hf8 == _T_110[9:0] ? 4'h1 : _GEN_3880; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3882 = 10'hf9 == _T_110[9:0] ? 4'h0 : _GEN_3881; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3883 = 10'hfa == _T_110[9:0] ? 4'ha : _GEN_3882; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3884 = 10'hfb == _T_110[9:0] ? 4'ha : _GEN_3883; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3885 = 10'hfc == _T_110[9:0] ? 4'ha : _GEN_3884; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3886 = 10'hfd == _T_110[9:0] ? 4'h3 : _GEN_3885; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3887 = 10'hfe == _T_110[9:0] ? 4'ha : _GEN_3886; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3888 = 10'hff == _T_110[9:0] ? 4'h0 : _GEN_3887; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3889 = 10'h100 == _T_110[9:0] ? 4'ha : _GEN_3888; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3890 = 10'h101 == _T_110[9:0] ? 4'h0 : _GEN_3889; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3891 = 10'h102 == _T_110[9:0] ? 4'h3 : _GEN_3890; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3892 = 10'h103 == _T_110[9:0] ? 4'ha : _GEN_3891; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3893 = 10'h104 == _T_110[9:0] ? 4'ha : _GEN_3892; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3894 = 10'h105 == _T_110[9:0] ? 4'ha : _GEN_3893; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3895 = 10'h106 == _T_110[9:0] ? 4'ha : _GEN_3894; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3896 = 10'h107 == _T_110[9:0] ? 4'ha : _GEN_3895; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3897 = 10'h108 == _T_110[9:0] ? 4'h1 : _GEN_3896; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3898 = 10'h109 == _T_110[9:0] ? 4'h0 : _GEN_3897; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3899 = 10'h10a == _T_110[9:0] ? 4'h0 : _GEN_3898; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3900 = 10'h10b == _T_110[9:0] ? 4'h0 : _GEN_3899; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3901 = 10'h10c == _T_110[9:0] ? 4'h0 : _GEN_3900; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3902 = 10'h10d == _T_110[9:0] ? 4'h0 : _GEN_3901; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3903 = 10'h10e == _T_110[9:0] ? 4'h0 : _GEN_3902; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3904 = 10'h10f == _T_110[9:0] ? 4'h0 : _GEN_3903; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3905 = 10'h110 == _T_110[9:0] ? 4'h0 : _GEN_3904; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3906 = 10'h111 == _T_110[9:0] ? 4'h0 : _GEN_3905; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3907 = 10'h112 == _T_110[9:0] ? 4'h0 : _GEN_3906; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3908 = 10'h113 == _T_110[9:0] ? 4'h0 : _GEN_3907; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3909 = 10'h114 == _T_110[9:0] ? 4'h0 : _GEN_3908; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3910 = 10'h115 == _T_110[9:0] ? 4'h0 : _GEN_3909; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3911 = 10'h116 == _T_110[9:0] ? 4'h1 : _GEN_3910; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3912 = 10'h117 == _T_110[9:0] ? 4'ha : _GEN_3911; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3913 = 10'h118 == _T_110[9:0] ? 4'ha : _GEN_3912; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3914 = 10'h119 == _T_110[9:0] ? 4'ha : _GEN_3913; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3915 = 10'h11a == _T_110[9:0] ? 4'h0 : _GEN_3914; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3916 = 10'h11b == _T_110[9:0] ? 4'ha : _GEN_3915; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3917 = 10'h11c == _T_110[9:0] ? 4'ha : _GEN_3916; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3918 = 10'h11d == _T_110[9:0] ? 4'h2 : _GEN_3917; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3919 = 10'h11e == _T_110[9:0] ? 4'h3 : _GEN_3918; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3920 = 10'h11f == _T_110[9:0] ? 4'h0 : _GEN_3919; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3921 = 10'h120 == _T_110[9:0] ? 4'ha : _GEN_3920; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3922 = 10'h121 == _T_110[9:0] ? 4'ha : _GEN_3921; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3923 = 10'h122 == _T_110[9:0] ? 4'h3 : _GEN_3922; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3924 = 10'h123 == _T_110[9:0] ? 4'ha : _GEN_3923; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3925 = 10'h124 == _T_110[9:0] ? 4'ha : _GEN_3924; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3926 = 10'h125 == _T_110[9:0] ? 4'ha : _GEN_3925; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3927 = 10'h126 == _T_110[9:0] ? 4'ha : _GEN_3926; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3928 = 10'h127 == _T_110[9:0] ? 4'h1 : _GEN_3927; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3929 = 10'h128 == _T_110[9:0] ? 4'h0 : _GEN_3928; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3930 = 10'h129 == _T_110[9:0] ? 4'ha : _GEN_3929; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3931 = 10'h12a == _T_110[9:0] ? 4'ha : _GEN_3930; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3932 = 10'h12b == _T_110[9:0] ? 4'h0 : _GEN_3931; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3933 = 10'h12c == _T_110[9:0] ? 4'h0 : _GEN_3932; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3934 = 10'h12d == _T_110[9:0] ? 4'h0 : _GEN_3933; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3935 = 10'h12e == _T_110[9:0] ? 4'h0 : _GEN_3934; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3936 = 10'h12f == _T_110[9:0] ? 4'h0 : _GEN_3935; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3937 = 10'h130 == _T_110[9:0] ? 4'h0 : _GEN_3936; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3938 = 10'h131 == _T_110[9:0] ? 4'h0 : _GEN_3937; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3939 = 10'h132 == _T_110[9:0] ? 4'h0 : _GEN_3938; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3940 = 10'h133 == _T_110[9:0] ? 4'h0 : _GEN_3939; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3941 = 10'h134 == _T_110[9:0] ? 4'ha : _GEN_3940; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3942 = 10'h135 == _T_110[9:0] ? 4'ha : _GEN_3941; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3943 = 10'h136 == _T_110[9:0] ? 4'h0 : _GEN_3942; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3944 = 10'h137 == _T_110[9:0] ? 4'h1 : _GEN_3943; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3945 = 10'h138 == _T_110[9:0] ? 4'ha : _GEN_3944; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3946 = 10'h139 == _T_110[9:0] ? 4'ha : _GEN_3945; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3947 = 10'h13a == _T_110[9:0] ? 4'ha : _GEN_3946; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3948 = 10'h13b == _T_110[9:0] ? 4'ha : _GEN_3947; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3949 = 10'h13c == _T_110[9:0] ? 4'ha : _GEN_3948; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3950 = 10'h13d == _T_110[9:0] ? 4'ha : _GEN_3949; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3951 = 10'h13e == _T_110[9:0] ? 4'h3 : _GEN_3950; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3952 = 10'h13f == _T_110[9:0] ? 4'h0 : _GEN_3951; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3953 = 10'h140 == _T_110[9:0] ? 4'ha : _GEN_3952; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3954 = 10'h141 == _T_110[9:0] ? 4'ha : _GEN_3953; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3955 = 10'h142 == _T_110[9:0] ? 4'h2 : _GEN_3954; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3956 = 10'h143 == _T_110[9:0] ? 4'h3 : _GEN_3955; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3957 = 10'h144 == _T_110[9:0] ? 4'ha : _GEN_3956; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3958 = 10'h145 == _T_110[9:0] ? 4'ha : _GEN_3957; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3959 = 10'h146 == _T_110[9:0] ? 4'h1 : _GEN_3958; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3960 = 10'h147 == _T_110[9:0] ? 4'h0 : _GEN_3959; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3961 = 10'h148 == _T_110[9:0] ? 4'ha : _GEN_3960; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3962 = 10'h149 == _T_110[9:0] ? 4'ha : _GEN_3961; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3963 = 10'h14a == _T_110[9:0] ? 4'ha : _GEN_3962; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3964 = 10'h14b == _T_110[9:0] ? 4'ha : _GEN_3963; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3965 = 10'h14c == _T_110[9:0] ? 4'ha : _GEN_3964; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3966 = 10'h14d == _T_110[9:0] ? 4'ha : _GEN_3965; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3967 = 10'h14e == _T_110[9:0] ? 4'ha : _GEN_3966; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3968 = 10'h14f == _T_110[9:0] ? 4'ha : _GEN_3967; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3969 = 10'h150 == _T_110[9:0] ? 4'ha : _GEN_3968; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3970 = 10'h151 == _T_110[9:0] ? 4'ha : _GEN_3969; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3971 = 10'h152 == _T_110[9:0] ? 4'ha : _GEN_3970; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3972 = 10'h153 == _T_110[9:0] ? 4'ha : _GEN_3971; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3973 = 10'h154 == _T_110[9:0] ? 4'ha : _GEN_3972; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3974 = 10'h155 == _T_110[9:0] ? 4'ha : _GEN_3973; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3975 = 10'h156 == _T_110[9:0] ? 4'ha : _GEN_3974; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3976 = 10'h157 == _T_110[9:0] ? 4'h0 : _GEN_3975; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3977 = 10'h158 == _T_110[9:0] ? 4'ha : _GEN_3976; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3978 = 10'h159 == _T_110[9:0] ? 4'ha : _GEN_3977; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3979 = 10'h15a == _T_110[9:0] ? 4'ha : _GEN_3978; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3980 = 10'h15b == _T_110[9:0] ? 4'ha : _GEN_3979; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3981 = 10'h15c == _T_110[9:0] ? 4'ha : _GEN_3980; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3982 = 10'h15d == _T_110[9:0] ? 4'h3 : _GEN_3981; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3983 = 10'h15e == _T_110[9:0] ? 4'h2 : _GEN_3982; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3984 = 10'h15f == _T_110[9:0] ? 4'h0 : _GEN_3983; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3985 = 10'h160 == _T_110[9:0] ? 4'ha : _GEN_3984; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3986 = 10'h161 == _T_110[9:0] ? 4'ha : _GEN_3985; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3987 = 10'h162 == _T_110[9:0] ? 4'ha : _GEN_3986; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3988 = 10'h163 == _T_110[9:0] ? 4'h2 : _GEN_3987; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3989 = 10'h164 == _T_110[9:0] ? 4'h3 : _GEN_3988; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3990 = 10'h165 == _T_110[9:0] ? 4'h1 : _GEN_3989; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3991 = 10'h166 == _T_110[9:0] ? 4'h0 : _GEN_3990; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3992 = 10'h167 == _T_110[9:0] ? 4'h0 : _GEN_3991; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3993 = 10'h168 == _T_110[9:0] ? 4'h5 : _GEN_3992; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3994 = 10'h169 == _T_110[9:0] ? 4'h3 : _GEN_3993; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3995 = 10'h16a == _T_110[9:0] ? 4'h5 : _GEN_3994; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3996 = 10'h16b == _T_110[9:0] ? 4'h5 : _GEN_3995; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3997 = 10'h16c == _T_110[9:0] ? 4'ha : _GEN_3996; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3998 = 10'h16d == _T_110[9:0] ? 4'ha : _GEN_3997; // @[Filter.scala 191:62]
  wire [3:0] _GEN_3999 = 10'h16e == _T_110[9:0] ? 4'ha : _GEN_3998; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4000 = 10'h16f == _T_110[9:0] ? 4'ha : _GEN_3999; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4001 = 10'h170 == _T_110[9:0] ? 4'ha : _GEN_4000; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4002 = 10'h171 == _T_110[9:0] ? 4'ha : _GEN_4001; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4003 = 10'h172 == _T_110[9:0] ? 4'ha : _GEN_4002; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4004 = 10'h173 == _T_110[9:0] ? 4'ha : _GEN_4003; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4005 = 10'h174 == _T_110[9:0] ? 4'ha : _GEN_4004; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4006 = 10'h175 == _T_110[9:0] ? 4'ha : _GEN_4005; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4007 = 10'h176 == _T_110[9:0] ? 4'h0 : _GEN_4006; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4008 = 10'h177 == _T_110[9:0] ? 4'h0 : _GEN_4007; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4009 = 10'h178 == _T_110[9:0] ? 4'h1 : _GEN_4008; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4010 = 10'h179 == _T_110[9:0] ? 4'ha : _GEN_4009; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4011 = 10'h17a == _T_110[9:0] ? 4'ha : _GEN_4010; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4012 = 10'h17b == _T_110[9:0] ? 4'ha : _GEN_4011; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4013 = 10'h17c == _T_110[9:0] ? 4'h3 : _GEN_4012; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4014 = 10'h17d == _T_110[9:0] ? 4'h2 : _GEN_4013; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4015 = 10'h17e == _T_110[9:0] ? 4'ha : _GEN_4014; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4016 = 10'h17f == _T_110[9:0] ? 4'h0 : _GEN_4015; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4017 = 10'h180 == _T_110[9:0] ? 4'h5 : _GEN_4016; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4018 = 10'h181 == _T_110[9:0] ? 4'h5 : _GEN_4017; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4019 = 10'h182 == _T_110[9:0] ? 4'h5 : _GEN_4018; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4020 = 10'h183 == _T_110[9:0] ? 4'h5 : _GEN_4019; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4021 = 10'h184 == _T_110[9:0] ? 4'h3 : _GEN_4020; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4022 = 10'h185 == _T_110[9:0] ? 4'h1 : _GEN_4021; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4023 = 10'h186 == _T_110[9:0] ? 4'hb : _GEN_4022; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4024 = 10'h187 == _T_110[9:0] ? 4'h0 : _GEN_4023; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4025 = 10'h188 == _T_110[9:0] ? 4'h5 : _GEN_4024; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4026 = 10'h189 == _T_110[9:0] ? 4'h5 : _GEN_4025; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4027 = 10'h18a == _T_110[9:0] ? 4'h5 : _GEN_4026; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4028 = 10'h18b == _T_110[9:0] ? 4'h5 : _GEN_4027; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4029 = 10'h18c == _T_110[9:0] ? 4'h5 : _GEN_4028; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4030 = 10'h18d == _T_110[9:0] ? 4'h5 : _GEN_4029; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4031 = 10'h18e == _T_110[9:0] ? 4'h5 : _GEN_4030; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4032 = 10'h18f == _T_110[9:0] ? 4'h5 : _GEN_4031; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4033 = 10'h190 == _T_110[9:0] ? 4'h5 : _GEN_4032; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4034 = 10'h191 == _T_110[9:0] ? 4'h5 : _GEN_4033; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4035 = 10'h192 == _T_110[9:0] ? 4'h3 : _GEN_4034; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4036 = 10'h193 == _T_110[9:0] ? 4'h5 : _GEN_4035; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4037 = 10'h194 == _T_110[9:0] ? 4'h5 : _GEN_4036; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4038 = 10'h195 == _T_110[9:0] ? 4'h5 : _GEN_4037; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4039 = 10'h196 == _T_110[9:0] ? 4'h0 : _GEN_4038; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4040 = 10'h197 == _T_110[9:0] ? 4'ha : _GEN_4039; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4041 = 10'h198 == _T_110[9:0] ? 4'h1 : _GEN_4040; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4042 = 10'h199 == _T_110[9:0] ? 4'ha : _GEN_4041; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4043 = 10'h19a == _T_110[9:0] ? 4'ha : _GEN_4042; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4044 = 10'h19b == _T_110[9:0] ? 4'ha : _GEN_4043; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4045 = 10'h19c == _T_110[9:0] ? 4'h3 : _GEN_4044; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4046 = 10'h19d == _T_110[9:0] ? 4'ha : _GEN_4045; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4047 = 10'h19e == _T_110[9:0] ? 4'ha : _GEN_4046; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4048 = 10'h19f == _T_110[9:0] ? 4'h0 : _GEN_4047; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4049 = 10'h1a0 == _T_110[9:0] ? 4'h5 : _GEN_4048; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4050 = 10'h1a1 == _T_110[9:0] ? 4'h5 : _GEN_4049; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4051 = 10'h1a2 == _T_110[9:0] ? 4'h3 : _GEN_4050; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4052 = 10'h1a3 == _T_110[9:0] ? 4'h5 : _GEN_4051; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4053 = 10'h1a4 == _T_110[9:0] ? 4'h3 : _GEN_4052; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4054 = 10'h1a5 == _T_110[9:0] ? 4'h0 : _GEN_4053; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4055 = 10'h1a6 == _T_110[9:0] ? 4'h5 : _GEN_4054; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4056 = 10'h1a7 == _T_110[9:0] ? 4'h0 : _GEN_4055; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4057 = 10'h1a8 == _T_110[9:0] ? 4'hb : _GEN_4056; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4058 = 10'h1a9 == _T_110[9:0] ? 4'h5 : _GEN_4057; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4059 = 10'h1aa == _T_110[9:0] ? 4'h5 : _GEN_4058; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4060 = 10'h1ab == _T_110[9:0] ? 4'h3 : _GEN_4059; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4061 = 10'h1ac == _T_110[9:0] ? 4'h5 : _GEN_4060; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4062 = 10'h1ad == _T_110[9:0] ? 4'h5 : _GEN_4061; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4063 = 10'h1ae == _T_110[9:0] ? 4'h5 : _GEN_4062; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4064 = 10'h1af == _T_110[9:0] ? 4'h5 : _GEN_4063; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4065 = 10'h1b0 == _T_110[9:0] ? 4'h5 : _GEN_4064; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4066 = 10'h1b1 == _T_110[9:0] ? 4'h5 : _GEN_4065; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4067 = 10'h1b2 == _T_110[9:0] ? 4'h5 : _GEN_4066; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4068 = 10'h1b3 == _T_110[9:0] ? 4'h5 : _GEN_4067; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4069 = 10'h1b4 == _T_110[9:0] ? 4'h5 : _GEN_4068; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4070 = 10'h1b5 == _T_110[9:0] ? 4'h5 : _GEN_4069; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4071 = 10'h1b6 == _T_110[9:0] ? 4'h0 : _GEN_4070; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4072 = 10'h1b7 == _T_110[9:0] ? 4'h5 : _GEN_4071; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4073 = 10'h1b8 == _T_110[9:0] ? 4'h0 : _GEN_4072; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4074 = 10'h1b9 == _T_110[9:0] ? 4'h5 : _GEN_4073; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4075 = 10'h1ba == _T_110[9:0] ? 4'h5 : _GEN_4074; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4076 = 10'h1bb == _T_110[9:0] ? 4'h5 : _GEN_4075; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4077 = 10'h1bc == _T_110[9:0] ? 4'h2 : _GEN_4076; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4078 = 10'h1bd == _T_110[9:0] ? 4'h3 : _GEN_4077; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4079 = 10'h1be == _T_110[9:0] ? 4'h5 : _GEN_4078; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4080 = 10'h1bf == _T_110[9:0] ? 4'h0 : _GEN_4079; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4081 = 10'h1c0 == _T_110[9:0] ? 4'h5 : _GEN_4080; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4082 = 10'h1c1 == _T_110[9:0] ? 4'h5 : _GEN_4081; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4083 = 10'h1c2 == _T_110[9:0] ? 4'h5 : _GEN_4082; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4084 = 10'h1c3 == _T_110[9:0] ? 4'h2 : _GEN_4083; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4085 = 10'h1c4 == _T_110[9:0] ? 4'h2 : _GEN_4084; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4086 = 10'h1c5 == _T_110[9:0] ? 4'h5 : _GEN_4085; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4087 = 10'h1c6 == _T_110[9:0] ? 4'h5 : _GEN_4086; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4088 = 10'h1c7 == _T_110[9:0] ? 4'h5 : _GEN_4087; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4089 = 10'h1c8 == _T_110[9:0] ? 4'h5 : _GEN_4088; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4090 = 10'h1c9 == _T_110[9:0] ? 4'hb : _GEN_4089; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4091 = 10'h1ca == _T_110[9:0] ? 4'hb : _GEN_4090; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4092 = 10'h1cb == _T_110[9:0] ? 4'hb : _GEN_4091; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4093 = 10'h1cc == _T_110[9:0] ? 4'hb : _GEN_4092; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4094 = 10'h1cd == _T_110[9:0] ? 4'hb : _GEN_4093; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4095 = 10'h1ce == _T_110[9:0] ? 4'hb : _GEN_4094; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4096 = 10'h1cf == _T_110[9:0] ? 4'hb : _GEN_4095; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4097 = 10'h1d0 == _T_110[9:0] ? 4'hb : _GEN_4096; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4098 = 10'h1d1 == _T_110[9:0] ? 4'hb : _GEN_4097; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4099 = 10'h1d2 == _T_110[9:0] ? 4'hb : _GEN_4098; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4100 = 10'h1d3 == _T_110[9:0] ? 4'hb : _GEN_4099; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4101 = 10'h1d4 == _T_110[9:0] ? 4'hb : _GEN_4100; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4102 = 10'h1d5 == _T_110[9:0] ? 4'hb : _GEN_4101; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4103 = 10'h1d6 == _T_110[9:0] ? 4'h5 : _GEN_4102; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4104 = 10'h1d7 == _T_110[9:0] ? 4'h5 : _GEN_4103; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4105 = 10'h1d8 == _T_110[9:0] ? 4'h5 : _GEN_4104; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4106 = 10'h1d9 == _T_110[9:0] ? 4'h5 : _GEN_4105; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4107 = 10'h1da == _T_110[9:0] ? 4'h5 : _GEN_4106; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4108 = 10'h1db == _T_110[9:0] ? 4'h5 : _GEN_4107; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4109 = 10'h1dc == _T_110[9:0] ? 4'h5 : _GEN_4108; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4110 = 10'h1dd == _T_110[9:0] ? 4'h3 : _GEN_4109; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4111 = 10'h1de == _T_110[9:0] ? 4'h5 : _GEN_4110; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4112 = 10'h1df == _T_110[9:0] ? 4'h0 : _GEN_4111; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4113 = 10'h1e0 == _T_110[9:0] ? 4'h3 : _GEN_4112; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4114 = 10'h1e1 == _T_110[9:0] ? 4'h5 : _GEN_4113; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4115 = 10'h1e2 == _T_110[9:0] ? 4'h2 : _GEN_4114; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4116 = 10'h1e3 == _T_110[9:0] ? 4'h2 : _GEN_4115; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4117 = 10'h1e4 == _T_110[9:0] ? 4'h5 : _GEN_4116; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4118 = 10'h1e5 == _T_110[9:0] ? 4'h5 : _GEN_4117; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4119 = 10'h1e6 == _T_110[9:0] ? 4'h5 : _GEN_4118; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4120 = 10'h1e7 == _T_110[9:0] ? 4'h5 : _GEN_4119; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4121 = 10'h1e8 == _T_110[9:0] ? 4'hb : _GEN_4120; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4122 = 10'h1e9 == _T_110[9:0] ? 4'h5 : _GEN_4121; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4123 = 10'h1ea == _T_110[9:0] ? 4'h5 : _GEN_4122; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4124 = 10'h1eb == _T_110[9:0] ? 4'hb : _GEN_4123; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4125 = 10'h1ec == _T_110[9:0] ? 4'h5 : _GEN_4124; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4126 = 10'h1ed == _T_110[9:0] ? 4'hb : _GEN_4125; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4127 = 10'h1ee == _T_110[9:0] ? 4'h5 : _GEN_4126; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4128 = 10'h1ef == _T_110[9:0] ? 4'hb : _GEN_4127; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4129 = 10'h1f0 == _T_110[9:0] ? 4'h5 : _GEN_4128; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4130 = 10'h1f1 == _T_110[9:0] ? 4'hb : _GEN_4129; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4131 = 10'h1f2 == _T_110[9:0] ? 4'hb : _GEN_4130; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4132 = 10'h1f3 == _T_110[9:0] ? 4'h5 : _GEN_4131; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4133 = 10'h1f4 == _T_110[9:0] ? 4'hb : _GEN_4132; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4134 = 10'h1f5 == _T_110[9:0] ? 4'hb : _GEN_4133; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4135 = 10'h1f6 == _T_110[9:0] ? 4'h5 : _GEN_4134; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4136 = 10'h1f7 == _T_110[9:0] ? 4'h5 : _GEN_4135; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4137 = 10'h1f8 == _T_110[9:0] ? 4'h5 : _GEN_4136; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4138 = 10'h1f9 == _T_110[9:0] ? 4'h5 : _GEN_4137; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4139 = 10'h1fa == _T_110[9:0] ? 4'h3 : _GEN_4138; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4140 = 10'h1fb == _T_110[9:0] ? 4'h5 : _GEN_4139; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4141 = 10'h1fc == _T_110[9:0] ? 4'h5 : _GEN_4140; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4142 = 10'h1fd == _T_110[9:0] ? 4'h2 : _GEN_4141; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4143 = 10'h1fe == _T_110[9:0] ? 4'h5 : _GEN_4142; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4144 = 10'h1ff == _T_110[9:0] ? 4'h0 : _GEN_4143; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4145 = 10'h200 == _T_110[9:0] ? 4'h5 : _GEN_4144; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4146 = 10'h201 == _T_110[9:0] ? 4'h5 : _GEN_4145; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4147 = 10'h202 == _T_110[9:0] ? 4'h3 : _GEN_4146; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4148 = 10'h203 == _T_110[9:0] ? 4'h5 : _GEN_4147; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4149 = 10'h204 == _T_110[9:0] ? 4'h5 : _GEN_4148; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4150 = 10'h205 == _T_110[9:0] ? 4'h5 : _GEN_4149; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4151 = 10'h206 == _T_110[9:0] ? 4'hb : _GEN_4150; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4152 = 10'h207 == _T_110[9:0] ? 4'hb : _GEN_4151; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4153 = 10'h208 == _T_110[9:0] ? 4'h5 : _GEN_4152; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4154 = 10'h209 == _T_110[9:0] ? 4'h5 : _GEN_4153; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4155 = 10'h20a == _T_110[9:0] ? 4'h5 : _GEN_4154; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4156 = 10'h20b == _T_110[9:0] ? 4'hb : _GEN_4155; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4157 = 10'h20c == _T_110[9:0] ? 4'h5 : _GEN_4156; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4158 = 10'h20d == _T_110[9:0] ? 4'hb : _GEN_4157; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4159 = 10'h20e == _T_110[9:0] ? 4'h5 : _GEN_4158; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4160 = 10'h20f == _T_110[9:0] ? 4'hb : _GEN_4159; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4161 = 10'h210 == _T_110[9:0] ? 4'h5 : _GEN_4160; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4162 = 10'h211 == _T_110[9:0] ? 4'h5 : _GEN_4161; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4163 = 10'h212 == _T_110[9:0] ? 4'hb : _GEN_4162; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4164 = 10'h213 == _T_110[9:0] ? 4'hb : _GEN_4163; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4165 = 10'h214 == _T_110[9:0] ? 4'hb : _GEN_4164; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4166 = 10'h215 == _T_110[9:0] ? 4'h5 : _GEN_4165; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4167 = 10'h216 == _T_110[9:0] ? 4'h5 : _GEN_4166; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4168 = 10'h217 == _T_110[9:0] ? 4'h5 : _GEN_4167; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4169 = 10'h218 == _T_110[9:0] ? 4'h5 : _GEN_4168; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4170 = 10'h219 == _T_110[9:0] ? 4'h5 : _GEN_4169; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4171 = 10'h21a == _T_110[9:0] ? 4'h5 : _GEN_4170; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4172 = 10'h21b == _T_110[9:0] ? 4'h5 : _GEN_4171; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4173 = 10'h21c == _T_110[9:0] ? 4'h3 : _GEN_4172; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4174 = 10'h21d == _T_110[9:0] ? 4'h2 : _GEN_4173; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4175 = 10'h21e == _T_110[9:0] ? 4'h5 : _GEN_4174; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4176 = 10'h21f == _T_110[9:0] ? 4'h0 : _GEN_4175; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4177 = 10'h220 == _T_110[9:0] ? 4'h0 : _GEN_4176; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4178 = 10'h221 == _T_110[9:0] ? 4'h0 : _GEN_4177; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4179 = 10'h222 == _T_110[9:0] ? 4'h0 : _GEN_4178; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4180 = 10'h223 == _T_110[9:0] ? 4'h0 : _GEN_4179; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4181 = 10'h224 == _T_110[9:0] ? 4'h0 : _GEN_4180; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4182 = 10'h225 == _T_110[9:0] ? 4'h0 : _GEN_4181; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4183 = 10'h226 == _T_110[9:0] ? 4'h0 : _GEN_4182; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4184 = 10'h227 == _T_110[9:0] ? 4'h0 : _GEN_4183; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4185 = 10'h228 == _T_110[9:0] ? 4'h0 : _GEN_4184; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4186 = 10'h229 == _T_110[9:0] ? 4'h0 : _GEN_4185; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4187 = 10'h22a == _T_110[9:0] ? 4'h0 : _GEN_4186; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4188 = 10'h22b == _T_110[9:0] ? 4'h0 : _GEN_4187; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4189 = 10'h22c == _T_110[9:0] ? 4'h0 : _GEN_4188; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4190 = 10'h22d == _T_110[9:0] ? 4'h0 : _GEN_4189; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4191 = 10'h22e == _T_110[9:0] ? 4'h0 : _GEN_4190; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4192 = 10'h22f == _T_110[9:0] ? 4'h0 : _GEN_4191; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4193 = 10'h230 == _T_110[9:0] ? 4'h0 : _GEN_4192; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4194 = 10'h231 == _T_110[9:0] ? 4'h0 : _GEN_4193; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4195 = 10'h232 == _T_110[9:0] ? 4'h0 : _GEN_4194; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4196 = 10'h233 == _T_110[9:0] ? 4'h0 : _GEN_4195; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4197 = 10'h234 == _T_110[9:0] ? 4'h0 : _GEN_4196; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4198 = 10'h235 == _T_110[9:0] ? 4'h0 : _GEN_4197; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4199 = 10'h236 == _T_110[9:0] ? 4'h0 : _GEN_4198; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4200 = 10'h237 == _T_110[9:0] ? 4'h0 : _GEN_4199; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4201 = 10'h238 == _T_110[9:0] ? 4'h0 : _GEN_4200; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4202 = 10'h239 == _T_110[9:0] ? 4'h0 : _GEN_4201; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4203 = 10'h23a == _T_110[9:0] ? 4'h0 : _GEN_4202; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4204 = 10'h23b == _T_110[9:0] ? 4'h0 : _GEN_4203; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4205 = 10'h23c == _T_110[9:0] ? 4'h0 : _GEN_4204; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4206 = 10'h23d == _T_110[9:0] ? 4'h0 : _GEN_4205; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4207 = 10'h23e == _T_110[9:0] ? 4'h0 : _GEN_4206; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4208 = 10'h23f == _T_110[9:0] ? 4'h0 : _GEN_4207; // @[Filter.scala 191:62]
  wire [4:0] _GEN_28310 = {{1'd0}, _GEN_4208}; // @[Filter.scala 191:62]
  wire [8:0] _T_112 = _GEN_28310 * 5'h14; // @[Filter.scala 191:62]
  wire [3:0] _GEN_4212 = 10'h3 == _T_110[9:0] ? 4'ha : 4'h3; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4213 = 10'h4 == _T_110[9:0] ? 4'h3 : _GEN_4212; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4214 = 10'h5 == _T_110[9:0] ? 4'h3 : _GEN_4213; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4215 = 10'h6 == _T_110[9:0] ? 4'h3 : _GEN_4214; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4216 = 10'h7 == _T_110[9:0] ? 4'h3 : _GEN_4215; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4217 = 10'h8 == _T_110[9:0] ? 4'h3 : _GEN_4216; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4218 = 10'h9 == _T_110[9:0] ? 4'h3 : _GEN_4217; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4219 = 10'ha == _T_110[9:0] ? 4'h3 : _GEN_4218; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4220 = 10'hb == _T_110[9:0] ? 4'h3 : _GEN_4219; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4221 = 10'hc == _T_110[9:0] ? 4'h5 : _GEN_4220; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4222 = 10'hd == _T_110[9:0] ? 4'h3 : _GEN_4221; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4223 = 10'he == _T_110[9:0] ? 4'h3 : _GEN_4222; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4224 = 10'hf == _T_110[9:0] ? 4'h3 : _GEN_4223; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4225 = 10'h10 == _T_110[9:0] ? 4'h3 : _GEN_4224; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4226 = 10'h11 == _T_110[9:0] ? 4'h3 : _GEN_4225; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4227 = 10'h12 == _T_110[9:0] ? 4'h3 : _GEN_4226; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4228 = 10'h13 == _T_110[9:0] ? 4'h3 : _GEN_4227; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4229 = 10'h14 == _T_110[9:0] ? 4'h3 : _GEN_4228; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4230 = 10'h15 == _T_110[9:0] ? 4'h3 : _GEN_4229; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4231 = 10'h16 == _T_110[9:0] ? 4'h3 : _GEN_4230; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4232 = 10'h17 == _T_110[9:0] ? 4'h3 : _GEN_4231; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4233 = 10'h18 == _T_110[9:0] ? 4'h3 : _GEN_4232; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4234 = 10'h19 == _T_110[9:0] ? 4'h3 : _GEN_4233; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4235 = 10'h1a == _T_110[9:0] ? 4'h3 : _GEN_4234; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4236 = 10'h1b == _T_110[9:0] ? 4'h3 : _GEN_4235; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4237 = 10'h1c == _T_110[9:0] ? 4'h3 : _GEN_4236; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4238 = 10'h1d == _T_110[9:0] ? 4'h3 : _GEN_4237; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4239 = 10'h1e == _T_110[9:0] ? 4'h3 : _GEN_4238; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4240 = 10'h1f == _T_110[9:0] ? 4'h0 : _GEN_4239; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4241 = 10'h20 == _T_110[9:0] ? 4'h3 : _GEN_4240; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4242 = 10'h21 == _T_110[9:0] ? 4'h5 : _GEN_4241; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4243 = 10'h22 == _T_110[9:0] ? 4'h3 : _GEN_4242; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4244 = 10'h23 == _T_110[9:0] ? 4'ha : _GEN_4243; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4245 = 10'h24 == _T_110[9:0] ? 4'h3 : _GEN_4244; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4246 = 10'h25 == _T_110[9:0] ? 4'h3 : _GEN_4245; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4247 = 10'h26 == _T_110[9:0] ? 4'h3 : _GEN_4246; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4248 = 10'h27 == _T_110[9:0] ? 4'h1 : _GEN_4247; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4249 = 10'h28 == _T_110[9:0] ? 4'h1 : _GEN_4248; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4250 = 10'h29 == _T_110[9:0] ? 4'h3 : _GEN_4249; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4251 = 10'h2a == _T_110[9:0] ? 4'h3 : _GEN_4250; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4252 = 10'h2b == _T_110[9:0] ? 4'h3 : _GEN_4251; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4253 = 10'h2c == _T_110[9:0] ? 4'h3 : _GEN_4252; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4254 = 10'h2d == _T_110[9:0] ? 4'h3 : _GEN_4253; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4255 = 10'h2e == _T_110[9:0] ? 4'h3 : _GEN_4254; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4256 = 10'h2f == _T_110[9:0] ? 4'h3 : _GEN_4255; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4257 = 10'h30 == _T_110[9:0] ? 4'h3 : _GEN_4256; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4258 = 10'h31 == _T_110[9:0] ? 4'h5 : _GEN_4257; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4259 = 10'h32 == _T_110[9:0] ? 4'h3 : _GEN_4258; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4260 = 10'h33 == _T_110[9:0] ? 4'h3 : _GEN_4259; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4261 = 10'h34 == _T_110[9:0] ? 4'h3 : _GEN_4260; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4262 = 10'h35 == _T_110[9:0] ? 4'h3 : _GEN_4261; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4263 = 10'h36 == _T_110[9:0] ? 4'h3 : _GEN_4262; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4264 = 10'h37 == _T_110[9:0] ? 4'h1 : _GEN_4263; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4265 = 10'h38 == _T_110[9:0] ? 4'h1 : _GEN_4264; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4266 = 10'h39 == _T_110[9:0] ? 4'h3 : _GEN_4265; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4267 = 10'h3a == _T_110[9:0] ? 4'h3 : _GEN_4266; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4268 = 10'h3b == _T_110[9:0] ? 4'h5 : _GEN_4267; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4269 = 10'h3c == _T_110[9:0] ? 4'h3 : _GEN_4268; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4270 = 10'h3d == _T_110[9:0] ? 4'ha : _GEN_4269; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4271 = 10'h3e == _T_110[9:0] ? 4'h3 : _GEN_4270; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4272 = 10'h3f == _T_110[9:0] ? 4'h0 : _GEN_4271; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4273 = 10'h40 == _T_110[9:0] ? 4'h3 : _GEN_4272; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4274 = 10'h41 == _T_110[9:0] ? 4'h3 : _GEN_4273; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4275 = 10'h42 == _T_110[9:0] ? 4'h3 : _GEN_4274; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4276 = 10'h43 == _T_110[9:0] ? 4'h7 : _GEN_4275; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4277 = 10'h44 == _T_110[9:0] ? 4'ha : _GEN_4276; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4278 = 10'h45 == _T_110[9:0] ? 4'h0 : _GEN_4277; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4279 = 10'h46 == _T_110[9:0] ? 4'h0 : _GEN_4278; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4280 = 10'h47 == _T_110[9:0] ? 4'h0 : _GEN_4279; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4281 = 10'h48 == _T_110[9:0] ? 4'h0 : _GEN_4280; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4282 = 10'h49 == _T_110[9:0] ? 4'h3 : _GEN_4281; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4283 = 10'h4a == _T_110[9:0] ? 4'h3 : _GEN_4282; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4284 = 10'h4b == _T_110[9:0] ? 4'h3 : _GEN_4283; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4285 = 10'h4c == _T_110[9:0] ? 4'h3 : _GEN_4284; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4286 = 10'h4d == _T_110[9:0] ? 4'h5 : _GEN_4285; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4287 = 10'h4e == _T_110[9:0] ? 4'h3 : _GEN_4286; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4288 = 10'h4f == _T_110[9:0] ? 4'h3 : _GEN_4287; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4289 = 10'h50 == _T_110[9:0] ? 4'h3 : _GEN_4288; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4290 = 10'h51 == _T_110[9:0] ? 4'h3 : _GEN_4289; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4291 = 10'h52 == _T_110[9:0] ? 4'h3 : _GEN_4290; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4292 = 10'h53 == _T_110[9:0] ? 4'h3 : _GEN_4291; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4293 = 10'h54 == _T_110[9:0] ? 4'h1 : _GEN_4292; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4294 = 10'h55 == _T_110[9:0] ? 4'h1 : _GEN_4293; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4295 = 10'h56 == _T_110[9:0] ? 4'h1 : _GEN_4294; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4296 = 10'h57 == _T_110[9:0] ? 4'h0 : _GEN_4295; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4297 = 10'h58 == _T_110[9:0] ? 4'h3 : _GEN_4296; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4298 = 10'h59 == _T_110[9:0] ? 4'h0 : _GEN_4297; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4299 = 10'h5a == _T_110[9:0] ? 4'h3 : _GEN_4298; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4300 = 10'h5b == _T_110[9:0] ? 4'h3 : _GEN_4299; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4301 = 10'h5c == _T_110[9:0] ? 4'h3 : _GEN_4300; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4302 = 10'h5d == _T_110[9:0] ? 4'ha : _GEN_4301; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4303 = 10'h5e == _T_110[9:0] ? 4'h3 : _GEN_4302; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4304 = 10'h5f == _T_110[9:0] ? 4'h0 : _GEN_4303; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4305 = 10'h60 == _T_110[9:0] ? 4'h3 : _GEN_4304; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4306 = 10'h61 == _T_110[9:0] ? 4'h3 : _GEN_4305; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4307 = 10'h62 == _T_110[9:0] ? 4'h3 : _GEN_4306; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4308 = 10'h63 == _T_110[9:0] ? 4'h3 : _GEN_4307; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4309 = 10'h64 == _T_110[9:0] ? 4'ha : _GEN_4308; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4310 = 10'h65 == _T_110[9:0] ? 4'h0 : _GEN_4309; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4311 = 10'h66 == _T_110[9:0] ? 4'h3 : _GEN_4310; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4312 = 10'h67 == _T_110[9:0] ? 4'h3 : _GEN_4311; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4313 = 10'h68 == _T_110[9:0] ? 4'h3 : _GEN_4312; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4314 = 10'h69 == _T_110[9:0] ? 4'h0 : _GEN_4313; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4315 = 10'h6a == _T_110[9:0] ? 4'h1 : _GEN_4314; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4316 = 10'h6b == _T_110[9:0] ? 4'h1 : _GEN_4315; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4317 = 10'h6c == _T_110[9:0] ? 4'h3 : _GEN_4316; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4318 = 10'h6d == _T_110[9:0] ? 4'h3 : _GEN_4317; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4319 = 10'h6e == _T_110[9:0] ? 4'h3 : _GEN_4318; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4320 = 10'h6f == _T_110[9:0] ? 4'h3 : _GEN_4319; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4321 = 10'h70 == _T_110[9:0] ? 4'h3 : _GEN_4320; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4322 = 10'h71 == _T_110[9:0] ? 4'h3 : _GEN_4321; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4323 = 10'h72 == _T_110[9:0] ? 4'h3 : _GEN_4322; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4324 = 10'h73 == _T_110[9:0] ? 4'h1 : _GEN_4323; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4325 = 10'h74 == _T_110[9:0] ? 4'h0 : _GEN_4324; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4326 = 10'h75 == _T_110[9:0] ? 4'h0 : _GEN_4325; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4327 = 10'h76 == _T_110[9:0] ? 4'h0 : _GEN_4326; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4328 = 10'h77 == _T_110[9:0] ? 4'h3 : _GEN_4327; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4329 = 10'h78 == _T_110[9:0] ? 4'h3 : _GEN_4328; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4330 = 10'h79 == _T_110[9:0] ? 4'h3 : _GEN_4329; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4331 = 10'h7a == _T_110[9:0] ? 4'h0 : _GEN_4330; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4332 = 10'h7b == _T_110[9:0] ? 4'h3 : _GEN_4331; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4333 = 10'h7c == _T_110[9:0] ? 4'h3 : _GEN_4332; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4334 = 10'h7d == _T_110[9:0] ? 4'h7 : _GEN_4333; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4335 = 10'h7e == _T_110[9:0] ? 4'ha : _GEN_4334; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4336 = 10'h7f == _T_110[9:0] ? 4'h0 : _GEN_4335; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4337 = 10'h80 == _T_110[9:0] ? 4'h3 : _GEN_4336; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4338 = 10'h81 == _T_110[9:0] ? 4'h3 : _GEN_4337; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4339 = 10'h82 == _T_110[9:0] ? 4'h1 : _GEN_4338; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4340 = 10'h83 == _T_110[9:0] ? 4'h0 : _GEN_4339; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4341 = 10'h84 == _T_110[9:0] ? 4'h7 : _GEN_4340; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4342 = 10'h85 == _T_110[9:0] ? 4'h1 : _GEN_4341; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4343 = 10'h86 == _T_110[9:0] ? 4'h1 : _GEN_4342; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4344 = 10'h87 == _T_110[9:0] ? 4'h3 : _GEN_4343; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4345 = 10'h88 == _T_110[9:0] ? 4'h3 : _GEN_4344; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4346 = 10'h89 == _T_110[9:0] ? 4'h0 : _GEN_4345; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4347 = 10'h8a == _T_110[9:0] ? 4'h0 : _GEN_4346; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4348 = 10'h8b == _T_110[9:0] ? 4'h1 : _GEN_4347; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4349 = 10'h8c == _T_110[9:0] ? 4'h1 : _GEN_4348; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4350 = 10'h8d == _T_110[9:0] ? 4'h1 : _GEN_4349; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4351 = 10'h8e == _T_110[9:0] ? 4'h1 : _GEN_4350; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4352 = 10'h8f == _T_110[9:0] ? 4'h1 : _GEN_4351; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4353 = 10'h90 == _T_110[9:0] ? 4'h1 : _GEN_4352; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4354 = 10'h91 == _T_110[9:0] ? 4'h1 : _GEN_4353; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4355 = 10'h92 == _T_110[9:0] ? 4'h1 : _GEN_4354; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4356 = 10'h93 == _T_110[9:0] ? 4'h0 : _GEN_4355; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4357 = 10'h94 == _T_110[9:0] ? 4'h0 : _GEN_4356; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4358 = 10'h95 == _T_110[9:0] ? 4'h3 : _GEN_4357; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4359 = 10'h96 == _T_110[9:0] ? 4'h3 : _GEN_4358; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4360 = 10'h97 == _T_110[9:0] ? 4'h3 : _GEN_4359; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4361 = 10'h98 == _T_110[9:0] ? 4'h1 : _GEN_4360; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4362 = 10'h99 == _T_110[9:0] ? 4'h0 : _GEN_4361; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4363 = 10'h9a == _T_110[9:0] ? 4'h1 : _GEN_4362; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4364 = 10'h9b == _T_110[9:0] ? 4'h1 : _GEN_4363; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4365 = 10'h9c == _T_110[9:0] ? 4'h3 : _GEN_4364; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4366 = 10'h9d == _T_110[9:0] ? 4'h3 : _GEN_4365; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4367 = 10'h9e == _T_110[9:0] ? 4'ha : _GEN_4366; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4368 = 10'h9f == _T_110[9:0] ? 4'h0 : _GEN_4367; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4369 = 10'ha0 == _T_110[9:0] ? 4'h3 : _GEN_4368; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4370 = 10'ha1 == _T_110[9:0] ? 4'h1 : _GEN_4369; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4371 = 10'ha2 == _T_110[9:0] ? 4'h0 : _GEN_4370; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4372 = 10'ha3 == _T_110[9:0] ? 4'ha : _GEN_4371; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4373 = 10'ha4 == _T_110[9:0] ? 4'h3 : _GEN_4372; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4374 = 10'ha5 == _T_110[9:0] ? 4'h3 : _GEN_4373; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4375 = 10'ha6 == _T_110[9:0] ? 4'h3 : _GEN_4374; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4376 = 10'ha7 == _T_110[9:0] ? 4'h0 : _GEN_4375; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4377 = 10'ha8 == _T_110[9:0] ? 4'h3 : _GEN_4376; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4378 = 10'ha9 == _T_110[9:0] ? 4'h1 : _GEN_4377; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4379 = 10'haa == _T_110[9:0] ? 4'h0 : _GEN_4378; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4380 = 10'hab == _T_110[9:0] ? 4'h0 : _GEN_4379; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4381 = 10'hac == _T_110[9:0] ? 4'h0 : _GEN_4380; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4382 = 10'had == _T_110[9:0] ? 4'h0 : _GEN_4381; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4383 = 10'hae == _T_110[9:0] ? 4'h0 : _GEN_4382; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4384 = 10'haf == _T_110[9:0] ? 4'h0 : _GEN_4383; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4385 = 10'hb0 == _T_110[9:0] ? 4'h0 : _GEN_4384; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4386 = 10'hb1 == _T_110[9:0] ? 4'h0 : _GEN_4385; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4387 = 10'hb2 == _T_110[9:0] ? 4'h0 : _GEN_4386; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4388 = 10'hb3 == _T_110[9:0] ? 4'h0 : _GEN_4387; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4389 = 10'hb4 == _T_110[9:0] ? 4'h1 : _GEN_4388; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4390 = 10'hb5 == _T_110[9:0] ? 4'h1 : _GEN_4389; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4391 = 10'hb6 == _T_110[9:0] ? 4'h3 : _GEN_4390; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4392 = 10'hb7 == _T_110[9:0] ? 4'h0 : _GEN_4391; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4393 = 10'hb8 == _T_110[9:0] ? 4'h3 : _GEN_4392; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4394 = 10'hb9 == _T_110[9:0] ? 4'h3 : _GEN_4393; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4395 = 10'hba == _T_110[9:0] ? 4'h3 : _GEN_4394; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4396 = 10'hbb == _T_110[9:0] ? 4'h0 : _GEN_4395; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4397 = 10'hbc == _T_110[9:0] ? 4'h3 : _GEN_4396; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4398 = 10'hbd == _T_110[9:0] ? 4'h3 : _GEN_4397; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4399 = 10'hbe == _T_110[9:0] ? 4'ha : _GEN_4398; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4400 = 10'hbf == _T_110[9:0] ? 4'h0 : _GEN_4399; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4401 = 10'hc0 == _T_110[9:0] ? 4'h3 : _GEN_4400; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4402 = 10'hc1 == _T_110[9:0] ? 4'h3 : _GEN_4401; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4403 = 10'hc2 == _T_110[9:0] ? 4'ha : _GEN_4402; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4404 = 10'hc3 == _T_110[9:0] ? 4'h7 : _GEN_4403; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4405 = 10'hc4 == _T_110[9:0] ? 4'h0 : _GEN_4404; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4406 = 10'hc5 == _T_110[9:0] ? 4'h0 : _GEN_4405; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4407 = 10'hc6 == _T_110[9:0] ? 4'h0 : _GEN_4406; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4408 = 10'hc7 == _T_110[9:0] ? 4'h3 : _GEN_4407; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4409 = 10'hc8 == _T_110[9:0] ? 4'h1 : _GEN_4408; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4410 = 10'hc9 == _T_110[9:0] ? 4'h0 : _GEN_4409; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4411 = 10'hca == _T_110[9:0] ? 4'h0 : _GEN_4410; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4412 = 10'hcb == _T_110[9:0] ? 4'h0 : _GEN_4411; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4413 = 10'hcc == _T_110[9:0] ? 4'h0 : _GEN_4412; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4414 = 10'hcd == _T_110[9:0] ? 4'h0 : _GEN_4413; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4415 = 10'hce == _T_110[9:0] ? 4'h0 : _GEN_4414; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4416 = 10'hcf == _T_110[9:0] ? 4'h0 : _GEN_4415; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4417 = 10'hd0 == _T_110[9:0] ? 4'h0 : _GEN_4416; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4418 = 10'hd1 == _T_110[9:0] ? 4'h0 : _GEN_4417; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4419 = 10'hd2 == _T_110[9:0] ? 4'h0 : _GEN_4418; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4420 = 10'hd3 == _T_110[9:0] ? 4'h0 : _GEN_4419; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4421 = 10'hd4 == _T_110[9:0] ? 4'h0 : _GEN_4420; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4422 = 10'hd5 == _T_110[9:0] ? 4'h0 : _GEN_4421; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4423 = 10'hd6 == _T_110[9:0] ? 4'h1 : _GEN_4422; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4424 = 10'hd7 == _T_110[9:0] ? 4'h3 : _GEN_4423; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4425 = 10'hd8 == _T_110[9:0] ? 4'h0 : _GEN_4424; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4426 = 10'hd9 == _T_110[9:0] ? 4'h3 : _GEN_4425; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4427 = 10'hda == _T_110[9:0] ? 4'h3 : _GEN_4426; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4428 = 10'hdb == _T_110[9:0] ? 4'h3 : _GEN_4427; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4429 = 10'hdc == _T_110[9:0] ? 4'h3 : _GEN_4428; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4430 = 10'hdd == _T_110[9:0] ? 4'ha : _GEN_4429; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4431 = 10'hde == _T_110[9:0] ? 4'h7 : _GEN_4430; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4432 = 10'hdf == _T_110[9:0] ? 4'h0 : _GEN_4431; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4433 = 10'he0 == _T_110[9:0] ? 4'h3 : _GEN_4432; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4434 = 10'he1 == _T_110[9:0] ? 4'h3 : _GEN_4433; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4435 = 10'he2 == _T_110[9:0] ? 4'ha : _GEN_4434; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4436 = 10'he3 == _T_110[9:0] ? 4'h3 : _GEN_4435; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4437 = 10'he4 == _T_110[9:0] ? 4'h3 : _GEN_4436; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4438 = 10'he5 == _T_110[9:0] ? 4'h3 : _GEN_4437; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4439 = 10'he6 == _T_110[9:0] ? 4'h3 : _GEN_4438; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4440 = 10'he7 == _T_110[9:0] ? 4'h1 : _GEN_4439; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4441 = 10'he8 == _T_110[9:0] ? 4'h1 : _GEN_4440; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4442 = 10'he9 == _T_110[9:0] ? 4'h1 : _GEN_4441; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4443 = 10'hea == _T_110[9:0] ? 4'h0 : _GEN_4442; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4444 = 10'heb == _T_110[9:0] ? 4'h0 : _GEN_4443; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4445 = 10'hec == _T_110[9:0] ? 4'h0 : _GEN_4444; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4446 = 10'hed == _T_110[9:0] ? 4'h0 : _GEN_4445; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4447 = 10'hee == _T_110[9:0] ? 4'h0 : _GEN_4446; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4448 = 10'hef == _T_110[9:0] ? 4'h0 : _GEN_4447; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4449 = 10'hf0 == _T_110[9:0] ? 4'h0 : _GEN_4448; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4450 = 10'hf1 == _T_110[9:0] ? 4'h0 : _GEN_4449; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4451 = 10'hf2 == _T_110[9:0] ? 4'h0 : _GEN_4450; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4452 = 10'hf3 == _T_110[9:0] ? 4'h0 : _GEN_4451; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4453 = 10'hf4 == _T_110[9:0] ? 4'h0 : _GEN_4452; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4454 = 10'hf5 == _T_110[9:0] ? 4'h1 : _GEN_4453; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4455 = 10'hf6 == _T_110[9:0] ? 4'h0 : _GEN_4454; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4456 = 10'hf7 == _T_110[9:0] ? 4'h0 : _GEN_4455; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4457 = 10'hf8 == _T_110[9:0] ? 4'h1 : _GEN_4456; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4458 = 10'hf9 == _T_110[9:0] ? 4'h0 : _GEN_4457; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4459 = 10'hfa == _T_110[9:0] ? 4'h3 : _GEN_4458; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4460 = 10'hfb == _T_110[9:0] ? 4'h3 : _GEN_4459; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4461 = 10'hfc == _T_110[9:0] ? 4'h3 : _GEN_4460; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4462 = 10'hfd == _T_110[9:0] ? 4'ha : _GEN_4461; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4463 = 10'hfe == _T_110[9:0] ? 4'h3 : _GEN_4462; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4464 = 10'hff == _T_110[9:0] ? 4'h0 : _GEN_4463; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4465 = 10'h100 == _T_110[9:0] ? 4'h3 : _GEN_4464; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4466 = 10'h101 == _T_110[9:0] ? 4'h0 : _GEN_4465; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4467 = 10'h102 == _T_110[9:0] ? 4'ha : _GEN_4466; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4468 = 10'h103 == _T_110[9:0] ? 4'h3 : _GEN_4467; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4469 = 10'h104 == _T_110[9:0] ? 4'h3 : _GEN_4468; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4470 = 10'h105 == _T_110[9:0] ? 4'h3 : _GEN_4469; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4471 = 10'h106 == _T_110[9:0] ? 4'h3 : _GEN_4470; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4472 = 10'h107 == _T_110[9:0] ? 4'h3 : _GEN_4471; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4473 = 10'h108 == _T_110[9:0] ? 4'h1 : _GEN_4472; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4474 = 10'h109 == _T_110[9:0] ? 4'h0 : _GEN_4473; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4475 = 10'h10a == _T_110[9:0] ? 4'h0 : _GEN_4474; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4476 = 10'h10b == _T_110[9:0] ? 4'h0 : _GEN_4475; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4477 = 10'h10c == _T_110[9:0] ? 4'h0 : _GEN_4476; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4478 = 10'h10d == _T_110[9:0] ? 4'h0 : _GEN_4477; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4479 = 10'h10e == _T_110[9:0] ? 4'h0 : _GEN_4478; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4480 = 10'h10f == _T_110[9:0] ? 4'h0 : _GEN_4479; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4481 = 10'h110 == _T_110[9:0] ? 4'h0 : _GEN_4480; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4482 = 10'h111 == _T_110[9:0] ? 4'h0 : _GEN_4481; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4483 = 10'h112 == _T_110[9:0] ? 4'h0 : _GEN_4482; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4484 = 10'h113 == _T_110[9:0] ? 4'h0 : _GEN_4483; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4485 = 10'h114 == _T_110[9:0] ? 4'h0 : _GEN_4484; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4486 = 10'h115 == _T_110[9:0] ? 4'h0 : _GEN_4485; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4487 = 10'h116 == _T_110[9:0] ? 4'h1 : _GEN_4486; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4488 = 10'h117 == _T_110[9:0] ? 4'h3 : _GEN_4487; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4489 = 10'h118 == _T_110[9:0] ? 4'h3 : _GEN_4488; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4490 = 10'h119 == _T_110[9:0] ? 4'h3 : _GEN_4489; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4491 = 10'h11a == _T_110[9:0] ? 4'h0 : _GEN_4490; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4492 = 10'h11b == _T_110[9:0] ? 4'h3 : _GEN_4491; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4493 = 10'h11c == _T_110[9:0] ? 4'h3 : _GEN_4492; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4494 = 10'h11d == _T_110[9:0] ? 4'h7 : _GEN_4493; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4495 = 10'h11e == _T_110[9:0] ? 4'ha : _GEN_4494; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4496 = 10'h11f == _T_110[9:0] ? 4'h0 : _GEN_4495; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4497 = 10'h120 == _T_110[9:0] ? 4'h3 : _GEN_4496; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4498 = 10'h121 == _T_110[9:0] ? 4'h3 : _GEN_4497; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4499 = 10'h122 == _T_110[9:0] ? 4'ha : _GEN_4498; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4500 = 10'h123 == _T_110[9:0] ? 4'h3 : _GEN_4499; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4501 = 10'h124 == _T_110[9:0] ? 4'h3 : _GEN_4500; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4502 = 10'h125 == _T_110[9:0] ? 4'h3 : _GEN_4501; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4503 = 10'h126 == _T_110[9:0] ? 4'h3 : _GEN_4502; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4504 = 10'h127 == _T_110[9:0] ? 4'h1 : _GEN_4503; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4505 = 10'h128 == _T_110[9:0] ? 4'h0 : _GEN_4504; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4506 = 10'h129 == _T_110[9:0] ? 4'h3 : _GEN_4505; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4507 = 10'h12a == _T_110[9:0] ? 4'h3 : _GEN_4506; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4508 = 10'h12b == _T_110[9:0] ? 4'h0 : _GEN_4507; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4509 = 10'h12c == _T_110[9:0] ? 4'h0 : _GEN_4508; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4510 = 10'h12d == _T_110[9:0] ? 4'h0 : _GEN_4509; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4511 = 10'h12e == _T_110[9:0] ? 4'h0 : _GEN_4510; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4512 = 10'h12f == _T_110[9:0] ? 4'h0 : _GEN_4511; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4513 = 10'h130 == _T_110[9:0] ? 4'h0 : _GEN_4512; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4514 = 10'h131 == _T_110[9:0] ? 4'h0 : _GEN_4513; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4515 = 10'h132 == _T_110[9:0] ? 4'h0 : _GEN_4514; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4516 = 10'h133 == _T_110[9:0] ? 4'h0 : _GEN_4515; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4517 = 10'h134 == _T_110[9:0] ? 4'h3 : _GEN_4516; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4518 = 10'h135 == _T_110[9:0] ? 4'h3 : _GEN_4517; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4519 = 10'h136 == _T_110[9:0] ? 4'h0 : _GEN_4518; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4520 = 10'h137 == _T_110[9:0] ? 4'h1 : _GEN_4519; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4521 = 10'h138 == _T_110[9:0] ? 4'h3 : _GEN_4520; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4522 = 10'h139 == _T_110[9:0] ? 4'h3 : _GEN_4521; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4523 = 10'h13a == _T_110[9:0] ? 4'h3 : _GEN_4522; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4524 = 10'h13b == _T_110[9:0] ? 4'h3 : _GEN_4523; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4525 = 10'h13c == _T_110[9:0] ? 4'h3 : _GEN_4524; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4526 = 10'h13d == _T_110[9:0] ? 4'h3 : _GEN_4525; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4527 = 10'h13e == _T_110[9:0] ? 4'ha : _GEN_4526; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4528 = 10'h13f == _T_110[9:0] ? 4'h0 : _GEN_4527; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4529 = 10'h140 == _T_110[9:0] ? 4'h5 : _GEN_4528; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4530 = 10'h141 == _T_110[9:0] ? 4'h3 : _GEN_4529; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4531 = 10'h142 == _T_110[9:0] ? 4'h7 : _GEN_4530; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4532 = 10'h143 == _T_110[9:0] ? 4'ha : _GEN_4531; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4533 = 10'h144 == _T_110[9:0] ? 4'h3 : _GEN_4532; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4534 = 10'h145 == _T_110[9:0] ? 4'h3 : _GEN_4533; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4535 = 10'h146 == _T_110[9:0] ? 4'h1 : _GEN_4534; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4536 = 10'h147 == _T_110[9:0] ? 4'h0 : _GEN_4535; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4537 = 10'h148 == _T_110[9:0] ? 4'h3 : _GEN_4536; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4538 = 10'h149 == _T_110[9:0] ? 4'h3 : _GEN_4537; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4539 = 10'h14a == _T_110[9:0] ? 4'h3 : _GEN_4538; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4540 = 10'h14b == _T_110[9:0] ? 4'h3 : _GEN_4539; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4541 = 10'h14c == _T_110[9:0] ? 4'h3 : _GEN_4540; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4542 = 10'h14d == _T_110[9:0] ? 4'h3 : _GEN_4541; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4543 = 10'h14e == _T_110[9:0] ? 4'h3 : _GEN_4542; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4544 = 10'h14f == _T_110[9:0] ? 4'h3 : _GEN_4543; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4545 = 10'h150 == _T_110[9:0] ? 4'h3 : _GEN_4544; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4546 = 10'h151 == _T_110[9:0] ? 4'h3 : _GEN_4545; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4547 = 10'h152 == _T_110[9:0] ? 4'h3 : _GEN_4546; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4548 = 10'h153 == _T_110[9:0] ? 4'h3 : _GEN_4547; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4549 = 10'h154 == _T_110[9:0] ? 4'h3 : _GEN_4548; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4550 = 10'h155 == _T_110[9:0] ? 4'h3 : _GEN_4549; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4551 = 10'h156 == _T_110[9:0] ? 4'h3 : _GEN_4550; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4552 = 10'h157 == _T_110[9:0] ? 4'h0 : _GEN_4551; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4553 = 10'h158 == _T_110[9:0] ? 4'h3 : _GEN_4552; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4554 = 10'h159 == _T_110[9:0] ? 4'h3 : _GEN_4553; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4555 = 10'h15a == _T_110[9:0] ? 4'h3 : _GEN_4554; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4556 = 10'h15b == _T_110[9:0] ? 4'h3 : _GEN_4555; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4557 = 10'h15c == _T_110[9:0] ? 4'h3 : _GEN_4556; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4558 = 10'h15d == _T_110[9:0] ? 4'ha : _GEN_4557; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4559 = 10'h15e == _T_110[9:0] ? 4'h7 : _GEN_4558; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4560 = 10'h15f == _T_110[9:0] ? 4'h0 : _GEN_4559; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4561 = 10'h160 == _T_110[9:0] ? 4'h3 : _GEN_4560; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4562 = 10'h161 == _T_110[9:0] ? 4'h3 : _GEN_4561; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4563 = 10'h162 == _T_110[9:0] ? 4'h3 : _GEN_4562; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4564 = 10'h163 == _T_110[9:0] ? 4'h7 : _GEN_4563; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4565 = 10'h164 == _T_110[9:0] ? 4'ha : _GEN_4564; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4566 = 10'h165 == _T_110[9:0] ? 4'h1 : _GEN_4565; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4567 = 10'h166 == _T_110[9:0] ? 4'h0 : _GEN_4566; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4568 = 10'h167 == _T_110[9:0] ? 4'h0 : _GEN_4567; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4569 = 10'h168 == _T_110[9:0] ? 4'hc : _GEN_4568; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4570 = 10'h169 == _T_110[9:0] ? 4'h9 : _GEN_4569; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4571 = 10'h16a == _T_110[9:0] ? 4'hc : _GEN_4570; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4572 = 10'h16b == _T_110[9:0] ? 4'hc : _GEN_4571; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4573 = 10'h16c == _T_110[9:0] ? 4'h3 : _GEN_4572; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4574 = 10'h16d == _T_110[9:0] ? 4'h3 : _GEN_4573; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4575 = 10'h16e == _T_110[9:0] ? 4'h3 : _GEN_4574; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4576 = 10'h16f == _T_110[9:0] ? 4'h3 : _GEN_4575; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4577 = 10'h170 == _T_110[9:0] ? 4'h5 : _GEN_4576; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4578 = 10'h171 == _T_110[9:0] ? 4'h3 : _GEN_4577; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4579 = 10'h172 == _T_110[9:0] ? 4'h3 : _GEN_4578; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4580 = 10'h173 == _T_110[9:0] ? 4'h3 : _GEN_4579; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4581 = 10'h174 == _T_110[9:0] ? 4'h3 : _GEN_4580; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4582 = 10'h175 == _T_110[9:0] ? 4'h3 : _GEN_4581; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4583 = 10'h176 == _T_110[9:0] ? 4'h0 : _GEN_4582; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4584 = 10'h177 == _T_110[9:0] ? 4'h0 : _GEN_4583; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4585 = 10'h178 == _T_110[9:0] ? 4'h1 : _GEN_4584; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4586 = 10'h179 == _T_110[9:0] ? 4'h3 : _GEN_4585; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4587 = 10'h17a == _T_110[9:0] ? 4'h5 : _GEN_4586; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4588 = 10'h17b == _T_110[9:0] ? 4'h3 : _GEN_4587; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4589 = 10'h17c == _T_110[9:0] ? 4'ha : _GEN_4588; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4590 = 10'h17d == _T_110[9:0] ? 4'h7 : _GEN_4589; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4591 = 10'h17e == _T_110[9:0] ? 4'h3 : _GEN_4590; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4592 = 10'h17f == _T_110[9:0] ? 4'h0 : _GEN_4591; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4593 = 10'h180 == _T_110[9:0] ? 4'hc : _GEN_4592; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4594 = 10'h181 == _T_110[9:0] ? 4'hc : _GEN_4593; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4595 = 10'h182 == _T_110[9:0] ? 4'hc : _GEN_4594; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4596 = 10'h183 == _T_110[9:0] ? 4'hc : _GEN_4595; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4597 = 10'h184 == _T_110[9:0] ? 4'ha : _GEN_4596; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4598 = 10'h185 == _T_110[9:0] ? 4'h1 : _GEN_4597; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4599 = 10'h186 == _T_110[9:0] ? 4'hc : _GEN_4598; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4600 = 10'h187 == _T_110[9:0] ? 4'h0 : _GEN_4599; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4601 = 10'h188 == _T_110[9:0] ? 4'hc : _GEN_4600; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4602 = 10'h189 == _T_110[9:0] ? 4'hc : _GEN_4601; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4603 = 10'h18a == _T_110[9:0] ? 4'hc : _GEN_4602; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4604 = 10'h18b == _T_110[9:0] ? 4'hc : _GEN_4603; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4605 = 10'h18c == _T_110[9:0] ? 4'hc : _GEN_4604; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4606 = 10'h18d == _T_110[9:0] ? 4'hc : _GEN_4605; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4607 = 10'h18e == _T_110[9:0] ? 4'hc : _GEN_4606; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4608 = 10'h18f == _T_110[9:0] ? 4'hc : _GEN_4607; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4609 = 10'h190 == _T_110[9:0] ? 4'hc : _GEN_4608; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4610 = 10'h191 == _T_110[9:0] ? 4'hc : _GEN_4609; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4611 = 10'h192 == _T_110[9:0] ? 4'h9 : _GEN_4610; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4612 = 10'h193 == _T_110[9:0] ? 4'hc : _GEN_4611; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4613 = 10'h194 == _T_110[9:0] ? 4'hc : _GEN_4612; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4614 = 10'h195 == _T_110[9:0] ? 4'hc : _GEN_4613; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4615 = 10'h196 == _T_110[9:0] ? 4'h0 : _GEN_4614; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4616 = 10'h197 == _T_110[9:0] ? 4'h3 : _GEN_4615; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4617 = 10'h198 == _T_110[9:0] ? 4'h1 : _GEN_4616; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4618 = 10'h199 == _T_110[9:0] ? 4'h3 : _GEN_4617; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4619 = 10'h19a == _T_110[9:0] ? 4'h3 : _GEN_4618; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4620 = 10'h19b == _T_110[9:0] ? 4'h3 : _GEN_4619; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4621 = 10'h19c == _T_110[9:0] ? 4'ha : _GEN_4620; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4622 = 10'h19d == _T_110[9:0] ? 4'h3 : _GEN_4621; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4623 = 10'h19e == _T_110[9:0] ? 4'h3 : _GEN_4622; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4624 = 10'h19f == _T_110[9:0] ? 4'h0 : _GEN_4623; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4625 = 10'h1a0 == _T_110[9:0] ? 4'hc : _GEN_4624; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4626 = 10'h1a1 == _T_110[9:0] ? 4'hc : _GEN_4625; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4627 = 10'h1a2 == _T_110[9:0] ? 4'h9 : _GEN_4626; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4628 = 10'h1a3 == _T_110[9:0] ? 4'hc : _GEN_4627; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4629 = 10'h1a4 == _T_110[9:0] ? 4'ha : _GEN_4628; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4630 = 10'h1a5 == _T_110[9:0] ? 4'h0 : _GEN_4629; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4631 = 10'h1a6 == _T_110[9:0] ? 4'hc : _GEN_4630; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4632 = 10'h1a7 == _T_110[9:0] ? 4'h0 : _GEN_4631; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4633 = 10'h1a8 == _T_110[9:0] ? 4'hc : _GEN_4632; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4634 = 10'h1a9 == _T_110[9:0] ? 4'hc : _GEN_4633; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4635 = 10'h1aa == _T_110[9:0] ? 4'hc : _GEN_4634; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4636 = 10'h1ab == _T_110[9:0] ? 4'h9 : _GEN_4635; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4637 = 10'h1ac == _T_110[9:0] ? 4'hc : _GEN_4636; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4638 = 10'h1ad == _T_110[9:0] ? 4'hc : _GEN_4637; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4639 = 10'h1ae == _T_110[9:0] ? 4'hc : _GEN_4638; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4640 = 10'h1af == _T_110[9:0] ? 4'hc : _GEN_4639; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4641 = 10'h1b0 == _T_110[9:0] ? 4'hc : _GEN_4640; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4642 = 10'h1b1 == _T_110[9:0] ? 4'hc : _GEN_4641; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4643 = 10'h1b2 == _T_110[9:0] ? 4'hc : _GEN_4642; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4644 = 10'h1b3 == _T_110[9:0] ? 4'hc : _GEN_4643; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4645 = 10'h1b4 == _T_110[9:0] ? 4'hc : _GEN_4644; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4646 = 10'h1b5 == _T_110[9:0] ? 4'hc : _GEN_4645; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4647 = 10'h1b6 == _T_110[9:0] ? 4'h0 : _GEN_4646; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4648 = 10'h1b7 == _T_110[9:0] ? 4'hc : _GEN_4647; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4649 = 10'h1b8 == _T_110[9:0] ? 4'h0 : _GEN_4648; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4650 = 10'h1b9 == _T_110[9:0] ? 4'hc : _GEN_4649; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4651 = 10'h1ba == _T_110[9:0] ? 4'hc : _GEN_4650; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4652 = 10'h1bb == _T_110[9:0] ? 4'hc : _GEN_4651; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4653 = 10'h1bc == _T_110[9:0] ? 4'h7 : _GEN_4652; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4654 = 10'h1bd == _T_110[9:0] ? 4'ha : _GEN_4653; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4655 = 10'h1be == _T_110[9:0] ? 4'hc : _GEN_4654; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4656 = 10'h1bf == _T_110[9:0] ? 4'h0 : _GEN_4655; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4657 = 10'h1c0 == _T_110[9:0] ? 4'hc : _GEN_4656; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4658 = 10'h1c1 == _T_110[9:0] ? 4'hc : _GEN_4657; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4659 = 10'h1c2 == _T_110[9:0] ? 4'hc : _GEN_4658; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4660 = 10'h1c3 == _T_110[9:0] ? 4'h7 : _GEN_4659; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4661 = 10'h1c4 == _T_110[9:0] ? 4'h7 : _GEN_4660; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4662 = 10'h1c5 == _T_110[9:0] ? 4'hc : _GEN_4661; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4663 = 10'h1c6 == _T_110[9:0] ? 4'hc : _GEN_4662; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4664 = 10'h1c7 == _T_110[9:0] ? 4'hc : _GEN_4663; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4665 = 10'h1c8 == _T_110[9:0] ? 4'hc : _GEN_4664; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4666 = 10'h1c9 == _T_110[9:0] ? 4'hc : _GEN_4665; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4667 = 10'h1ca == _T_110[9:0] ? 4'hc : _GEN_4666; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4668 = 10'h1cb == _T_110[9:0] ? 4'hc : _GEN_4667; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4669 = 10'h1cc == _T_110[9:0] ? 4'hc : _GEN_4668; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4670 = 10'h1cd == _T_110[9:0] ? 4'hc : _GEN_4669; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4671 = 10'h1ce == _T_110[9:0] ? 4'hc : _GEN_4670; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4672 = 10'h1cf == _T_110[9:0] ? 4'hc : _GEN_4671; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4673 = 10'h1d0 == _T_110[9:0] ? 4'hc : _GEN_4672; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4674 = 10'h1d1 == _T_110[9:0] ? 4'hc : _GEN_4673; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4675 = 10'h1d2 == _T_110[9:0] ? 4'hc : _GEN_4674; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4676 = 10'h1d3 == _T_110[9:0] ? 4'hc : _GEN_4675; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4677 = 10'h1d4 == _T_110[9:0] ? 4'hc : _GEN_4676; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4678 = 10'h1d5 == _T_110[9:0] ? 4'hc : _GEN_4677; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4679 = 10'h1d6 == _T_110[9:0] ? 4'hc : _GEN_4678; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4680 = 10'h1d7 == _T_110[9:0] ? 4'hc : _GEN_4679; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4681 = 10'h1d8 == _T_110[9:0] ? 4'hc : _GEN_4680; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4682 = 10'h1d9 == _T_110[9:0] ? 4'hc : _GEN_4681; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4683 = 10'h1da == _T_110[9:0] ? 4'hc : _GEN_4682; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4684 = 10'h1db == _T_110[9:0] ? 4'hc : _GEN_4683; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4685 = 10'h1dc == _T_110[9:0] ? 4'hc : _GEN_4684; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4686 = 10'h1dd == _T_110[9:0] ? 4'ha : _GEN_4685; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4687 = 10'h1de == _T_110[9:0] ? 4'hc : _GEN_4686; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4688 = 10'h1df == _T_110[9:0] ? 4'h0 : _GEN_4687; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4689 = 10'h1e0 == _T_110[9:0] ? 4'h9 : _GEN_4688; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4690 = 10'h1e1 == _T_110[9:0] ? 4'hc : _GEN_4689; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4691 = 10'h1e2 == _T_110[9:0] ? 4'h7 : _GEN_4690; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4692 = 10'h1e3 == _T_110[9:0] ? 4'h7 : _GEN_4691; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4693 = 10'h1e4 == _T_110[9:0] ? 4'hc : _GEN_4692; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4694 = 10'h1e5 == _T_110[9:0] ? 4'hc : _GEN_4693; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4695 = 10'h1e6 == _T_110[9:0] ? 4'hc : _GEN_4694; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4696 = 10'h1e7 == _T_110[9:0] ? 4'hc : _GEN_4695; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4697 = 10'h1e8 == _T_110[9:0] ? 4'hc : _GEN_4696; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4698 = 10'h1e9 == _T_110[9:0] ? 4'hc : _GEN_4697; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4699 = 10'h1ea == _T_110[9:0] ? 4'hc : _GEN_4698; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4700 = 10'h1eb == _T_110[9:0] ? 4'hc : _GEN_4699; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4701 = 10'h1ec == _T_110[9:0] ? 4'hc : _GEN_4700; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4702 = 10'h1ed == _T_110[9:0] ? 4'hc : _GEN_4701; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4703 = 10'h1ee == _T_110[9:0] ? 4'hc : _GEN_4702; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4704 = 10'h1ef == _T_110[9:0] ? 4'hc : _GEN_4703; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4705 = 10'h1f0 == _T_110[9:0] ? 4'hc : _GEN_4704; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4706 = 10'h1f1 == _T_110[9:0] ? 4'hc : _GEN_4705; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4707 = 10'h1f2 == _T_110[9:0] ? 4'hc : _GEN_4706; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4708 = 10'h1f3 == _T_110[9:0] ? 4'hc : _GEN_4707; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4709 = 10'h1f4 == _T_110[9:0] ? 4'hc : _GEN_4708; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4710 = 10'h1f5 == _T_110[9:0] ? 4'hc : _GEN_4709; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4711 = 10'h1f6 == _T_110[9:0] ? 4'hc : _GEN_4710; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4712 = 10'h1f7 == _T_110[9:0] ? 4'hc : _GEN_4711; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4713 = 10'h1f8 == _T_110[9:0] ? 4'hc : _GEN_4712; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4714 = 10'h1f9 == _T_110[9:0] ? 4'hc : _GEN_4713; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4715 = 10'h1fa == _T_110[9:0] ? 4'h9 : _GEN_4714; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4716 = 10'h1fb == _T_110[9:0] ? 4'hc : _GEN_4715; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4717 = 10'h1fc == _T_110[9:0] ? 4'hc : _GEN_4716; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4718 = 10'h1fd == _T_110[9:0] ? 4'h7 : _GEN_4717; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4719 = 10'h1fe == _T_110[9:0] ? 4'hc : _GEN_4718; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4720 = 10'h1ff == _T_110[9:0] ? 4'h0 : _GEN_4719; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4721 = 10'h200 == _T_110[9:0] ? 4'hc : _GEN_4720; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4722 = 10'h201 == _T_110[9:0] ? 4'hc : _GEN_4721; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4723 = 10'h202 == _T_110[9:0] ? 4'ha : _GEN_4722; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4724 = 10'h203 == _T_110[9:0] ? 4'hc : _GEN_4723; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4725 = 10'h204 == _T_110[9:0] ? 4'hc : _GEN_4724; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4726 = 10'h205 == _T_110[9:0] ? 4'hc : _GEN_4725; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4727 = 10'h206 == _T_110[9:0] ? 4'hc : _GEN_4726; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4728 = 10'h207 == _T_110[9:0] ? 4'hc : _GEN_4727; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4729 = 10'h208 == _T_110[9:0] ? 4'hc : _GEN_4728; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4730 = 10'h209 == _T_110[9:0] ? 4'hc : _GEN_4729; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4731 = 10'h20a == _T_110[9:0] ? 4'hc : _GEN_4730; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4732 = 10'h20b == _T_110[9:0] ? 4'hc : _GEN_4731; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4733 = 10'h20c == _T_110[9:0] ? 4'hc : _GEN_4732; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4734 = 10'h20d == _T_110[9:0] ? 4'hc : _GEN_4733; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4735 = 10'h20e == _T_110[9:0] ? 4'hc : _GEN_4734; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4736 = 10'h20f == _T_110[9:0] ? 4'hc : _GEN_4735; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4737 = 10'h210 == _T_110[9:0] ? 4'hc : _GEN_4736; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4738 = 10'h211 == _T_110[9:0] ? 4'hc : _GEN_4737; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4739 = 10'h212 == _T_110[9:0] ? 4'hc : _GEN_4738; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4740 = 10'h213 == _T_110[9:0] ? 4'hc : _GEN_4739; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4741 = 10'h214 == _T_110[9:0] ? 4'hc : _GEN_4740; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4742 = 10'h215 == _T_110[9:0] ? 4'hc : _GEN_4741; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4743 = 10'h216 == _T_110[9:0] ? 4'hc : _GEN_4742; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4744 = 10'h217 == _T_110[9:0] ? 4'hc : _GEN_4743; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4745 = 10'h218 == _T_110[9:0] ? 4'hc : _GEN_4744; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4746 = 10'h219 == _T_110[9:0] ? 4'hc : _GEN_4745; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4747 = 10'h21a == _T_110[9:0] ? 4'hc : _GEN_4746; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4748 = 10'h21b == _T_110[9:0] ? 4'hc : _GEN_4747; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4749 = 10'h21c == _T_110[9:0] ? 4'ha : _GEN_4748; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4750 = 10'h21d == _T_110[9:0] ? 4'h7 : _GEN_4749; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4751 = 10'h21e == _T_110[9:0] ? 4'hc : _GEN_4750; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4752 = 10'h21f == _T_110[9:0] ? 4'h0 : _GEN_4751; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4753 = 10'h220 == _T_110[9:0] ? 4'h0 : _GEN_4752; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4754 = 10'h221 == _T_110[9:0] ? 4'h0 : _GEN_4753; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4755 = 10'h222 == _T_110[9:0] ? 4'h0 : _GEN_4754; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4756 = 10'h223 == _T_110[9:0] ? 4'h0 : _GEN_4755; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4757 = 10'h224 == _T_110[9:0] ? 4'h0 : _GEN_4756; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4758 = 10'h225 == _T_110[9:0] ? 4'h0 : _GEN_4757; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4759 = 10'h226 == _T_110[9:0] ? 4'h0 : _GEN_4758; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4760 = 10'h227 == _T_110[9:0] ? 4'h0 : _GEN_4759; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4761 = 10'h228 == _T_110[9:0] ? 4'h0 : _GEN_4760; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4762 = 10'h229 == _T_110[9:0] ? 4'h0 : _GEN_4761; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4763 = 10'h22a == _T_110[9:0] ? 4'h0 : _GEN_4762; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4764 = 10'h22b == _T_110[9:0] ? 4'h0 : _GEN_4763; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4765 = 10'h22c == _T_110[9:0] ? 4'h0 : _GEN_4764; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4766 = 10'h22d == _T_110[9:0] ? 4'h0 : _GEN_4765; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4767 = 10'h22e == _T_110[9:0] ? 4'h0 : _GEN_4766; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4768 = 10'h22f == _T_110[9:0] ? 4'h0 : _GEN_4767; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4769 = 10'h230 == _T_110[9:0] ? 4'h0 : _GEN_4768; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4770 = 10'h231 == _T_110[9:0] ? 4'h0 : _GEN_4769; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4771 = 10'h232 == _T_110[9:0] ? 4'h0 : _GEN_4770; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4772 = 10'h233 == _T_110[9:0] ? 4'h0 : _GEN_4771; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4773 = 10'h234 == _T_110[9:0] ? 4'h0 : _GEN_4772; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4774 = 10'h235 == _T_110[9:0] ? 4'h0 : _GEN_4773; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4775 = 10'h236 == _T_110[9:0] ? 4'h0 : _GEN_4774; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4776 = 10'h237 == _T_110[9:0] ? 4'h0 : _GEN_4775; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4777 = 10'h238 == _T_110[9:0] ? 4'h0 : _GEN_4776; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4778 = 10'h239 == _T_110[9:0] ? 4'h0 : _GEN_4777; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4779 = 10'h23a == _T_110[9:0] ? 4'h0 : _GEN_4778; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4780 = 10'h23b == _T_110[9:0] ? 4'h0 : _GEN_4779; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4781 = 10'h23c == _T_110[9:0] ? 4'h0 : _GEN_4780; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4782 = 10'h23d == _T_110[9:0] ? 4'h0 : _GEN_4781; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4783 = 10'h23e == _T_110[9:0] ? 4'h0 : _GEN_4782; // @[Filter.scala 191:102]
  wire [3:0] _GEN_4784 = 10'h23f == _T_110[9:0] ? 4'h0 : _GEN_4783; // @[Filter.scala 191:102]
  wire [6:0] _GEN_28312 = {{3'd0}, _GEN_4784}; // @[Filter.scala 191:102]
  wire [10:0] _T_117 = _GEN_28312 * 7'h46; // @[Filter.scala 191:102]
  wire [10:0] _GEN_28313 = {{2'd0}, _T_112}; // @[Filter.scala 191:69]
  wire [10:0] _T_119 = _GEN_28313 + _T_117; // @[Filter.scala 191:69]
  wire [3:0] _GEN_4816 = 10'h1f == _T_110[9:0] ? 4'h0 : 4'h3; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4817 = 10'h20 == _T_110[9:0] ? 4'h3 : _GEN_4816; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4818 = 10'h21 == _T_110[9:0] ? 4'h3 : _GEN_4817; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4819 = 10'h22 == _T_110[9:0] ? 4'h3 : _GEN_4818; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4820 = 10'h23 == _T_110[9:0] ? 4'h3 : _GEN_4819; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4821 = 10'h24 == _T_110[9:0] ? 4'h3 : _GEN_4820; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4822 = 10'h25 == _T_110[9:0] ? 4'h3 : _GEN_4821; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4823 = 10'h26 == _T_110[9:0] ? 4'h3 : _GEN_4822; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4824 = 10'h27 == _T_110[9:0] ? 4'h9 : _GEN_4823; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4825 = 10'h28 == _T_110[9:0] ? 4'h9 : _GEN_4824; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4826 = 10'h29 == _T_110[9:0] ? 4'h3 : _GEN_4825; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4827 = 10'h2a == _T_110[9:0] ? 4'h3 : _GEN_4826; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4828 = 10'h2b == _T_110[9:0] ? 4'h3 : _GEN_4827; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4829 = 10'h2c == _T_110[9:0] ? 4'h3 : _GEN_4828; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4830 = 10'h2d == _T_110[9:0] ? 4'h3 : _GEN_4829; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4831 = 10'h2e == _T_110[9:0] ? 4'h3 : _GEN_4830; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4832 = 10'h2f == _T_110[9:0] ? 4'h3 : _GEN_4831; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4833 = 10'h30 == _T_110[9:0] ? 4'h3 : _GEN_4832; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4834 = 10'h31 == _T_110[9:0] ? 4'h3 : _GEN_4833; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4835 = 10'h32 == _T_110[9:0] ? 4'h3 : _GEN_4834; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4836 = 10'h33 == _T_110[9:0] ? 4'h3 : _GEN_4835; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4837 = 10'h34 == _T_110[9:0] ? 4'h3 : _GEN_4836; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4838 = 10'h35 == _T_110[9:0] ? 4'h3 : _GEN_4837; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4839 = 10'h36 == _T_110[9:0] ? 4'h3 : _GEN_4838; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4840 = 10'h37 == _T_110[9:0] ? 4'h9 : _GEN_4839; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4841 = 10'h38 == _T_110[9:0] ? 4'h9 : _GEN_4840; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4842 = 10'h39 == _T_110[9:0] ? 4'h3 : _GEN_4841; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4843 = 10'h3a == _T_110[9:0] ? 4'h3 : _GEN_4842; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4844 = 10'h3b == _T_110[9:0] ? 4'h3 : _GEN_4843; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4845 = 10'h3c == _T_110[9:0] ? 4'h3 : _GEN_4844; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4846 = 10'h3d == _T_110[9:0] ? 4'h3 : _GEN_4845; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4847 = 10'h3e == _T_110[9:0] ? 4'h3 : _GEN_4846; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4848 = 10'h3f == _T_110[9:0] ? 4'h0 : _GEN_4847; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4849 = 10'h40 == _T_110[9:0] ? 4'h3 : _GEN_4848; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4850 = 10'h41 == _T_110[9:0] ? 4'h3 : _GEN_4849; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4851 = 10'h42 == _T_110[9:0] ? 4'h3 : _GEN_4850; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4852 = 10'h43 == _T_110[9:0] ? 4'h2 : _GEN_4851; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4853 = 10'h44 == _T_110[9:0] ? 4'h3 : _GEN_4852; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4854 = 10'h45 == _T_110[9:0] ? 4'hf : _GEN_4853; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4855 = 10'h46 == _T_110[9:0] ? 4'hf : _GEN_4854; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4856 = 10'h47 == _T_110[9:0] ? 4'hf : _GEN_4855; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4857 = 10'h48 == _T_110[9:0] ? 4'hf : _GEN_4856; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4858 = 10'h49 == _T_110[9:0] ? 4'h3 : _GEN_4857; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4859 = 10'h4a == _T_110[9:0] ? 4'h3 : _GEN_4858; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4860 = 10'h4b == _T_110[9:0] ? 4'h3 : _GEN_4859; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4861 = 10'h4c == _T_110[9:0] ? 4'h3 : _GEN_4860; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4862 = 10'h4d == _T_110[9:0] ? 4'h3 : _GEN_4861; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4863 = 10'h4e == _T_110[9:0] ? 4'h3 : _GEN_4862; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4864 = 10'h4f == _T_110[9:0] ? 4'h3 : _GEN_4863; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4865 = 10'h50 == _T_110[9:0] ? 4'h3 : _GEN_4864; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4866 = 10'h51 == _T_110[9:0] ? 4'h3 : _GEN_4865; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4867 = 10'h52 == _T_110[9:0] ? 4'h3 : _GEN_4866; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4868 = 10'h53 == _T_110[9:0] ? 4'h3 : _GEN_4867; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4869 = 10'h54 == _T_110[9:0] ? 4'h9 : _GEN_4868; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4870 = 10'h55 == _T_110[9:0] ? 4'h9 : _GEN_4869; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4871 = 10'h56 == _T_110[9:0] ? 4'h9 : _GEN_4870; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4872 = 10'h57 == _T_110[9:0] ? 4'hf : _GEN_4871; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4873 = 10'h58 == _T_110[9:0] ? 4'h3 : _GEN_4872; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4874 = 10'h59 == _T_110[9:0] ? 4'hf : _GEN_4873; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4875 = 10'h5a == _T_110[9:0] ? 4'h3 : _GEN_4874; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4876 = 10'h5b == _T_110[9:0] ? 4'h3 : _GEN_4875; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4877 = 10'h5c == _T_110[9:0] ? 4'h3 : _GEN_4876; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4878 = 10'h5d == _T_110[9:0] ? 4'h3 : _GEN_4877; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4879 = 10'h5e == _T_110[9:0] ? 4'h3 : _GEN_4878; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4880 = 10'h5f == _T_110[9:0] ? 4'h0 : _GEN_4879; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4881 = 10'h60 == _T_110[9:0] ? 4'h3 : _GEN_4880; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4882 = 10'h61 == _T_110[9:0] ? 4'h3 : _GEN_4881; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4883 = 10'h62 == _T_110[9:0] ? 4'h3 : _GEN_4882; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4884 = 10'h63 == _T_110[9:0] ? 4'h3 : _GEN_4883; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4885 = 10'h64 == _T_110[9:0] ? 4'h3 : _GEN_4884; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4886 = 10'h65 == _T_110[9:0] ? 4'hf : _GEN_4885; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4887 = 10'h66 == _T_110[9:0] ? 4'h3 : _GEN_4886; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4888 = 10'h67 == _T_110[9:0] ? 4'h3 : _GEN_4887; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4889 = 10'h68 == _T_110[9:0] ? 4'h3 : _GEN_4888; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4890 = 10'h69 == _T_110[9:0] ? 4'hf : _GEN_4889; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4891 = 10'h6a == _T_110[9:0] ? 4'h9 : _GEN_4890; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4892 = 10'h6b == _T_110[9:0] ? 4'h9 : _GEN_4891; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4893 = 10'h6c == _T_110[9:0] ? 4'h3 : _GEN_4892; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4894 = 10'h6d == _T_110[9:0] ? 4'h3 : _GEN_4893; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4895 = 10'h6e == _T_110[9:0] ? 4'h3 : _GEN_4894; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4896 = 10'h6f == _T_110[9:0] ? 4'h3 : _GEN_4895; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4897 = 10'h70 == _T_110[9:0] ? 4'h3 : _GEN_4896; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4898 = 10'h71 == _T_110[9:0] ? 4'h3 : _GEN_4897; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4899 = 10'h72 == _T_110[9:0] ? 4'h3 : _GEN_4898; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4900 = 10'h73 == _T_110[9:0] ? 4'h9 : _GEN_4899; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4901 = 10'h74 == _T_110[9:0] ? 4'hf : _GEN_4900; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4902 = 10'h75 == _T_110[9:0] ? 4'hf : _GEN_4901; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4903 = 10'h76 == _T_110[9:0] ? 4'hf : _GEN_4902; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4904 = 10'h77 == _T_110[9:0] ? 4'h3 : _GEN_4903; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4905 = 10'h78 == _T_110[9:0] ? 4'h3 : _GEN_4904; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4906 = 10'h79 == _T_110[9:0] ? 4'h3 : _GEN_4905; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4907 = 10'h7a == _T_110[9:0] ? 4'hf : _GEN_4906; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4908 = 10'h7b == _T_110[9:0] ? 4'h3 : _GEN_4907; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4909 = 10'h7c == _T_110[9:0] ? 4'h3 : _GEN_4908; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4910 = 10'h7d == _T_110[9:0] ? 4'h2 : _GEN_4909; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4911 = 10'h7e == _T_110[9:0] ? 4'h3 : _GEN_4910; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4912 = 10'h7f == _T_110[9:0] ? 4'h0 : _GEN_4911; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4913 = 10'h80 == _T_110[9:0] ? 4'h3 : _GEN_4912; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4914 = 10'h81 == _T_110[9:0] ? 4'h3 : _GEN_4913; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4915 = 10'h82 == _T_110[9:0] ? 4'h9 : _GEN_4914; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4916 = 10'h83 == _T_110[9:0] ? 4'hf : _GEN_4915; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4917 = 10'h84 == _T_110[9:0] ? 4'h2 : _GEN_4916; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4918 = 10'h85 == _T_110[9:0] ? 4'h9 : _GEN_4917; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4919 = 10'h86 == _T_110[9:0] ? 4'h9 : _GEN_4918; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4920 = 10'h87 == _T_110[9:0] ? 4'h3 : _GEN_4919; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4921 = 10'h88 == _T_110[9:0] ? 4'h3 : _GEN_4920; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4922 = 10'h89 == _T_110[9:0] ? 4'hf : _GEN_4921; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4923 = 10'h8a == _T_110[9:0] ? 4'hf : _GEN_4922; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4924 = 10'h8b == _T_110[9:0] ? 4'h9 : _GEN_4923; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4925 = 10'h8c == _T_110[9:0] ? 4'h9 : _GEN_4924; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4926 = 10'h8d == _T_110[9:0] ? 4'h9 : _GEN_4925; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4927 = 10'h8e == _T_110[9:0] ? 4'h9 : _GEN_4926; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4928 = 10'h8f == _T_110[9:0] ? 4'h9 : _GEN_4927; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4929 = 10'h90 == _T_110[9:0] ? 4'h9 : _GEN_4928; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4930 = 10'h91 == _T_110[9:0] ? 4'h9 : _GEN_4929; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4931 = 10'h92 == _T_110[9:0] ? 4'h9 : _GEN_4930; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4932 = 10'h93 == _T_110[9:0] ? 4'hf : _GEN_4931; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4933 = 10'h94 == _T_110[9:0] ? 4'hf : _GEN_4932; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4934 = 10'h95 == _T_110[9:0] ? 4'h3 : _GEN_4933; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4935 = 10'h96 == _T_110[9:0] ? 4'h3 : _GEN_4934; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4936 = 10'h97 == _T_110[9:0] ? 4'h3 : _GEN_4935; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4937 = 10'h98 == _T_110[9:0] ? 4'h9 : _GEN_4936; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4938 = 10'h99 == _T_110[9:0] ? 4'hf : _GEN_4937; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4939 = 10'h9a == _T_110[9:0] ? 4'h9 : _GEN_4938; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4940 = 10'h9b == _T_110[9:0] ? 4'h9 : _GEN_4939; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4941 = 10'h9c == _T_110[9:0] ? 4'h3 : _GEN_4940; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4942 = 10'h9d == _T_110[9:0] ? 4'h3 : _GEN_4941; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4943 = 10'h9e == _T_110[9:0] ? 4'h3 : _GEN_4942; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4944 = 10'h9f == _T_110[9:0] ? 4'h0 : _GEN_4943; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4945 = 10'ha0 == _T_110[9:0] ? 4'h3 : _GEN_4944; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4946 = 10'ha1 == _T_110[9:0] ? 4'h9 : _GEN_4945; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4947 = 10'ha2 == _T_110[9:0] ? 4'hf : _GEN_4946; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4948 = 10'ha3 == _T_110[9:0] ? 4'h3 : _GEN_4947; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4949 = 10'ha4 == _T_110[9:0] ? 4'h3 : _GEN_4948; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4950 = 10'ha5 == _T_110[9:0] ? 4'h3 : _GEN_4949; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4951 = 10'ha6 == _T_110[9:0] ? 4'h3 : _GEN_4950; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4952 = 10'ha7 == _T_110[9:0] ? 4'hf : _GEN_4951; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4953 = 10'ha8 == _T_110[9:0] ? 4'h3 : _GEN_4952; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4954 = 10'ha9 == _T_110[9:0] ? 4'h9 : _GEN_4953; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4955 = 10'haa == _T_110[9:0] ? 4'hf : _GEN_4954; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4956 = 10'hab == _T_110[9:0] ? 4'hf : _GEN_4955; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4957 = 10'hac == _T_110[9:0] ? 4'hf : _GEN_4956; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4958 = 10'had == _T_110[9:0] ? 4'hf : _GEN_4957; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4959 = 10'hae == _T_110[9:0] ? 4'hf : _GEN_4958; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4960 = 10'haf == _T_110[9:0] ? 4'hf : _GEN_4959; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4961 = 10'hb0 == _T_110[9:0] ? 4'hf : _GEN_4960; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4962 = 10'hb1 == _T_110[9:0] ? 4'hf : _GEN_4961; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4963 = 10'hb2 == _T_110[9:0] ? 4'hf : _GEN_4962; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4964 = 10'hb3 == _T_110[9:0] ? 4'hf : _GEN_4963; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4965 = 10'hb4 == _T_110[9:0] ? 4'h9 : _GEN_4964; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4966 = 10'hb5 == _T_110[9:0] ? 4'h9 : _GEN_4965; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4967 = 10'hb6 == _T_110[9:0] ? 4'h3 : _GEN_4966; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4968 = 10'hb7 == _T_110[9:0] ? 4'hf : _GEN_4967; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4969 = 10'hb8 == _T_110[9:0] ? 4'h3 : _GEN_4968; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4970 = 10'hb9 == _T_110[9:0] ? 4'h3 : _GEN_4969; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4971 = 10'hba == _T_110[9:0] ? 4'h3 : _GEN_4970; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4972 = 10'hbb == _T_110[9:0] ? 4'hf : _GEN_4971; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4973 = 10'hbc == _T_110[9:0] ? 4'h3 : _GEN_4972; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4974 = 10'hbd == _T_110[9:0] ? 4'h3 : _GEN_4973; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4975 = 10'hbe == _T_110[9:0] ? 4'h3 : _GEN_4974; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4976 = 10'hbf == _T_110[9:0] ? 4'h0 : _GEN_4975; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4977 = 10'hc0 == _T_110[9:0] ? 4'h3 : _GEN_4976; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4978 = 10'hc1 == _T_110[9:0] ? 4'h3 : _GEN_4977; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4979 = 10'hc2 == _T_110[9:0] ? 4'h3 : _GEN_4978; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4980 = 10'hc3 == _T_110[9:0] ? 4'h2 : _GEN_4979; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4981 = 10'hc4 == _T_110[9:0] ? 4'hf : _GEN_4980; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4982 = 10'hc5 == _T_110[9:0] ? 4'hf : _GEN_4981; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4983 = 10'hc6 == _T_110[9:0] ? 4'hf : _GEN_4982; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4984 = 10'hc7 == _T_110[9:0] ? 4'h3 : _GEN_4983; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4985 = 10'hc8 == _T_110[9:0] ? 4'h9 : _GEN_4984; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4986 = 10'hc9 == _T_110[9:0] ? 4'hf : _GEN_4985; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4987 = 10'hca == _T_110[9:0] ? 4'hf : _GEN_4986; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4988 = 10'hcb == _T_110[9:0] ? 4'hf : _GEN_4987; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4989 = 10'hcc == _T_110[9:0] ? 4'hf : _GEN_4988; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4990 = 10'hcd == _T_110[9:0] ? 4'hf : _GEN_4989; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4991 = 10'hce == _T_110[9:0] ? 4'hf : _GEN_4990; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4992 = 10'hcf == _T_110[9:0] ? 4'hf : _GEN_4991; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4993 = 10'hd0 == _T_110[9:0] ? 4'hf : _GEN_4992; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4994 = 10'hd1 == _T_110[9:0] ? 4'hf : _GEN_4993; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4995 = 10'hd2 == _T_110[9:0] ? 4'hf : _GEN_4994; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4996 = 10'hd3 == _T_110[9:0] ? 4'hf : _GEN_4995; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4997 = 10'hd4 == _T_110[9:0] ? 4'hf : _GEN_4996; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4998 = 10'hd5 == _T_110[9:0] ? 4'hf : _GEN_4997; // @[Filter.scala 191:142]
  wire [3:0] _GEN_4999 = 10'hd6 == _T_110[9:0] ? 4'h9 : _GEN_4998; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5000 = 10'hd7 == _T_110[9:0] ? 4'h3 : _GEN_4999; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5001 = 10'hd8 == _T_110[9:0] ? 4'hf : _GEN_5000; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5002 = 10'hd9 == _T_110[9:0] ? 4'h3 : _GEN_5001; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5003 = 10'hda == _T_110[9:0] ? 4'h3 : _GEN_5002; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5004 = 10'hdb == _T_110[9:0] ? 4'h3 : _GEN_5003; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5005 = 10'hdc == _T_110[9:0] ? 4'h3 : _GEN_5004; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5006 = 10'hdd == _T_110[9:0] ? 4'h3 : _GEN_5005; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5007 = 10'hde == _T_110[9:0] ? 4'h2 : _GEN_5006; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5008 = 10'hdf == _T_110[9:0] ? 4'h0 : _GEN_5007; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5009 = 10'he0 == _T_110[9:0] ? 4'h3 : _GEN_5008; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5010 = 10'he1 == _T_110[9:0] ? 4'h3 : _GEN_5009; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5011 = 10'he2 == _T_110[9:0] ? 4'h3 : _GEN_5010; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5012 = 10'he3 == _T_110[9:0] ? 4'h3 : _GEN_5011; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5013 = 10'he4 == _T_110[9:0] ? 4'h3 : _GEN_5012; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5014 = 10'he5 == _T_110[9:0] ? 4'h3 : _GEN_5013; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5015 = 10'he6 == _T_110[9:0] ? 4'h3 : _GEN_5014; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5016 = 10'he7 == _T_110[9:0] ? 4'h9 : _GEN_5015; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5017 = 10'he8 == _T_110[9:0] ? 4'h9 : _GEN_5016; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5018 = 10'he9 == _T_110[9:0] ? 4'h9 : _GEN_5017; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5019 = 10'hea == _T_110[9:0] ? 4'hf : _GEN_5018; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5020 = 10'heb == _T_110[9:0] ? 4'hf : _GEN_5019; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5021 = 10'hec == _T_110[9:0] ? 4'hf : _GEN_5020; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5022 = 10'hed == _T_110[9:0] ? 4'hf : _GEN_5021; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5023 = 10'hee == _T_110[9:0] ? 4'hf : _GEN_5022; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5024 = 10'hef == _T_110[9:0] ? 4'hf : _GEN_5023; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5025 = 10'hf0 == _T_110[9:0] ? 4'hf : _GEN_5024; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5026 = 10'hf1 == _T_110[9:0] ? 4'hf : _GEN_5025; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5027 = 10'hf2 == _T_110[9:0] ? 4'hf : _GEN_5026; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5028 = 10'hf3 == _T_110[9:0] ? 4'hf : _GEN_5027; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5029 = 10'hf4 == _T_110[9:0] ? 4'hf : _GEN_5028; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5030 = 10'hf5 == _T_110[9:0] ? 4'h9 : _GEN_5029; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5031 = 10'hf6 == _T_110[9:0] ? 4'hf : _GEN_5030; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5032 = 10'hf7 == _T_110[9:0] ? 4'hf : _GEN_5031; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5033 = 10'hf8 == _T_110[9:0] ? 4'h9 : _GEN_5032; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5034 = 10'hf9 == _T_110[9:0] ? 4'hf : _GEN_5033; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5035 = 10'hfa == _T_110[9:0] ? 4'h3 : _GEN_5034; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5036 = 10'hfb == _T_110[9:0] ? 4'h3 : _GEN_5035; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5037 = 10'hfc == _T_110[9:0] ? 4'h3 : _GEN_5036; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5038 = 10'hfd == _T_110[9:0] ? 4'h3 : _GEN_5037; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5039 = 10'hfe == _T_110[9:0] ? 4'h3 : _GEN_5038; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5040 = 10'hff == _T_110[9:0] ? 4'h0 : _GEN_5039; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5041 = 10'h100 == _T_110[9:0] ? 4'h3 : _GEN_5040; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5042 = 10'h101 == _T_110[9:0] ? 4'hf : _GEN_5041; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5043 = 10'h102 == _T_110[9:0] ? 4'h3 : _GEN_5042; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5044 = 10'h103 == _T_110[9:0] ? 4'h3 : _GEN_5043; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5045 = 10'h104 == _T_110[9:0] ? 4'h3 : _GEN_5044; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5046 = 10'h105 == _T_110[9:0] ? 4'h3 : _GEN_5045; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5047 = 10'h106 == _T_110[9:0] ? 4'h3 : _GEN_5046; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5048 = 10'h107 == _T_110[9:0] ? 4'h3 : _GEN_5047; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5049 = 10'h108 == _T_110[9:0] ? 4'h9 : _GEN_5048; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5050 = 10'h109 == _T_110[9:0] ? 4'hf : _GEN_5049; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5051 = 10'h10a == _T_110[9:0] ? 4'hf : _GEN_5050; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5052 = 10'h10b == _T_110[9:0] ? 4'hf : _GEN_5051; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5053 = 10'h10c == _T_110[9:0] ? 4'hf : _GEN_5052; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5054 = 10'h10d == _T_110[9:0] ? 4'h0 : _GEN_5053; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5055 = 10'h10e == _T_110[9:0] ? 4'hf : _GEN_5054; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5056 = 10'h10f == _T_110[9:0] ? 4'hf : _GEN_5055; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5057 = 10'h110 == _T_110[9:0] ? 4'hf : _GEN_5056; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5058 = 10'h111 == _T_110[9:0] ? 4'h0 : _GEN_5057; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5059 = 10'h112 == _T_110[9:0] ? 4'hf : _GEN_5058; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5060 = 10'h113 == _T_110[9:0] ? 4'hf : _GEN_5059; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5061 = 10'h114 == _T_110[9:0] ? 4'hf : _GEN_5060; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5062 = 10'h115 == _T_110[9:0] ? 4'hf : _GEN_5061; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5063 = 10'h116 == _T_110[9:0] ? 4'h9 : _GEN_5062; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5064 = 10'h117 == _T_110[9:0] ? 4'h3 : _GEN_5063; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5065 = 10'h118 == _T_110[9:0] ? 4'h3 : _GEN_5064; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5066 = 10'h119 == _T_110[9:0] ? 4'h3 : _GEN_5065; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5067 = 10'h11a == _T_110[9:0] ? 4'hf : _GEN_5066; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5068 = 10'h11b == _T_110[9:0] ? 4'h3 : _GEN_5067; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5069 = 10'h11c == _T_110[9:0] ? 4'h3 : _GEN_5068; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5070 = 10'h11d == _T_110[9:0] ? 4'h2 : _GEN_5069; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5071 = 10'h11e == _T_110[9:0] ? 4'h3 : _GEN_5070; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5072 = 10'h11f == _T_110[9:0] ? 4'h0 : _GEN_5071; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5073 = 10'h120 == _T_110[9:0] ? 4'h3 : _GEN_5072; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5074 = 10'h121 == _T_110[9:0] ? 4'h3 : _GEN_5073; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5075 = 10'h122 == _T_110[9:0] ? 4'h3 : _GEN_5074; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5076 = 10'h123 == _T_110[9:0] ? 4'h3 : _GEN_5075; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5077 = 10'h124 == _T_110[9:0] ? 4'h3 : _GEN_5076; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5078 = 10'h125 == _T_110[9:0] ? 4'h3 : _GEN_5077; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5079 = 10'h126 == _T_110[9:0] ? 4'h3 : _GEN_5078; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5080 = 10'h127 == _T_110[9:0] ? 4'h9 : _GEN_5079; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5081 = 10'h128 == _T_110[9:0] ? 4'hf : _GEN_5080; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5082 = 10'h129 == _T_110[9:0] ? 4'h3 : _GEN_5081; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5083 = 10'h12a == _T_110[9:0] ? 4'h3 : _GEN_5082; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5084 = 10'h12b == _T_110[9:0] ? 4'hf : _GEN_5083; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5085 = 10'h12c == _T_110[9:0] ? 4'hf : _GEN_5084; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5086 = 10'h12d == _T_110[9:0] ? 4'hf : _GEN_5085; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5087 = 10'h12e == _T_110[9:0] ? 4'hf : _GEN_5086; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5088 = 10'h12f == _T_110[9:0] ? 4'hf : _GEN_5087; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5089 = 10'h130 == _T_110[9:0] ? 4'hf : _GEN_5088; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5090 = 10'h131 == _T_110[9:0] ? 4'hf : _GEN_5089; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5091 = 10'h132 == _T_110[9:0] ? 4'hf : _GEN_5090; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5092 = 10'h133 == _T_110[9:0] ? 4'hf : _GEN_5091; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5093 = 10'h134 == _T_110[9:0] ? 4'h3 : _GEN_5092; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5094 = 10'h135 == _T_110[9:0] ? 4'h3 : _GEN_5093; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5095 = 10'h136 == _T_110[9:0] ? 4'hf : _GEN_5094; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5096 = 10'h137 == _T_110[9:0] ? 4'h9 : _GEN_5095; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5097 = 10'h138 == _T_110[9:0] ? 4'h3 : _GEN_5096; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5098 = 10'h139 == _T_110[9:0] ? 4'h3 : _GEN_5097; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5099 = 10'h13a == _T_110[9:0] ? 4'h3 : _GEN_5098; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5100 = 10'h13b == _T_110[9:0] ? 4'h3 : _GEN_5099; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5101 = 10'h13c == _T_110[9:0] ? 4'h3 : _GEN_5100; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5102 = 10'h13d == _T_110[9:0] ? 4'h3 : _GEN_5101; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5103 = 10'h13e == _T_110[9:0] ? 4'h3 : _GEN_5102; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5104 = 10'h13f == _T_110[9:0] ? 4'h0 : _GEN_5103; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5105 = 10'h140 == _T_110[9:0] ? 4'h3 : _GEN_5104; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5106 = 10'h141 == _T_110[9:0] ? 4'h3 : _GEN_5105; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5107 = 10'h142 == _T_110[9:0] ? 4'h2 : _GEN_5106; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5108 = 10'h143 == _T_110[9:0] ? 4'h3 : _GEN_5107; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5109 = 10'h144 == _T_110[9:0] ? 4'h3 : _GEN_5108; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5110 = 10'h145 == _T_110[9:0] ? 4'h3 : _GEN_5109; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5111 = 10'h146 == _T_110[9:0] ? 4'h9 : _GEN_5110; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5112 = 10'h147 == _T_110[9:0] ? 4'hf : _GEN_5111; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5113 = 10'h148 == _T_110[9:0] ? 4'h3 : _GEN_5112; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5114 = 10'h149 == _T_110[9:0] ? 4'h3 : _GEN_5113; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5115 = 10'h14a == _T_110[9:0] ? 4'h3 : _GEN_5114; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5116 = 10'h14b == _T_110[9:0] ? 4'h3 : _GEN_5115; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5117 = 10'h14c == _T_110[9:0] ? 4'h3 : _GEN_5116; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5118 = 10'h14d == _T_110[9:0] ? 4'h3 : _GEN_5117; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5119 = 10'h14e == _T_110[9:0] ? 4'h3 : _GEN_5118; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5120 = 10'h14f == _T_110[9:0] ? 4'h3 : _GEN_5119; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5121 = 10'h150 == _T_110[9:0] ? 4'h3 : _GEN_5120; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5122 = 10'h151 == _T_110[9:0] ? 4'h3 : _GEN_5121; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5123 = 10'h152 == _T_110[9:0] ? 4'h3 : _GEN_5122; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5124 = 10'h153 == _T_110[9:0] ? 4'h3 : _GEN_5123; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5125 = 10'h154 == _T_110[9:0] ? 4'h3 : _GEN_5124; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5126 = 10'h155 == _T_110[9:0] ? 4'h3 : _GEN_5125; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5127 = 10'h156 == _T_110[9:0] ? 4'h3 : _GEN_5126; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5128 = 10'h157 == _T_110[9:0] ? 4'hf : _GEN_5127; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5129 = 10'h158 == _T_110[9:0] ? 4'h3 : _GEN_5128; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5130 = 10'h159 == _T_110[9:0] ? 4'h3 : _GEN_5129; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5131 = 10'h15a == _T_110[9:0] ? 4'h3 : _GEN_5130; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5132 = 10'h15b == _T_110[9:0] ? 4'h3 : _GEN_5131; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5133 = 10'h15c == _T_110[9:0] ? 4'h3 : _GEN_5132; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5134 = 10'h15d == _T_110[9:0] ? 4'h3 : _GEN_5133; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5135 = 10'h15e == _T_110[9:0] ? 4'h2 : _GEN_5134; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5136 = 10'h15f == _T_110[9:0] ? 4'h0 : _GEN_5135; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5137 = 10'h160 == _T_110[9:0] ? 4'h3 : _GEN_5136; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5138 = 10'h161 == _T_110[9:0] ? 4'h3 : _GEN_5137; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5139 = 10'h162 == _T_110[9:0] ? 4'h3 : _GEN_5138; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5140 = 10'h163 == _T_110[9:0] ? 4'h2 : _GEN_5139; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5141 = 10'h164 == _T_110[9:0] ? 4'h3 : _GEN_5140; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5142 = 10'h165 == _T_110[9:0] ? 4'h9 : _GEN_5141; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5143 = 10'h166 == _T_110[9:0] ? 4'hf : _GEN_5142; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5144 = 10'h167 == _T_110[9:0] ? 4'hf : _GEN_5143; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5145 = 10'h168 == _T_110[9:0] ? 4'hd : _GEN_5144; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5146 = 10'h169 == _T_110[9:0] ? 4'h9 : _GEN_5145; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5147 = 10'h16a == _T_110[9:0] ? 4'hd : _GEN_5146; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5148 = 10'h16b == _T_110[9:0] ? 4'hd : _GEN_5147; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5149 = 10'h16c == _T_110[9:0] ? 4'h3 : _GEN_5148; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5150 = 10'h16d == _T_110[9:0] ? 4'h3 : _GEN_5149; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5151 = 10'h16e == _T_110[9:0] ? 4'h3 : _GEN_5150; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5152 = 10'h16f == _T_110[9:0] ? 4'h3 : _GEN_5151; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5153 = 10'h170 == _T_110[9:0] ? 4'h3 : _GEN_5152; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5154 = 10'h171 == _T_110[9:0] ? 4'h3 : _GEN_5153; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5155 = 10'h172 == _T_110[9:0] ? 4'h3 : _GEN_5154; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5156 = 10'h173 == _T_110[9:0] ? 4'h3 : _GEN_5155; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5157 = 10'h174 == _T_110[9:0] ? 4'h3 : _GEN_5156; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5158 = 10'h175 == _T_110[9:0] ? 4'h3 : _GEN_5157; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5159 = 10'h176 == _T_110[9:0] ? 4'hf : _GEN_5158; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5160 = 10'h177 == _T_110[9:0] ? 4'hf : _GEN_5159; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5161 = 10'h178 == _T_110[9:0] ? 4'h9 : _GEN_5160; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5162 = 10'h179 == _T_110[9:0] ? 4'h3 : _GEN_5161; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5163 = 10'h17a == _T_110[9:0] ? 4'h3 : _GEN_5162; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5164 = 10'h17b == _T_110[9:0] ? 4'h3 : _GEN_5163; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5165 = 10'h17c == _T_110[9:0] ? 4'h3 : _GEN_5164; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5166 = 10'h17d == _T_110[9:0] ? 4'h2 : _GEN_5165; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5167 = 10'h17e == _T_110[9:0] ? 4'h3 : _GEN_5166; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5168 = 10'h17f == _T_110[9:0] ? 4'h0 : _GEN_5167; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5169 = 10'h180 == _T_110[9:0] ? 4'hd : _GEN_5168; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5170 = 10'h181 == _T_110[9:0] ? 4'hd : _GEN_5169; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5171 = 10'h182 == _T_110[9:0] ? 4'hd : _GEN_5170; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5172 = 10'h183 == _T_110[9:0] ? 4'hd : _GEN_5171; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5173 = 10'h184 == _T_110[9:0] ? 4'h3 : _GEN_5172; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5174 = 10'h185 == _T_110[9:0] ? 4'h9 : _GEN_5173; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5175 = 10'h186 == _T_110[9:0] ? 4'hb : _GEN_5174; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5176 = 10'h187 == _T_110[9:0] ? 4'hf : _GEN_5175; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5177 = 10'h188 == _T_110[9:0] ? 4'hd : _GEN_5176; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5178 = 10'h189 == _T_110[9:0] ? 4'hd : _GEN_5177; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5179 = 10'h18a == _T_110[9:0] ? 4'hd : _GEN_5178; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5180 = 10'h18b == _T_110[9:0] ? 4'hd : _GEN_5179; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5181 = 10'h18c == _T_110[9:0] ? 4'hd : _GEN_5180; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5182 = 10'h18d == _T_110[9:0] ? 4'hd : _GEN_5181; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5183 = 10'h18e == _T_110[9:0] ? 4'hd : _GEN_5182; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5184 = 10'h18f == _T_110[9:0] ? 4'hd : _GEN_5183; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5185 = 10'h190 == _T_110[9:0] ? 4'hd : _GEN_5184; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5186 = 10'h191 == _T_110[9:0] ? 4'hd : _GEN_5185; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5187 = 10'h192 == _T_110[9:0] ? 4'h9 : _GEN_5186; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5188 = 10'h193 == _T_110[9:0] ? 4'hd : _GEN_5187; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5189 = 10'h194 == _T_110[9:0] ? 4'hd : _GEN_5188; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5190 = 10'h195 == _T_110[9:0] ? 4'hd : _GEN_5189; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5191 = 10'h196 == _T_110[9:0] ? 4'hf : _GEN_5190; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5192 = 10'h197 == _T_110[9:0] ? 4'h3 : _GEN_5191; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5193 = 10'h198 == _T_110[9:0] ? 4'h9 : _GEN_5192; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5194 = 10'h199 == _T_110[9:0] ? 4'h3 : _GEN_5193; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5195 = 10'h19a == _T_110[9:0] ? 4'h3 : _GEN_5194; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5196 = 10'h19b == _T_110[9:0] ? 4'h3 : _GEN_5195; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5197 = 10'h19c == _T_110[9:0] ? 4'h3 : _GEN_5196; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5198 = 10'h19d == _T_110[9:0] ? 4'h3 : _GEN_5197; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5199 = 10'h19e == _T_110[9:0] ? 4'h3 : _GEN_5198; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5200 = 10'h19f == _T_110[9:0] ? 4'h0 : _GEN_5199; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5201 = 10'h1a0 == _T_110[9:0] ? 4'hd : _GEN_5200; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5202 = 10'h1a1 == _T_110[9:0] ? 4'hd : _GEN_5201; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5203 = 10'h1a2 == _T_110[9:0] ? 4'h9 : _GEN_5202; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5204 = 10'h1a3 == _T_110[9:0] ? 4'hd : _GEN_5203; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5205 = 10'h1a4 == _T_110[9:0] ? 4'h3 : _GEN_5204; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5206 = 10'h1a5 == _T_110[9:0] ? 4'hf : _GEN_5205; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5207 = 10'h1a6 == _T_110[9:0] ? 4'hd : _GEN_5206; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5208 = 10'h1a7 == _T_110[9:0] ? 4'hf : _GEN_5207; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5209 = 10'h1a8 == _T_110[9:0] ? 4'hb : _GEN_5208; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5210 = 10'h1a9 == _T_110[9:0] ? 4'hd : _GEN_5209; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5211 = 10'h1aa == _T_110[9:0] ? 4'hd : _GEN_5210; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5212 = 10'h1ab == _T_110[9:0] ? 4'h9 : _GEN_5211; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5213 = 10'h1ac == _T_110[9:0] ? 4'hd : _GEN_5212; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5214 = 10'h1ad == _T_110[9:0] ? 4'hd : _GEN_5213; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5215 = 10'h1ae == _T_110[9:0] ? 4'hd : _GEN_5214; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5216 = 10'h1af == _T_110[9:0] ? 4'hd : _GEN_5215; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5217 = 10'h1b0 == _T_110[9:0] ? 4'hd : _GEN_5216; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5218 = 10'h1b1 == _T_110[9:0] ? 4'hd : _GEN_5217; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5219 = 10'h1b2 == _T_110[9:0] ? 4'hd : _GEN_5218; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5220 = 10'h1b3 == _T_110[9:0] ? 4'hd : _GEN_5219; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5221 = 10'h1b4 == _T_110[9:0] ? 4'hd : _GEN_5220; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5222 = 10'h1b5 == _T_110[9:0] ? 4'hd : _GEN_5221; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5223 = 10'h1b6 == _T_110[9:0] ? 4'hf : _GEN_5222; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5224 = 10'h1b7 == _T_110[9:0] ? 4'hd : _GEN_5223; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5225 = 10'h1b8 == _T_110[9:0] ? 4'hf : _GEN_5224; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5226 = 10'h1b9 == _T_110[9:0] ? 4'hd : _GEN_5225; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5227 = 10'h1ba == _T_110[9:0] ? 4'hd : _GEN_5226; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5228 = 10'h1bb == _T_110[9:0] ? 4'hd : _GEN_5227; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5229 = 10'h1bc == _T_110[9:0] ? 4'h2 : _GEN_5228; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5230 = 10'h1bd == _T_110[9:0] ? 4'h3 : _GEN_5229; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5231 = 10'h1be == _T_110[9:0] ? 4'hd : _GEN_5230; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5232 = 10'h1bf == _T_110[9:0] ? 4'h0 : _GEN_5231; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5233 = 10'h1c0 == _T_110[9:0] ? 4'hd : _GEN_5232; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5234 = 10'h1c1 == _T_110[9:0] ? 4'hd : _GEN_5233; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5235 = 10'h1c2 == _T_110[9:0] ? 4'hd : _GEN_5234; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5236 = 10'h1c3 == _T_110[9:0] ? 4'h2 : _GEN_5235; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5237 = 10'h1c4 == _T_110[9:0] ? 4'h2 : _GEN_5236; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5238 = 10'h1c5 == _T_110[9:0] ? 4'hd : _GEN_5237; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5239 = 10'h1c6 == _T_110[9:0] ? 4'hd : _GEN_5238; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5240 = 10'h1c7 == _T_110[9:0] ? 4'hd : _GEN_5239; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5241 = 10'h1c8 == _T_110[9:0] ? 4'hd : _GEN_5240; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5242 = 10'h1c9 == _T_110[9:0] ? 4'hb : _GEN_5241; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5243 = 10'h1ca == _T_110[9:0] ? 4'hb : _GEN_5242; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5244 = 10'h1cb == _T_110[9:0] ? 4'hb : _GEN_5243; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5245 = 10'h1cc == _T_110[9:0] ? 4'hb : _GEN_5244; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5246 = 10'h1cd == _T_110[9:0] ? 4'hb : _GEN_5245; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5247 = 10'h1ce == _T_110[9:0] ? 4'hb : _GEN_5246; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5248 = 10'h1cf == _T_110[9:0] ? 4'hb : _GEN_5247; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5249 = 10'h1d0 == _T_110[9:0] ? 4'hb : _GEN_5248; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5250 = 10'h1d1 == _T_110[9:0] ? 4'hb : _GEN_5249; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5251 = 10'h1d2 == _T_110[9:0] ? 4'hb : _GEN_5250; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5252 = 10'h1d3 == _T_110[9:0] ? 4'hb : _GEN_5251; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5253 = 10'h1d4 == _T_110[9:0] ? 4'hb : _GEN_5252; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5254 = 10'h1d5 == _T_110[9:0] ? 4'hb : _GEN_5253; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5255 = 10'h1d6 == _T_110[9:0] ? 4'hd : _GEN_5254; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5256 = 10'h1d7 == _T_110[9:0] ? 4'hd : _GEN_5255; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5257 = 10'h1d8 == _T_110[9:0] ? 4'hd : _GEN_5256; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5258 = 10'h1d9 == _T_110[9:0] ? 4'hd : _GEN_5257; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5259 = 10'h1da == _T_110[9:0] ? 4'hd : _GEN_5258; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5260 = 10'h1db == _T_110[9:0] ? 4'hd : _GEN_5259; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5261 = 10'h1dc == _T_110[9:0] ? 4'hd : _GEN_5260; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5262 = 10'h1dd == _T_110[9:0] ? 4'h3 : _GEN_5261; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5263 = 10'h1de == _T_110[9:0] ? 4'hd : _GEN_5262; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5264 = 10'h1df == _T_110[9:0] ? 4'h0 : _GEN_5263; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5265 = 10'h1e0 == _T_110[9:0] ? 4'h9 : _GEN_5264; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5266 = 10'h1e1 == _T_110[9:0] ? 4'hd : _GEN_5265; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5267 = 10'h1e2 == _T_110[9:0] ? 4'h2 : _GEN_5266; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5268 = 10'h1e3 == _T_110[9:0] ? 4'h2 : _GEN_5267; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5269 = 10'h1e4 == _T_110[9:0] ? 4'hd : _GEN_5268; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5270 = 10'h1e5 == _T_110[9:0] ? 4'hd : _GEN_5269; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5271 = 10'h1e6 == _T_110[9:0] ? 4'hd : _GEN_5270; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5272 = 10'h1e7 == _T_110[9:0] ? 4'hd : _GEN_5271; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5273 = 10'h1e8 == _T_110[9:0] ? 4'hb : _GEN_5272; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5274 = 10'h1e9 == _T_110[9:0] ? 4'hd : _GEN_5273; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5275 = 10'h1ea == _T_110[9:0] ? 4'hd : _GEN_5274; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5276 = 10'h1eb == _T_110[9:0] ? 4'hb : _GEN_5275; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5277 = 10'h1ec == _T_110[9:0] ? 4'hd : _GEN_5276; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5278 = 10'h1ed == _T_110[9:0] ? 4'hb : _GEN_5277; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5279 = 10'h1ee == _T_110[9:0] ? 4'hd : _GEN_5278; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5280 = 10'h1ef == _T_110[9:0] ? 4'hb : _GEN_5279; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5281 = 10'h1f0 == _T_110[9:0] ? 4'hd : _GEN_5280; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5282 = 10'h1f1 == _T_110[9:0] ? 4'hb : _GEN_5281; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5283 = 10'h1f2 == _T_110[9:0] ? 4'hb : _GEN_5282; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5284 = 10'h1f3 == _T_110[9:0] ? 4'hd : _GEN_5283; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5285 = 10'h1f4 == _T_110[9:0] ? 4'hb : _GEN_5284; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5286 = 10'h1f5 == _T_110[9:0] ? 4'hb : _GEN_5285; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5287 = 10'h1f6 == _T_110[9:0] ? 4'hd : _GEN_5286; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5288 = 10'h1f7 == _T_110[9:0] ? 4'hd : _GEN_5287; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5289 = 10'h1f8 == _T_110[9:0] ? 4'hd : _GEN_5288; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5290 = 10'h1f9 == _T_110[9:0] ? 4'hd : _GEN_5289; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5291 = 10'h1fa == _T_110[9:0] ? 4'h9 : _GEN_5290; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5292 = 10'h1fb == _T_110[9:0] ? 4'hd : _GEN_5291; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5293 = 10'h1fc == _T_110[9:0] ? 4'hd : _GEN_5292; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5294 = 10'h1fd == _T_110[9:0] ? 4'h2 : _GEN_5293; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5295 = 10'h1fe == _T_110[9:0] ? 4'hd : _GEN_5294; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5296 = 10'h1ff == _T_110[9:0] ? 4'h0 : _GEN_5295; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5297 = 10'h200 == _T_110[9:0] ? 4'hd : _GEN_5296; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5298 = 10'h201 == _T_110[9:0] ? 4'hd : _GEN_5297; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5299 = 10'h202 == _T_110[9:0] ? 4'h3 : _GEN_5298; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5300 = 10'h203 == _T_110[9:0] ? 4'hd : _GEN_5299; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5301 = 10'h204 == _T_110[9:0] ? 4'hd : _GEN_5300; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5302 = 10'h205 == _T_110[9:0] ? 4'hd : _GEN_5301; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5303 = 10'h206 == _T_110[9:0] ? 4'hb : _GEN_5302; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5304 = 10'h207 == _T_110[9:0] ? 4'hb : _GEN_5303; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5305 = 10'h208 == _T_110[9:0] ? 4'hd : _GEN_5304; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5306 = 10'h209 == _T_110[9:0] ? 4'hd : _GEN_5305; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5307 = 10'h20a == _T_110[9:0] ? 4'hd : _GEN_5306; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5308 = 10'h20b == _T_110[9:0] ? 4'hb : _GEN_5307; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5309 = 10'h20c == _T_110[9:0] ? 4'hd : _GEN_5308; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5310 = 10'h20d == _T_110[9:0] ? 4'hb : _GEN_5309; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5311 = 10'h20e == _T_110[9:0] ? 4'hd : _GEN_5310; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5312 = 10'h20f == _T_110[9:0] ? 4'hb : _GEN_5311; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5313 = 10'h210 == _T_110[9:0] ? 4'hd : _GEN_5312; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5314 = 10'h211 == _T_110[9:0] ? 4'hd : _GEN_5313; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5315 = 10'h212 == _T_110[9:0] ? 4'hb : _GEN_5314; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5316 = 10'h213 == _T_110[9:0] ? 4'hb : _GEN_5315; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5317 = 10'h214 == _T_110[9:0] ? 4'hb : _GEN_5316; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5318 = 10'h215 == _T_110[9:0] ? 4'hd : _GEN_5317; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5319 = 10'h216 == _T_110[9:0] ? 4'hd : _GEN_5318; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5320 = 10'h217 == _T_110[9:0] ? 4'hd : _GEN_5319; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5321 = 10'h218 == _T_110[9:0] ? 4'hd : _GEN_5320; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5322 = 10'h219 == _T_110[9:0] ? 4'hd : _GEN_5321; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5323 = 10'h21a == _T_110[9:0] ? 4'hd : _GEN_5322; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5324 = 10'h21b == _T_110[9:0] ? 4'hd : _GEN_5323; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5325 = 10'h21c == _T_110[9:0] ? 4'h3 : _GEN_5324; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5326 = 10'h21d == _T_110[9:0] ? 4'h2 : _GEN_5325; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5327 = 10'h21e == _T_110[9:0] ? 4'hd : _GEN_5326; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5328 = 10'h21f == _T_110[9:0] ? 4'h0 : _GEN_5327; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5329 = 10'h220 == _T_110[9:0] ? 4'h0 : _GEN_5328; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5330 = 10'h221 == _T_110[9:0] ? 4'h0 : _GEN_5329; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5331 = 10'h222 == _T_110[9:0] ? 4'h0 : _GEN_5330; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5332 = 10'h223 == _T_110[9:0] ? 4'h0 : _GEN_5331; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5333 = 10'h224 == _T_110[9:0] ? 4'h0 : _GEN_5332; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5334 = 10'h225 == _T_110[9:0] ? 4'h0 : _GEN_5333; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5335 = 10'h226 == _T_110[9:0] ? 4'h0 : _GEN_5334; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5336 = 10'h227 == _T_110[9:0] ? 4'h0 : _GEN_5335; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5337 = 10'h228 == _T_110[9:0] ? 4'h0 : _GEN_5336; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5338 = 10'h229 == _T_110[9:0] ? 4'h0 : _GEN_5337; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5339 = 10'h22a == _T_110[9:0] ? 4'h0 : _GEN_5338; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5340 = 10'h22b == _T_110[9:0] ? 4'h0 : _GEN_5339; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5341 = 10'h22c == _T_110[9:0] ? 4'h0 : _GEN_5340; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5342 = 10'h22d == _T_110[9:0] ? 4'h0 : _GEN_5341; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5343 = 10'h22e == _T_110[9:0] ? 4'h0 : _GEN_5342; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5344 = 10'h22f == _T_110[9:0] ? 4'h0 : _GEN_5343; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5345 = 10'h230 == _T_110[9:0] ? 4'h0 : _GEN_5344; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5346 = 10'h231 == _T_110[9:0] ? 4'h0 : _GEN_5345; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5347 = 10'h232 == _T_110[9:0] ? 4'h0 : _GEN_5346; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5348 = 10'h233 == _T_110[9:0] ? 4'h0 : _GEN_5347; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5349 = 10'h234 == _T_110[9:0] ? 4'h0 : _GEN_5348; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5350 = 10'h235 == _T_110[9:0] ? 4'h0 : _GEN_5349; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5351 = 10'h236 == _T_110[9:0] ? 4'h0 : _GEN_5350; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5352 = 10'h237 == _T_110[9:0] ? 4'h0 : _GEN_5351; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5353 = 10'h238 == _T_110[9:0] ? 4'h0 : _GEN_5352; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5354 = 10'h239 == _T_110[9:0] ? 4'h0 : _GEN_5353; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5355 = 10'h23a == _T_110[9:0] ? 4'h0 : _GEN_5354; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5356 = 10'h23b == _T_110[9:0] ? 4'h0 : _GEN_5355; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5357 = 10'h23c == _T_110[9:0] ? 4'h0 : _GEN_5356; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5358 = 10'h23d == _T_110[9:0] ? 4'h0 : _GEN_5357; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5359 = 10'h23e == _T_110[9:0] ? 4'h0 : _GEN_5358; // @[Filter.scala 191:142]
  wire [3:0] _GEN_5360 = 10'h23f == _T_110[9:0] ? 4'h0 : _GEN_5359; // @[Filter.scala 191:142]
  wire [7:0] _T_124 = _GEN_5360 * 4'ha; // @[Filter.scala 191:142]
  wire [10:0] _GEN_28315 = {{3'd0}, _T_124}; // @[Filter.scala 191:109]
  wire [10:0] _T_126 = _T_119 + _GEN_28315; // @[Filter.scala 191:109]
  wire [10:0] _T_127 = _T_126 / 11'h64; // @[Filter.scala 191:150]
  wire  _T_129 = _T_100 >= 6'h20; // @[Filter.scala 194:31]
  wire  _T_133 = _T_107 >= 32'h12; // @[Filter.scala 194:63]
  wire  _T_134 = _T_129 | _T_133; // @[Filter.scala 194:58]
  wire [10:0] _GEN_5937 = io_SPI_distort ? _T_127 : {{7'd0}, _GEN_4208}; // @[Filter.scala 196:35]
  wire [10:0] _GEN_5938 = _T_134 ? 11'h0 : _GEN_5937; // @[Filter.scala 194:80]
  wire [10:0] _GEN_6515 = io_SPI_distort ? _T_127 : {{7'd0}, _GEN_4784}; // @[Filter.scala 196:35]
  wire [10:0] _GEN_6516 = _T_134 ? 11'h0 : _GEN_6515; // @[Filter.scala 194:80]
  wire [10:0] _GEN_7093 = io_SPI_distort ? _T_127 : {{7'd0}, _GEN_5360}; // @[Filter.scala 196:35]
  wire [10:0] _GEN_7094 = _T_134 ? 11'h0 : _GEN_7093; // @[Filter.scala 194:80]
  wire [31:0] _T_162 = pixelIndex + 32'h2; // @[Filter.scala 189:31]
  wire [31:0] _GEN_2 = _T_162 % 32'h20; // @[Filter.scala 189:38]
  wire [5:0] _T_163 = _GEN_2[5:0]; // @[Filter.scala 189:38]
  wire [5:0] _T_165 = _T_163 + _GEN_28295; // @[Filter.scala 189:53]
  wire [5:0] _T_167 = _T_165 - 6'h1; // @[Filter.scala 189:69]
  wire [31:0] _T_170 = _T_162 / 32'h20; // @[Filter.scala 190:38]
  wire [31:0] _T_172 = _T_170 + _GEN_28296; // @[Filter.scala 190:53]
  wire [31:0] _T_174 = _T_172 - 32'h1; // @[Filter.scala 190:69]
  wire [37:0] _T_175 = _T_174 * 32'h20; // @[Filter.scala 191:42]
  wire [37:0] _GEN_28321 = {{32'd0}, _T_167}; // @[Filter.scala 191:57]
  wire [37:0] _T_177 = _T_175 + _GEN_28321; // @[Filter.scala 191:57]
  wire [3:0] _GEN_7098 = 10'h3 == _T_177[9:0] ? 4'h3 : 4'ha; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7099 = 10'h4 == _T_177[9:0] ? 4'ha : _GEN_7098; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7100 = 10'h5 == _T_177[9:0] ? 4'ha : _GEN_7099; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7101 = 10'h6 == _T_177[9:0] ? 4'ha : _GEN_7100; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7102 = 10'h7 == _T_177[9:0] ? 4'ha : _GEN_7101; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7103 = 10'h8 == _T_177[9:0] ? 4'ha : _GEN_7102; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7104 = 10'h9 == _T_177[9:0] ? 4'ha : _GEN_7103; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7105 = 10'ha == _T_177[9:0] ? 4'ha : _GEN_7104; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7106 = 10'hb == _T_177[9:0] ? 4'ha : _GEN_7105; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7107 = 10'hc == _T_177[9:0] ? 4'ha : _GEN_7106; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7108 = 10'hd == _T_177[9:0] ? 4'ha : _GEN_7107; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7109 = 10'he == _T_177[9:0] ? 4'ha : _GEN_7108; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7110 = 10'hf == _T_177[9:0] ? 4'ha : _GEN_7109; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7111 = 10'h10 == _T_177[9:0] ? 4'ha : _GEN_7110; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7112 = 10'h11 == _T_177[9:0] ? 4'ha : _GEN_7111; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7113 = 10'h12 == _T_177[9:0] ? 4'ha : _GEN_7112; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7114 = 10'h13 == _T_177[9:0] ? 4'ha : _GEN_7113; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7115 = 10'h14 == _T_177[9:0] ? 4'ha : _GEN_7114; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7116 = 10'h15 == _T_177[9:0] ? 4'ha : _GEN_7115; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7117 = 10'h16 == _T_177[9:0] ? 4'ha : _GEN_7116; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7118 = 10'h17 == _T_177[9:0] ? 4'ha : _GEN_7117; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7119 = 10'h18 == _T_177[9:0] ? 4'ha : _GEN_7118; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7120 = 10'h19 == _T_177[9:0] ? 4'ha : _GEN_7119; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7121 = 10'h1a == _T_177[9:0] ? 4'ha : _GEN_7120; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7122 = 10'h1b == _T_177[9:0] ? 4'ha : _GEN_7121; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7123 = 10'h1c == _T_177[9:0] ? 4'ha : _GEN_7122; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7124 = 10'h1d == _T_177[9:0] ? 4'ha : _GEN_7123; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7125 = 10'h1e == _T_177[9:0] ? 4'ha : _GEN_7124; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7126 = 10'h1f == _T_177[9:0] ? 4'h0 : _GEN_7125; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7127 = 10'h20 == _T_177[9:0] ? 4'ha : _GEN_7126; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7128 = 10'h21 == _T_177[9:0] ? 4'ha : _GEN_7127; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7129 = 10'h22 == _T_177[9:0] ? 4'ha : _GEN_7128; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7130 = 10'h23 == _T_177[9:0] ? 4'h3 : _GEN_7129; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7131 = 10'h24 == _T_177[9:0] ? 4'ha : _GEN_7130; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7132 = 10'h25 == _T_177[9:0] ? 4'ha : _GEN_7131; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7133 = 10'h26 == _T_177[9:0] ? 4'ha : _GEN_7132; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7134 = 10'h27 == _T_177[9:0] ? 4'h1 : _GEN_7133; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7135 = 10'h28 == _T_177[9:0] ? 4'h1 : _GEN_7134; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7136 = 10'h29 == _T_177[9:0] ? 4'ha : _GEN_7135; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7137 = 10'h2a == _T_177[9:0] ? 4'ha : _GEN_7136; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7138 = 10'h2b == _T_177[9:0] ? 4'ha : _GEN_7137; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7139 = 10'h2c == _T_177[9:0] ? 4'ha : _GEN_7138; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7140 = 10'h2d == _T_177[9:0] ? 4'ha : _GEN_7139; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7141 = 10'h2e == _T_177[9:0] ? 4'ha : _GEN_7140; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7142 = 10'h2f == _T_177[9:0] ? 4'ha : _GEN_7141; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7143 = 10'h30 == _T_177[9:0] ? 4'ha : _GEN_7142; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7144 = 10'h31 == _T_177[9:0] ? 4'ha : _GEN_7143; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7145 = 10'h32 == _T_177[9:0] ? 4'ha : _GEN_7144; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7146 = 10'h33 == _T_177[9:0] ? 4'ha : _GEN_7145; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7147 = 10'h34 == _T_177[9:0] ? 4'ha : _GEN_7146; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7148 = 10'h35 == _T_177[9:0] ? 4'ha : _GEN_7147; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7149 = 10'h36 == _T_177[9:0] ? 4'ha : _GEN_7148; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7150 = 10'h37 == _T_177[9:0] ? 4'h1 : _GEN_7149; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7151 = 10'h38 == _T_177[9:0] ? 4'h1 : _GEN_7150; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7152 = 10'h39 == _T_177[9:0] ? 4'ha : _GEN_7151; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7153 = 10'h3a == _T_177[9:0] ? 4'ha : _GEN_7152; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7154 = 10'h3b == _T_177[9:0] ? 4'ha : _GEN_7153; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7155 = 10'h3c == _T_177[9:0] ? 4'ha : _GEN_7154; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7156 = 10'h3d == _T_177[9:0] ? 4'h3 : _GEN_7155; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7157 = 10'h3e == _T_177[9:0] ? 4'ha : _GEN_7156; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7158 = 10'h3f == _T_177[9:0] ? 4'h0 : _GEN_7157; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7159 = 10'h40 == _T_177[9:0] ? 4'ha : _GEN_7158; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7160 = 10'h41 == _T_177[9:0] ? 4'ha : _GEN_7159; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7161 = 10'h42 == _T_177[9:0] ? 4'ha : _GEN_7160; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7162 = 10'h43 == _T_177[9:0] ? 4'h2 : _GEN_7161; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7163 = 10'h44 == _T_177[9:0] ? 4'h3 : _GEN_7162; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7164 = 10'h45 == _T_177[9:0] ? 4'h0 : _GEN_7163; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7165 = 10'h46 == _T_177[9:0] ? 4'h0 : _GEN_7164; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7166 = 10'h47 == _T_177[9:0] ? 4'h0 : _GEN_7165; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7167 = 10'h48 == _T_177[9:0] ? 4'h0 : _GEN_7166; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7168 = 10'h49 == _T_177[9:0] ? 4'ha : _GEN_7167; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7169 = 10'h4a == _T_177[9:0] ? 4'ha : _GEN_7168; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7170 = 10'h4b == _T_177[9:0] ? 4'ha : _GEN_7169; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7171 = 10'h4c == _T_177[9:0] ? 4'ha : _GEN_7170; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7172 = 10'h4d == _T_177[9:0] ? 4'ha : _GEN_7171; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7173 = 10'h4e == _T_177[9:0] ? 4'ha : _GEN_7172; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7174 = 10'h4f == _T_177[9:0] ? 4'ha : _GEN_7173; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7175 = 10'h50 == _T_177[9:0] ? 4'ha : _GEN_7174; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7176 = 10'h51 == _T_177[9:0] ? 4'ha : _GEN_7175; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7177 = 10'h52 == _T_177[9:0] ? 4'ha : _GEN_7176; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7178 = 10'h53 == _T_177[9:0] ? 4'ha : _GEN_7177; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7179 = 10'h54 == _T_177[9:0] ? 4'h1 : _GEN_7178; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7180 = 10'h55 == _T_177[9:0] ? 4'h1 : _GEN_7179; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7181 = 10'h56 == _T_177[9:0] ? 4'h1 : _GEN_7180; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7182 = 10'h57 == _T_177[9:0] ? 4'h0 : _GEN_7181; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7183 = 10'h58 == _T_177[9:0] ? 4'ha : _GEN_7182; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7184 = 10'h59 == _T_177[9:0] ? 4'h0 : _GEN_7183; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7185 = 10'h5a == _T_177[9:0] ? 4'ha : _GEN_7184; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7186 = 10'h5b == _T_177[9:0] ? 4'ha : _GEN_7185; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7187 = 10'h5c == _T_177[9:0] ? 4'ha : _GEN_7186; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7188 = 10'h5d == _T_177[9:0] ? 4'h3 : _GEN_7187; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7189 = 10'h5e == _T_177[9:0] ? 4'ha : _GEN_7188; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7190 = 10'h5f == _T_177[9:0] ? 4'h0 : _GEN_7189; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7191 = 10'h60 == _T_177[9:0] ? 4'ha : _GEN_7190; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7192 = 10'h61 == _T_177[9:0] ? 4'ha : _GEN_7191; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7193 = 10'h62 == _T_177[9:0] ? 4'ha : _GEN_7192; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7194 = 10'h63 == _T_177[9:0] ? 4'ha : _GEN_7193; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7195 = 10'h64 == _T_177[9:0] ? 4'h3 : _GEN_7194; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7196 = 10'h65 == _T_177[9:0] ? 4'h0 : _GEN_7195; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7197 = 10'h66 == _T_177[9:0] ? 4'ha : _GEN_7196; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7198 = 10'h67 == _T_177[9:0] ? 4'ha : _GEN_7197; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7199 = 10'h68 == _T_177[9:0] ? 4'ha : _GEN_7198; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7200 = 10'h69 == _T_177[9:0] ? 4'h0 : _GEN_7199; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7201 = 10'h6a == _T_177[9:0] ? 4'h1 : _GEN_7200; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7202 = 10'h6b == _T_177[9:0] ? 4'h1 : _GEN_7201; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7203 = 10'h6c == _T_177[9:0] ? 4'ha : _GEN_7202; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7204 = 10'h6d == _T_177[9:0] ? 4'ha : _GEN_7203; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7205 = 10'h6e == _T_177[9:0] ? 4'ha : _GEN_7204; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7206 = 10'h6f == _T_177[9:0] ? 4'ha : _GEN_7205; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7207 = 10'h70 == _T_177[9:0] ? 4'ha : _GEN_7206; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7208 = 10'h71 == _T_177[9:0] ? 4'ha : _GEN_7207; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7209 = 10'h72 == _T_177[9:0] ? 4'ha : _GEN_7208; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7210 = 10'h73 == _T_177[9:0] ? 4'h1 : _GEN_7209; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7211 = 10'h74 == _T_177[9:0] ? 4'h0 : _GEN_7210; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7212 = 10'h75 == _T_177[9:0] ? 4'h0 : _GEN_7211; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7213 = 10'h76 == _T_177[9:0] ? 4'h0 : _GEN_7212; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7214 = 10'h77 == _T_177[9:0] ? 4'ha : _GEN_7213; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7215 = 10'h78 == _T_177[9:0] ? 4'ha : _GEN_7214; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7216 = 10'h79 == _T_177[9:0] ? 4'ha : _GEN_7215; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7217 = 10'h7a == _T_177[9:0] ? 4'h0 : _GEN_7216; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7218 = 10'h7b == _T_177[9:0] ? 4'ha : _GEN_7217; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7219 = 10'h7c == _T_177[9:0] ? 4'ha : _GEN_7218; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7220 = 10'h7d == _T_177[9:0] ? 4'h2 : _GEN_7219; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7221 = 10'h7e == _T_177[9:0] ? 4'h3 : _GEN_7220; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7222 = 10'h7f == _T_177[9:0] ? 4'h0 : _GEN_7221; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7223 = 10'h80 == _T_177[9:0] ? 4'ha : _GEN_7222; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7224 = 10'h81 == _T_177[9:0] ? 4'ha : _GEN_7223; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7225 = 10'h82 == _T_177[9:0] ? 4'h1 : _GEN_7224; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7226 = 10'h83 == _T_177[9:0] ? 4'h0 : _GEN_7225; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7227 = 10'h84 == _T_177[9:0] ? 4'h2 : _GEN_7226; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7228 = 10'h85 == _T_177[9:0] ? 4'h1 : _GEN_7227; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7229 = 10'h86 == _T_177[9:0] ? 4'h1 : _GEN_7228; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7230 = 10'h87 == _T_177[9:0] ? 4'ha : _GEN_7229; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7231 = 10'h88 == _T_177[9:0] ? 4'ha : _GEN_7230; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7232 = 10'h89 == _T_177[9:0] ? 4'h0 : _GEN_7231; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7233 = 10'h8a == _T_177[9:0] ? 4'h0 : _GEN_7232; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7234 = 10'h8b == _T_177[9:0] ? 4'h1 : _GEN_7233; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7235 = 10'h8c == _T_177[9:0] ? 4'h1 : _GEN_7234; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7236 = 10'h8d == _T_177[9:0] ? 4'h1 : _GEN_7235; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7237 = 10'h8e == _T_177[9:0] ? 4'h1 : _GEN_7236; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7238 = 10'h8f == _T_177[9:0] ? 4'h1 : _GEN_7237; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7239 = 10'h90 == _T_177[9:0] ? 4'h1 : _GEN_7238; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7240 = 10'h91 == _T_177[9:0] ? 4'h1 : _GEN_7239; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7241 = 10'h92 == _T_177[9:0] ? 4'h1 : _GEN_7240; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7242 = 10'h93 == _T_177[9:0] ? 4'h0 : _GEN_7241; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7243 = 10'h94 == _T_177[9:0] ? 4'h0 : _GEN_7242; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7244 = 10'h95 == _T_177[9:0] ? 4'ha : _GEN_7243; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7245 = 10'h96 == _T_177[9:0] ? 4'ha : _GEN_7244; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7246 = 10'h97 == _T_177[9:0] ? 4'ha : _GEN_7245; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7247 = 10'h98 == _T_177[9:0] ? 4'h1 : _GEN_7246; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7248 = 10'h99 == _T_177[9:0] ? 4'h0 : _GEN_7247; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7249 = 10'h9a == _T_177[9:0] ? 4'h1 : _GEN_7248; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7250 = 10'h9b == _T_177[9:0] ? 4'h1 : _GEN_7249; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7251 = 10'h9c == _T_177[9:0] ? 4'ha : _GEN_7250; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7252 = 10'h9d == _T_177[9:0] ? 4'ha : _GEN_7251; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7253 = 10'h9e == _T_177[9:0] ? 4'h3 : _GEN_7252; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7254 = 10'h9f == _T_177[9:0] ? 4'h0 : _GEN_7253; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7255 = 10'ha0 == _T_177[9:0] ? 4'ha : _GEN_7254; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7256 = 10'ha1 == _T_177[9:0] ? 4'h1 : _GEN_7255; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7257 = 10'ha2 == _T_177[9:0] ? 4'h0 : _GEN_7256; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7258 = 10'ha3 == _T_177[9:0] ? 4'h3 : _GEN_7257; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7259 = 10'ha4 == _T_177[9:0] ? 4'ha : _GEN_7258; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7260 = 10'ha5 == _T_177[9:0] ? 4'ha : _GEN_7259; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7261 = 10'ha6 == _T_177[9:0] ? 4'ha : _GEN_7260; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7262 = 10'ha7 == _T_177[9:0] ? 4'h0 : _GEN_7261; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7263 = 10'ha8 == _T_177[9:0] ? 4'ha : _GEN_7262; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7264 = 10'ha9 == _T_177[9:0] ? 4'h1 : _GEN_7263; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7265 = 10'haa == _T_177[9:0] ? 4'h0 : _GEN_7264; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7266 = 10'hab == _T_177[9:0] ? 4'h0 : _GEN_7265; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7267 = 10'hac == _T_177[9:0] ? 4'h0 : _GEN_7266; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7268 = 10'had == _T_177[9:0] ? 4'h0 : _GEN_7267; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7269 = 10'hae == _T_177[9:0] ? 4'h0 : _GEN_7268; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7270 = 10'haf == _T_177[9:0] ? 4'h0 : _GEN_7269; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7271 = 10'hb0 == _T_177[9:0] ? 4'h0 : _GEN_7270; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7272 = 10'hb1 == _T_177[9:0] ? 4'h0 : _GEN_7271; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7273 = 10'hb2 == _T_177[9:0] ? 4'h0 : _GEN_7272; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7274 = 10'hb3 == _T_177[9:0] ? 4'h0 : _GEN_7273; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7275 = 10'hb4 == _T_177[9:0] ? 4'h1 : _GEN_7274; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7276 = 10'hb5 == _T_177[9:0] ? 4'h1 : _GEN_7275; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7277 = 10'hb6 == _T_177[9:0] ? 4'ha : _GEN_7276; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7278 = 10'hb7 == _T_177[9:0] ? 4'h0 : _GEN_7277; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7279 = 10'hb8 == _T_177[9:0] ? 4'ha : _GEN_7278; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7280 = 10'hb9 == _T_177[9:0] ? 4'ha : _GEN_7279; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7281 = 10'hba == _T_177[9:0] ? 4'ha : _GEN_7280; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7282 = 10'hbb == _T_177[9:0] ? 4'h0 : _GEN_7281; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7283 = 10'hbc == _T_177[9:0] ? 4'ha : _GEN_7282; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7284 = 10'hbd == _T_177[9:0] ? 4'ha : _GEN_7283; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7285 = 10'hbe == _T_177[9:0] ? 4'h3 : _GEN_7284; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7286 = 10'hbf == _T_177[9:0] ? 4'h0 : _GEN_7285; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7287 = 10'hc0 == _T_177[9:0] ? 4'ha : _GEN_7286; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7288 = 10'hc1 == _T_177[9:0] ? 4'ha : _GEN_7287; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7289 = 10'hc2 == _T_177[9:0] ? 4'h3 : _GEN_7288; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7290 = 10'hc3 == _T_177[9:0] ? 4'h2 : _GEN_7289; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7291 = 10'hc4 == _T_177[9:0] ? 4'h0 : _GEN_7290; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7292 = 10'hc5 == _T_177[9:0] ? 4'h0 : _GEN_7291; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7293 = 10'hc6 == _T_177[9:0] ? 4'h0 : _GEN_7292; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7294 = 10'hc7 == _T_177[9:0] ? 4'ha : _GEN_7293; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7295 = 10'hc8 == _T_177[9:0] ? 4'h1 : _GEN_7294; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7296 = 10'hc9 == _T_177[9:0] ? 4'h0 : _GEN_7295; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7297 = 10'hca == _T_177[9:0] ? 4'h0 : _GEN_7296; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7298 = 10'hcb == _T_177[9:0] ? 4'h0 : _GEN_7297; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7299 = 10'hcc == _T_177[9:0] ? 4'h0 : _GEN_7298; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7300 = 10'hcd == _T_177[9:0] ? 4'h0 : _GEN_7299; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7301 = 10'hce == _T_177[9:0] ? 4'h0 : _GEN_7300; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7302 = 10'hcf == _T_177[9:0] ? 4'h0 : _GEN_7301; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7303 = 10'hd0 == _T_177[9:0] ? 4'h0 : _GEN_7302; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7304 = 10'hd1 == _T_177[9:0] ? 4'h0 : _GEN_7303; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7305 = 10'hd2 == _T_177[9:0] ? 4'h0 : _GEN_7304; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7306 = 10'hd3 == _T_177[9:0] ? 4'h0 : _GEN_7305; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7307 = 10'hd4 == _T_177[9:0] ? 4'h0 : _GEN_7306; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7308 = 10'hd5 == _T_177[9:0] ? 4'h0 : _GEN_7307; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7309 = 10'hd6 == _T_177[9:0] ? 4'h1 : _GEN_7308; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7310 = 10'hd7 == _T_177[9:0] ? 4'ha : _GEN_7309; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7311 = 10'hd8 == _T_177[9:0] ? 4'h0 : _GEN_7310; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7312 = 10'hd9 == _T_177[9:0] ? 4'ha : _GEN_7311; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7313 = 10'hda == _T_177[9:0] ? 4'ha : _GEN_7312; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7314 = 10'hdb == _T_177[9:0] ? 4'ha : _GEN_7313; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7315 = 10'hdc == _T_177[9:0] ? 4'ha : _GEN_7314; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7316 = 10'hdd == _T_177[9:0] ? 4'h3 : _GEN_7315; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7317 = 10'hde == _T_177[9:0] ? 4'h2 : _GEN_7316; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7318 = 10'hdf == _T_177[9:0] ? 4'h0 : _GEN_7317; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7319 = 10'he0 == _T_177[9:0] ? 4'ha : _GEN_7318; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7320 = 10'he1 == _T_177[9:0] ? 4'ha : _GEN_7319; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7321 = 10'he2 == _T_177[9:0] ? 4'h3 : _GEN_7320; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7322 = 10'he3 == _T_177[9:0] ? 4'ha : _GEN_7321; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7323 = 10'he4 == _T_177[9:0] ? 4'ha : _GEN_7322; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7324 = 10'he5 == _T_177[9:0] ? 4'ha : _GEN_7323; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7325 = 10'he6 == _T_177[9:0] ? 4'ha : _GEN_7324; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7326 = 10'he7 == _T_177[9:0] ? 4'h1 : _GEN_7325; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7327 = 10'he8 == _T_177[9:0] ? 4'h1 : _GEN_7326; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7328 = 10'he9 == _T_177[9:0] ? 4'h1 : _GEN_7327; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7329 = 10'hea == _T_177[9:0] ? 4'h0 : _GEN_7328; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7330 = 10'heb == _T_177[9:0] ? 4'h0 : _GEN_7329; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7331 = 10'hec == _T_177[9:0] ? 4'h0 : _GEN_7330; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7332 = 10'hed == _T_177[9:0] ? 4'h0 : _GEN_7331; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7333 = 10'hee == _T_177[9:0] ? 4'h0 : _GEN_7332; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7334 = 10'hef == _T_177[9:0] ? 4'h0 : _GEN_7333; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7335 = 10'hf0 == _T_177[9:0] ? 4'h0 : _GEN_7334; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7336 = 10'hf1 == _T_177[9:0] ? 4'h0 : _GEN_7335; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7337 = 10'hf2 == _T_177[9:0] ? 4'h0 : _GEN_7336; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7338 = 10'hf3 == _T_177[9:0] ? 4'h0 : _GEN_7337; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7339 = 10'hf4 == _T_177[9:0] ? 4'h0 : _GEN_7338; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7340 = 10'hf5 == _T_177[9:0] ? 4'h1 : _GEN_7339; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7341 = 10'hf6 == _T_177[9:0] ? 4'h0 : _GEN_7340; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7342 = 10'hf7 == _T_177[9:0] ? 4'h0 : _GEN_7341; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7343 = 10'hf8 == _T_177[9:0] ? 4'h1 : _GEN_7342; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7344 = 10'hf9 == _T_177[9:0] ? 4'h0 : _GEN_7343; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7345 = 10'hfa == _T_177[9:0] ? 4'ha : _GEN_7344; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7346 = 10'hfb == _T_177[9:0] ? 4'ha : _GEN_7345; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7347 = 10'hfc == _T_177[9:0] ? 4'ha : _GEN_7346; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7348 = 10'hfd == _T_177[9:0] ? 4'h3 : _GEN_7347; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7349 = 10'hfe == _T_177[9:0] ? 4'ha : _GEN_7348; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7350 = 10'hff == _T_177[9:0] ? 4'h0 : _GEN_7349; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7351 = 10'h100 == _T_177[9:0] ? 4'ha : _GEN_7350; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7352 = 10'h101 == _T_177[9:0] ? 4'h0 : _GEN_7351; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7353 = 10'h102 == _T_177[9:0] ? 4'h3 : _GEN_7352; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7354 = 10'h103 == _T_177[9:0] ? 4'ha : _GEN_7353; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7355 = 10'h104 == _T_177[9:0] ? 4'ha : _GEN_7354; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7356 = 10'h105 == _T_177[9:0] ? 4'ha : _GEN_7355; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7357 = 10'h106 == _T_177[9:0] ? 4'ha : _GEN_7356; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7358 = 10'h107 == _T_177[9:0] ? 4'ha : _GEN_7357; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7359 = 10'h108 == _T_177[9:0] ? 4'h1 : _GEN_7358; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7360 = 10'h109 == _T_177[9:0] ? 4'h0 : _GEN_7359; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7361 = 10'h10a == _T_177[9:0] ? 4'h0 : _GEN_7360; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7362 = 10'h10b == _T_177[9:0] ? 4'h0 : _GEN_7361; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7363 = 10'h10c == _T_177[9:0] ? 4'h0 : _GEN_7362; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7364 = 10'h10d == _T_177[9:0] ? 4'h0 : _GEN_7363; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7365 = 10'h10e == _T_177[9:0] ? 4'h0 : _GEN_7364; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7366 = 10'h10f == _T_177[9:0] ? 4'h0 : _GEN_7365; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7367 = 10'h110 == _T_177[9:0] ? 4'h0 : _GEN_7366; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7368 = 10'h111 == _T_177[9:0] ? 4'h0 : _GEN_7367; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7369 = 10'h112 == _T_177[9:0] ? 4'h0 : _GEN_7368; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7370 = 10'h113 == _T_177[9:0] ? 4'h0 : _GEN_7369; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7371 = 10'h114 == _T_177[9:0] ? 4'h0 : _GEN_7370; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7372 = 10'h115 == _T_177[9:0] ? 4'h0 : _GEN_7371; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7373 = 10'h116 == _T_177[9:0] ? 4'h1 : _GEN_7372; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7374 = 10'h117 == _T_177[9:0] ? 4'ha : _GEN_7373; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7375 = 10'h118 == _T_177[9:0] ? 4'ha : _GEN_7374; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7376 = 10'h119 == _T_177[9:0] ? 4'ha : _GEN_7375; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7377 = 10'h11a == _T_177[9:0] ? 4'h0 : _GEN_7376; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7378 = 10'h11b == _T_177[9:0] ? 4'ha : _GEN_7377; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7379 = 10'h11c == _T_177[9:0] ? 4'ha : _GEN_7378; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7380 = 10'h11d == _T_177[9:0] ? 4'h2 : _GEN_7379; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7381 = 10'h11e == _T_177[9:0] ? 4'h3 : _GEN_7380; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7382 = 10'h11f == _T_177[9:0] ? 4'h0 : _GEN_7381; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7383 = 10'h120 == _T_177[9:0] ? 4'ha : _GEN_7382; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7384 = 10'h121 == _T_177[9:0] ? 4'ha : _GEN_7383; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7385 = 10'h122 == _T_177[9:0] ? 4'h3 : _GEN_7384; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7386 = 10'h123 == _T_177[9:0] ? 4'ha : _GEN_7385; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7387 = 10'h124 == _T_177[9:0] ? 4'ha : _GEN_7386; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7388 = 10'h125 == _T_177[9:0] ? 4'ha : _GEN_7387; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7389 = 10'h126 == _T_177[9:0] ? 4'ha : _GEN_7388; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7390 = 10'h127 == _T_177[9:0] ? 4'h1 : _GEN_7389; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7391 = 10'h128 == _T_177[9:0] ? 4'h0 : _GEN_7390; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7392 = 10'h129 == _T_177[9:0] ? 4'ha : _GEN_7391; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7393 = 10'h12a == _T_177[9:0] ? 4'ha : _GEN_7392; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7394 = 10'h12b == _T_177[9:0] ? 4'h0 : _GEN_7393; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7395 = 10'h12c == _T_177[9:0] ? 4'h0 : _GEN_7394; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7396 = 10'h12d == _T_177[9:0] ? 4'h0 : _GEN_7395; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7397 = 10'h12e == _T_177[9:0] ? 4'h0 : _GEN_7396; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7398 = 10'h12f == _T_177[9:0] ? 4'h0 : _GEN_7397; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7399 = 10'h130 == _T_177[9:0] ? 4'h0 : _GEN_7398; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7400 = 10'h131 == _T_177[9:0] ? 4'h0 : _GEN_7399; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7401 = 10'h132 == _T_177[9:0] ? 4'h0 : _GEN_7400; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7402 = 10'h133 == _T_177[9:0] ? 4'h0 : _GEN_7401; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7403 = 10'h134 == _T_177[9:0] ? 4'ha : _GEN_7402; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7404 = 10'h135 == _T_177[9:0] ? 4'ha : _GEN_7403; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7405 = 10'h136 == _T_177[9:0] ? 4'h0 : _GEN_7404; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7406 = 10'h137 == _T_177[9:0] ? 4'h1 : _GEN_7405; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7407 = 10'h138 == _T_177[9:0] ? 4'ha : _GEN_7406; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7408 = 10'h139 == _T_177[9:0] ? 4'ha : _GEN_7407; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7409 = 10'h13a == _T_177[9:0] ? 4'ha : _GEN_7408; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7410 = 10'h13b == _T_177[9:0] ? 4'ha : _GEN_7409; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7411 = 10'h13c == _T_177[9:0] ? 4'ha : _GEN_7410; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7412 = 10'h13d == _T_177[9:0] ? 4'ha : _GEN_7411; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7413 = 10'h13e == _T_177[9:0] ? 4'h3 : _GEN_7412; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7414 = 10'h13f == _T_177[9:0] ? 4'h0 : _GEN_7413; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7415 = 10'h140 == _T_177[9:0] ? 4'ha : _GEN_7414; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7416 = 10'h141 == _T_177[9:0] ? 4'ha : _GEN_7415; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7417 = 10'h142 == _T_177[9:0] ? 4'h2 : _GEN_7416; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7418 = 10'h143 == _T_177[9:0] ? 4'h3 : _GEN_7417; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7419 = 10'h144 == _T_177[9:0] ? 4'ha : _GEN_7418; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7420 = 10'h145 == _T_177[9:0] ? 4'ha : _GEN_7419; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7421 = 10'h146 == _T_177[9:0] ? 4'h1 : _GEN_7420; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7422 = 10'h147 == _T_177[9:0] ? 4'h0 : _GEN_7421; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7423 = 10'h148 == _T_177[9:0] ? 4'ha : _GEN_7422; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7424 = 10'h149 == _T_177[9:0] ? 4'ha : _GEN_7423; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7425 = 10'h14a == _T_177[9:0] ? 4'ha : _GEN_7424; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7426 = 10'h14b == _T_177[9:0] ? 4'ha : _GEN_7425; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7427 = 10'h14c == _T_177[9:0] ? 4'ha : _GEN_7426; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7428 = 10'h14d == _T_177[9:0] ? 4'ha : _GEN_7427; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7429 = 10'h14e == _T_177[9:0] ? 4'ha : _GEN_7428; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7430 = 10'h14f == _T_177[9:0] ? 4'ha : _GEN_7429; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7431 = 10'h150 == _T_177[9:0] ? 4'ha : _GEN_7430; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7432 = 10'h151 == _T_177[9:0] ? 4'ha : _GEN_7431; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7433 = 10'h152 == _T_177[9:0] ? 4'ha : _GEN_7432; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7434 = 10'h153 == _T_177[9:0] ? 4'ha : _GEN_7433; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7435 = 10'h154 == _T_177[9:0] ? 4'ha : _GEN_7434; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7436 = 10'h155 == _T_177[9:0] ? 4'ha : _GEN_7435; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7437 = 10'h156 == _T_177[9:0] ? 4'ha : _GEN_7436; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7438 = 10'h157 == _T_177[9:0] ? 4'h0 : _GEN_7437; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7439 = 10'h158 == _T_177[9:0] ? 4'ha : _GEN_7438; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7440 = 10'h159 == _T_177[9:0] ? 4'ha : _GEN_7439; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7441 = 10'h15a == _T_177[9:0] ? 4'ha : _GEN_7440; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7442 = 10'h15b == _T_177[9:0] ? 4'ha : _GEN_7441; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7443 = 10'h15c == _T_177[9:0] ? 4'ha : _GEN_7442; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7444 = 10'h15d == _T_177[9:0] ? 4'h3 : _GEN_7443; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7445 = 10'h15e == _T_177[9:0] ? 4'h2 : _GEN_7444; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7446 = 10'h15f == _T_177[9:0] ? 4'h0 : _GEN_7445; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7447 = 10'h160 == _T_177[9:0] ? 4'ha : _GEN_7446; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7448 = 10'h161 == _T_177[9:0] ? 4'ha : _GEN_7447; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7449 = 10'h162 == _T_177[9:0] ? 4'ha : _GEN_7448; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7450 = 10'h163 == _T_177[9:0] ? 4'h2 : _GEN_7449; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7451 = 10'h164 == _T_177[9:0] ? 4'h3 : _GEN_7450; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7452 = 10'h165 == _T_177[9:0] ? 4'h1 : _GEN_7451; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7453 = 10'h166 == _T_177[9:0] ? 4'h0 : _GEN_7452; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7454 = 10'h167 == _T_177[9:0] ? 4'h0 : _GEN_7453; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7455 = 10'h168 == _T_177[9:0] ? 4'h5 : _GEN_7454; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7456 = 10'h169 == _T_177[9:0] ? 4'h3 : _GEN_7455; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7457 = 10'h16a == _T_177[9:0] ? 4'h5 : _GEN_7456; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7458 = 10'h16b == _T_177[9:0] ? 4'h5 : _GEN_7457; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7459 = 10'h16c == _T_177[9:0] ? 4'ha : _GEN_7458; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7460 = 10'h16d == _T_177[9:0] ? 4'ha : _GEN_7459; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7461 = 10'h16e == _T_177[9:0] ? 4'ha : _GEN_7460; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7462 = 10'h16f == _T_177[9:0] ? 4'ha : _GEN_7461; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7463 = 10'h170 == _T_177[9:0] ? 4'ha : _GEN_7462; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7464 = 10'h171 == _T_177[9:0] ? 4'ha : _GEN_7463; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7465 = 10'h172 == _T_177[9:0] ? 4'ha : _GEN_7464; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7466 = 10'h173 == _T_177[9:0] ? 4'ha : _GEN_7465; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7467 = 10'h174 == _T_177[9:0] ? 4'ha : _GEN_7466; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7468 = 10'h175 == _T_177[9:0] ? 4'ha : _GEN_7467; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7469 = 10'h176 == _T_177[9:0] ? 4'h0 : _GEN_7468; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7470 = 10'h177 == _T_177[9:0] ? 4'h0 : _GEN_7469; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7471 = 10'h178 == _T_177[9:0] ? 4'h1 : _GEN_7470; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7472 = 10'h179 == _T_177[9:0] ? 4'ha : _GEN_7471; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7473 = 10'h17a == _T_177[9:0] ? 4'ha : _GEN_7472; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7474 = 10'h17b == _T_177[9:0] ? 4'ha : _GEN_7473; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7475 = 10'h17c == _T_177[9:0] ? 4'h3 : _GEN_7474; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7476 = 10'h17d == _T_177[9:0] ? 4'h2 : _GEN_7475; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7477 = 10'h17e == _T_177[9:0] ? 4'ha : _GEN_7476; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7478 = 10'h17f == _T_177[9:0] ? 4'h0 : _GEN_7477; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7479 = 10'h180 == _T_177[9:0] ? 4'h5 : _GEN_7478; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7480 = 10'h181 == _T_177[9:0] ? 4'h5 : _GEN_7479; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7481 = 10'h182 == _T_177[9:0] ? 4'h5 : _GEN_7480; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7482 = 10'h183 == _T_177[9:0] ? 4'h5 : _GEN_7481; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7483 = 10'h184 == _T_177[9:0] ? 4'h3 : _GEN_7482; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7484 = 10'h185 == _T_177[9:0] ? 4'h1 : _GEN_7483; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7485 = 10'h186 == _T_177[9:0] ? 4'hb : _GEN_7484; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7486 = 10'h187 == _T_177[9:0] ? 4'h0 : _GEN_7485; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7487 = 10'h188 == _T_177[9:0] ? 4'h5 : _GEN_7486; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7488 = 10'h189 == _T_177[9:0] ? 4'h5 : _GEN_7487; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7489 = 10'h18a == _T_177[9:0] ? 4'h5 : _GEN_7488; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7490 = 10'h18b == _T_177[9:0] ? 4'h5 : _GEN_7489; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7491 = 10'h18c == _T_177[9:0] ? 4'h5 : _GEN_7490; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7492 = 10'h18d == _T_177[9:0] ? 4'h5 : _GEN_7491; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7493 = 10'h18e == _T_177[9:0] ? 4'h5 : _GEN_7492; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7494 = 10'h18f == _T_177[9:0] ? 4'h5 : _GEN_7493; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7495 = 10'h190 == _T_177[9:0] ? 4'h5 : _GEN_7494; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7496 = 10'h191 == _T_177[9:0] ? 4'h5 : _GEN_7495; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7497 = 10'h192 == _T_177[9:0] ? 4'h3 : _GEN_7496; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7498 = 10'h193 == _T_177[9:0] ? 4'h5 : _GEN_7497; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7499 = 10'h194 == _T_177[9:0] ? 4'h5 : _GEN_7498; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7500 = 10'h195 == _T_177[9:0] ? 4'h5 : _GEN_7499; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7501 = 10'h196 == _T_177[9:0] ? 4'h0 : _GEN_7500; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7502 = 10'h197 == _T_177[9:0] ? 4'ha : _GEN_7501; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7503 = 10'h198 == _T_177[9:0] ? 4'h1 : _GEN_7502; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7504 = 10'h199 == _T_177[9:0] ? 4'ha : _GEN_7503; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7505 = 10'h19a == _T_177[9:0] ? 4'ha : _GEN_7504; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7506 = 10'h19b == _T_177[9:0] ? 4'ha : _GEN_7505; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7507 = 10'h19c == _T_177[9:0] ? 4'h3 : _GEN_7506; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7508 = 10'h19d == _T_177[9:0] ? 4'ha : _GEN_7507; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7509 = 10'h19e == _T_177[9:0] ? 4'ha : _GEN_7508; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7510 = 10'h19f == _T_177[9:0] ? 4'h0 : _GEN_7509; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7511 = 10'h1a0 == _T_177[9:0] ? 4'h5 : _GEN_7510; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7512 = 10'h1a1 == _T_177[9:0] ? 4'h5 : _GEN_7511; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7513 = 10'h1a2 == _T_177[9:0] ? 4'h3 : _GEN_7512; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7514 = 10'h1a3 == _T_177[9:0] ? 4'h5 : _GEN_7513; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7515 = 10'h1a4 == _T_177[9:0] ? 4'h3 : _GEN_7514; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7516 = 10'h1a5 == _T_177[9:0] ? 4'h0 : _GEN_7515; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7517 = 10'h1a6 == _T_177[9:0] ? 4'h5 : _GEN_7516; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7518 = 10'h1a7 == _T_177[9:0] ? 4'h0 : _GEN_7517; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7519 = 10'h1a8 == _T_177[9:0] ? 4'hb : _GEN_7518; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7520 = 10'h1a9 == _T_177[9:0] ? 4'h5 : _GEN_7519; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7521 = 10'h1aa == _T_177[9:0] ? 4'h5 : _GEN_7520; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7522 = 10'h1ab == _T_177[9:0] ? 4'h3 : _GEN_7521; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7523 = 10'h1ac == _T_177[9:0] ? 4'h5 : _GEN_7522; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7524 = 10'h1ad == _T_177[9:0] ? 4'h5 : _GEN_7523; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7525 = 10'h1ae == _T_177[9:0] ? 4'h5 : _GEN_7524; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7526 = 10'h1af == _T_177[9:0] ? 4'h5 : _GEN_7525; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7527 = 10'h1b0 == _T_177[9:0] ? 4'h5 : _GEN_7526; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7528 = 10'h1b1 == _T_177[9:0] ? 4'h5 : _GEN_7527; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7529 = 10'h1b2 == _T_177[9:0] ? 4'h5 : _GEN_7528; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7530 = 10'h1b3 == _T_177[9:0] ? 4'h5 : _GEN_7529; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7531 = 10'h1b4 == _T_177[9:0] ? 4'h5 : _GEN_7530; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7532 = 10'h1b5 == _T_177[9:0] ? 4'h5 : _GEN_7531; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7533 = 10'h1b6 == _T_177[9:0] ? 4'h0 : _GEN_7532; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7534 = 10'h1b7 == _T_177[9:0] ? 4'h5 : _GEN_7533; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7535 = 10'h1b8 == _T_177[9:0] ? 4'h0 : _GEN_7534; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7536 = 10'h1b9 == _T_177[9:0] ? 4'h5 : _GEN_7535; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7537 = 10'h1ba == _T_177[9:0] ? 4'h5 : _GEN_7536; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7538 = 10'h1bb == _T_177[9:0] ? 4'h5 : _GEN_7537; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7539 = 10'h1bc == _T_177[9:0] ? 4'h2 : _GEN_7538; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7540 = 10'h1bd == _T_177[9:0] ? 4'h3 : _GEN_7539; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7541 = 10'h1be == _T_177[9:0] ? 4'h5 : _GEN_7540; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7542 = 10'h1bf == _T_177[9:0] ? 4'h0 : _GEN_7541; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7543 = 10'h1c0 == _T_177[9:0] ? 4'h5 : _GEN_7542; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7544 = 10'h1c1 == _T_177[9:0] ? 4'h5 : _GEN_7543; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7545 = 10'h1c2 == _T_177[9:0] ? 4'h5 : _GEN_7544; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7546 = 10'h1c3 == _T_177[9:0] ? 4'h2 : _GEN_7545; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7547 = 10'h1c4 == _T_177[9:0] ? 4'h2 : _GEN_7546; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7548 = 10'h1c5 == _T_177[9:0] ? 4'h5 : _GEN_7547; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7549 = 10'h1c6 == _T_177[9:0] ? 4'h5 : _GEN_7548; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7550 = 10'h1c7 == _T_177[9:0] ? 4'h5 : _GEN_7549; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7551 = 10'h1c8 == _T_177[9:0] ? 4'h5 : _GEN_7550; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7552 = 10'h1c9 == _T_177[9:0] ? 4'hb : _GEN_7551; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7553 = 10'h1ca == _T_177[9:0] ? 4'hb : _GEN_7552; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7554 = 10'h1cb == _T_177[9:0] ? 4'hb : _GEN_7553; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7555 = 10'h1cc == _T_177[9:0] ? 4'hb : _GEN_7554; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7556 = 10'h1cd == _T_177[9:0] ? 4'hb : _GEN_7555; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7557 = 10'h1ce == _T_177[9:0] ? 4'hb : _GEN_7556; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7558 = 10'h1cf == _T_177[9:0] ? 4'hb : _GEN_7557; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7559 = 10'h1d0 == _T_177[9:0] ? 4'hb : _GEN_7558; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7560 = 10'h1d1 == _T_177[9:0] ? 4'hb : _GEN_7559; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7561 = 10'h1d2 == _T_177[9:0] ? 4'hb : _GEN_7560; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7562 = 10'h1d3 == _T_177[9:0] ? 4'hb : _GEN_7561; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7563 = 10'h1d4 == _T_177[9:0] ? 4'hb : _GEN_7562; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7564 = 10'h1d5 == _T_177[9:0] ? 4'hb : _GEN_7563; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7565 = 10'h1d6 == _T_177[9:0] ? 4'h5 : _GEN_7564; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7566 = 10'h1d7 == _T_177[9:0] ? 4'h5 : _GEN_7565; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7567 = 10'h1d8 == _T_177[9:0] ? 4'h5 : _GEN_7566; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7568 = 10'h1d9 == _T_177[9:0] ? 4'h5 : _GEN_7567; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7569 = 10'h1da == _T_177[9:0] ? 4'h5 : _GEN_7568; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7570 = 10'h1db == _T_177[9:0] ? 4'h5 : _GEN_7569; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7571 = 10'h1dc == _T_177[9:0] ? 4'h5 : _GEN_7570; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7572 = 10'h1dd == _T_177[9:0] ? 4'h3 : _GEN_7571; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7573 = 10'h1de == _T_177[9:0] ? 4'h5 : _GEN_7572; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7574 = 10'h1df == _T_177[9:0] ? 4'h0 : _GEN_7573; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7575 = 10'h1e0 == _T_177[9:0] ? 4'h3 : _GEN_7574; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7576 = 10'h1e1 == _T_177[9:0] ? 4'h5 : _GEN_7575; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7577 = 10'h1e2 == _T_177[9:0] ? 4'h2 : _GEN_7576; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7578 = 10'h1e3 == _T_177[9:0] ? 4'h2 : _GEN_7577; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7579 = 10'h1e4 == _T_177[9:0] ? 4'h5 : _GEN_7578; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7580 = 10'h1e5 == _T_177[9:0] ? 4'h5 : _GEN_7579; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7581 = 10'h1e6 == _T_177[9:0] ? 4'h5 : _GEN_7580; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7582 = 10'h1e7 == _T_177[9:0] ? 4'h5 : _GEN_7581; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7583 = 10'h1e8 == _T_177[9:0] ? 4'hb : _GEN_7582; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7584 = 10'h1e9 == _T_177[9:0] ? 4'h5 : _GEN_7583; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7585 = 10'h1ea == _T_177[9:0] ? 4'h5 : _GEN_7584; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7586 = 10'h1eb == _T_177[9:0] ? 4'hb : _GEN_7585; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7587 = 10'h1ec == _T_177[9:0] ? 4'h5 : _GEN_7586; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7588 = 10'h1ed == _T_177[9:0] ? 4'hb : _GEN_7587; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7589 = 10'h1ee == _T_177[9:0] ? 4'h5 : _GEN_7588; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7590 = 10'h1ef == _T_177[9:0] ? 4'hb : _GEN_7589; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7591 = 10'h1f0 == _T_177[9:0] ? 4'h5 : _GEN_7590; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7592 = 10'h1f1 == _T_177[9:0] ? 4'hb : _GEN_7591; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7593 = 10'h1f2 == _T_177[9:0] ? 4'hb : _GEN_7592; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7594 = 10'h1f3 == _T_177[9:0] ? 4'h5 : _GEN_7593; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7595 = 10'h1f4 == _T_177[9:0] ? 4'hb : _GEN_7594; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7596 = 10'h1f5 == _T_177[9:0] ? 4'hb : _GEN_7595; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7597 = 10'h1f6 == _T_177[9:0] ? 4'h5 : _GEN_7596; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7598 = 10'h1f7 == _T_177[9:0] ? 4'h5 : _GEN_7597; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7599 = 10'h1f8 == _T_177[9:0] ? 4'h5 : _GEN_7598; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7600 = 10'h1f9 == _T_177[9:0] ? 4'h5 : _GEN_7599; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7601 = 10'h1fa == _T_177[9:0] ? 4'h3 : _GEN_7600; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7602 = 10'h1fb == _T_177[9:0] ? 4'h5 : _GEN_7601; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7603 = 10'h1fc == _T_177[9:0] ? 4'h5 : _GEN_7602; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7604 = 10'h1fd == _T_177[9:0] ? 4'h2 : _GEN_7603; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7605 = 10'h1fe == _T_177[9:0] ? 4'h5 : _GEN_7604; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7606 = 10'h1ff == _T_177[9:0] ? 4'h0 : _GEN_7605; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7607 = 10'h200 == _T_177[9:0] ? 4'h5 : _GEN_7606; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7608 = 10'h201 == _T_177[9:0] ? 4'h5 : _GEN_7607; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7609 = 10'h202 == _T_177[9:0] ? 4'h3 : _GEN_7608; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7610 = 10'h203 == _T_177[9:0] ? 4'h5 : _GEN_7609; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7611 = 10'h204 == _T_177[9:0] ? 4'h5 : _GEN_7610; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7612 = 10'h205 == _T_177[9:0] ? 4'h5 : _GEN_7611; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7613 = 10'h206 == _T_177[9:0] ? 4'hb : _GEN_7612; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7614 = 10'h207 == _T_177[9:0] ? 4'hb : _GEN_7613; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7615 = 10'h208 == _T_177[9:0] ? 4'h5 : _GEN_7614; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7616 = 10'h209 == _T_177[9:0] ? 4'h5 : _GEN_7615; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7617 = 10'h20a == _T_177[9:0] ? 4'h5 : _GEN_7616; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7618 = 10'h20b == _T_177[9:0] ? 4'hb : _GEN_7617; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7619 = 10'h20c == _T_177[9:0] ? 4'h5 : _GEN_7618; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7620 = 10'h20d == _T_177[9:0] ? 4'hb : _GEN_7619; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7621 = 10'h20e == _T_177[9:0] ? 4'h5 : _GEN_7620; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7622 = 10'h20f == _T_177[9:0] ? 4'hb : _GEN_7621; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7623 = 10'h210 == _T_177[9:0] ? 4'h5 : _GEN_7622; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7624 = 10'h211 == _T_177[9:0] ? 4'h5 : _GEN_7623; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7625 = 10'h212 == _T_177[9:0] ? 4'hb : _GEN_7624; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7626 = 10'h213 == _T_177[9:0] ? 4'hb : _GEN_7625; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7627 = 10'h214 == _T_177[9:0] ? 4'hb : _GEN_7626; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7628 = 10'h215 == _T_177[9:0] ? 4'h5 : _GEN_7627; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7629 = 10'h216 == _T_177[9:0] ? 4'h5 : _GEN_7628; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7630 = 10'h217 == _T_177[9:0] ? 4'h5 : _GEN_7629; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7631 = 10'h218 == _T_177[9:0] ? 4'h5 : _GEN_7630; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7632 = 10'h219 == _T_177[9:0] ? 4'h5 : _GEN_7631; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7633 = 10'h21a == _T_177[9:0] ? 4'h5 : _GEN_7632; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7634 = 10'h21b == _T_177[9:0] ? 4'h5 : _GEN_7633; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7635 = 10'h21c == _T_177[9:0] ? 4'h3 : _GEN_7634; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7636 = 10'h21d == _T_177[9:0] ? 4'h2 : _GEN_7635; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7637 = 10'h21e == _T_177[9:0] ? 4'h5 : _GEN_7636; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7638 = 10'h21f == _T_177[9:0] ? 4'h0 : _GEN_7637; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7639 = 10'h220 == _T_177[9:0] ? 4'h0 : _GEN_7638; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7640 = 10'h221 == _T_177[9:0] ? 4'h0 : _GEN_7639; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7641 = 10'h222 == _T_177[9:0] ? 4'h0 : _GEN_7640; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7642 = 10'h223 == _T_177[9:0] ? 4'h0 : _GEN_7641; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7643 = 10'h224 == _T_177[9:0] ? 4'h0 : _GEN_7642; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7644 = 10'h225 == _T_177[9:0] ? 4'h0 : _GEN_7643; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7645 = 10'h226 == _T_177[9:0] ? 4'h0 : _GEN_7644; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7646 = 10'h227 == _T_177[9:0] ? 4'h0 : _GEN_7645; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7647 = 10'h228 == _T_177[9:0] ? 4'h0 : _GEN_7646; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7648 = 10'h229 == _T_177[9:0] ? 4'h0 : _GEN_7647; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7649 = 10'h22a == _T_177[9:0] ? 4'h0 : _GEN_7648; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7650 = 10'h22b == _T_177[9:0] ? 4'h0 : _GEN_7649; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7651 = 10'h22c == _T_177[9:0] ? 4'h0 : _GEN_7650; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7652 = 10'h22d == _T_177[9:0] ? 4'h0 : _GEN_7651; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7653 = 10'h22e == _T_177[9:0] ? 4'h0 : _GEN_7652; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7654 = 10'h22f == _T_177[9:0] ? 4'h0 : _GEN_7653; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7655 = 10'h230 == _T_177[9:0] ? 4'h0 : _GEN_7654; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7656 = 10'h231 == _T_177[9:0] ? 4'h0 : _GEN_7655; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7657 = 10'h232 == _T_177[9:0] ? 4'h0 : _GEN_7656; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7658 = 10'h233 == _T_177[9:0] ? 4'h0 : _GEN_7657; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7659 = 10'h234 == _T_177[9:0] ? 4'h0 : _GEN_7658; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7660 = 10'h235 == _T_177[9:0] ? 4'h0 : _GEN_7659; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7661 = 10'h236 == _T_177[9:0] ? 4'h0 : _GEN_7660; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7662 = 10'h237 == _T_177[9:0] ? 4'h0 : _GEN_7661; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7663 = 10'h238 == _T_177[9:0] ? 4'h0 : _GEN_7662; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7664 = 10'h239 == _T_177[9:0] ? 4'h0 : _GEN_7663; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7665 = 10'h23a == _T_177[9:0] ? 4'h0 : _GEN_7664; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7666 = 10'h23b == _T_177[9:0] ? 4'h0 : _GEN_7665; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7667 = 10'h23c == _T_177[9:0] ? 4'h0 : _GEN_7666; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7668 = 10'h23d == _T_177[9:0] ? 4'h0 : _GEN_7667; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7669 = 10'h23e == _T_177[9:0] ? 4'h0 : _GEN_7668; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7670 = 10'h23f == _T_177[9:0] ? 4'h0 : _GEN_7669; // @[Filter.scala 191:62]
  wire [4:0] _GEN_28322 = {{1'd0}, _GEN_7670}; // @[Filter.scala 191:62]
  wire [8:0] _T_179 = _GEN_28322 * 5'h14; // @[Filter.scala 191:62]
  wire [3:0] _GEN_7674 = 10'h3 == _T_177[9:0] ? 4'ha : 4'h3; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7675 = 10'h4 == _T_177[9:0] ? 4'h3 : _GEN_7674; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7676 = 10'h5 == _T_177[9:0] ? 4'h3 : _GEN_7675; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7677 = 10'h6 == _T_177[9:0] ? 4'h3 : _GEN_7676; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7678 = 10'h7 == _T_177[9:0] ? 4'h3 : _GEN_7677; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7679 = 10'h8 == _T_177[9:0] ? 4'h3 : _GEN_7678; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7680 = 10'h9 == _T_177[9:0] ? 4'h3 : _GEN_7679; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7681 = 10'ha == _T_177[9:0] ? 4'h3 : _GEN_7680; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7682 = 10'hb == _T_177[9:0] ? 4'h3 : _GEN_7681; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7683 = 10'hc == _T_177[9:0] ? 4'h5 : _GEN_7682; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7684 = 10'hd == _T_177[9:0] ? 4'h3 : _GEN_7683; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7685 = 10'he == _T_177[9:0] ? 4'h3 : _GEN_7684; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7686 = 10'hf == _T_177[9:0] ? 4'h3 : _GEN_7685; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7687 = 10'h10 == _T_177[9:0] ? 4'h3 : _GEN_7686; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7688 = 10'h11 == _T_177[9:0] ? 4'h3 : _GEN_7687; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7689 = 10'h12 == _T_177[9:0] ? 4'h3 : _GEN_7688; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7690 = 10'h13 == _T_177[9:0] ? 4'h3 : _GEN_7689; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7691 = 10'h14 == _T_177[9:0] ? 4'h3 : _GEN_7690; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7692 = 10'h15 == _T_177[9:0] ? 4'h3 : _GEN_7691; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7693 = 10'h16 == _T_177[9:0] ? 4'h3 : _GEN_7692; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7694 = 10'h17 == _T_177[9:0] ? 4'h3 : _GEN_7693; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7695 = 10'h18 == _T_177[9:0] ? 4'h3 : _GEN_7694; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7696 = 10'h19 == _T_177[9:0] ? 4'h3 : _GEN_7695; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7697 = 10'h1a == _T_177[9:0] ? 4'h3 : _GEN_7696; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7698 = 10'h1b == _T_177[9:0] ? 4'h3 : _GEN_7697; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7699 = 10'h1c == _T_177[9:0] ? 4'h3 : _GEN_7698; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7700 = 10'h1d == _T_177[9:0] ? 4'h3 : _GEN_7699; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7701 = 10'h1e == _T_177[9:0] ? 4'h3 : _GEN_7700; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7702 = 10'h1f == _T_177[9:0] ? 4'h0 : _GEN_7701; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7703 = 10'h20 == _T_177[9:0] ? 4'h3 : _GEN_7702; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7704 = 10'h21 == _T_177[9:0] ? 4'h5 : _GEN_7703; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7705 = 10'h22 == _T_177[9:0] ? 4'h3 : _GEN_7704; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7706 = 10'h23 == _T_177[9:0] ? 4'ha : _GEN_7705; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7707 = 10'h24 == _T_177[9:0] ? 4'h3 : _GEN_7706; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7708 = 10'h25 == _T_177[9:0] ? 4'h3 : _GEN_7707; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7709 = 10'h26 == _T_177[9:0] ? 4'h3 : _GEN_7708; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7710 = 10'h27 == _T_177[9:0] ? 4'h1 : _GEN_7709; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7711 = 10'h28 == _T_177[9:0] ? 4'h1 : _GEN_7710; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7712 = 10'h29 == _T_177[9:0] ? 4'h3 : _GEN_7711; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7713 = 10'h2a == _T_177[9:0] ? 4'h3 : _GEN_7712; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7714 = 10'h2b == _T_177[9:0] ? 4'h3 : _GEN_7713; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7715 = 10'h2c == _T_177[9:0] ? 4'h3 : _GEN_7714; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7716 = 10'h2d == _T_177[9:0] ? 4'h3 : _GEN_7715; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7717 = 10'h2e == _T_177[9:0] ? 4'h3 : _GEN_7716; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7718 = 10'h2f == _T_177[9:0] ? 4'h3 : _GEN_7717; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7719 = 10'h30 == _T_177[9:0] ? 4'h3 : _GEN_7718; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7720 = 10'h31 == _T_177[9:0] ? 4'h5 : _GEN_7719; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7721 = 10'h32 == _T_177[9:0] ? 4'h3 : _GEN_7720; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7722 = 10'h33 == _T_177[9:0] ? 4'h3 : _GEN_7721; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7723 = 10'h34 == _T_177[9:0] ? 4'h3 : _GEN_7722; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7724 = 10'h35 == _T_177[9:0] ? 4'h3 : _GEN_7723; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7725 = 10'h36 == _T_177[9:0] ? 4'h3 : _GEN_7724; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7726 = 10'h37 == _T_177[9:0] ? 4'h1 : _GEN_7725; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7727 = 10'h38 == _T_177[9:0] ? 4'h1 : _GEN_7726; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7728 = 10'h39 == _T_177[9:0] ? 4'h3 : _GEN_7727; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7729 = 10'h3a == _T_177[9:0] ? 4'h3 : _GEN_7728; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7730 = 10'h3b == _T_177[9:0] ? 4'h5 : _GEN_7729; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7731 = 10'h3c == _T_177[9:0] ? 4'h3 : _GEN_7730; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7732 = 10'h3d == _T_177[9:0] ? 4'ha : _GEN_7731; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7733 = 10'h3e == _T_177[9:0] ? 4'h3 : _GEN_7732; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7734 = 10'h3f == _T_177[9:0] ? 4'h0 : _GEN_7733; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7735 = 10'h40 == _T_177[9:0] ? 4'h3 : _GEN_7734; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7736 = 10'h41 == _T_177[9:0] ? 4'h3 : _GEN_7735; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7737 = 10'h42 == _T_177[9:0] ? 4'h3 : _GEN_7736; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7738 = 10'h43 == _T_177[9:0] ? 4'h7 : _GEN_7737; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7739 = 10'h44 == _T_177[9:0] ? 4'ha : _GEN_7738; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7740 = 10'h45 == _T_177[9:0] ? 4'h0 : _GEN_7739; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7741 = 10'h46 == _T_177[9:0] ? 4'h0 : _GEN_7740; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7742 = 10'h47 == _T_177[9:0] ? 4'h0 : _GEN_7741; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7743 = 10'h48 == _T_177[9:0] ? 4'h0 : _GEN_7742; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7744 = 10'h49 == _T_177[9:0] ? 4'h3 : _GEN_7743; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7745 = 10'h4a == _T_177[9:0] ? 4'h3 : _GEN_7744; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7746 = 10'h4b == _T_177[9:0] ? 4'h3 : _GEN_7745; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7747 = 10'h4c == _T_177[9:0] ? 4'h3 : _GEN_7746; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7748 = 10'h4d == _T_177[9:0] ? 4'h5 : _GEN_7747; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7749 = 10'h4e == _T_177[9:0] ? 4'h3 : _GEN_7748; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7750 = 10'h4f == _T_177[9:0] ? 4'h3 : _GEN_7749; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7751 = 10'h50 == _T_177[9:0] ? 4'h3 : _GEN_7750; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7752 = 10'h51 == _T_177[9:0] ? 4'h3 : _GEN_7751; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7753 = 10'h52 == _T_177[9:0] ? 4'h3 : _GEN_7752; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7754 = 10'h53 == _T_177[9:0] ? 4'h3 : _GEN_7753; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7755 = 10'h54 == _T_177[9:0] ? 4'h1 : _GEN_7754; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7756 = 10'h55 == _T_177[9:0] ? 4'h1 : _GEN_7755; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7757 = 10'h56 == _T_177[9:0] ? 4'h1 : _GEN_7756; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7758 = 10'h57 == _T_177[9:0] ? 4'h0 : _GEN_7757; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7759 = 10'h58 == _T_177[9:0] ? 4'h3 : _GEN_7758; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7760 = 10'h59 == _T_177[9:0] ? 4'h0 : _GEN_7759; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7761 = 10'h5a == _T_177[9:0] ? 4'h3 : _GEN_7760; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7762 = 10'h5b == _T_177[9:0] ? 4'h3 : _GEN_7761; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7763 = 10'h5c == _T_177[9:0] ? 4'h3 : _GEN_7762; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7764 = 10'h5d == _T_177[9:0] ? 4'ha : _GEN_7763; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7765 = 10'h5e == _T_177[9:0] ? 4'h3 : _GEN_7764; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7766 = 10'h5f == _T_177[9:0] ? 4'h0 : _GEN_7765; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7767 = 10'h60 == _T_177[9:0] ? 4'h3 : _GEN_7766; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7768 = 10'h61 == _T_177[9:0] ? 4'h3 : _GEN_7767; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7769 = 10'h62 == _T_177[9:0] ? 4'h3 : _GEN_7768; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7770 = 10'h63 == _T_177[9:0] ? 4'h3 : _GEN_7769; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7771 = 10'h64 == _T_177[9:0] ? 4'ha : _GEN_7770; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7772 = 10'h65 == _T_177[9:0] ? 4'h0 : _GEN_7771; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7773 = 10'h66 == _T_177[9:0] ? 4'h3 : _GEN_7772; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7774 = 10'h67 == _T_177[9:0] ? 4'h3 : _GEN_7773; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7775 = 10'h68 == _T_177[9:0] ? 4'h3 : _GEN_7774; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7776 = 10'h69 == _T_177[9:0] ? 4'h0 : _GEN_7775; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7777 = 10'h6a == _T_177[9:0] ? 4'h1 : _GEN_7776; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7778 = 10'h6b == _T_177[9:0] ? 4'h1 : _GEN_7777; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7779 = 10'h6c == _T_177[9:0] ? 4'h3 : _GEN_7778; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7780 = 10'h6d == _T_177[9:0] ? 4'h3 : _GEN_7779; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7781 = 10'h6e == _T_177[9:0] ? 4'h3 : _GEN_7780; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7782 = 10'h6f == _T_177[9:0] ? 4'h3 : _GEN_7781; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7783 = 10'h70 == _T_177[9:0] ? 4'h3 : _GEN_7782; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7784 = 10'h71 == _T_177[9:0] ? 4'h3 : _GEN_7783; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7785 = 10'h72 == _T_177[9:0] ? 4'h3 : _GEN_7784; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7786 = 10'h73 == _T_177[9:0] ? 4'h1 : _GEN_7785; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7787 = 10'h74 == _T_177[9:0] ? 4'h0 : _GEN_7786; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7788 = 10'h75 == _T_177[9:0] ? 4'h0 : _GEN_7787; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7789 = 10'h76 == _T_177[9:0] ? 4'h0 : _GEN_7788; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7790 = 10'h77 == _T_177[9:0] ? 4'h3 : _GEN_7789; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7791 = 10'h78 == _T_177[9:0] ? 4'h3 : _GEN_7790; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7792 = 10'h79 == _T_177[9:0] ? 4'h3 : _GEN_7791; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7793 = 10'h7a == _T_177[9:0] ? 4'h0 : _GEN_7792; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7794 = 10'h7b == _T_177[9:0] ? 4'h3 : _GEN_7793; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7795 = 10'h7c == _T_177[9:0] ? 4'h3 : _GEN_7794; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7796 = 10'h7d == _T_177[9:0] ? 4'h7 : _GEN_7795; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7797 = 10'h7e == _T_177[9:0] ? 4'ha : _GEN_7796; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7798 = 10'h7f == _T_177[9:0] ? 4'h0 : _GEN_7797; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7799 = 10'h80 == _T_177[9:0] ? 4'h3 : _GEN_7798; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7800 = 10'h81 == _T_177[9:0] ? 4'h3 : _GEN_7799; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7801 = 10'h82 == _T_177[9:0] ? 4'h1 : _GEN_7800; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7802 = 10'h83 == _T_177[9:0] ? 4'h0 : _GEN_7801; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7803 = 10'h84 == _T_177[9:0] ? 4'h7 : _GEN_7802; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7804 = 10'h85 == _T_177[9:0] ? 4'h1 : _GEN_7803; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7805 = 10'h86 == _T_177[9:0] ? 4'h1 : _GEN_7804; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7806 = 10'h87 == _T_177[9:0] ? 4'h3 : _GEN_7805; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7807 = 10'h88 == _T_177[9:0] ? 4'h3 : _GEN_7806; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7808 = 10'h89 == _T_177[9:0] ? 4'h0 : _GEN_7807; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7809 = 10'h8a == _T_177[9:0] ? 4'h0 : _GEN_7808; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7810 = 10'h8b == _T_177[9:0] ? 4'h1 : _GEN_7809; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7811 = 10'h8c == _T_177[9:0] ? 4'h1 : _GEN_7810; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7812 = 10'h8d == _T_177[9:0] ? 4'h1 : _GEN_7811; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7813 = 10'h8e == _T_177[9:0] ? 4'h1 : _GEN_7812; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7814 = 10'h8f == _T_177[9:0] ? 4'h1 : _GEN_7813; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7815 = 10'h90 == _T_177[9:0] ? 4'h1 : _GEN_7814; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7816 = 10'h91 == _T_177[9:0] ? 4'h1 : _GEN_7815; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7817 = 10'h92 == _T_177[9:0] ? 4'h1 : _GEN_7816; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7818 = 10'h93 == _T_177[9:0] ? 4'h0 : _GEN_7817; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7819 = 10'h94 == _T_177[9:0] ? 4'h0 : _GEN_7818; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7820 = 10'h95 == _T_177[9:0] ? 4'h3 : _GEN_7819; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7821 = 10'h96 == _T_177[9:0] ? 4'h3 : _GEN_7820; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7822 = 10'h97 == _T_177[9:0] ? 4'h3 : _GEN_7821; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7823 = 10'h98 == _T_177[9:0] ? 4'h1 : _GEN_7822; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7824 = 10'h99 == _T_177[9:0] ? 4'h0 : _GEN_7823; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7825 = 10'h9a == _T_177[9:0] ? 4'h1 : _GEN_7824; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7826 = 10'h9b == _T_177[9:0] ? 4'h1 : _GEN_7825; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7827 = 10'h9c == _T_177[9:0] ? 4'h3 : _GEN_7826; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7828 = 10'h9d == _T_177[9:0] ? 4'h3 : _GEN_7827; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7829 = 10'h9e == _T_177[9:0] ? 4'ha : _GEN_7828; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7830 = 10'h9f == _T_177[9:0] ? 4'h0 : _GEN_7829; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7831 = 10'ha0 == _T_177[9:0] ? 4'h3 : _GEN_7830; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7832 = 10'ha1 == _T_177[9:0] ? 4'h1 : _GEN_7831; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7833 = 10'ha2 == _T_177[9:0] ? 4'h0 : _GEN_7832; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7834 = 10'ha3 == _T_177[9:0] ? 4'ha : _GEN_7833; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7835 = 10'ha4 == _T_177[9:0] ? 4'h3 : _GEN_7834; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7836 = 10'ha5 == _T_177[9:0] ? 4'h3 : _GEN_7835; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7837 = 10'ha6 == _T_177[9:0] ? 4'h3 : _GEN_7836; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7838 = 10'ha7 == _T_177[9:0] ? 4'h0 : _GEN_7837; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7839 = 10'ha8 == _T_177[9:0] ? 4'h3 : _GEN_7838; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7840 = 10'ha9 == _T_177[9:0] ? 4'h1 : _GEN_7839; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7841 = 10'haa == _T_177[9:0] ? 4'h0 : _GEN_7840; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7842 = 10'hab == _T_177[9:0] ? 4'h0 : _GEN_7841; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7843 = 10'hac == _T_177[9:0] ? 4'h0 : _GEN_7842; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7844 = 10'had == _T_177[9:0] ? 4'h0 : _GEN_7843; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7845 = 10'hae == _T_177[9:0] ? 4'h0 : _GEN_7844; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7846 = 10'haf == _T_177[9:0] ? 4'h0 : _GEN_7845; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7847 = 10'hb0 == _T_177[9:0] ? 4'h0 : _GEN_7846; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7848 = 10'hb1 == _T_177[9:0] ? 4'h0 : _GEN_7847; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7849 = 10'hb2 == _T_177[9:0] ? 4'h0 : _GEN_7848; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7850 = 10'hb3 == _T_177[9:0] ? 4'h0 : _GEN_7849; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7851 = 10'hb4 == _T_177[9:0] ? 4'h1 : _GEN_7850; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7852 = 10'hb5 == _T_177[9:0] ? 4'h1 : _GEN_7851; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7853 = 10'hb6 == _T_177[9:0] ? 4'h3 : _GEN_7852; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7854 = 10'hb7 == _T_177[9:0] ? 4'h0 : _GEN_7853; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7855 = 10'hb8 == _T_177[9:0] ? 4'h3 : _GEN_7854; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7856 = 10'hb9 == _T_177[9:0] ? 4'h3 : _GEN_7855; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7857 = 10'hba == _T_177[9:0] ? 4'h3 : _GEN_7856; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7858 = 10'hbb == _T_177[9:0] ? 4'h0 : _GEN_7857; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7859 = 10'hbc == _T_177[9:0] ? 4'h3 : _GEN_7858; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7860 = 10'hbd == _T_177[9:0] ? 4'h3 : _GEN_7859; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7861 = 10'hbe == _T_177[9:0] ? 4'ha : _GEN_7860; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7862 = 10'hbf == _T_177[9:0] ? 4'h0 : _GEN_7861; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7863 = 10'hc0 == _T_177[9:0] ? 4'h3 : _GEN_7862; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7864 = 10'hc1 == _T_177[9:0] ? 4'h3 : _GEN_7863; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7865 = 10'hc2 == _T_177[9:0] ? 4'ha : _GEN_7864; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7866 = 10'hc3 == _T_177[9:0] ? 4'h7 : _GEN_7865; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7867 = 10'hc4 == _T_177[9:0] ? 4'h0 : _GEN_7866; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7868 = 10'hc5 == _T_177[9:0] ? 4'h0 : _GEN_7867; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7869 = 10'hc6 == _T_177[9:0] ? 4'h0 : _GEN_7868; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7870 = 10'hc7 == _T_177[9:0] ? 4'h3 : _GEN_7869; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7871 = 10'hc8 == _T_177[9:0] ? 4'h1 : _GEN_7870; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7872 = 10'hc9 == _T_177[9:0] ? 4'h0 : _GEN_7871; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7873 = 10'hca == _T_177[9:0] ? 4'h0 : _GEN_7872; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7874 = 10'hcb == _T_177[9:0] ? 4'h0 : _GEN_7873; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7875 = 10'hcc == _T_177[9:0] ? 4'h0 : _GEN_7874; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7876 = 10'hcd == _T_177[9:0] ? 4'h0 : _GEN_7875; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7877 = 10'hce == _T_177[9:0] ? 4'h0 : _GEN_7876; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7878 = 10'hcf == _T_177[9:0] ? 4'h0 : _GEN_7877; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7879 = 10'hd0 == _T_177[9:0] ? 4'h0 : _GEN_7878; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7880 = 10'hd1 == _T_177[9:0] ? 4'h0 : _GEN_7879; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7881 = 10'hd2 == _T_177[9:0] ? 4'h0 : _GEN_7880; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7882 = 10'hd3 == _T_177[9:0] ? 4'h0 : _GEN_7881; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7883 = 10'hd4 == _T_177[9:0] ? 4'h0 : _GEN_7882; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7884 = 10'hd5 == _T_177[9:0] ? 4'h0 : _GEN_7883; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7885 = 10'hd6 == _T_177[9:0] ? 4'h1 : _GEN_7884; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7886 = 10'hd7 == _T_177[9:0] ? 4'h3 : _GEN_7885; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7887 = 10'hd8 == _T_177[9:0] ? 4'h0 : _GEN_7886; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7888 = 10'hd9 == _T_177[9:0] ? 4'h3 : _GEN_7887; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7889 = 10'hda == _T_177[9:0] ? 4'h3 : _GEN_7888; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7890 = 10'hdb == _T_177[9:0] ? 4'h3 : _GEN_7889; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7891 = 10'hdc == _T_177[9:0] ? 4'h3 : _GEN_7890; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7892 = 10'hdd == _T_177[9:0] ? 4'ha : _GEN_7891; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7893 = 10'hde == _T_177[9:0] ? 4'h7 : _GEN_7892; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7894 = 10'hdf == _T_177[9:0] ? 4'h0 : _GEN_7893; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7895 = 10'he0 == _T_177[9:0] ? 4'h3 : _GEN_7894; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7896 = 10'he1 == _T_177[9:0] ? 4'h3 : _GEN_7895; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7897 = 10'he2 == _T_177[9:0] ? 4'ha : _GEN_7896; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7898 = 10'he3 == _T_177[9:0] ? 4'h3 : _GEN_7897; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7899 = 10'he4 == _T_177[9:0] ? 4'h3 : _GEN_7898; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7900 = 10'he5 == _T_177[9:0] ? 4'h3 : _GEN_7899; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7901 = 10'he6 == _T_177[9:0] ? 4'h3 : _GEN_7900; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7902 = 10'he7 == _T_177[9:0] ? 4'h1 : _GEN_7901; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7903 = 10'he8 == _T_177[9:0] ? 4'h1 : _GEN_7902; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7904 = 10'he9 == _T_177[9:0] ? 4'h1 : _GEN_7903; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7905 = 10'hea == _T_177[9:0] ? 4'h0 : _GEN_7904; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7906 = 10'heb == _T_177[9:0] ? 4'h0 : _GEN_7905; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7907 = 10'hec == _T_177[9:0] ? 4'h0 : _GEN_7906; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7908 = 10'hed == _T_177[9:0] ? 4'h0 : _GEN_7907; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7909 = 10'hee == _T_177[9:0] ? 4'h0 : _GEN_7908; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7910 = 10'hef == _T_177[9:0] ? 4'h0 : _GEN_7909; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7911 = 10'hf0 == _T_177[9:0] ? 4'h0 : _GEN_7910; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7912 = 10'hf1 == _T_177[9:0] ? 4'h0 : _GEN_7911; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7913 = 10'hf2 == _T_177[9:0] ? 4'h0 : _GEN_7912; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7914 = 10'hf3 == _T_177[9:0] ? 4'h0 : _GEN_7913; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7915 = 10'hf4 == _T_177[9:0] ? 4'h0 : _GEN_7914; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7916 = 10'hf5 == _T_177[9:0] ? 4'h1 : _GEN_7915; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7917 = 10'hf6 == _T_177[9:0] ? 4'h0 : _GEN_7916; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7918 = 10'hf7 == _T_177[9:0] ? 4'h0 : _GEN_7917; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7919 = 10'hf8 == _T_177[9:0] ? 4'h1 : _GEN_7918; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7920 = 10'hf9 == _T_177[9:0] ? 4'h0 : _GEN_7919; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7921 = 10'hfa == _T_177[9:0] ? 4'h3 : _GEN_7920; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7922 = 10'hfb == _T_177[9:0] ? 4'h3 : _GEN_7921; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7923 = 10'hfc == _T_177[9:0] ? 4'h3 : _GEN_7922; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7924 = 10'hfd == _T_177[9:0] ? 4'ha : _GEN_7923; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7925 = 10'hfe == _T_177[9:0] ? 4'h3 : _GEN_7924; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7926 = 10'hff == _T_177[9:0] ? 4'h0 : _GEN_7925; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7927 = 10'h100 == _T_177[9:0] ? 4'h3 : _GEN_7926; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7928 = 10'h101 == _T_177[9:0] ? 4'h0 : _GEN_7927; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7929 = 10'h102 == _T_177[9:0] ? 4'ha : _GEN_7928; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7930 = 10'h103 == _T_177[9:0] ? 4'h3 : _GEN_7929; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7931 = 10'h104 == _T_177[9:0] ? 4'h3 : _GEN_7930; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7932 = 10'h105 == _T_177[9:0] ? 4'h3 : _GEN_7931; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7933 = 10'h106 == _T_177[9:0] ? 4'h3 : _GEN_7932; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7934 = 10'h107 == _T_177[9:0] ? 4'h3 : _GEN_7933; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7935 = 10'h108 == _T_177[9:0] ? 4'h1 : _GEN_7934; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7936 = 10'h109 == _T_177[9:0] ? 4'h0 : _GEN_7935; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7937 = 10'h10a == _T_177[9:0] ? 4'h0 : _GEN_7936; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7938 = 10'h10b == _T_177[9:0] ? 4'h0 : _GEN_7937; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7939 = 10'h10c == _T_177[9:0] ? 4'h0 : _GEN_7938; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7940 = 10'h10d == _T_177[9:0] ? 4'h0 : _GEN_7939; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7941 = 10'h10e == _T_177[9:0] ? 4'h0 : _GEN_7940; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7942 = 10'h10f == _T_177[9:0] ? 4'h0 : _GEN_7941; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7943 = 10'h110 == _T_177[9:0] ? 4'h0 : _GEN_7942; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7944 = 10'h111 == _T_177[9:0] ? 4'h0 : _GEN_7943; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7945 = 10'h112 == _T_177[9:0] ? 4'h0 : _GEN_7944; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7946 = 10'h113 == _T_177[9:0] ? 4'h0 : _GEN_7945; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7947 = 10'h114 == _T_177[9:0] ? 4'h0 : _GEN_7946; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7948 = 10'h115 == _T_177[9:0] ? 4'h0 : _GEN_7947; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7949 = 10'h116 == _T_177[9:0] ? 4'h1 : _GEN_7948; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7950 = 10'h117 == _T_177[9:0] ? 4'h3 : _GEN_7949; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7951 = 10'h118 == _T_177[9:0] ? 4'h3 : _GEN_7950; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7952 = 10'h119 == _T_177[9:0] ? 4'h3 : _GEN_7951; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7953 = 10'h11a == _T_177[9:0] ? 4'h0 : _GEN_7952; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7954 = 10'h11b == _T_177[9:0] ? 4'h3 : _GEN_7953; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7955 = 10'h11c == _T_177[9:0] ? 4'h3 : _GEN_7954; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7956 = 10'h11d == _T_177[9:0] ? 4'h7 : _GEN_7955; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7957 = 10'h11e == _T_177[9:0] ? 4'ha : _GEN_7956; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7958 = 10'h11f == _T_177[9:0] ? 4'h0 : _GEN_7957; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7959 = 10'h120 == _T_177[9:0] ? 4'h3 : _GEN_7958; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7960 = 10'h121 == _T_177[9:0] ? 4'h3 : _GEN_7959; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7961 = 10'h122 == _T_177[9:0] ? 4'ha : _GEN_7960; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7962 = 10'h123 == _T_177[9:0] ? 4'h3 : _GEN_7961; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7963 = 10'h124 == _T_177[9:0] ? 4'h3 : _GEN_7962; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7964 = 10'h125 == _T_177[9:0] ? 4'h3 : _GEN_7963; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7965 = 10'h126 == _T_177[9:0] ? 4'h3 : _GEN_7964; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7966 = 10'h127 == _T_177[9:0] ? 4'h1 : _GEN_7965; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7967 = 10'h128 == _T_177[9:0] ? 4'h0 : _GEN_7966; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7968 = 10'h129 == _T_177[9:0] ? 4'h3 : _GEN_7967; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7969 = 10'h12a == _T_177[9:0] ? 4'h3 : _GEN_7968; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7970 = 10'h12b == _T_177[9:0] ? 4'h0 : _GEN_7969; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7971 = 10'h12c == _T_177[9:0] ? 4'h0 : _GEN_7970; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7972 = 10'h12d == _T_177[9:0] ? 4'h0 : _GEN_7971; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7973 = 10'h12e == _T_177[9:0] ? 4'h0 : _GEN_7972; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7974 = 10'h12f == _T_177[9:0] ? 4'h0 : _GEN_7973; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7975 = 10'h130 == _T_177[9:0] ? 4'h0 : _GEN_7974; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7976 = 10'h131 == _T_177[9:0] ? 4'h0 : _GEN_7975; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7977 = 10'h132 == _T_177[9:0] ? 4'h0 : _GEN_7976; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7978 = 10'h133 == _T_177[9:0] ? 4'h0 : _GEN_7977; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7979 = 10'h134 == _T_177[9:0] ? 4'h3 : _GEN_7978; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7980 = 10'h135 == _T_177[9:0] ? 4'h3 : _GEN_7979; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7981 = 10'h136 == _T_177[9:0] ? 4'h0 : _GEN_7980; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7982 = 10'h137 == _T_177[9:0] ? 4'h1 : _GEN_7981; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7983 = 10'h138 == _T_177[9:0] ? 4'h3 : _GEN_7982; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7984 = 10'h139 == _T_177[9:0] ? 4'h3 : _GEN_7983; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7985 = 10'h13a == _T_177[9:0] ? 4'h3 : _GEN_7984; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7986 = 10'h13b == _T_177[9:0] ? 4'h3 : _GEN_7985; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7987 = 10'h13c == _T_177[9:0] ? 4'h3 : _GEN_7986; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7988 = 10'h13d == _T_177[9:0] ? 4'h3 : _GEN_7987; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7989 = 10'h13e == _T_177[9:0] ? 4'ha : _GEN_7988; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7990 = 10'h13f == _T_177[9:0] ? 4'h0 : _GEN_7989; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7991 = 10'h140 == _T_177[9:0] ? 4'h5 : _GEN_7990; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7992 = 10'h141 == _T_177[9:0] ? 4'h3 : _GEN_7991; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7993 = 10'h142 == _T_177[9:0] ? 4'h7 : _GEN_7992; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7994 = 10'h143 == _T_177[9:0] ? 4'ha : _GEN_7993; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7995 = 10'h144 == _T_177[9:0] ? 4'h3 : _GEN_7994; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7996 = 10'h145 == _T_177[9:0] ? 4'h3 : _GEN_7995; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7997 = 10'h146 == _T_177[9:0] ? 4'h1 : _GEN_7996; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7998 = 10'h147 == _T_177[9:0] ? 4'h0 : _GEN_7997; // @[Filter.scala 191:102]
  wire [3:0] _GEN_7999 = 10'h148 == _T_177[9:0] ? 4'h3 : _GEN_7998; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8000 = 10'h149 == _T_177[9:0] ? 4'h3 : _GEN_7999; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8001 = 10'h14a == _T_177[9:0] ? 4'h3 : _GEN_8000; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8002 = 10'h14b == _T_177[9:0] ? 4'h3 : _GEN_8001; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8003 = 10'h14c == _T_177[9:0] ? 4'h3 : _GEN_8002; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8004 = 10'h14d == _T_177[9:0] ? 4'h3 : _GEN_8003; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8005 = 10'h14e == _T_177[9:0] ? 4'h3 : _GEN_8004; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8006 = 10'h14f == _T_177[9:0] ? 4'h3 : _GEN_8005; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8007 = 10'h150 == _T_177[9:0] ? 4'h3 : _GEN_8006; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8008 = 10'h151 == _T_177[9:0] ? 4'h3 : _GEN_8007; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8009 = 10'h152 == _T_177[9:0] ? 4'h3 : _GEN_8008; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8010 = 10'h153 == _T_177[9:0] ? 4'h3 : _GEN_8009; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8011 = 10'h154 == _T_177[9:0] ? 4'h3 : _GEN_8010; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8012 = 10'h155 == _T_177[9:0] ? 4'h3 : _GEN_8011; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8013 = 10'h156 == _T_177[9:0] ? 4'h3 : _GEN_8012; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8014 = 10'h157 == _T_177[9:0] ? 4'h0 : _GEN_8013; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8015 = 10'h158 == _T_177[9:0] ? 4'h3 : _GEN_8014; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8016 = 10'h159 == _T_177[9:0] ? 4'h3 : _GEN_8015; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8017 = 10'h15a == _T_177[9:0] ? 4'h3 : _GEN_8016; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8018 = 10'h15b == _T_177[9:0] ? 4'h3 : _GEN_8017; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8019 = 10'h15c == _T_177[9:0] ? 4'h3 : _GEN_8018; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8020 = 10'h15d == _T_177[9:0] ? 4'ha : _GEN_8019; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8021 = 10'h15e == _T_177[9:0] ? 4'h7 : _GEN_8020; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8022 = 10'h15f == _T_177[9:0] ? 4'h0 : _GEN_8021; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8023 = 10'h160 == _T_177[9:0] ? 4'h3 : _GEN_8022; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8024 = 10'h161 == _T_177[9:0] ? 4'h3 : _GEN_8023; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8025 = 10'h162 == _T_177[9:0] ? 4'h3 : _GEN_8024; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8026 = 10'h163 == _T_177[9:0] ? 4'h7 : _GEN_8025; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8027 = 10'h164 == _T_177[9:0] ? 4'ha : _GEN_8026; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8028 = 10'h165 == _T_177[9:0] ? 4'h1 : _GEN_8027; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8029 = 10'h166 == _T_177[9:0] ? 4'h0 : _GEN_8028; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8030 = 10'h167 == _T_177[9:0] ? 4'h0 : _GEN_8029; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8031 = 10'h168 == _T_177[9:0] ? 4'hc : _GEN_8030; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8032 = 10'h169 == _T_177[9:0] ? 4'h9 : _GEN_8031; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8033 = 10'h16a == _T_177[9:0] ? 4'hc : _GEN_8032; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8034 = 10'h16b == _T_177[9:0] ? 4'hc : _GEN_8033; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8035 = 10'h16c == _T_177[9:0] ? 4'h3 : _GEN_8034; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8036 = 10'h16d == _T_177[9:0] ? 4'h3 : _GEN_8035; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8037 = 10'h16e == _T_177[9:0] ? 4'h3 : _GEN_8036; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8038 = 10'h16f == _T_177[9:0] ? 4'h3 : _GEN_8037; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8039 = 10'h170 == _T_177[9:0] ? 4'h5 : _GEN_8038; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8040 = 10'h171 == _T_177[9:0] ? 4'h3 : _GEN_8039; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8041 = 10'h172 == _T_177[9:0] ? 4'h3 : _GEN_8040; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8042 = 10'h173 == _T_177[9:0] ? 4'h3 : _GEN_8041; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8043 = 10'h174 == _T_177[9:0] ? 4'h3 : _GEN_8042; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8044 = 10'h175 == _T_177[9:0] ? 4'h3 : _GEN_8043; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8045 = 10'h176 == _T_177[9:0] ? 4'h0 : _GEN_8044; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8046 = 10'h177 == _T_177[9:0] ? 4'h0 : _GEN_8045; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8047 = 10'h178 == _T_177[9:0] ? 4'h1 : _GEN_8046; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8048 = 10'h179 == _T_177[9:0] ? 4'h3 : _GEN_8047; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8049 = 10'h17a == _T_177[9:0] ? 4'h5 : _GEN_8048; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8050 = 10'h17b == _T_177[9:0] ? 4'h3 : _GEN_8049; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8051 = 10'h17c == _T_177[9:0] ? 4'ha : _GEN_8050; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8052 = 10'h17d == _T_177[9:0] ? 4'h7 : _GEN_8051; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8053 = 10'h17e == _T_177[9:0] ? 4'h3 : _GEN_8052; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8054 = 10'h17f == _T_177[9:0] ? 4'h0 : _GEN_8053; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8055 = 10'h180 == _T_177[9:0] ? 4'hc : _GEN_8054; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8056 = 10'h181 == _T_177[9:0] ? 4'hc : _GEN_8055; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8057 = 10'h182 == _T_177[9:0] ? 4'hc : _GEN_8056; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8058 = 10'h183 == _T_177[9:0] ? 4'hc : _GEN_8057; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8059 = 10'h184 == _T_177[9:0] ? 4'ha : _GEN_8058; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8060 = 10'h185 == _T_177[9:0] ? 4'h1 : _GEN_8059; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8061 = 10'h186 == _T_177[9:0] ? 4'hc : _GEN_8060; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8062 = 10'h187 == _T_177[9:0] ? 4'h0 : _GEN_8061; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8063 = 10'h188 == _T_177[9:0] ? 4'hc : _GEN_8062; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8064 = 10'h189 == _T_177[9:0] ? 4'hc : _GEN_8063; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8065 = 10'h18a == _T_177[9:0] ? 4'hc : _GEN_8064; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8066 = 10'h18b == _T_177[9:0] ? 4'hc : _GEN_8065; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8067 = 10'h18c == _T_177[9:0] ? 4'hc : _GEN_8066; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8068 = 10'h18d == _T_177[9:0] ? 4'hc : _GEN_8067; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8069 = 10'h18e == _T_177[9:0] ? 4'hc : _GEN_8068; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8070 = 10'h18f == _T_177[9:0] ? 4'hc : _GEN_8069; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8071 = 10'h190 == _T_177[9:0] ? 4'hc : _GEN_8070; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8072 = 10'h191 == _T_177[9:0] ? 4'hc : _GEN_8071; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8073 = 10'h192 == _T_177[9:0] ? 4'h9 : _GEN_8072; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8074 = 10'h193 == _T_177[9:0] ? 4'hc : _GEN_8073; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8075 = 10'h194 == _T_177[9:0] ? 4'hc : _GEN_8074; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8076 = 10'h195 == _T_177[9:0] ? 4'hc : _GEN_8075; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8077 = 10'h196 == _T_177[9:0] ? 4'h0 : _GEN_8076; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8078 = 10'h197 == _T_177[9:0] ? 4'h3 : _GEN_8077; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8079 = 10'h198 == _T_177[9:0] ? 4'h1 : _GEN_8078; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8080 = 10'h199 == _T_177[9:0] ? 4'h3 : _GEN_8079; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8081 = 10'h19a == _T_177[9:0] ? 4'h3 : _GEN_8080; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8082 = 10'h19b == _T_177[9:0] ? 4'h3 : _GEN_8081; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8083 = 10'h19c == _T_177[9:0] ? 4'ha : _GEN_8082; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8084 = 10'h19d == _T_177[9:0] ? 4'h3 : _GEN_8083; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8085 = 10'h19e == _T_177[9:0] ? 4'h3 : _GEN_8084; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8086 = 10'h19f == _T_177[9:0] ? 4'h0 : _GEN_8085; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8087 = 10'h1a0 == _T_177[9:0] ? 4'hc : _GEN_8086; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8088 = 10'h1a1 == _T_177[9:0] ? 4'hc : _GEN_8087; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8089 = 10'h1a2 == _T_177[9:0] ? 4'h9 : _GEN_8088; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8090 = 10'h1a3 == _T_177[9:0] ? 4'hc : _GEN_8089; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8091 = 10'h1a4 == _T_177[9:0] ? 4'ha : _GEN_8090; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8092 = 10'h1a5 == _T_177[9:0] ? 4'h0 : _GEN_8091; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8093 = 10'h1a6 == _T_177[9:0] ? 4'hc : _GEN_8092; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8094 = 10'h1a7 == _T_177[9:0] ? 4'h0 : _GEN_8093; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8095 = 10'h1a8 == _T_177[9:0] ? 4'hc : _GEN_8094; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8096 = 10'h1a9 == _T_177[9:0] ? 4'hc : _GEN_8095; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8097 = 10'h1aa == _T_177[9:0] ? 4'hc : _GEN_8096; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8098 = 10'h1ab == _T_177[9:0] ? 4'h9 : _GEN_8097; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8099 = 10'h1ac == _T_177[9:0] ? 4'hc : _GEN_8098; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8100 = 10'h1ad == _T_177[9:0] ? 4'hc : _GEN_8099; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8101 = 10'h1ae == _T_177[9:0] ? 4'hc : _GEN_8100; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8102 = 10'h1af == _T_177[9:0] ? 4'hc : _GEN_8101; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8103 = 10'h1b0 == _T_177[9:0] ? 4'hc : _GEN_8102; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8104 = 10'h1b1 == _T_177[9:0] ? 4'hc : _GEN_8103; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8105 = 10'h1b2 == _T_177[9:0] ? 4'hc : _GEN_8104; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8106 = 10'h1b3 == _T_177[9:0] ? 4'hc : _GEN_8105; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8107 = 10'h1b4 == _T_177[9:0] ? 4'hc : _GEN_8106; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8108 = 10'h1b5 == _T_177[9:0] ? 4'hc : _GEN_8107; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8109 = 10'h1b6 == _T_177[9:0] ? 4'h0 : _GEN_8108; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8110 = 10'h1b7 == _T_177[9:0] ? 4'hc : _GEN_8109; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8111 = 10'h1b8 == _T_177[9:0] ? 4'h0 : _GEN_8110; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8112 = 10'h1b9 == _T_177[9:0] ? 4'hc : _GEN_8111; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8113 = 10'h1ba == _T_177[9:0] ? 4'hc : _GEN_8112; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8114 = 10'h1bb == _T_177[9:0] ? 4'hc : _GEN_8113; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8115 = 10'h1bc == _T_177[9:0] ? 4'h7 : _GEN_8114; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8116 = 10'h1bd == _T_177[9:0] ? 4'ha : _GEN_8115; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8117 = 10'h1be == _T_177[9:0] ? 4'hc : _GEN_8116; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8118 = 10'h1bf == _T_177[9:0] ? 4'h0 : _GEN_8117; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8119 = 10'h1c0 == _T_177[9:0] ? 4'hc : _GEN_8118; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8120 = 10'h1c1 == _T_177[9:0] ? 4'hc : _GEN_8119; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8121 = 10'h1c2 == _T_177[9:0] ? 4'hc : _GEN_8120; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8122 = 10'h1c3 == _T_177[9:0] ? 4'h7 : _GEN_8121; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8123 = 10'h1c4 == _T_177[9:0] ? 4'h7 : _GEN_8122; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8124 = 10'h1c5 == _T_177[9:0] ? 4'hc : _GEN_8123; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8125 = 10'h1c6 == _T_177[9:0] ? 4'hc : _GEN_8124; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8126 = 10'h1c7 == _T_177[9:0] ? 4'hc : _GEN_8125; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8127 = 10'h1c8 == _T_177[9:0] ? 4'hc : _GEN_8126; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8128 = 10'h1c9 == _T_177[9:0] ? 4'hc : _GEN_8127; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8129 = 10'h1ca == _T_177[9:0] ? 4'hc : _GEN_8128; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8130 = 10'h1cb == _T_177[9:0] ? 4'hc : _GEN_8129; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8131 = 10'h1cc == _T_177[9:0] ? 4'hc : _GEN_8130; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8132 = 10'h1cd == _T_177[9:0] ? 4'hc : _GEN_8131; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8133 = 10'h1ce == _T_177[9:0] ? 4'hc : _GEN_8132; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8134 = 10'h1cf == _T_177[9:0] ? 4'hc : _GEN_8133; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8135 = 10'h1d0 == _T_177[9:0] ? 4'hc : _GEN_8134; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8136 = 10'h1d1 == _T_177[9:0] ? 4'hc : _GEN_8135; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8137 = 10'h1d2 == _T_177[9:0] ? 4'hc : _GEN_8136; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8138 = 10'h1d3 == _T_177[9:0] ? 4'hc : _GEN_8137; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8139 = 10'h1d4 == _T_177[9:0] ? 4'hc : _GEN_8138; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8140 = 10'h1d5 == _T_177[9:0] ? 4'hc : _GEN_8139; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8141 = 10'h1d6 == _T_177[9:0] ? 4'hc : _GEN_8140; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8142 = 10'h1d7 == _T_177[9:0] ? 4'hc : _GEN_8141; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8143 = 10'h1d8 == _T_177[9:0] ? 4'hc : _GEN_8142; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8144 = 10'h1d9 == _T_177[9:0] ? 4'hc : _GEN_8143; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8145 = 10'h1da == _T_177[9:0] ? 4'hc : _GEN_8144; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8146 = 10'h1db == _T_177[9:0] ? 4'hc : _GEN_8145; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8147 = 10'h1dc == _T_177[9:0] ? 4'hc : _GEN_8146; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8148 = 10'h1dd == _T_177[9:0] ? 4'ha : _GEN_8147; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8149 = 10'h1de == _T_177[9:0] ? 4'hc : _GEN_8148; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8150 = 10'h1df == _T_177[9:0] ? 4'h0 : _GEN_8149; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8151 = 10'h1e0 == _T_177[9:0] ? 4'h9 : _GEN_8150; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8152 = 10'h1e1 == _T_177[9:0] ? 4'hc : _GEN_8151; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8153 = 10'h1e2 == _T_177[9:0] ? 4'h7 : _GEN_8152; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8154 = 10'h1e3 == _T_177[9:0] ? 4'h7 : _GEN_8153; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8155 = 10'h1e4 == _T_177[9:0] ? 4'hc : _GEN_8154; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8156 = 10'h1e5 == _T_177[9:0] ? 4'hc : _GEN_8155; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8157 = 10'h1e6 == _T_177[9:0] ? 4'hc : _GEN_8156; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8158 = 10'h1e7 == _T_177[9:0] ? 4'hc : _GEN_8157; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8159 = 10'h1e8 == _T_177[9:0] ? 4'hc : _GEN_8158; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8160 = 10'h1e9 == _T_177[9:0] ? 4'hc : _GEN_8159; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8161 = 10'h1ea == _T_177[9:0] ? 4'hc : _GEN_8160; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8162 = 10'h1eb == _T_177[9:0] ? 4'hc : _GEN_8161; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8163 = 10'h1ec == _T_177[9:0] ? 4'hc : _GEN_8162; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8164 = 10'h1ed == _T_177[9:0] ? 4'hc : _GEN_8163; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8165 = 10'h1ee == _T_177[9:0] ? 4'hc : _GEN_8164; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8166 = 10'h1ef == _T_177[9:0] ? 4'hc : _GEN_8165; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8167 = 10'h1f0 == _T_177[9:0] ? 4'hc : _GEN_8166; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8168 = 10'h1f1 == _T_177[9:0] ? 4'hc : _GEN_8167; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8169 = 10'h1f2 == _T_177[9:0] ? 4'hc : _GEN_8168; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8170 = 10'h1f3 == _T_177[9:0] ? 4'hc : _GEN_8169; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8171 = 10'h1f4 == _T_177[9:0] ? 4'hc : _GEN_8170; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8172 = 10'h1f5 == _T_177[9:0] ? 4'hc : _GEN_8171; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8173 = 10'h1f6 == _T_177[9:0] ? 4'hc : _GEN_8172; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8174 = 10'h1f7 == _T_177[9:0] ? 4'hc : _GEN_8173; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8175 = 10'h1f8 == _T_177[9:0] ? 4'hc : _GEN_8174; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8176 = 10'h1f9 == _T_177[9:0] ? 4'hc : _GEN_8175; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8177 = 10'h1fa == _T_177[9:0] ? 4'h9 : _GEN_8176; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8178 = 10'h1fb == _T_177[9:0] ? 4'hc : _GEN_8177; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8179 = 10'h1fc == _T_177[9:0] ? 4'hc : _GEN_8178; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8180 = 10'h1fd == _T_177[9:0] ? 4'h7 : _GEN_8179; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8181 = 10'h1fe == _T_177[9:0] ? 4'hc : _GEN_8180; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8182 = 10'h1ff == _T_177[9:0] ? 4'h0 : _GEN_8181; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8183 = 10'h200 == _T_177[9:0] ? 4'hc : _GEN_8182; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8184 = 10'h201 == _T_177[9:0] ? 4'hc : _GEN_8183; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8185 = 10'h202 == _T_177[9:0] ? 4'ha : _GEN_8184; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8186 = 10'h203 == _T_177[9:0] ? 4'hc : _GEN_8185; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8187 = 10'h204 == _T_177[9:0] ? 4'hc : _GEN_8186; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8188 = 10'h205 == _T_177[9:0] ? 4'hc : _GEN_8187; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8189 = 10'h206 == _T_177[9:0] ? 4'hc : _GEN_8188; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8190 = 10'h207 == _T_177[9:0] ? 4'hc : _GEN_8189; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8191 = 10'h208 == _T_177[9:0] ? 4'hc : _GEN_8190; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8192 = 10'h209 == _T_177[9:0] ? 4'hc : _GEN_8191; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8193 = 10'h20a == _T_177[9:0] ? 4'hc : _GEN_8192; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8194 = 10'h20b == _T_177[9:0] ? 4'hc : _GEN_8193; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8195 = 10'h20c == _T_177[9:0] ? 4'hc : _GEN_8194; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8196 = 10'h20d == _T_177[9:0] ? 4'hc : _GEN_8195; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8197 = 10'h20e == _T_177[9:0] ? 4'hc : _GEN_8196; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8198 = 10'h20f == _T_177[9:0] ? 4'hc : _GEN_8197; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8199 = 10'h210 == _T_177[9:0] ? 4'hc : _GEN_8198; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8200 = 10'h211 == _T_177[9:0] ? 4'hc : _GEN_8199; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8201 = 10'h212 == _T_177[9:0] ? 4'hc : _GEN_8200; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8202 = 10'h213 == _T_177[9:0] ? 4'hc : _GEN_8201; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8203 = 10'h214 == _T_177[9:0] ? 4'hc : _GEN_8202; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8204 = 10'h215 == _T_177[9:0] ? 4'hc : _GEN_8203; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8205 = 10'h216 == _T_177[9:0] ? 4'hc : _GEN_8204; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8206 = 10'h217 == _T_177[9:0] ? 4'hc : _GEN_8205; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8207 = 10'h218 == _T_177[9:0] ? 4'hc : _GEN_8206; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8208 = 10'h219 == _T_177[9:0] ? 4'hc : _GEN_8207; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8209 = 10'h21a == _T_177[9:0] ? 4'hc : _GEN_8208; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8210 = 10'h21b == _T_177[9:0] ? 4'hc : _GEN_8209; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8211 = 10'h21c == _T_177[9:0] ? 4'ha : _GEN_8210; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8212 = 10'h21d == _T_177[9:0] ? 4'h7 : _GEN_8211; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8213 = 10'h21e == _T_177[9:0] ? 4'hc : _GEN_8212; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8214 = 10'h21f == _T_177[9:0] ? 4'h0 : _GEN_8213; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8215 = 10'h220 == _T_177[9:0] ? 4'h0 : _GEN_8214; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8216 = 10'h221 == _T_177[9:0] ? 4'h0 : _GEN_8215; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8217 = 10'h222 == _T_177[9:0] ? 4'h0 : _GEN_8216; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8218 = 10'h223 == _T_177[9:0] ? 4'h0 : _GEN_8217; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8219 = 10'h224 == _T_177[9:0] ? 4'h0 : _GEN_8218; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8220 = 10'h225 == _T_177[9:0] ? 4'h0 : _GEN_8219; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8221 = 10'h226 == _T_177[9:0] ? 4'h0 : _GEN_8220; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8222 = 10'h227 == _T_177[9:0] ? 4'h0 : _GEN_8221; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8223 = 10'h228 == _T_177[9:0] ? 4'h0 : _GEN_8222; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8224 = 10'h229 == _T_177[9:0] ? 4'h0 : _GEN_8223; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8225 = 10'h22a == _T_177[9:0] ? 4'h0 : _GEN_8224; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8226 = 10'h22b == _T_177[9:0] ? 4'h0 : _GEN_8225; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8227 = 10'h22c == _T_177[9:0] ? 4'h0 : _GEN_8226; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8228 = 10'h22d == _T_177[9:0] ? 4'h0 : _GEN_8227; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8229 = 10'h22e == _T_177[9:0] ? 4'h0 : _GEN_8228; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8230 = 10'h22f == _T_177[9:0] ? 4'h0 : _GEN_8229; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8231 = 10'h230 == _T_177[9:0] ? 4'h0 : _GEN_8230; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8232 = 10'h231 == _T_177[9:0] ? 4'h0 : _GEN_8231; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8233 = 10'h232 == _T_177[9:0] ? 4'h0 : _GEN_8232; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8234 = 10'h233 == _T_177[9:0] ? 4'h0 : _GEN_8233; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8235 = 10'h234 == _T_177[9:0] ? 4'h0 : _GEN_8234; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8236 = 10'h235 == _T_177[9:0] ? 4'h0 : _GEN_8235; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8237 = 10'h236 == _T_177[9:0] ? 4'h0 : _GEN_8236; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8238 = 10'h237 == _T_177[9:0] ? 4'h0 : _GEN_8237; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8239 = 10'h238 == _T_177[9:0] ? 4'h0 : _GEN_8238; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8240 = 10'h239 == _T_177[9:0] ? 4'h0 : _GEN_8239; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8241 = 10'h23a == _T_177[9:0] ? 4'h0 : _GEN_8240; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8242 = 10'h23b == _T_177[9:0] ? 4'h0 : _GEN_8241; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8243 = 10'h23c == _T_177[9:0] ? 4'h0 : _GEN_8242; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8244 = 10'h23d == _T_177[9:0] ? 4'h0 : _GEN_8243; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8245 = 10'h23e == _T_177[9:0] ? 4'h0 : _GEN_8244; // @[Filter.scala 191:102]
  wire [3:0] _GEN_8246 = 10'h23f == _T_177[9:0] ? 4'h0 : _GEN_8245; // @[Filter.scala 191:102]
  wire [6:0] _GEN_28324 = {{3'd0}, _GEN_8246}; // @[Filter.scala 191:102]
  wire [10:0] _T_184 = _GEN_28324 * 7'h46; // @[Filter.scala 191:102]
  wire [10:0] _GEN_28325 = {{2'd0}, _T_179}; // @[Filter.scala 191:69]
  wire [10:0] _T_186 = _GEN_28325 + _T_184; // @[Filter.scala 191:69]
  wire [3:0] _GEN_8278 = 10'h1f == _T_177[9:0] ? 4'h0 : 4'h3; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8279 = 10'h20 == _T_177[9:0] ? 4'h3 : _GEN_8278; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8280 = 10'h21 == _T_177[9:0] ? 4'h3 : _GEN_8279; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8281 = 10'h22 == _T_177[9:0] ? 4'h3 : _GEN_8280; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8282 = 10'h23 == _T_177[9:0] ? 4'h3 : _GEN_8281; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8283 = 10'h24 == _T_177[9:0] ? 4'h3 : _GEN_8282; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8284 = 10'h25 == _T_177[9:0] ? 4'h3 : _GEN_8283; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8285 = 10'h26 == _T_177[9:0] ? 4'h3 : _GEN_8284; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8286 = 10'h27 == _T_177[9:0] ? 4'h9 : _GEN_8285; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8287 = 10'h28 == _T_177[9:0] ? 4'h9 : _GEN_8286; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8288 = 10'h29 == _T_177[9:0] ? 4'h3 : _GEN_8287; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8289 = 10'h2a == _T_177[9:0] ? 4'h3 : _GEN_8288; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8290 = 10'h2b == _T_177[9:0] ? 4'h3 : _GEN_8289; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8291 = 10'h2c == _T_177[9:0] ? 4'h3 : _GEN_8290; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8292 = 10'h2d == _T_177[9:0] ? 4'h3 : _GEN_8291; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8293 = 10'h2e == _T_177[9:0] ? 4'h3 : _GEN_8292; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8294 = 10'h2f == _T_177[9:0] ? 4'h3 : _GEN_8293; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8295 = 10'h30 == _T_177[9:0] ? 4'h3 : _GEN_8294; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8296 = 10'h31 == _T_177[9:0] ? 4'h3 : _GEN_8295; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8297 = 10'h32 == _T_177[9:0] ? 4'h3 : _GEN_8296; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8298 = 10'h33 == _T_177[9:0] ? 4'h3 : _GEN_8297; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8299 = 10'h34 == _T_177[9:0] ? 4'h3 : _GEN_8298; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8300 = 10'h35 == _T_177[9:0] ? 4'h3 : _GEN_8299; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8301 = 10'h36 == _T_177[9:0] ? 4'h3 : _GEN_8300; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8302 = 10'h37 == _T_177[9:0] ? 4'h9 : _GEN_8301; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8303 = 10'h38 == _T_177[9:0] ? 4'h9 : _GEN_8302; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8304 = 10'h39 == _T_177[9:0] ? 4'h3 : _GEN_8303; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8305 = 10'h3a == _T_177[9:0] ? 4'h3 : _GEN_8304; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8306 = 10'h3b == _T_177[9:0] ? 4'h3 : _GEN_8305; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8307 = 10'h3c == _T_177[9:0] ? 4'h3 : _GEN_8306; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8308 = 10'h3d == _T_177[9:0] ? 4'h3 : _GEN_8307; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8309 = 10'h3e == _T_177[9:0] ? 4'h3 : _GEN_8308; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8310 = 10'h3f == _T_177[9:0] ? 4'h0 : _GEN_8309; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8311 = 10'h40 == _T_177[9:0] ? 4'h3 : _GEN_8310; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8312 = 10'h41 == _T_177[9:0] ? 4'h3 : _GEN_8311; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8313 = 10'h42 == _T_177[9:0] ? 4'h3 : _GEN_8312; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8314 = 10'h43 == _T_177[9:0] ? 4'h2 : _GEN_8313; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8315 = 10'h44 == _T_177[9:0] ? 4'h3 : _GEN_8314; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8316 = 10'h45 == _T_177[9:0] ? 4'hf : _GEN_8315; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8317 = 10'h46 == _T_177[9:0] ? 4'hf : _GEN_8316; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8318 = 10'h47 == _T_177[9:0] ? 4'hf : _GEN_8317; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8319 = 10'h48 == _T_177[9:0] ? 4'hf : _GEN_8318; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8320 = 10'h49 == _T_177[9:0] ? 4'h3 : _GEN_8319; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8321 = 10'h4a == _T_177[9:0] ? 4'h3 : _GEN_8320; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8322 = 10'h4b == _T_177[9:0] ? 4'h3 : _GEN_8321; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8323 = 10'h4c == _T_177[9:0] ? 4'h3 : _GEN_8322; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8324 = 10'h4d == _T_177[9:0] ? 4'h3 : _GEN_8323; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8325 = 10'h4e == _T_177[9:0] ? 4'h3 : _GEN_8324; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8326 = 10'h4f == _T_177[9:0] ? 4'h3 : _GEN_8325; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8327 = 10'h50 == _T_177[9:0] ? 4'h3 : _GEN_8326; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8328 = 10'h51 == _T_177[9:0] ? 4'h3 : _GEN_8327; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8329 = 10'h52 == _T_177[9:0] ? 4'h3 : _GEN_8328; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8330 = 10'h53 == _T_177[9:0] ? 4'h3 : _GEN_8329; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8331 = 10'h54 == _T_177[9:0] ? 4'h9 : _GEN_8330; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8332 = 10'h55 == _T_177[9:0] ? 4'h9 : _GEN_8331; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8333 = 10'h56 == _T_177[9:0] ? 4'h9 : _GEN_8332; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8334 = 10'h57 == _T_177[9:0] ? 4'hf : _GEN_8333; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8335 = 10'h58 == _T_177[9:0] ? 4'h3 : _GEN_8334; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8336 = 10'h59 == _T_177[9:0] ? 4'hf : _GEN_8335; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8337 = 10'h5a == _T_177[9:0] ? 4'h3 : _GEN_8336; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8338 = 10'h5b == _T_177[9:0] ? 4'h3 : _GEN_8337; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8339 = 10'h5c == _T_177[9:0] ? 4'h3 : _GEN_8338; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8340 = 10'h5d == _T_177[9:0] ? 4'h3 : _GEN_8339; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8341 = 10'h5e == _T_177[9:0] ? 4'h3 : _GEN_8340; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8342 = 10'h5f == _T_177[9:0] ? 4'h0 : _GEN_8341; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8343 = 10'h60 == _T_177[9:0] ? 4'h3 : _GEN_8342; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8344 = 10'h61 == _T_177[9:0] ? 4'h3 : _GEN_8343; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8345 = 10'h62 == _T_177[9:0] ? 4'h3 : _GEN_8344; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8346 = 10'h63 == _T_177[9:0] ? 4'h3 : _GEN_8345; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8347 = 10'h64 == _T_177[9:0] ? 4'h3 : _GEN_8346; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8348 = 10'h65 == _T_177[9:0] ? 4'hf : _GEN_8347; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8349 = 10'h66 == _T_177[9:0] ? 4'h3 : _GEN_8348; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8350 = 10'h67 == _T_177[9:0] ? 4'h3 : _GEN_8349; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8351 = 10'h68 == _T_177[9:0] ? 4'h3 : _GEN_8350; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8352 = 10'h69 == _T_177[9:0] ? 4'hf : _GEN_8351; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8353 = 10'h6a == _T_177[9:0] ? 4'h9 : _GEN_8352; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8354 = 10'h6b == _T_177[9:0] ? 4'h9 : _GEN_8353; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8355 = 10'h6c == _T_177[9:0] ? 4'h3 : _GEN_8354; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8356 = 10'h6d == _T_177[9:0] ? 4'h3 : _GEN_8355; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8357 = 10'h6e == _T_177[9:0] ? 4'h3 : _GEN_8356; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8358 = 10'h6f == _T_177[9:0] ? 4'h3 : _GEN_8357; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8359 = 10'h70 == _T_177[9:0] ? 4'h3 : _GEN_8358; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8360 = 10'h71 == _T_177[9:0] ? 4'h3 : _GEN_8359; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8361 = 10'h72 == _T_177[9:0] ? 4'h3 : _GEN_8360; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8362 = 10'h73 == _T_177[9:0] ? 4'h9 : _GEN_8361; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8363 = 10'h74 == _T_177[9:0] ? 4'hf : _GEN_8362; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8364 = 10'h75 == _T_177[9:0] ? 4'hf : _GEN_8363; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8365 = 10'h76 == _T_177[9:0] ? 4'hf : _GEN_8364; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8366 = 10'h77 == _T_177[9:0] ? 4'h3 : _GEN_8365; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8367 = 10'h78 == _T_177[9:0] ? 4'h3 : _GEN_8366; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8368 = 10'h79 == _T_177[9:0] ? 4'h3 : _GEN_8367; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8369 = 10'h7a == _T_177[9:0] ? 4'hf : _GEN_8368; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8370 = 10'h7b == _T_177[9:0] ? 4'h3 : _GEN_8369; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8371 = 10'h7c == _T_177[9:0] ? 4'h3 : _GEN_8370; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8372 = 10'h7d == _T_177[9:0] ? 4'h2 : _GEN_8371; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8373 = 10'h7e == _T_177[9:0] ? 4'h3 : _GEN_8372; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8374 = 10'h7f == _T_177[9:0] ? 4'h0 : _GEN_8373; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8375 = 10'h80 == _T_177[9:0] ? 4'h3 : _GEN_8374; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8376 = 10'h81 == _T_177[9:0] ? 4'h3 : _GEN_8375; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8377 = 10'h82 == _T_177[9:0] ? 4'h9 : _GEN_8376; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8378 = 10'h83 == _T_177[9:0] ? 4'hf : _GEN_8377; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8379 = 10'h84 == _T_177[9:0] ? 4'h2 : _GEN_8378; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8380 = 10'h85 == _T_177[9:0] ? 4'h9 : _GEN_8379; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8381 = 10'h86 == _T_177[9:0] ? 4'h9 : _GEN_8380; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8382 = 10'h87 == _T_177[9:0] ? 4'h3 : _GEN_8381; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8383 = 10'h88 == _T_177[9:0] ? 4'h3 : _GEN_8382; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8384 = 10'h89 == _T_177[9:0] ? 4'hf : _GEN_8383; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8385 = 10'h8a == _T_177[9:0] ? 4'hf : _GEN_8384; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8386 = 10'h8b == _T_177[9:0] ? 4'h9 : _GEN_8385; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8387 = 10'h8c == _T_177[9:0] ? 4'h9 : _GEN_8386; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8388 = 10'h8d == _T_177[9:0] ? 4'h9 : _GEN_8387; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8389 = 10'h8e == _T_177[9:0] ? 4'h9 : _GEN_8388; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8390 = 10'h8f == _T_177[9:0] ? 4'h9 : _GEN_8389; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8391 = 10'h90 == _T_177[9:0] ? 4'h9 : _GEN_8390; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8392 = 10'h91 == _T_177[9:0] ? 4'h9 : _GEN_8391; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8393 = 10'h92 == _T_177[9:0] ? 4'h9 : _GEN_8392; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8394 = 10'h93 == _T_177[9:0] ? 4'hf : _GEN_8393; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8395 = 10'h94 == _T_177[9:0] ? 4'hf : _GEN_8394; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8396 = 10'h95 == _T_177[9:0] ? 4'h3 : _GEN_8395; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8397 = 10'h96 == _T_177[9:0] ? 4'h3 : _GEN_8396; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8398 = 10'h97 == _T_177[9:0] ? 4'h3 : _GEN_8397; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8399 = 10'h98 == _T_177[9:0] ? 4'h9 : _GEN_8398; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8400 = 10'h99 == _T_177[9:0] ? 4'hf : _GEN_8399; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8401 = 10'h9a == _T_177[9:0] ? 4'h9 : _GEN_8400; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8402 = 10'h9b == _T_177[9:0] ? 4'h9 : _GEN_8401; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8403 = 10'h9c == _T_177[9:0] ? 4'h3 : _GEN_8402; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8404 = 10'h9d == _T_177[9:0] ? 4'h3 : _GEN_8403; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8405 = 10'h9e == _T_177[9:0] ? 4'h3 : _GEN_8404; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8406 = 10'h9f == _T_177[9:0] ? 4'h0 : _GEN_8405; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8407 = 10'ha0 == _T_177[9:0] ? 4'h3 : _GEN_8406; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8408 = 10'ha1 == _T_177[9:0] ? 4'h9 : _GEN_8407; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8409 = 10'ha2 == _T_177[9:0] ? 4'hf : _GEN_8408; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8410 = 10'ha3 == _T_177[9:0] ? 4'h3 : _GEN_8409; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8411 = 10'ha4 == _T_177[9:0] ? 4'h3 : _GEN_8410; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8412 = 10'ha5 == _T_177[9:0] ? 4'h3 : _GEN_8411; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8413 = 10'ha6 == _T_177[9:0] ? 4'h3 : _GEN_8412; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8414 = 10'ha7 == _T_177[9:0] ? 4'hf : _GEN_8413; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8415 = 10'ha8 == _T_177[9:0] ? 4'h3 : _GEN_8414; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8416 = 10'ha9 == _T_177[9:0] ? 4'h9 : _GEN_8415; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8417 = 10'haa == _T_177[9:0] ? 4'hf : _GEN_8416; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8418 = 10'hab == _T_177[9:0] ? 4'hf : _GEN_8417; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8419 = 10'hac == _T_177[9:0] ? 4'hf : _GEN_8418; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8420 = 10'had == _T_177[9:0] ? 4'hf : _GEN_8419; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8421 = 10'hae == _T_177[9:0] ? 4'hf : _GEN_8420; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8422 = 10'haf == _T_177[9:0] ? 4'hf : _GEN_8421; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8423 = 10'hb0 == _T_177[9:0] ? 4'hf : _GEN_8422; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8424 = 10'hb1 == _T_177[9:0] ? 4'hf : _GEN_8423; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8425 = 10'hb2 == _T_177[9:0] ? 4'hf : _GEN_8424; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8426 = 10'hb3 == _T_177[9:0] ? 4'hf : _GEN_8425; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8427 = 10'hb4 == _T_177[9:0] ? 4'h9 : _GEN_8426; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8428 = 10'hb5 == _T_177[9:0] ? 4'h9 : _GEN_8427; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8429 = 10'hb6 == _T_177[9:0] ? 4'h3 : _GEN_8428; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8430 = 10'hb7 == _T_177[9:0] ? 4'hf : _GEN_8429; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8431 = 10'hb8 == _T_177[9:0] ? 4'h3 : _GEN_8430; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8432 = 10'hb9 == _T_177[9:0] ? 4'h3 : _GEN_8431; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8433 = 10'hba == _T_177[9:0] ? 4'h3 : _GEN_8432; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8434 = 10'hbb == _T_177[9:0] ? 4'hf : _GEN_8433; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8435 = 10'hbc == _T_177[9:0] ? 4'h3 : _GEN_8434; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8436 = 10'hbd == _T_177[9:0] ? 4'h3 : _GEN_8435; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8437 = 10'hbe == _T_177[9:0] ? 4'h3 : _GEN_8436; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8438 = 10'hbf == _T_177[9:0] ? 4'h0 : _GEN_8437; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8439 = 10'hc0 == _T_177[9:0] ? 4'h3 : _GEN_8438; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8440 = 10'hc1 == _T_177[9:0] ? 4'h3 : _GEN_8439; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8441 = 10'hc2 == _T_177[9:0] ? 4'h3 : _GEN_8440; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8442 = 10'hc3 == _T_177[9:0] ? 4'h2 : _GEN_8441; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8443 = 10'hc4 == _T_177[9:0] ? 4'hf : _GEN_8442; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8444 = 10'hc5 == _T_177[9:0] ? 4'hf : _GEN_8443; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8445 = 10'hc6 == _T_177[9:0] ? 4'hf : _GEN_8444; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8446 = 10'hc7 == _T_177[9:0] ? 4'h3 : _GEN_8445; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8447 = 10'hc8 == _T_177[9:0] ? 4'h9 : _GEN_8446; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8448 = 10'hc9 == _T_177[9:0] ? 4'hf : _GEN_8447; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8449 = 10'hca == _T_177[9:0] ? 4'hf : _GEN_8448; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8450 = 10'hcb == _T_177[9:0] ? 4'hf : _GEN_8449; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8451 = 10'hcc == _T_177[9:0] ? 4'hf : _GEN_8450; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8452 = 10'hcd == _T_177[9:0] ? 4'hf : _GEN_8451; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8453 = 10'hce == _T_177[9:0] ? 4'hf : _GEN_8452; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8454 = 10'hcf == _T_177[9:0] ? 4'hf : _GEN_8453; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8455 = 10'hd0 == _T_177[9:0] ? 4'hf : _GEN_8454; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8456 = 10'hd1 == _T_177[9:0] ? 4'hf : _GEN_8455; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8457 = 10'hd2 == _T_177[9:0] ? 4'hf : _GEN_8456; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8458 = 10'hd3 == _T_177[9:0] ? 4'hf : _GEN_8457; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8459 = 10'hd4 == _T_177[9:0] ? 4'hf : _GEN_8458; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8460 = 10'hd5 == _T_177[9:0] ? 4'hf : _GEN_8459; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8461 = 10'hd6 == _T_177[9:0] ? 4'h9 : _GEN_8460; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8462 = 10'hd7 == _T_177[9:0] ? 4'h3 : _GEN_8461; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8463 = 10'hd8 == _T_177[9:0] ? 4'hf : _GEN_8462; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8464 = 10'hd9 == _T_177[9:0] ? 4'h3 : _GEN_8463; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8465 = 10'hda == _T_177[9:0] ? 4'h3 : _GEN_8464; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8466 = 10'hdb == _T_177[9:0] ? 4'h3 : _GEN_8465; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8467 = 10'hdc == _T_177[9:0] ? 4'h3 : _GEN_8466; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8468 = 10'hdd == _T_177[9:0] ? 4'h3 : _GEN_8467; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8469 = 10'hde == _T_177[9:0] ? 4'h2 : _GEN_8468; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8470 = 10'hdf == _T_177[9:0] ? 4'h0 : _GEN_8469; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8471 = 10'he0 == _T_177[9:0] ? 4'h3 : _GEN_8470; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8472 = 10'he1 == _T_177[9:0] ? 4'h3 : _GEN_8471; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8473 = 10'he2 == _T_177[9:0] ? 4'h3 : _GEN_8472; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8474 = 10'he3 == _T_177[9:0] ? 4'h3 : _GEN_8473; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8475 = 10'he4 == _T_177[9:0] ? 4'h3 : _GEN_8474; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8476 = 10'he5 == _T_177[9:0] ? 4'h3 : _GEN_8475; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8477 = 10'he6 == _T_177[9:0] ? 4'h3 : _GEN_8476; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8478 = 10'he7 == _T_177[9:0] ? 4'h9 : _GEN_8477; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8479 = 10'he8 == _T_177[9:0] ? 4'h9 : _GEN_8478; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8480 = 10'he9 == _T_177[9:0] ? 4'h9 : _GEN_8479; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8481 = 10'hea == _T_177[9:0] ? 4'hf : _GEN_8480; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8482 = 10'heb == _T_177[9:0] ? 4'hf : _GEN_8481; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8483 = 10'hec == _T_177[9:0] ? 4'hf : _GEN_8482; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8484 = 10'hed == _T_177[9:0] ? 4'hf : _GEN_8483; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8485 = 10'hee == _T_177[9:0] ? 4'hf : _GEN_8484; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8486 = 10'hef == _T_177[9:0] ? 4'hf : _GEN_8485; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8487 = 10'hf0 == _T_177[9:0] ? 4'hf : _GEN_8486; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8488 = 10'hf1 == _T_177[9:0] ? 4'hf : _GEN_8487; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8489 = 10'hf2 == _T_177[9:0] ? 4'hf : _GEN_8488; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8490 = 10'hf3 == _T_177[9:0] ? 4'hf : _GEN_8489; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8491 = 10'hf4 == _T_177[9:0] ? 4'hf : _GEN_8490; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8492 = 10'hf5 == _T_177[9:0] ? 4'h9 : _GEN_8491; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8493 = 10'hf6 == _T_177[9:0] ? 4'hf : _GEN_8492; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8494 = 10'hf7 == _T_177[9:0] ? 4'hf : _GEN_8493; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8495 = 10'hf8 == _T_177[9:0] ? 4'h9 : _GEN_8494; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8496 = 10'hf9 == _T_177[9:0] ? 4'hf : _GEN_8495; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8497 = 10'hfa == _T_177[9:0] ? 4'h3 : _GEN_8496; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8498 = 10'hfb == _T_177[9:0] ? 4'h3 : _GEN_8497; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8499 = 10'hfc == _T_177[9:0] ? 4'h3 : _GEN_8498; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8500 = 10'hfd == _T_177[9:0] ? 4'h3 : _GEN_8499; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8501 = 10'hfe == _T_177[9:0] ? 4'h3 : _GEN_8500; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8502 = 10'hff == _T_177[9:0] ? 4'h0 : _GEN_8501; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8503 = 10'h100 == _T_177[9:0] ? 4'h3 : _GEN_8502; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8504 = 10'h101 == _T_177[9:0] ? 4'hf : _GEN_8503; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8505 = 10'h102 == _T_177[9:0] ? 4'h3 : _GEN_8504; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8506 = 10'h103 == _T_177[9:0] ? 4'h3 : _GEN_8505; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8507 = 10'h104 == _T_177[9:0] ? 4'h3 : _GEN_8506; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8508 = 10'h105 == _T_177[9:0] ? 4'h3 : _GEN_8507; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8509 = 10'h106 == _T_177[9:0] ? 4'h3 : _GEN_8508; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8510 = 10'h107 == _T_177[9:0] ? 4'h3 : _GEN_8509; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8511 = 10'h108 == _T_177[9:0] ? 4'h9 : _GEN_8510; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8512 = 10'h109 == _T_177[9:0] ? 4'hf : _GEN_8511; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8513 = 10'h10a == _T_177[9:0] ? 4'hf : _GEN_8512; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8514 = 10'h10b == _T_177[9:0] ? 4'hf : _GEN_8513; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8515 = 10'h10c == _T_177[9:0] ? 4'hf : _GEN_8514; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8516 = 10'h10d == _T_177[9:0] ? 4'h0 : _GEN_8515; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8517 = 10'h10e == _T_177[9:0] ? 4'hf : _GEN_8516; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8518 = 10'h10f == _T_177[9:0] ? 4'hf : _GEN_8517; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8519 = 10'h110 == _T_177[9:0] ? 4'hf : _GEN_8518; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8520 = 10'h111 == _T_177[9:0] ? 4'h0 : _GEN_8519; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8521 = 10'h112 == _T_177[9:0] ? 4'hf : _GEN_8520; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8522 = 10'h113 == _T_177[9:0] ? 4'hf : _GEN_8521; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8523 = 10'h114 == _T_177[9:0] ? 4'hf : _GEN_8522; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8524 = 10'h115 == _T_177[9:0] ? 4'hf : _GEN_8523; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8525 = 10'h116 == _T_177[9:0] ? 4'h9 : _GEN_8524; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8526 = 10'h117 == _T_177[9:0] ? 4'h3 : _GEN_8525; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8527 = 10'h118 == _T_177[9:0] ? 4'h3 : _GEN_8526; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8528 = 10'h119 == _T_177[9:0] ? 4'h3 : _GEN_8527; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8529 = 10'h11a == _T_177[9:0] ? 4'hf : _GEN_8528; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8530 = 10'h11b == _T_177[9:0] ? 4'h3 : _GEN_8529; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8531 = 10'h11c == _T_177[9:0] ? 4'h3 : _GEN_8530; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8532 = 10'h11d == _T_177[9:0] ? 4'h2 : _GEN_8531; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8533 = 10'h11e == _T_177[9:0] ? 4'h3 : _GEN_8532; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8534 = 10'h11f == _T_177[9:0] ? 4'h0 : _GEN_8533; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8535 = 10'h120 == _T_177[9:0] ? 4'h3 : _GEN_8534; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8536 = 10'h121 == _T_177[9:0] ? 4'h3 : _GEN_8535; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8537 = 10'h122 == _T_177[9:0] ? 4'h3 : _GEN_8536; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8538 = 10'h123 == _T_177[9:0] ? 4'h3 : _GEN_8537; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8539 = 10'h124 == _T_177[9:0] ? 4'h3 : _GEN_8538; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8540 = 10'h125 == _T_177[9:0] ? 4'h3 : _GEN_8539; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8541 = 10'h126 == _T_177[9:0] ? 4'h3 : _GEN_8540; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8542 = 10'h127 == _T_177[9:0] ? 4'h9 : _GEN_8541; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8543 = 10'h128 == _T_177[9:0] ? 4'hf : _GEN_8542; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8544 = 10'h129 == _T_177[9:0] ? 4'h3 : _GEN_8543; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8545 = 10'h12a == _T_177[9:0] ? 4'h3 : _GEN_8544; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8546 = 10'h12b == _T_177[9:0] ? 4'hf : _GEN_8545; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8547 = 10'h12c == _T_177[9:0] ? 4'hf : _GEN_8546; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8548 = 10'h12d == _T_177[9:0] ? 4'hf : _GEN_8547; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8549 = 10'h12e == _T_177[9:0] ? 4'hf : _GEN_8548; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8550 = 10'h12f == _T_177[9:0] ? 4'hf : _GEN_8549; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8551 = 10'h130 == _T_177[9:0] ? 4'hf : _GEN_8550; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8552 = 10'h131 == _T_177[9:0] ? 4'hf : _GEN_8551; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8553 = 10'h132 == _T_177[9:0] ? 4'hf : _GEN_8552; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8554 = 10'h133 == _T_177[9:0] ? 4'hf : _GEN_8553; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8555 = 10'h134 == _T_177[9:0] ? 4'h3 : _GEN_8554; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8556 = 10'h135 == _T_177[9:0] ? 4'h3 : _GEN_8555; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8557 = 10'h136 == _T_177[9:0] ? 4'hf : _GEN_8556; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8558 = 10'h137 == _T_177[9:0] ? 4'h9 : _GEN_8557; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8559 = 10'h138 == _T_177[9:0] ? 4'h3 : _GEN_8558; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8560 = 10'h139 == _T_177[9:0] ? 4'h3 : _GEN_8559; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8561 = 10'h13a == _T_177[9:0] ? 4'h3 : _GEN_8560; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8562 = 10'h13b == _T_177[9:0] ? 4'h3 : _GEN_8561; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8563 = 10'h13c == _T_177[9:0] ? 4'h3 : _GEN_8562; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8564 = 10'h13d == _T_177[9:0] ? 4'h3 : _GEN_8563; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8565 = 10'h13e == _T_177[9:0] ? 4'h3 : _GEN_8564; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8566 = 10'h13f == _T_177[9:0] ? 4'h0 : _GEN_8565; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8567 = 10'h140 == _T_177[9:0] ? 4'h3 : _GEN_8566; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8568 = 10'h141 == _T_177[9:0] ? 4'h3 : _GEN_8567; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8569 = 10'h142 == _T_177[9:0] ? 4'h2 : _GEN_8568; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8570 = 10'h143 == _T_177[9:0] ? 4'h3 : _GEN_8569; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8571 = 10'h144 == _T_177[9:0] ? 4'h3 : _GEN_8570; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8572 = 10'h145 == _T_177[9:0] ? 4'h3 : _GEN_8571; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8573 = 10'h146 == _T_177[9:0] ? 4'h9 : _GEN_8572; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8574 = 10'h147 == _T_177[9:0] ? 4'hf : _GEN_8573; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8575 = 10'h148 == _T_177[9:0] ? 4'h3 : _GEN_8574; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8576 = 10'h149 == _T_177[9:0] ? 4'h3 : _GEN_8575; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8577 = 10'h14a == _T_177[9:0] ? 4'h3 : _GEN_8576; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8578 = 10'h14b == _T_177[9:0] ? 4'h3 : _GEN_8577; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8579 = 10'h14c == _T_177[9:0] ? 4'h3 : _GEN_8578; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8580 = 10'h14d == _T_177[9:0] ? 4'h3 : _GEN_8579; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8581 = 10'h14e == _T_177[9:0] ? 4'h3 : _GEN_8580; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8582 = 10'h14f == _T_177[9:0] ? 4'h3 : _GEN_8581; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8583 = 10'h150 == _T_177[9:0] ? 4'h3 : _GEN_8582; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8584 = 10'h151 == _T_177[9:0] ? 4'h3 : _GEN_8583; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8585 = 10'h152 == _T_177[9:0] ? 4'h3 : _GEN_8584; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8586 = 10'h153 == _T_177[9:0] ? 4'h3 : _GEN_8585; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8587 = 10'h154 == _T_177[9:0] ? 4'h3 : _GEN_8586; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8588 = 10'h155 == _T_177[9:0] ? 4'h3 : _GEN_8587; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8589 = 10'h156 == _T_177[9:0] ? 4'h3 : _GEN_8588; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8590 = 10'h157 == _T_177[9:0] ? 4'hf : _GEN_8589; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8591 = 10'h158 == _T_177[9:0] ? 4'h3 : _GEN_8590; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8592 = 10'h159 == _T_177[9:0] ? 4'h3 : _GEN_8591; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8593 = 10'h15a == _T_177[9:0] ? 4'h3 : _GEN_8592; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8594 = 10'h15b == _T_177[9:0] ? 4'h3 : _GEN_8593; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8595 = 10'h15c == _T_177[9:0] ? 4'h3 : _GEN_8594; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8596 = 10'h15d == _T_177[9:0] ? 4'h3 : _GEN_8595; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8597 = 10'h15e == _T_177[9:0] ? 4'h2 : _GEN_8596; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8598 = 10'h15f == _T_177[9:0] ? 4'h0 : _GEN_8597; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8599 = 10'h160 == _T_177[9:0] ? 4'h3 : _GEN_8598; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8600 = 10'h161 == _T_177[9:0] ? 4'h3 : _GEN_8599; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8601 = 10'h162 == _T_177[9:0] ? 4'h3 : _GEN_8600; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8602 = 10'h163 == _T_177[9:0] ? 4'h2 : _GEN_8601; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8603 = 10'h164 == _T_177[9:0] ? 4'h3 : _GEN_8602; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8604 = 10'h165 == _T_177[9:0] ? 4'h9 : _GEN_8603; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8605 = 10'h166 == _T_177[9:0] ? 4'hf : _GEN_8604; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8606 = 10'h167 == _T_177[9:0] ? 4'hf : _GEN_8605; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8607 = 10'h168 == _T_177[9:0] ? 4'hd : _GEN_8606; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8608 = 10'h169 == _T_177[9:0] ? 4'h9 : _GEN_8607; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8609 = 10'h16a == _T_177[9:0] ? 4'hd : _GEN_8608; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8610 = 10'h16b == _T_177[9:0] ? 4'hd : _GEN_8609; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8611 = 10'h16c == _T_177[9:0] ? 4'h3 : _GEN_8610; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8612 = 10'h16d == _T_177[9:0] ? 4'h3 : _GEN_8611; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8613 = 10'h16e == _T_177[9:0] ? 4'h3 : _GEN_8612; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8614 = 10'h16f == _T_177[9:0] ? 4'h3 : _GEN_8613; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8615 = 10'h170 == _T_177[9:0] ? 4'h3 : _GEN_8614; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8616 = 10'h171 == _T_177[9:0] ? 4'h3 : _GEN_8615; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8617 = 10'h172 == _T_177[9:0] ? 4'h3 : _GEN_8616; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8618 = 10'h173 == _T_177[9:0] ? 4'h3 : _GEN_8617; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8619 = 10'h174 == _T_177[9:0] ? 4'h3 : _GEN_8618; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8620 = 10'h175 == _T_177[9:0] ? 4'h3 : _GEN_8619; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8621 = 10'h176 == _T_177[9:0] ? 4'hf : _GEN_8620; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8622 = 10'h177 == _T_177[9:0] ? 4'hf : _GEN_8621; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8623 = 10'h178 == _T_177[9:0] ? 4'h9 : _GEN_8622; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8624 = 10'h179 == _T_177[9:0] ? 4'h3 : _GEN_8623; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8625 = 10'h17a == _T_177[9:0] ? 4'h3 : _GEN_8624; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8626 = 10'h17b == _T_177[9:0] ? 4'h3 : _GEN_8625; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8627 = 10'h17c == _T_177[9:0] ? 4'h3 : _GEN_8626; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8628 = 10'h17d == _T_177[9:0] ? 4'h2 : _GEN_8627; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8629 = 10'h17e == _T_177[9:0] ? 4'h3 : _GEN_8628; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8630 = 10'h17f == _T_177[9:0] ? 4'h0 : _GEN_8629; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8631 = 10'h180 == _T_177[9:0] ? 4'hd : _GEN_8630; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8632 = 10'h181 == _T_177[9:0] ? 4'hd : _GEN_8631; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8633 = 10'h182 == _T_177[9:0] ? 4'hd : _GEN_8632; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8634 = 10'h183 == _T_177[9:0] ? 4'hd : _GEN_8633; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8635 = 10'h184 == _T_177[9:0] ? 4'h3 : _GEN_8634; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8636 = 10'h185 == _T_177[9:0] ? 4'h9 : _GEN_8635; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8637 = 10'h186 == _T_177[9:0] ? 4'hb : _GEN_8636; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8638 = 10'h187 == _T_177[9:0] ? 4'hf : _GEN_8637; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8639 = 10'h188 == _T_177[9:0] ? 4'hd : _GEN_8638; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8640 = 10'h189 == _T_177[9:0] ? 4'hd : _GEN_8639; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8641 = 10'h18a == _T_177[9:0] ? 4'hd : _GEN_8640; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8642 = 10'h18b == _T_177[9:0] ? 4'hd : _GEN_8641; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8643 = 10'h18c == _T_177[9:0] ? 4'hd : _GEN_8642; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8644 = 10'h18d == _T_177[9:0] ? 4'hd : _GEN_8643; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8645 = 10'h18e == _T_177[9:0] ? 4'hd : _GEN_8644; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8646 = 10'h18f == _T_177[9:0] ? 4'hd : _GEN_8645; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8647 = 10'h190 == _T_177[9:0] ? 4'hd : _GEN_8646; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8648 = 10'h191 == _T_177[9:0] ? 4'hd : _GEN_8647; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8649 = 10'h192 == _T_177[9:0] ? 4'h9 : _GEN_8648; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8650 = 10'h193 == _T_177[9:0] ? 4'hd : _GEN_8649; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8651 = 10'h194 == _T_177[9:0] ? 4'hd : _GEN_8650; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8652 = 10'h195 == _T_177[9:0] ? 4'hd : _GEN_8651; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8653 = 10'h196 == _T_177[9:0] ? 4'hf : _GEN_8652; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8654 = 10'h197 == _T_177[9:0] ? 4'h3 : _GEN_8653; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8655 = 10'h198 == _T_177[9:0] ? 4'h9 : _GEN_8654; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8656 = 10'h199 == _T_177[9:0] ? 4'h3 : _GEN_8655; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8657 = 10'h19a == _T_177[9:0] ? 4'h3 : _GEN_8656; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8658 = 10'h19b == _T_177[9:0] ? 4'h3 : _GEN_8657; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8659 = 10'h19c == _T_177[9:0] ? 4'h3 : _GEN_8658; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8660 = 10'h19d == _T_177[9:0] ? 4'h3 : _GEN_8659; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8661 = 10'h19e == _T_177[9:0] ? 4'h3 : _GEN_8660; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8662 = 10'h19f == _T_177[9:0] ? 4'h0 : _GEN_8661; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8663 = 10'h1a0 == _T_177[9:0] ? 4'hd : _GEN_8662; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8664 = 10'h1a1 == _T_177[9:0] ? 4'hd : _GEN_8663; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8665 = 10'h1a2 == _T_177[9:0] ? 4'h9 : _GEN_8664; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8666 = 10'h1a3 == _T_177[9:0] ? 4'hd : _GEN_8665; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8667 = 10'h1a4 == _T_177[9:0] ? 4'h3 : _GEN_8666; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8668 = 10'h1a5 == _T_177[9:0] ? 4'hf : _GEN_8667; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8669 = 10'h1a6 == _T_177[9:0] ? 4'hd : _GEN_8668; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8670 = 10'h1a7 == _T_177[9:0] ? 4'hf : _GEN_8669; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8671 = 10'h1a8 == _T_177[9:0] ? 4'hb : _GEN_8670; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8672 = 10'h1a9 == _T_177[9:0] ? 4'hd : _GEN_8671; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8673 = 10'h1aa == _T_177[9:0] ? 4'hd : _GEN_8672; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8674 = 10'h1ab == _T_177[9:0] ? 4'h9 : _GEN_8673; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8675 = 10'h1ac == _T_177[9:0] ? 4'hd : _GEN_8674; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8676 = 10'h1ad == _T_177[9:0] ? 4'hd : _GEN_8675; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8677 = 10'h1ae == _T_177[9:0] ? 4'hd : _GEN_8676; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8678 = 10'h1af == _T_177[9:0] ? 4'hd : _GEN_8677; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8679 = 10'h1b0 == _T_177[9:0] ? 4'hd : _GEN_8678; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8680 = 10'h1b1 == _T_177[9:0] ? 4'hd : _GEN_8679; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8681 = 10'h1b2 == _T_177[9:0] ? 4'hd : _GEN_8680; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8682 = 10'h1b3 == _T_177[9:0] ? 4'hd : _GEN_8681; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8683 = 10'h1b4 == _T_177[9:0] ? 4'hd : _GEN_8682; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8684 = 10'h1b5 == _T_177[9:0] ? 4'hd : _GEN_8683; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8685 = 10'h1b6 == _T_177[9:0] ? 4'hf : _GEN_8684; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8686 = 10'h1b7 == _T_177[9:0] ? 4'hd : _GEN_8685; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8687 = 10'h1b8 == _T_177[9:0] ? 4'hf : _GEN_8686; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8688 = 10'h1b9 == _T_177[9:0] ? 4'hd : _GEN_8687; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8689 = 10'h1ba == _T_177[9:0] ? 4'hd : _GEN_8688; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8690 = 10'h1bb == _T_177[9:0] ? 4'hd : _GEN_8689; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8691 = 10'h1bc == _T_177[9:0] ? 4'h2 : _GEN_8690; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8692 = 10'h1bd == _T_177[9:0] ? 4'h3 : _GEN_8691; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8693 = 10'h1be == _T_177[9:0] ? 4'hd : _GEN_8692; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8694 = 10'h1bf == _T_177[9:0] ? 4'h0 : _GEN_8693; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8695 = 10'h1c0 == _T_177[9:0] ? 4'hd : _GEN_8694; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8696 = 10'h1c1 == _T_177[9:0] ? 4'hd : _GEN_8695; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8697 = 10'h1c2 == _T_177[9:0] ? 4'hd : _GEN_8696; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8698 = 10'h1c3 == _T_177[9:0] ? 4'h2 : _GEN_8697; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8699 = 10'h1c4 == _T_177[9:0] ? 4'h2 : _GEN_8698; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8700 = 10'h1c5 == _T_177[9:0] ? 4'hd : _GEN_8699; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8701 = 10'h1c6 == _T_177[9:0] ? 4'hd : _GEN_8700; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8702 = 10'h1c7 == _T_177[9:0] ? 4'hd : _GEN_8701; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8703 = 10'h1c8 == _T_177[9:0] ? 4'hd : _GEN_8702; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8704 = 10'h1c9 == _T_177[9:0] ? 4'hb : _GEN_8703; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8705 = 10'h1ca == _T_177[9:0] ? 4'hb : _GEN_8704; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8706 = 10'h1cb == _T_177[9:0] ? 4'hb : _GEN_8705; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8707 = 10'h1cc == _T_177[9:0] ? 4'hb : _GEN_8706; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8708 = 10'h1cd == _T_177[9:0] ? 4'hb : _GEN_8707; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8709 = 10'h1ce == _T_177[9:0] ? 4'hb : _GEN_8708; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8710 = 10'h1cf == _T_177[9:0] ? 4'hb : _GEN_8709; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8711 = 10'h1d0 == _T_177[9:0] ? 4'hb : _GEN_8710; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8712 = 10'h1d1 == _T_177[9:0] ? 4'hb : _GEN_8711; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8713 = 10'h1d2 == _T_177[9:0] ? 4'hb : _GEN_8712; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8714 = 10'h1d3 == _T_177[9:0] ? 4'hb : _GEN_8713; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8715 = 10'h1d4 == _T_177[9:0] ? 4'hb : _GEN_8714; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8716 = 10'h1d5 == _T_177[9:0] ? 4'hb : _GEN_8715; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8717 = 10'h1d6 == _T_177[9:0] ? 4'hd : _GEN_8716; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8718 = 10'h1d7 == _T_177[9:0] ? 4'hd : _GEN_8717; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8719 = 10'h1d8 == _T_177[9:0] ? 4'hd : _GEN_8718; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8720 = 10'h1d9 == _T_177[9:0] ? 4'hd : _GEN_8719; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8721 = 10'h1da == _T_177[9:0] ? 4'hd : _GEN_8720; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8722 = 10'h1db == _T_177[9:0] ? 4'hd : _GEN_8721; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8723 = 10'h1dc == _T_177[9:0] ? 4'hd : _GEN_8722; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8724 = 10'h1dd == _T_177[9:0] ? 4'h3 : _GEN_8723; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8725 = 10'h1de == _T_177[9:0] ? 4'hd : _GEN_8724; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8726 = 10'h1df == _T_177[9:0] ? 4'h0 : _GEN_8725; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8727 = 10'h1e0 == _T_177[9:0] ? 4'h9 : _GEN_8726; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8728 = 10'h1e1 == _T_177[9:0] ? 4'hd : _GEN_8727; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8729 = 10'h1e2 == _T_177[9:0] ? 4'h2 : _GEN_8728; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8730 = 10'h1e3 == _T_177[9:0] ? 4'h2 : _GEN_8729; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8731 = 10'h1e4 == _T_177[9:0] ? 4'hd : _GEN_8730; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8732 = 10'h1e5 == _T_177[9:0] ? 4'hd : _GEN_8731; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8733 = 10'h1e6 == _T_177[9:0] ? 4'hd : _GEN_8732; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8734 = 10'h1e7 == _T_177[9:0] ? 4'hd : _GEN_8733; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8735 = 10'h1e8 == _T_177[9:0] ? 4'hb : _GEN_8734; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8736 = 10'h1e9 == _T_177[9:0] ? 4'hd : _GEN_8735; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8737 = 10'h1ea == _T_177[9:0] ? 4'hd : _GEN_8736; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8738 = 10'h1eb == _T_177[9:0] ? 4'hb : _GEN_8737; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8739 = 10'h1ec == _T_177[9:0] ? 4'hd : _GEN_8738; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8740 = 10'h1ed == _T_177[9:0] ? 4'hb : _GEN_8739; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8741 = 10'h1ee == _T_177[9:0] ? 4'hd : _GEN_8740; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8742 = 10'h1ef == _T_177[9:0] ? 4'hb : _GEN_8741; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8743 = 10'h1f0 == _T_177[9:0] ? 4'hd : _GEN_8742; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8744 = 10'h1f1 == _T_177[9:0] ? 4'hb : _GEN_8743; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8745 = 10'h1f2 == _T_177[9:0] ? 4'hb : _GEN_8744; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8746 = 10'h1f3 == _T_177[9:0] ? 4'hd : _GEN_8745; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8747 = 10'h1f4 == _T_177[9:0] ? 4'hb : _GEN_8746; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8748 = 10'h1f5 == _T_177[9:0] ? 4'hb : _GEN_8747; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8749 = 10'h1f6 == _T_177[9:0] ? 4'hd : _GEN_8748; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8750 = 10'h1f7 == _T_177[9:0] ? 4'hd : _GEN_8749; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8751 = 10'h1f8 == _T_177[9:0] ? 4'hd : _GEN_8750; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8752 = 10'h1f9 == _T_177[9:0] ? 4'hd : _GEN_8751; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8753 = 10'h1fa == _T_177[9:0] ? 4'h9 : _GEN_8752; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8754 = 10'h1fb == _T_177[9:0] ? 4'hd : _GEN_8753; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8755 = 10'h1fc == _T_177[9:0] ? 4'hd : _GEN_8754; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8756 = 10'h1fd == _T_177[9:0] ? 4'h2 : _GEN_8755; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8757 = 10'h1fe == _T_177[9:0] ? 4'hd : _GEN_8756; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8758 = 10'h1ff == _T_177[9:0] ? 4'h0 : _GEN_8757; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8759 = 10'h200 == _T_177[9:0] ? 4'hd : _GEN_8758; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8760 = 10'h201 == _T_177[9:0] ? 4'hd : _GEN_8759; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8761 = 10'h202 == _T_177[9:0] ? 4'h3 : _GEN_8760; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8762 = 10'h203 == _T_177[9:0] ? 4'hd : _GEN_8761; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8763 = 10'h204 == _T_177[9:0] ? 4'hd : _GEN_8762; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8764 = 10'h205 == _T_177[9:0] ? 4'hd : _GEN_8763; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8765 = 10'h206 == _T_177[9:0] ? 4'hb : _GEN_8764; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8766 = 10'h207 == _T_177[9:0] ? 4'hb : _GEN_8765; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8767 = 10'h208 == _T_177[9:0] ? 4'hd : _GEN_8766; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8768 = 10'h209 == _T_177[9:0] ? 4'hd : _GEN_8767; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8769 = 10'h20a == _T_177[9:0] ? 4'hd : _GEN_8768; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8770 = 10'h20b == _T_177[9:0] ? 4'hb : _GEN_8769; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8771 = 10'h20c == _T_177[9:0] ? 4'hd : _GEN_8770; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8772 = 10'h20d == _T_177[9:0] ? 4'hb : _GEN_8771; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8773 = 10'h20e == _T_177[9:0] ? 4'hd : _GEN_8772; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8774 = 10'h20f == _T_177[9:0] ? 4'hb : _GEN_8773; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8775 = 10'h210 == _T_177[9:0] ? 4'hd : _GEN_8774; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8776 = 10'h211 == _T_177[9:0] ? 4'hd : _GEN_8775; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8777 = 10'h212 == _T_177[9:0] ? 4'hb : _GEN_8776; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8778 = 10'h213 == _T_177[9:0] ? 4'hb : _GEN_8777; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8779 = 10'h214 == _T_177[9:0] ? 4'hb : _GEN_8778; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8780 = 10'h215 == _T_177[9:0] ? 4'hd : _GEN_8779; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8781 = 10'h216 == _T_177[9:0] ? 4'hd : _GEN_8780; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8782 = 10'h217 == _T_177[9:0] ? 4'hd : _GEN_8781; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8783 = 10'h218 == _T_177[9:0] ? 4'hd : _GEN_8782; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8784 = 10'h219 == _T_177[9:0] ? 4'hd : _GEN_8783; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8785 = 10'h21a == _T_177[9:0] ? 4'hd : _GEN_8784; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8786 = 10'h21b == _T_177[9:0] ? 4'hd : _GEN_8785; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8787 = 10'h21c == _T_177[9:0] ? 4'h3 : _GEN_8786; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8788 = 10'h21d == _T_177[9:0] ? 4'h2 : _GEN_8787; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8789 = 10'h21e == _T_177[9:0] ? 4'hd : _GEN_8788; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8790 = 10'h21f == _T_177[9:0] ? 4'h0 : _GEN_8789; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8791 = 10'h220 == _T_177[9:0] ? 4'h0 : _GEN_8790; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8792 = 10'h221 == _T_177[9:0] ? 4'h0 : _GEN_8791; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8793 = 10'h222 == _T_177[9:0] ? 4'h0 : _GEN_8792; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8794 = 10'h223 == _T_177[9:0] ? 4'h0 : _GEN_8793; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8795 = 10'h224 == _T_177[9:0] ? 4'h0 : _GEN_8794; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8796 = 10'h225 == _T_177[9:0] ? 4'h0 : _GEN_8795; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8797 = 10'h226 == _T_177[9:0] ? 4'h0 : _GEN_8796; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8798 = 10'h227 == _T_177[9:0] ? 4'h0 : _GEN_8797; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8799 = 10'h228 == _T_177[9:0] ? 4'h0 : _GEN_8798; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8800 = 10'h229 == _T_177[9:0] ? 4'h0 : _GEN_8799; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8801 = 10'h22a == _T_177[9:0] ? 4'h0 : _GEN_8800; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8802 = 10'h22b == _T_177[9:0] ? 4'h0 : _GEN_8801; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8803 = 10'h22c == _T_177[9:0] ? 4'h0 : _GEN_8802; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8804 = 10'h22d == _T_177[9:0] ? 4'h0 : _GEN_8803; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8805 = 10'h22e == _T_177[9:0] ? 4'h0 : _GEN_8804; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8806 = 10'h22f == _T_177[9:0] ? 4'h0 : _GEN_8805; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8807 = 10'h230 == _T_177[9:0] ? 4'h0 : _GEN_8806; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8808 = 10'h231 == _T_177[9:0] ? 4'h0 : _GEN_8807; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8809 = 10'h232 == _T_177[9:0] ? 4'h0 : _GEN_8808; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8810 = 10'h233 == _T_177[9:0] ? 4'h0 : _GEN_8809; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8811 = 10'h234 == _T_177[9:0] ? 4'h0 : _GEN_8810; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8812 = 10'h235 == _T_177[9:0] ? 4'h0 : _GEN_8811; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8813 = 10'h236 == _T_177[9:0] ? 4'h0 : _GEN_8812; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8814 = 10'h237 == _T_177[9:0] ? 4'h0 : _GEN_8813; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8815 = 10'h238 == _T_177[9:0] ? 4'h0 : _GEN_8814; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8816 = 10'h239 == _T_177[9:0] ? 4'h0 : _GEN_8815; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8817 = 10'h23a == _T_177[9:0] ? 4'h0 : _GEN_8816; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8818 = 10'h23b == _T_177[9:0] ? 4'h0 : _GEN_8817; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8819 = 10'h23c == _T_177[9:0] ? 4'h0 : _GEN_8818; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8820 = 10'h23d == _T_177[9:0] ? 4'h0 : _GEN_8819; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8821 = 10'h23e == _T_177[9:0] ? 4'h0 : _GEN_8820; // @[Filter.scala 191:142]
  wire [3:0] _GEN_8822 = 10'h23f == _T_177[9:0] ? 4'h0 : _GEN_8821; // @[Filter.scala 191:142]
  wire [7:0] _T_191 = _GEN_8822 * 4'ha; // @[Filter.scala 191:142]
  wire [10:0] _GEN_28327 = {{3'd0}, _T_191}; // @[Filter.scala 191:109]
  wire [10:0] _T_193 = _T_186 + _GEN_28327; // @[Filter.scala 191:109]
  wire [10:0] _T_194 = _T_193 / 11'h64; // @[Filter.scala 191:150]
  wire  _T_196 = _T_167 >= 6'h20; // @[Filter.scala 194:31]
  wire  _T_200 = _T_174 >= 32'h12; // @[Filter.scala 194:63]
  wire  _T_201 = _T_196 | _T_200; // @[Filter.scala 194:58]
  wire [10:0] _GEN_9399 = io_SPI_distort ? _T_194 : {{7'd0}, _GEN_7670}; // @[Filter.scala 196:35]
  wire [10:0] _GEN_9400 = _T_201 ? 11'h0 : _GEN_9399; // @[Filter.scala 194:80]
  wire [10:0] _GEN_9977 = io_SPI_distort ? _T_194 : {{7'd0}, _GEN_8246}; // @[Filter.scala 196:35]
  wire [10:0] _GEN_9978 = _T_201 ? 11'h0 : _GEN_9977; // @[Filter.scala 194:80]
  wire [10:0] _GEN_10555 = io_SPI_distort ? _T_194 : {{7'd0}, _GEN_8822}; // @[Filter.scala 196:35]
  wire [10:0] _GEN_10556 = _T_201 ? 11'h0 : _GEN_10555; // @[Filter.scala 194:80]
  wire [31:0] _T_229 = pixelIndex + 32'h3; // @[Filter.scala 189:31]
  wire [31:0] _GEN_3 = _T_229 % 32'h20; // @[Filter.scala 189:38]
  wire [5:0] _T_230 = _GEN_3[5:0]; // @[Filter.scala 189:38]
  wire [5:0] _T_232 = _T_230 + _GEN_28295; // @[Filter.scala 189:53]
  wire [5:0] _T_234 = _T_232 - 6'h1; // @[Filter.scala 189:69]
  wire [31:0] _T_237 = _T_229 / 32'h20; // @[Filter.scala 190:38]
  wire [31:0] _T_239 = _T_237 + _GEN_28296; // @[Filter.scala 190:53]
  wire [31:0] _T_241 = _T_239 - 32'h1; // @[Filter.scala 190:69]
  wire [37:0] _T_242 = _T_241 * 32'h20; // @[Filter.scala 191:42]
  wire [37:0] _GEN_28333 = {{32'd0}, _T_234}; // @[Filter.scala 191:57]
  wire [37:0] _T_244 = _T_242 + _GEN_28333; // @[Filter.scala 191:57]
  wire [3:0] _GEN_10560 = 10'h3 == _T_244[9:0] ? 4'h3 : 4'ha; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10561 = 10'h4 == _T_244[9:0] ? 4'ha : _GEN_10560; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10562 = 10'h5 == _T_244[9:0] ? 4'ha : _GEN_10561; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10563 = 10'h6 == _T_244[9:0] ? 4'ha : _GEN_10562; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10564 = 10'h7 == _T_244[9:0] ? 4'ha : _GEN_10563; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10565 = 10'h8 == _T_244[9:0] ? 4'ha : _GEN_10564; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10566 = 10'h9 == _T_244[9:0] ? 4'ha : _GEN_10565; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10567 = 10'ha == _T_244[9:0] ? 4'ha : _GEN_10566; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10568 = 10'hb == _T_244[9:0] ? 4'ha : _GEN_10567; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10569 = 10'hc == _T_244[9:0] ? 4'ha : _GEN_10568; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10570 = 10'hd == _T_244[9:0] ? 4'ha : _GEN_10569; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10571 = 10'he == _T_244[9:0] ? 4'ha : _GEN_10570; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10572 = 10'hf == _T_244[9:0] ? 4'ha : _GEN_10571; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10573 = 10'h10 == _T_244[9:0] ? 4'ha : _GEN_10572; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10574 = 10'h11 == _T_244[9:0] ? 4'ha : _GEN_10573; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10575 = 10'h12 == _T_244[9:0] ? 4'ha : _GEN_10574; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10576 = 10'h13 == _T_244[9:0] ? 4'ha : _GEN_10575; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10577 = 10'h14 == _T_244[9:0] ? 4'ha : _GEN_10576; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10578 = 10'h15 == _T_244[9:0] ? 4'ha : _GEN_10577; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10579 = 10'h16 == _T_244[9:0] ? 4'ha : _GEN_10578; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10580 = 10'h17 == _T_244[9:0] ? 4'ha : _GEN_10579; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10581 = 10'h18 == _T_244[9:0] ? 4'ha : _GEN_10580; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10582 = 10'h19 == _T_244[9:0] ? 4'ha : _GEN_10581; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10583 = 10'h1a == _T_244[9:0] ? 4'ha : _GEN_10582; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10584 = 10'h1b == _T_244[9:0] ? 4'ha : _GEN_10583; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10585 = 10'h1c == _T_244[9:0] ? 4'ha : _GEN_10584; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10586 = 10'h1d == _T_244[9:0] ? 4'ha : _GEN_10585; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10587 = 10'h1e == _T_244[9:0] ? 4'ha : _GEN_10586; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10588 = 10'h1f == _T_244[9:0] ? 4'h0 : _GEN_10587; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10589 = 10'h20 == _T_244[9:0] ? 4'ha : _GEN_10588; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10590 = 10'h21 == _T_244[9:0] ? 4'ha : _GEN_10589; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10591 = 10'h22 == _T_244[9:0] ? 4'ha : _GEN_10590; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10592 = 10'h23 == _T_244[9:0] ? 4'h3 : _GEN_10591; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10593 = 10'h24 == _T_244[9:0] ? 4'ha : _GEN_10592; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10594 = 10'h25 == _T_244[9:0] ? 4'ha : _GEN_10593; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10595 = 10'h26 == _T_244[9:0] ? 4'ha : _GEN_10594; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10596 = 10'h27 == _T_244[9:0] ? 4'h1 : _GEN_10595; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10597 = 10'h28 == _T_244[9:0] ? 4'h1 : _GEN_10596; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10598 = 10'h29 == _T_244[9:0] ? 4'ha : _GEN_10597; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10599 = 10'h2a == _T_244[9:0] ? 4'ha : _GEN_10598; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10600 = 10'h2b == _T_244[9:0] ? 4'ha : _GEN_10599; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10601 = 10'h2c == _T_244[9:0] ? 4'ha : _GEN_10600; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10602 = 10'h2d == _T_244[9:0] ? 4'ha : _GEN_10601; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10603 = 10'h2e == _T_244[9:0] ? 4'ha : _GEN_10602; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10604 = 10'h2f == _T_244[9:0] ? 4'ha : _GEN_10603; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10605 = 10'h30 == _T_244[9:0] ? 4'ha : _GEN_10604; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10606 = 10'h31 == _T_244[9:0] ? 4'ha : _GEN_10605; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10607 = 10'h32 == _T_244[9:0] ? 4'ha : _GEN_10606; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10608 = 10'h33 == _T_244[9:0] ? 4'ha : _GEN_10607; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10609 = 10'h34 == _T_244[9:0] ? 4'ha : _GEN_10608; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10610 = 10'h35 == _T_244[9:0] ? 4'ha : _GEN_10609; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10611 = 10'h36 == _T_244[9:0] ? 4'ha : _GEN_10610; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10612 = 10'h37 == _T_244[9:0] ? 4'h1 : _GEN_10611; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10613 = 10'h38 == _T_244[9:0] ? 4'h1 : _GEN_10612; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10614 = 10'h39 == _T_244[9:0] ? 4'ha : _GEN_10613; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10615 = 10'h3a == _T_244[9:0] ? 4'ha : _GEN_10614; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10616 = 10'h3b == _T_244[9:0] ? 4'ha : _GEN_10615; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10617 = 10'h3c == _T_244[9:0] ? 4'ha : _GEN_10616; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10618 = 10'h3d == _T_244[9:0] ? 4'h3 : _GEN_10617; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10619 = 10'h3e == _T_244[9:0] ? 4'ha : _GEN_10618; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10620 = 10'h3f == _T_244[9:0] ? 4'h0 : _GEN_10619; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10621 = 10'h40 == _T_244[9:0] ? 4'ha : _GEN_10620; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10622 = 10'h41 == _T_244[9:0] ? 4'ha : _GEN_10621; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10623 = 10'h42 == _T_244[9:0] ? 4'ha : _GEN_10622; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10624 = 10'h43 == _T_244[9:0] ? 4'h2 : _GEN_10623; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10625 = 10'h44 == _T_244[9:0] ? 4'h3 : _GEN_10624; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10626 = 10'h45 == _T_244[9:0] ? 4'h0 : _GEN_10625; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10627 = 10'h46 == _T_244[9:0] ? 4'h0 : _GEN_10626; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10628 = 10'h47 == _T_244[9:0] ? 4'h0 : _GEN_10627; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10629 = 10'h48 == _T_244[9:0] ? 4'h0 : _GEN_10628; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10630 = 10'h49 == _T_244[9:0] ? 4'ha : _GEN_10629; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10631 = 10'h4a == _T_244[9:0] ? 4'ha : _GEN_10630; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10632 = 10'h4b == _T_244[9:0] ? 4'ha : _GEN_10631; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10633 = 10'h4c == _T_244[9:0] ? 4'ha : _GEN_10632; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10634 = 10'h4d == _T_244[9:0] ? 4'ha : _GEN_10633; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10635 = 10'h4e == _T_244[9:0] ? 4'ha : _GEN_10634; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10636 = 10'h4f == _T_244[9:0] ? 4'ha : _GEN_10635; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10637 = 10'h50 == _T_244[9:0] ? 4'ha : _GEN_10636; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10638 = 10'h51 == _T_244[9:0] ? 4'ha : _GEN_10637; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10639 = 10'h52 == _T_244[9:0] ? 4'ha : _GEN_10638; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10640 = 10'h53 == _T_244[9:0] ? 4'ha : _GEN_10639; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10641 = 10'h54 == _T_244[9:0] ? 4'h1 : _GEN_10640; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10642 = 10'h55 == _T_244[9:0] ? 4'h1 : _GEN_10641; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10643 = 10'h56 == _T_244[9:0] ? 4'h1 : _GEN_10642; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10644 = 10'h57 == _T_244[9:0] ? 4'h0 : _GEN_10643; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10645 = 10'h58 == _T_244[9:0] ? 4'ha : _GEN_10644; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10646 = 10'h59 == _T_244[9:0] ? 4'h0 : _GEN_10645; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10647 = 10'h5a == _T_244[9:0] ? 4'ha : _GEN_10646; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10648 = 10'h5b == _T_244[9:0] ? 4'ha : _GEN_10647; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10649 = 10'h5c == _T_244[9:0] ? 4'ha : _GEN_10648; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10650 = 10'h5d == _T_244[9:0] ? 4'h3 : _GEN_10649; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10651 = 10'h5e == _T_244[9:0] ? 4'ha : _GEN_10650; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10652 = 10'h5f == _T_244[9:0] ? 4'h0 : _GEN_10651; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10653 = 10'h60 == _T_244[9:0] ? 4'ha : _GEN_10652; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10654 = 10'h61 == _T_244[9:0] ? 4'ha : _GEN_10653; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10655 = 10'h62 == _T_244[9:0] ? 4'ha : _GEN_10654; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10656 = 10'h63 == _T_244[9:0] ? 4'ha : _GEN_10655; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10657 = 10'h64 == _T_244[9:0] ? 4'h3 : _GEN_10656; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10658 = 10'h65 == _T_244[9:0] ? 4'h0 : _GEN_10657; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10659 = 10'h66 == _T_244[9:0] ? 4'ha : _GEN_10658; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10660 = 10'h67 == _T_244[9:0] ? 4'ha : _GEN_10659; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10661 = 10'h68 == _T_244[9:0] ? 4'ha : _GEN_10660; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10662 = 10'h69 == _T_244[9:0] ? 4'h0 : _GEN_10661; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10663 = 10'h6a == _T_244[9:0] ? 4'h1 : _GEN_10662; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10664 = 10'h6b == _T_244[9:0] ? 4'h1 : _GEN_10663; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10665 = 10'h6c == _T_244[9:0] ? 4'ha : _GEN_10664; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10666 = 10'h6d == _T_244[9:0] ? 4'ha : _GEN_10665; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10667 = 10'h6e == _T_244[9:0] ? 4'ha : _GEN_10666; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10668 = 10'h6f == _T_244[9:0] ? 4'ha : _GEN_10667; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10669 = 10'h70 == _T_244[9:0] ? 4'ha : _GEN_10668; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10670 = 10'h71 == _T_244[9:0] ? 4'ha : _GEN_10669; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10671 = 10'h72 == _T_244[9:0] ? 4'ha : _GEN_10670; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10672 = 10'h73 == _T_244[9:0] ? 4'h1 : _GEN_10671; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10673 = 10'h74 == _T_244[9:0] ? 4'h0 : _GEN_10672; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10674 = 10'h75 == _T_244[9:0] ? 4'h0 : _GEN_10673; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10675 = 10'h76 == _T_244[9:0] ? 4'h0 : _GEN_10674; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10676 = 10'h77 == _T_244[9:0] ? 4'ha : _GEN_10675; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10677 = 10'h78 == _T_244[9:0] ? 4'ha : _GEN_10676; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10678 = 10'h79 == _T_244[9:0] ? 4'ha : _GEN_10677; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10679 = 10'h7a == _T_244[9:0] ? 4'h0 : _GEN_10678; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10680 = 10'h7b == _T_244[9:0] ? 4'ha : _GEN_10679; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10681 = 10'h7c == _T_244[9:0] ? 4'ha : _GEN_10680; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10682 = 10'h7d == _T_244[9:0] ? 4'h2 : _GEN_10681; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10683 = 10'h7e == _T_244[9:0] ? 4'h3 : _GEN_10682; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10684 = 10'h7f == _T_244[9:0] ? 4'h0 : _GEN_10683; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10685 = 10'h80 == _T_244[9:0] ? 4'ha : _GEN_10684; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10686 = 10'h81 == _T_244[9:0] ? 4'ha : _GEN_10685; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10687 = 10'h82 == _T_244[9:0] ? 4'h1 : _GEN_10686; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10688 = 10'h83 == _T_244[9:0] ? 4'h0 : _GEN_10687; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10689 = 10'h84 == _T_244[9:0] ? 4'h2 : _GEN_10688; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10690 = 10'h85 == _T_244[9:0] ? 4'h1 : _GEN_10689; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10691 = 10'h86 == _T_244[9:0] ? 4'h1 : _GEN_10690; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10692 = 10'h87 == _T_244[9:0] ? 4'ha : _GEN_10691; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10693 = 10'h88 == _T_244[9:0] ? 4'ha : _GEN_10692; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10694 = 10'h89 == _T_244[9:0] ? 4'h0 : _GEN_10693; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10695 = 10'h8a == _T_244[9:0] ? 4'h0 : _GEN_10694; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10696 = 10'h8b == _T_244[9:0] ? 4'h1 : _GEN_10695; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10697 = 10'h8c == _T_244[9:0] ? 4'h1 : _GEN_10696; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10698 = 10'h8d == _T_244[9:0] ? 4'h1 : _GEN_10697; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10699 = 10'h8e == _T_244[9:0] ? 4'h1 : _GEN_10698; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10700 = 10'h8f == _T_244[9:0] ? 4'h1 : _GEN_10699; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10701 = 10'h90 == _T_244[9:0] ? 4'h1 : _GEN_10700; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10702 = 10'h91 == _T_244[9:0] ? 4'h1 : _GEN_10701; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10703 = 10'h92 == _T_244[9:0] ? 4'h1 : _GEN_10702; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10704 = 10'h93 == _T_244[9:0] ? 4'h0 : _GEN_10703; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10705 = 10'h94 == _T_244[9:0] ? 4'h0 : _GEN_10704; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10706 = 10'h95 == _T_244[9:0] ? 4'ha : _GEN_10705; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10707 = 10'h96 == _T_244[9:0] ? 4'ha : _GEN_10706; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10708 = 10'h97 == _T_244[9:0] ? 4'ha : _GEN_10707; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10709 = 10'h98 == _T_244[9:0] ? 4'h1 : _GEN_10708; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10710 = 10'h99 == _T_244[9:0] ? 4'h0 : _GEN_10709; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10711 = 10'h9a == _T_244[9:0] ? 4'h1 : _GEN_10710; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10712 = 10'h9b == _T_244[9:0] ? 4'h1 : _GEN_10711; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10713 = 10'h9c == _T_244[9:0] ? 4'ha : _GEN_10712; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10714 = 10'h9d == _T_244[9:0] ? 4'ha : _GEN_10713; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10715 = 10'h9e == _T_244[9:0] ? 4'h3 : _GEN_10714; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10716 = 10'h9f == _T_244[9:0] ? 4'h0 : _GEN_10715; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10717 = 10'ha0 == _T_244[9:0] ? 4'ha : _GEN_10716; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10718 = 10'ha1 == _T_244[9:0] ? 4'h1 : _GEN_10717; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10719 = 10'ha2 == _T_244[9:0] ? 4'h0 : _GEN_10718; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10720 = 10'ha3 == _T_244[9:0] ? 4'h3 : _GEN_10719; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10721 = 10'ha4 == _T_244[9:0] ? 4'ha : _GEN_10720; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10722 = 10'ha5 == _T_244[9:0] ? 4'ha : _GEN_10721; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10723 = 10'ha6 == _T_244[9:0] ? 4'ha : _GEN_10722; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10724 = 10'ha7 == _T_244[9:0] ? 4'h0 : _GEN_10723; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10725 = 10'ha8 == _T_244[9:0] ? 4'ha : _GEN_10724; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10726 = 10'ha9 == _T_244[9:0] ? 4'h1 : _GEN_10725; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10727 = 10'haa == _T_244[9:0] ? 4'h0 : _GEN_10726; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10728 = 10'hab == _T_244[9:0] ? 4'h0 : _GEN_10727; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10729 = 10'hac == _T_244[9:0] ? 4'h0 : _GEN_10728; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10730 = 10'had == _T_244[9:0] ? 4'h0 : _GEN_10729; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10731 = 10'hae == _T_244[9:0] ? 4'h0 : _GEN_10730; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10732 = 10'haf == _T_244[9:0] ? 4'h0 : _GEN_10731; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10733 = 10'hb0 == _T_244[9:0] ? 4'h0 : _GEN_10732; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10734 = 10'hb1 == _T_244[9:0] ? 4'h0 : _GEN_10733; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10735 = 10'hb2 == _T_244[9:0] ? 4'h0 : _GEN_10734; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10736 = 10'hb3 == _T_244[9:0] ? 4'h0 : _GEN_10735; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10737 = 10'hb4 == _T_244[9:0] ? 4'h1 : _GEN_10736; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10738 = 10'hb5 == _T_244[9:0] ? 4'h1 : _GEN_10737; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10739 = 10'hb6 == _T_244[9:0] ? 4'ha : _GEN_10738; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10740 = 10'hb7 == _T_244[9:0] ? 4'h0 : _GEN_10739; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10741 = 10'hb8 == _T_244[9:0] ? 4'ha : _GEN_10740; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10742 = 10'hb9 == _T_244[9:0] ? 4'ha : _GEN_10741; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10743 = 10'hba == _T_244[9:0] ? 4'ha : _GEN_10742; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10744 = 10'hbb == _T_244[9:0] ? 4'h0 : _GEN_10743; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10745 = 10'hbc == _T_244[9:0] ? 4'ha : _GEN_10744; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10746 = 10'hbd == _T_244[9:0] ? 4'ha : _GEN_10745; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10747 = 10'hbe == _T_244[9:0] ? 4'h3 : _GEN_10746; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10748 = 10'hbf == _T_244[9:0] ? 4'h0 : _GEN_10747; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10749 = 10'hc0 == _T_244[9:0] ? 4'ha : _GEN_10748; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10750 = 10'hc1 == _T_244[9:0] ? 4'ha : _GEN_10749; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10751 = 10'hc2 == _T_244[9:0] ? 4'h3 : _GEN_10750; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10752 = 10'hc3 == _T_244[9:0] ? 4'h2 : _GEN_10751; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10753 = 10'hc4 == _T_244[9:0] ? 4'h0 : _GEN_10752; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10754 = 10'hc5 == _T_244[9:0] ? 4'h0 : _GEN_10753; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10755 = 10'hc6 == _T_244[9:0] ? 4'h0 : _GEN_10754; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10756 = 10'hc7 == _T_244[9:0] ? 4'ha : _GEN_10755; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10757 = 10'hc8 == _T_244[9:0] ? 4'h1 : _GEN_10756; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10758 = 10'hc9 == _T_244[9:0] ? 4'h0 : _GEN_10757; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10759 = 10'hca == _T_244[9:0] ? 4'h0 : _GEN_10758; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10760 = 10'hcb == _T_244[9:0] ? 4'h0 : _GEN_10759; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10761 = 10'hcc == _T_244[9:0] ? 4'h0 : _GEN_10760; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10762 = 10'hcd == _T_244[9:0] ? 4'h0 : _GEN_10761; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10763 = 10'hce == _T_244[9:0] ? 4'h0 : _GEN_10762; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10764 = 10'hcf == _T_244[9:0] ? 4'h0 : _GEN_10763; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10765 = 10'hd0 == _T_244[9:0] ? 4'h0 : _GEN_10764; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10766 = 10'hd1 == _T_244[9:0] ? 4'h0 : _GEN_10765; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10767 = 10'hd2 == _T_244[9:0] ? 4'h0 : _GEN_10766; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10768 = 10'hd3 == _T_244[9:0] ? 4'h0 : _GEN_10767; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10769 = 10'hd4 == _T_244[9:0] ? 4'h0 : _GEN_10768; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10770 = 10'hd5 == _T_244[9:0] ? 4'h0 : _GEN_10769; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10771 = 10'hd6 == _T_244[9:0] ? 4'h1 : _GEN_10770; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10772 = 10'hd7 == _T_244[9:0] ? 4'ha : _GEN_10771; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10773 = 10'hd8 == _T_244[9:0] ? 4'h0 : _GEN_10772; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10774 = 10'hd9 == _T_244[9:0] ? 4'ha : _GEN_10773; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10775 = 10'hda == _T_244[9:0] ? 4'ha : _GEN_10774; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10776 = 10'hdb == _T_244[9:0] ? 4'ha : _GEN_10775; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10777 = 10'hdc == _T_244[9:0] ? 4'ha : _GEN_10776; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10778 = 10'hdd == _T_244[9:0] ? 4'h3 : _GEN_10777; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10779 = 10'hde == _T_244[9:0] ? 4'h2 : _GEN_10778; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10780 = 10'hdf == _T_244[9:0] ? 4'h0 : _GEN_10779; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10781 = 10'he0 == _T_244[9:0] ? 4'ha : _GEN_10780; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10782 = 10'he1 == _T_244[9:0] ? 4'ha : _GEN_10781; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10783 = 10'he2 == _T_244[9:0] ? 4'h3 : _GEN_10782; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10784 = 10'he3 == _T_244[9:0] ? 4'ha : _GEN_10783; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10785 = 10'he4 == _T_244[9:0] ? 4'ha : _GEN_10784; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10786 = 10'he5 == _T_244[9:0] ? 4'ha : _GEN_10785; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10787 = 10'he6 == _T_244[9:0] ? 4'ha : _GEN_10786; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10788 = 10'he7 == _T_244[9:0] ? 4'h1 : _GEN_10787; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10789 = 10'he8 == _T_244[9:0] ? 4'h1 : _GEN_10788; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10790 = 10'he9 == _T_244[9:0] ? 4'h1 : _GEN_10789; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10791 = 10'hea == _T_244[9:0] ? 4'h0 : _GEN_10790; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10792 = 10'heb == _T_244[9:0] ? 4'h0 : _GEN_10791; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10793 = 10'hec == _T_244[9:0] ? 4'h0 : _GEN_10792; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10794 = 10'hed == _T_244[9:0] ? 4'h0 : _GEN_10793; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10795 = 10'hee == _T_244[9:0] ? 4'h0 : _GEN_10794; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10796 = 10'hef == _T_244[9:0] ? 4'h0 : _GEN_10795; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10797 = 10'hf0 == _T_244[9:0] ? 4'h0 : _GEN_10796; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10798 = 10'hf1 == _T_244[9:0] ? 4'h0 : _GEN_10797; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10799 = 10'hf2 == _T_244[9:0] ? 4'h0 : _GEN_10798; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10800 = 10'hf3 == _T_244[9:0] ? 4'h0 : _GEN_10799; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10801 = 10'hf4 == _T_244[9:0] ? 4'h0 : _GEN_10800; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10802 = 10'hf5 == _T_244[9:0] ? 4'h1 : _GEN_10801; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10803 = 10'hf6 == _T_244[9:0] ? 4'h0 : _GEN_10802; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10804 = 10'hf7 == _T_244[9:0] ? 4'h0 : _GEN_10803; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10805 = 10'hf8 == _T_244[9:0] ? 4'h1 : _GEN_10804; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10806 = 10'hf9 == _T_244[9:0] ? 4'h0 : _GEN_10805; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10807 = 10'hfa == _T_244[9:0] ? 4'ha : _GEN_10806; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10808 = 10'hfb == _T_244[9:0] ? 4'ha : _GEN_10807; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10809 = 10'hfc == _T_244[9:0] ? 4'ha : _GEN_10808; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10810 = 10'hfd == _T_244[9:0] ? 4'h3 : _GEN_10809; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10811 = 10'hfe == _T_244[9:0] ? 4'ha : _GEN_10810; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10812 = 10'hff == _T_244[9:0] ? 4'h0 : _GEN_10811; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10813 = 10'h100 == _T_244[9:0] ? 4'ha : _GEN_10812; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10814 = 10'h101 == _T_244[9:0] ? 4'h0 : _GEN_10813; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10815 = 10'h102 == _T_244[9:0] ? 4'h3 : _GEN_10814; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10816 = 10'h103 == _T_244[9:0] ? 4'ha : _GEN_10815; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10817 = 10'h104 == _T_244[9:0] ? 4'ha : _GEN_10816; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10818 = 10'h105 == _T_244[9:0] ? 4'ha : _GEN_10817; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10819 = 10'h106 == _T_244[9:0] ? 4'ha : _GEN_10818; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10820 = 10'h107 == _T_244[9:0] ? 4'ha : _GEN_10819; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10821 = 10'h108 == _T_244[9:0] ? 4'h1 : _GEN_10820; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10822 = 10'h109 == _T_244[9:0] ? 4'h0 : _GEN_10821; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10823 = 10'h10a == _T_244[9:0] ? 4'h0 : _GEN_10822; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10824 = 10'h10b == _T_244[9:0] ? 4'h0 : _GEN_10823; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10825 = 10'h10c == _T_244[9:0] ? 4'h0 : _GEN_10824; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10826 = 10'h10d == _T_244[9:0] ? 4'h0 : _GEN_10825; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10827 = 10'h10e == _T_244[9:0] ? 4'h0 : _GEN_10826; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10828 = 10'h10f == _T_244[9:0] ? 4'h0 : _GEN_10827; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10829 = 10'h110 == _T_244[9:0] ? 4'h0 : _GEN_10828; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10830 = 10'h111 == _T_244[9:0] ? 4'h0 : _GEN_10829; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10831 = 10'h112 == _T_244[9:0] ? 4'h0 : _GEN_10830; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10832 = 10'h113 == _T_244[9:0] ? 4'h0 : _GEN_10831; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10833 = 10'h114 == _T_244[9:0] ? 4'h0 : _GEN_10832; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10834 = 10'h115 == _T_244[9:0] ? 4'h0 : _GEN_10833; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10835 = 10'h116 == _T_244[9:0] ? 4'h1 : _GEN_10834; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10836 = 10'h117 == _T_244[9:0] ? 4'ha : _GEN_10835; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10837 = 10'h118 == _T_244[9:0] ? 4'ha : _GEN_10836; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10838 = 10'h119 == _T_244[9:0] ? 4'ha : _GEN_10837; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10839 = 10'h11a == _T_244[9:0] ? 4'h0 : _GEN_10838; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10840 = 10'h11b == _T_244[9:0] ? 4'ha : _GEN_10839; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10841 = 10'h11c == _T_244[9:0] ? 4'ha : _GEN_10840; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10842 = 10'h11d == _T_244[9:0] ? 4'h2 : _GEN_10841; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10843 = 10'h11e == _T_244[9:0] ? 4'h3 : _GEN_10842; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10844 = 10'h11f == _T_244[9:0] ? 4'h0 : _GEN_10843; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10845 = 10'h120 == _T_244[9:0] ? 4'ha : _GEN_10844; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10846 = 10'h121 == _T_244[9:0] ? 4'ha : _GEN_10845; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10847 = 10'h122 == _T_244[9:0] ? 4'h3 : _GEN_10846; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10848 = 10'h123 == _T_244[9:0] ? 4'ha : _GEN_10847; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10849 = 10'h124 == _T_244[9:0] ? 4'ha : _GEN_10848; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10850 = 10'h125 == _T_244[9:0] ? 4'ha : _GEN_10849; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10851 = 10'h126 == _T_244[9:0] ? 4'ha : _GEN_10850; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10852 = 10'h127 == _T_244[9:0] ? 4'h1 : _GEN_10851; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10853 = 10'h128 == _T_244[9:0] ? 4'h0 : _GEN_10852; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10854 = 10'h129 == _T_244[9:0] ? 4'ha : _GEN_10853; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10855 = 10'h12a == _T_244[9:0] ? 4'ha : _GEN_10854; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10856 = 10'h12b == _T_244[9:0] ? 4'h0 : _GEN_10855; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10857 = 10'h12c == _T_244[9:0] ? 4'h0 : _GEN_10856; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10858 = 10'h12d == _T_244[9:0] ? 4'h0 : _GEN_10857; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10859 = 10'h12e == _T_244[9:0] ? 4'h0 : _GEN_10858; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10860 = 10'h12f == _T_244[9:0] ? 4'h0 : _GEN_10859; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10861 = 10'h130 == _T_244[9:0] ? 4'h0 : _GEN_10860; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10862 = 10'h131 == _T_244[9:0] ? 4'h0 : _GEN_10861; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10863 = 10'h132 == _T_244[9:0] ? 4'h0 : _GEN_10862; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10864 = 10'h133 == _T_244[9:0] ? 4'h0 : _GEN_10863; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10865 = 10'h134 == _T_244[9:0] ? 4'ha : _GEN_10864; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10866 = 10'h135 == _T_244[9:0] ? 4'ha : _GEN_10865; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10867 = 10'h136 == _T_244[9:0] ? 4'h0 : _GEN_10866; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10868 = 10'h137 == _T_244[9:0] ? 4'h1 : _GEN_10867; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10869 = 10'h138 == _T_244[9:0] ? 4'ha : _GEN_10868; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10870 = 10'h139 == _T_244[9:0] ? 4'ha : _GEN_10869; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10871 = 10'h13a == _T_244[9:0] ? 4'ha : _GEN_10870; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10872 = 10'h13b == _T_244[9:0] ? 4'ha : _GEN_10871; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10873 = 10'h13c == _T_244[9:0] ? 4'ha : _GEN_10872; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10874 = 10'h13d == _T_244[9:0] ? 4'ha : _GEN_10873; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10875 = 10'h13e == _T_244[9:0] ? 4'h3 : _GEN_10874; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10876 = 10'h13f == _T_244[9:0] ? 4'h0 : _GEN_10875; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10877 = 10'h140 == _T_244[9:0] ? 4'ha : _GEN_10876; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10878 = 10'h141 == _T_244[9:0] ? 4'ha : _GEN_10877; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10879 = 10'h142 == _T_244[9:0] ? 4'h2 : _GEN_10878; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10880 = 10'h143 == _T_244[9:0] ? 4'h3 : _GEN_10879; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10881 = 10'h144 == _T_244[9:0] ? 4'ha : _GEN_10880; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10882 = 10'h145 == _T_244[9:0] ? 4'ha : _GEN_10881; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10883 = 10'h146 == _T_244[9:0] ? 4'h1 : _GEN_10882; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10884 = 10'h147 == _T_244[9:0] ? 4'h0 : _GEN_10883; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10885 = 10'h148 == _T_244[9:0] ? 4'ha : _GEN_10884; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10886 = 10'h149 == _T_244[9:0] ? 4'ha : _GEN_10885; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10887 = 10'h14a == _T_244[9:0] ? 4'ha : _GEN_10886; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10888 = 10'h14b == _T_244[9:0] ? 4'ha : _GEN_10887; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10889 = 10'h14c == _T_244[9:0] ? 4'ha : _GEN_10888; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10890 = 10'h14d == _T_244[9:0] ? 4'ha : _GEN_10889; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10891 = 10'h14e == _T_244[9:0] ? 4'ha : _GEN_10890; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10892 = 10'h14f == _T_244[9:0] ? 4'ha : _GEN_10891; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10893 = 10'h150 == _T_244[9:0] ? 4'ha : _GEN_10892; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10894 = 10'h151 == _T_244[9:0] ? 4'ha : _GEN_10893; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10895 = 10'h152 == _T_244[9:0] ? 4'ha : _GEN_10894; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10896 = 10'h153 == _T_244[9:0] ? 4'ha : _GEN_10895; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10897 = 10'h154 == _T_244[9:0] ? 4'ha : _GEN_10896; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10898 = 10'h155 == _T_244[9:0] ? 4'ha : _GEN_10897; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10899 = 10'h156 == _T_244[9:0] ? 4'ha : _GEN_10898; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10900 = 10'h157 == _T_244[9:0] ? 4'h0 : _GEN_10899; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10901 = 10'h158 == _T_244[9:0] ? 4'ha : _GEN_10900; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10902 = 10'h159 == _T_244[9:0] ? 4'ha : _GEN_10901; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10903 = 10'h15a == _T_244[9:0] ? 4'ha : _GEN_10902; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10904 = 10'h15b == _T_244[9:0] ? 4'ha : _GEN_10903; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10905 = 10'h15c == _T_244[9:0] ? 4'ha : _GEN_10904; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10906 = 10'h15d == _T_244[9:0] ? 4'h3 : _GEN_10905; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10907 = 10'h15e == _T_244[9:0] ? 4'h2 : _GEN_10906; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10908 = 10'h15f == _T_244[9:0] ? 4'h0 : _GEN_10907; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10909 = 10'h160 == _T_244[9:0] ? 4'ha : _GEN_10908; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10910 = 10'h161 == _T_244[9:0] ? 4'ha : _GEN_10909; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10911 = 10'h162 == _T_244[9:0] ? 4'ha : _GEN_10910; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10912 = 10'h163 == _T_244[9:0] ? 4'h2 : _GEN_10911; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10913 = 10'h164 == _T_244[9:0] ? 4'h3 : _GEN_10912; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10914 = 10'h165 == _T_244[9:0] ? 4'h1 : _GEN_10913; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10915 = 10'h166 == _T_244[9:0] ? 4'h0 : _GEN_10914; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10916 = 10'h167 == _T_244[9:0] ? 4'h0 : _GEN_10915; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10917 = 10'h168 == _T_244[9:0] ? 4'h5 : _GEN_10916; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10918 = 10'h169 == _T_244[9:0] ? 4'h3 : _GEN_10917; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10919 = 10'h16a == _T_244[9:0] ? 4'h5 : _GEN_10918; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10920 = 10'h16b == _T_244[9:0] ? 4'h5 : _GEN_10919; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10921 = 10'h16c == _T_244[9:0] ? 4'ha : _GEN_10920; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10922 = 10'h16d == _T_244[9:0] ? 4'ha : _GEN_10921; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10923 = 10'h16e == _T_244[9:0] ? 4'ha : _GEN_10922; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10924 = 10'h16f == _T_244[9:0] ? 4'ha : _GEN_10923; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10925 = 10'h170 == _T_244[9:0] ? 4'ha : _GEN_10924; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10926 = 10'h171 == _T_244[9:0] ? 4'ha : _GEN_10925; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10927 = 10'h172 == _T_244[9:0] ? 4'ha : _GEN_10926; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10928 = 10'h173 == _T_244[9:0] ? 4'ha : _GEN_10927; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10929 = 10'h174 == _T_244[9:0] ? 4'ha : _GEN_10928; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10930 = 10'h175 == _T_244[9:0] ? 4'ha : _GEN_10929; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10931 = 10'h176 == _T_244[9:0] ? 4'h0 : _GEN_10930; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10932 = 10'h177 == _T_244[9:0] ? 4'h0 : _GEN_10931; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10933 = 10'h178 == _T_244[9:0] ? 4'h1 : _GEN_10932; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10934 = 10'h179 == _T_244[9:0] ? 4'ha : _GEN_10933; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10935 = 10'h17a == _T_244[9:0] ? 4'ha : _GEN_10934; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10936 = 10'h17b == _T_244[9:0] ? 4'ha : _GEN_10935; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10937 = 10'h17c == _T_244[9:0] ? 4'h3 : _GEN_10936; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10938 = 10'h17d == _T_244[9:0] ? 4'h2 : _GEN_10937; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10939 = 10'h17e == _T_244[9:0] ? 4'ha : _GEN_10938; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10940 = 10'h17f == _T_244[9:0] ? 4'h0 : _GEN_10939; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10941 = 10'h180 == _T_244[9:0] ? 4'h5 : _GEN_10940; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10942 = 10'h181 == _T_244[9:0] ? 4'h5 : _GEN_10941; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10943 = 10'h182 == _T_244[9:0] ? 4'h5 : _GEN_10942; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10944 = 10'h183 == _T_244[9:0] ? 4'h5 : _GEN_10943; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10945 = 10'h184 == _T_244[9:0] ? 4'h3 : _GEN_10944; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10946 = 10'h185 == _T_244[9:0] ? 4'h1 : _GEN_10945; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10947 = 10'h186 == _T_244[9:0] ? 4'hb : _GEN_10946; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10948 = 10'h187 == _T_244[9:0] ? 4'h0 : _GEN_10947; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10949 = 10'h188 == _T_244[9:0] ? 4'h5 : _GEN_10948; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10950 = 10'h189 == _T_244[9:0] ? 4'h5 : _GEN_10949; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10951 = 10'h18a == _T_244[9:0] ? 4'h5 : _GEN_10950; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10952 = 10'h18b == _T_244[9:0] ? 4'h5 : _GEN_10951; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10953 = 10'h18c == _T_244[9:0] ? 4'h5 : _GEN_10952; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10954 = 10'h18d == _T_244[9:0] ? 4'h5 : _GEN_10953; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10955 = 10'h18e == _T_244[9:0] ? 4'h5 : _GEN_10954; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10956 = 10'h18f == _T_244[9:0] ? 4'h5 : _GEN_10955; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10957 = 10'h190 == _T_244[9:0] ? 4'h5 : _GEN_10956; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10958 = 10'h191 == _T_244[9:0] ? 4'h5 : _GEN_10957; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10959 = 10'h192 == _T_244[9:0] ? 4'h3 : _GEN_10958; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10960 = 10'h193 == _T_244[9:0] ? 4'h5 : _GEN_10959; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10961 = 10'h194 == _T_244[9:0] ? 4'h5 : _GEN_10960; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10962 = 10'h195 == _T_244[9:0] ? 4'h5 : _GEN_10961; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10963 = 10'h196 == _T_244[9:0] ? 4'h0 : _GEN_10962; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10964 = 10'h197 == _T_244[9:0] ? 4'ha : _GEN_10963; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10965 = 10'h198 == _T_244[9:0] ? 4'h1 : _GEN_10964; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10966 = 10'h199 == _T_244[9:0] ? 4'ha : _GEN_10965; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10967 = 10'h19a == _T_244[9:0] ? 4'ha : _GEN_10966; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10968 = 10'h19b == _T_244[9:0] ? 4'ha : _GEN_10967; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10969 = 10'h19c == _T_244[9:0] ? 4'h3 : _GEN_10968; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10970 = 10'h19d == _T_244[9:0] ? 4'ha : _GEN_10969; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10971 = 10'h19e == _T_244[9:0] ? 4'ha : _GEN_10970; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10972 = 10'h19f == _T_244[9:0] ? 4'h0 : _GEN_10971; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10973 = 10'h1a0 == _T_244[9:0] ? 4'h5 : _GEN_10972; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10974 = 10'h1a1 == _T_244[9:0] ? 4'h5 : _GEN_10973; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10975 = 10'h1a2 == _T_244[9:0] ? 4'h3 : _GEN_10974; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10976 = 10'h1a3 == _T_244[9:0] ? 4'h5 : _GEN_10975; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10977 = 10'h1a4 == _T_244[9:0] ? 4'h3 : _GEN_10976; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10978 = 10'h1a5 == _T_244[9:0] ? 4'h0 : _GEN_10977; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10979 = 10'h1a6 == _T_244[9:0] ? 4'h5 : _GEN_10978; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10980 = 10'h1a7 == _T_244[9:0] ? 4'h0 : _GEN_10979; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10981 = 10'h1a8 == _T_244[9:0] ? 4'hb : _GEN_10980; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10982 = 10'h1a9 == _T_244[9:0] ? 4'h5 : _GEN_10981; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10983 = 10'h1aa == _T_244[9:0] ? 4'h5 : _GEN_10982; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10984 = 10'h1ab == _T_244[9:0] ? 4'h3 : _GEN_10983; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10985 = 10'h1ac == _T_244[9:0] ? 4'h5 : _GEN_10984; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10986 = 10'h1ad == _T_244[9:0] ? 4'h5 : _GEN_10985; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10987 = 10'h1ae == _T_244[9:0] ? 4'h5 : _GEN_10986; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10988 = 10'h1af == _T_244[9:0] ? 4'h5 : _GEN_10987; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10989 = 10'h1b0 == _T_244[9:0] ? 4'h5 : _GEN_10988; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10990 = 10'h1b1 == _T_244[9:0] ? 4'h5 : _GEN_10989; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10991 = 10'h1b2 == _T_244[9:0] ? 4'h5 : _GEN_10990; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10992 = 10'h1b3 == _T_244[9:0] ? 4'h5 : _GEN_10991; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10993 = 10'h1b4 == _T_244[9:0] ? 4'h5 : _GEN_10992; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10994 = 10'h1b5 == _T_244[9:0] ? 4'h5 : _GEN_10993; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10995 = 10'h1b6 == _T_244[9:0] ? 4'h0 : _GEN_10994; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10996 = 10'h1b7 == _T_244[9:0] ? 4'h5 : _GEN_10995; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10997 = 10'h1b8 == _T_244[9:0] ? 4'h0 : _GEN_10996; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10998 = 10'h1b9 == _T_244[9:0] ? 4'h5 : _GEN_10997; // @[Filter.scala 191:62]
  wire [3:0] _GEN_10999 = 10'h1ba == _T_244[9:0] ? 4'h5 : _GEN_10998; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11000 = 10'h1bb == _T_244[9:0] ? 4'h5 : _GEN_10999; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11001 = 10'h1bc == _T_244[9:0] ? 4'h2 : _GEN_11000; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11002 = 10'h1bd == _T_244[9:0] ? 4'h3 : _GEN_11001; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11003 = 10'h1be == _T_244[9:0] ? 4'h5 : _GEN_11002; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11004 = 10'h1bf == _T_244[9:0] ? 4'h0 : _GEN_11003; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11005 = 10'h1c0 == _T_244[9:0] ? 4'h5 : _GEN_11004; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11006 = 10'h1c1 == _T_244[9:0] ? 4'h5 : _GEN_11005; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11007 = 10'h1c2 == _T_244[9:0] ? 4'h5 : _GEN_11006; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11008 = 10'h1c3 == _T_244[9:0] ? 4'h2 : _GEN_11007; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11009 = 10'h1c4 == _T_244[9:0] ? 4'h2 : _GEN_11008; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11010 = 10'h1c5 == _T_244[9:0] ? 4'h5 : _GEN_11009; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11011 = 10'h1c6 == _T_244[9:0] ? 4'h5 : _GEN_11010; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11012 = 10'h1c7 == _T_244[9:0] ? 4'h5 : _GEN_11011; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11013 = 10'h1c8 == _T_244[9:0] ? 4'h5 : _GEN_11012; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11014 = 10'h1c9 == _T_244[9:0] ? 4'hb : _GEN_11013; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11015 = 10'h1ca == _T_244[9:0] ? 4'hb : _GEN_11014; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11016 = 10'h1cb == _T_244[9:0] ? 4'hb : _GEN_11015; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11017 = 10'h1cc == _T_244[9:0] ? 4'hb : _GEN_11016; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11018 = 10'h1cd == _T_244[9:0] ? 4'hb : _GEN_11017; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11019 = 10'h1ce == _T_244[9:0] ? 4'hb : _GEN_11018; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11020 = 10'h1cf == _T_244[9:0] ? 4'hb : _GEN_11019; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11021 = 10'h1d0 == _T_244[9:0] ? 4'hb : _GEN_11020; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11022 = 10'h1d1 == _T_244[9:0] ? 4'hb : _GEN_11021; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11023 = 10'h1d2 == _T_244[9:0] ? 4'hb : _GEN_11022; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11024 = 10'h1d3 == _T_244[9:0] ? 4'hb : _GEN_11023; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11025 = 10'h1d4 == _T_244[9:0] ? 4'hb : _GEN_11024; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11026 = 10'h1d5 == _T_244[9:0] ? 4'hb : _GEN_11025; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11027 = 10'h1d6 == _T_244[9:0] ? 4'h5 : _GEN_11026; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11028 = 10'h1d7 == _T_244[9:0] ? 4'h5 : _GEN_11027; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11029 = 10'h1d8 == _T_244[9:0] ? 4'h5 : _GEN_11028; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11030 = 10'h1d9 == _T_244[9:0] ? 4'h5 : _GEN_11029; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11031 = 10'h1da == _T_244[9:0] ? 4'h5 : _GEN_11030; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11032 = 10'h1db == _T_244[9:0] ? 4'h5 : _GEN_11031; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11033 = 10'h1dc == _T_244[9:0] ? 4'h5 : _GEN_11032; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11034 = 10'h1dd == _T_244[9:0] ? 4'h3 : _GEN_11033; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11035 = 10'h1de == _T_244[9:0] ? 4'h5 : _GEN_11034; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11036 = 10'h1df == _T_244[9:0] ? 4'h0 : _GEN_11035; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11037 = 10'h1e0 == _T_244[9:0] ? 4'h3 : _GEN_11036; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11038 = 10'h1e1 == _T_244[9:0] ? 4'h5 : _GEN_11037; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11039 = 10'h1e2 == _T_244[9:0] ? 4'h2 : _GEN_11038; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11040 = 10'h1e3 == _T_244[9:0] ? 4'h2 : _GEN_11039; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11041 = 10'h1e4 == _T_244[9:0] ? 4'h5 : _GEN_11040; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11042 = 10'h1e5 == _T_244[9:0] ? 4'h5 : _GEN_11041; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11043 = 10'h1e6 == _T_244[9:0] ? 4'h5 : _GEN_11042; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11044 = 10'h1e7 == _T_244[9:0] ? 4'h5 : _GEN_11043; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11045 = 10'h1e8 == _T_244[9:0] ? 4'hb : _GEN_11044; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11046 = 10'h1e9 == _T_244[9:0] ? 4'h5 : _GEN_11045; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11047 = 10'h1ea == _T_244[9:0] ? 4'h5 : _GEN_11046; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11048 = 10'h1eb == _T_244[9:0] ? 4'hb : _GEN_11047; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11049 = 10'h1ec == _T_244[9:0] ? 4'h5 : _GEN_11048; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11050 = 10'h1ed == _T_244[9:0] ? 4'hb : _GEN_11049; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11051 = 10'h1ee == _T_244[9:0] ? 4'h5 : _GEN_11050; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11052 = 10'h1ef == _T_244[9:0] ? 4'hb : _GEN_11051; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11053 = 10'h1f0 == _T_244[9:0] ? 4'h5 : _GEN_11052; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11054 = 10'h1f1 == _T_244[9:0] ? 4'hb : _GEN_11053; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11055 = 10'h1f2 == _T_244[9:0] ? 4'hb : _GEN_11054; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11056 = 10'h1f3 == _T_244[9:0] ? 4'h5 : _GEN_11055; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11057 = 10'h1f4 == _T_244[9:0] ? 4'hb : _GEN_11056; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11058 = 10'h1f5 == _T_244[9:0] ? 4'hb : _GEN_11057; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11059 = 10'h1f6 == _T_244[9:0] ? 4'h5 : _GEN_11058; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11060 = 10'h1f7 == _T_244[9:0] ? 4'h5 : _GEN_11059; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11061 = 10'h1f8 == _T_244[9:0] ? 4'h5 : _GEN_11060; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11062 = 10'h1f9 == _T_244[9:0] ? 4'h5 : _GEN_11061; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11063 = 10'h1fa == _T_244[9:0] ? 4'h3 : _GEN_11062; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11064 = 10'h1fb == _T_244[9:0] ? 4'h5 : _GEN_11063; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11065 = 10'h1fc == _T_244[9:0] ? 4'h5 : _GEN_11064; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11066 = 10'h1fd == _T_244[9:0] ? 4'h2 : _GEN_11065; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11067 = 10'h1fe == _T_244[9:0] ? 4'h5 : _GEN_11066; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11068 = 10'h1ff == _T_244[9:0] ? 4'h0 : _GEN_11067; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11069 = 10'h200 == _T_244[9:0] ? 4'h5 : _GEN_11068; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11070 = 10'h201 == _T_244[9:0] ? 4'h5 : _GEN_11069; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11071 = 10'h202 == _T_244[9:0] ? 4'h3 : _GEN_11070; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11072 = 10'h203 == _T_244[9:0] ? 4'h5 : _GEN_11071; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11073 = 10'h204 == _T_244[9:0] ? 4'h5 : _GEN_11072; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11074 = 10'h205 == _T_244[9:0] ? 4'h5 : _GEN_11073; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11075 = 10'h206 == _T_244[9:0] ? 4'hb : _GEN_11074; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11076 = 10'h207 == _T_244[9:0] ? 4'hb : _GEN_11075; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11077 = 10'h208 == _T_244[9:0] ? 4'h5 : _GEN_11076; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11078 = 10'h209 == _T_244[9:0] ? 4'h5 : _GEN_11077; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11079 = 10'h20a == _T_244[9:0] ? 4'h5 : _GEN_11078; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11080 = 10'h20b == _T_244[9:0] ? 4'hb : _GEN_11079; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11081 = 10'h20c == _T_244[9:0] ? 4'h5 : _GEN_11080; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11082 = 10'h20d == _T_244[9:0] ? 4'hb : _GEN_11081; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11083 = 10'h20e == _T_244[9:0] ? 4'h5 : _GEN_11082; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11084 = 10'h20f == _T_244[9:0] ? 4'hb : _GEN_11083; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11085 = 10'h210 == _T_244[9:0] ? 4'h5 : _GEN_11084; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11086 = 10'h211 == _T_244[9:0] ? 4'h5 : _GEN_11085; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11087 = 10'h212 == _T_244[9:0] ? 4'hb : _GEN_11086; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11088 = 10'h213 == _T_244[9:0] ? 4'hb : _GEN_11087; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11089 = 10'h214 == _T_244[9:0] ? 4'hb : _GEN_11088; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11090 = 10'h215 == _T_244[9:0] ? 4'h5 : _GEN_11089; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11091 = 10'h216 == _T_244[9:0] ? 4'h5 : _GEN_11090; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11092 = 10'h217 == _T_244[9:0] ? 4'h5 : _GEN_11091; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11093 = 10'h218 == _T_244[9:0] ? 4'h5 : _GEN_11092; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11094 = 10'h219 == _T_244[9:0] ? 4'h5 : _GEN_11093; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11095 = 10'h21a == _T_244[9:0] ? 4'h5 : _GEN_11094; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11096 = 10'h21b == _T_244[9:0] ? 4'h5 : _GEN_11095; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11097 = 10'h21c == _T_244[9:0] ? 4'h3 : _GEN_11096; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11098 = 10'h21d == _T_244[9:0] ? 4'h2 : _GEN_11097; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11099 = 10'h21e == _T_244[9:0] ? 4'h5 : _GEN_11098; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11100 = 10'h21f == _T_244[9:0] ? 4'h0 : _GEN_11099; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11101 = 10'h220 == _T_244[9:0] ? 4'h0 : _GEN_11100; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11102 = 10'h221 == _T_244[9:0] ? 4'h0 : _GEN_11101; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11103 = 10'h222 == _T_244[9:0] ? 4'h0 : _GEN_11102; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11104 = 10'h223 == _T_244[9:0] ? 4'h0 : _GEN_11103; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11105 = 10'h224 == _T_244[9:0] ? 4'h0 : _GEN_11104; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11106 = 10'h225 == _T_244[9:0] ? 4'h0 : _GEN_11105; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11107 = 10'h226 == _T_244[9:0] ? 4'h0 : _GEN_11106; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11108 = 10'h227 == _T_244[9:0] ? 4'h0 : _GEN_11107; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11109 = 10'h228 == _T_244[9:0] ? 4'h0 : _GEN_11108; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11110 = 10'h229 == _T_244[9:0] ? 4'h0 : _GEN_11109; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11111 = 10'h22a == _T_244[9:0] ? 4'h0 : _GEN_11110; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11112 = 10'h22b == _T_244[9:0] ? 4'h0 : _GEN_11111; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11113 = 10'h22c == _T_244[9:0] ? 4'h0 : _GEN_11112; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11114 = 10'h22d == _T_244[9:0] ? 4'h0 : _GEN_11113; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11115 = 10'h22e == _T_244[9:0] ? 4'h0 : _GEN_11114; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11116 = 10'h22f == _T_244[9:0] ? 4'h0 : _GEN_11115; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11117 = 10'h230 == _T_244[9:0] ? 4'h0 : _GEN_11116; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11118 = 10'h231 == _T_244[9:0] ? 4'h0 : _GEN_11117; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11119 = 10'h232 == _T_244[9:0] ? 4'h0 : _GEN_11118; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11120 = 10'h233 == _T_244[9:0] ? 4'h0 : _GEN_11119; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11121 = 10'h234 == _T_244[9:0] ? 4'h0 : _GEN_11120; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11122 = 10'h235 == _T_244[9:0] ? 4'h0 : _GEN_11121; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11123 = 10'h236 == _T_244[9:0] ? 4'h0 : _GEN_11122; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11124 = 10'h237 == _T_244[9:0] ? 4'h0 : _GEN_11123; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11125 = 10'h238 == _T_244[9:0] ? 4'h0 : _GEN_11124; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11126 = 10'h239 == _T_244[9:0] ? 4'h0 : _GEN_11125; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11127 = 10'h23a == _T_244[9:0] ? 4'h0 : _GEN_11126; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11128 = 10'h23b == _T_244[9:0] ? 4'h0 : _GEN_11127; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11129 = 10'h23c == _T_244[9:0] ? 4'h0 : _GEN_11128; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11130 = 10'h23d == _T_244[9:0] ? 4'h0 : _GEN_11129; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11131 = 10'h23e == _T_244[9:0] ? 4'h0 : _GEN_11130; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11132 = 10'h23f == _T_244[9:0] ? 4'h0 : _GEN_11131; // @[Filter.scala 191:62]
  wire [4:0] _GEN_28334 = {{1'd0}, _GEN_11132}; // @[Filter.scala 191:62]
  wire [8:0] _T_246 = _GEN_28334 * 5'h14; // @[Filter.scala 191:62]
  wire [3:0] _GEN_11136 = 10'h3 == _T_244[9:0] ? 4'ha : 4'h3; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11137 = 10'h4 == _T_244[9:0] ? 4'h3 : _GEN_11136; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11138 = 10'h5 == _T_244[9:0] ? 4'h3 : _GEN_11137; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11139 = 10'h6 == _T_244[9:0] ? 4'h3 : _GEN_11138; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11140 = 10'h7 == _T_244[9:0] ? 4'h3 : _GEN_11139; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11141 = 10'h8 == _T_244[9:0] ? 4'h3 : _GEN_11140; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11142 = 10'h9 == _T_244[9:0] ? 4'h3 : _GEN_11141; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11143 = 10'ha == _T_244[9:0] ? 4'h3 : _GEN_11142; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11144 = 10'hb == _T_244[9:0] ? 4'h3 : _GEN_11143; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11145 = 10'hc == _T_244[9:0] ? 4'h5 : _GEN_11144; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11146 = 10'hd == _T_244[9:0] ? 4'h3 : _GEN_11145; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11147 = 10'he == _T_244[9:0] ? 4'h3 : _GEN_11146; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11148 = 10'hf == _T_244[9:0] ? 4'h3 : _GEN_11147; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11149 = 10'h10 == _T_244[9:0] ? 4'h3 : _GEN_11148; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11150 = 10'h11 == _T_244[9:0] ? 4'h3 : _GEN_11149; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11151 = 10'h12 == _T_244[9:0] ? 4'h3 : _GEN_11150; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11152 = 10'h13 == _T_244[9:0] ? 4'h3 : _GEN_11151; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11153 = 10'h14 == _T_244[9:0] ? 4'h3 : _GEN_11152; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11154 = 10'h15 == _T_244[9:0] ? 4'h3 : _GEN_11153; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11155 = 10'h16 == _T_244[9:0] ? 4'h3 : _GEN_11154; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11156 = 10'h17 == _T_244[9:0] ? 4'h3 : _GEN_11155; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11157 = 10'h18 == _T_244[9:0] ? 4'h3 : _GEN_11156; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11158 = 10'h19 == _T_244[9:0] ? 4'h3 : _GEN_11157; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11159 = 10'h1a == _T_244[9:0] ? 4'h3 : _GEN_11158; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11160 = 10'h1b == _T_244[9:0] ? 4'h3 : _GEN_11159; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11161 = 10'h1c == _T_244[9:0] ? 4'h3 : _GEN_11160; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11162 = 10'h1d == _T_244[9:0] ? 4'h3 : _GEN_11161; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11163 = 10'h1e == _T_244[9:0] ? 4'h3 : _GEN_11162; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11164 = 10'h1f == _T_244[9:0] ? 4'h0 : _GEN_11163; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11165 = 10'h20 == _T_244[9:0] ? 4'h3 : _GEN_11164; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11166 = 10'h21 == _T_244[9:0] ? 4'h5 : _GEN_11165; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11167 = 10'h22 == _T_244[9:0] ? 4'h3 : _GEN_11166; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11168 = 10'h23 == _T_244[9:0] ? 4'ha : _GEN_11167; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11169 = 10'h24 == _T_244[9:0] ? 4'h3 : _GEN_11168; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11170 = 10'h25 == _T_244[9:0] ? 4'h3 : _GEN_11169; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11171 = 10'h26 == _T_244[9:0] ? 4'h3 : _GEN_11170; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11172 = 10'h27 == _T_244[9:0] ? 4'h1 : _GEN_11171; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11173 = 10'h28 == _T_244[9:0] ? 4'h1 : _GEN_11172; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11174 = 10'h29 == _T_244[9:0] ? 4'h3 : _GEN_11173; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11175 = 10'h2a == _T_244[9:0] ? 4'h3 : _GEN_11174; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11176 = 10'h2b == _T_244[9:0] ? 4'h3 : _GEN_11175; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11177 = 10'h2c == _T_244[9:0] ? 4'h3 : _GEN_11176; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11178 = 10'h2d == _T_244[9:0] ? 4'h3 : _GEN_11177; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11179 = 10'h2e == _T_244[9:0] ? 4'h3 : _GEN_11178; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11180 = 10'h2f == _T_244[9:0] ? 4'h3 : _GEN_11179; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11181 = 10'h30 == _T_244[9:0] ? 4'h3 : _GEN_11180; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11182 = 10'h31 == _T_244[9:0] ? 4'h5 : _GEN_11181; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11183 = 10'h32 == _T_244[9:0] ? 4'h3 : _GEN_11182; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11184 = 10'h33 == _T_244[9:0] ? 4'h3 : _GEN_11183; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11185 = 10'h34 == _T_244[9:0] ? 4'h3 : _GEN_11184; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11186 = 10'h35 == _T_244[9:0] ? 4'h3 : _GEN_11185; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11187 = 10'h36 == _T_244[9:0] ? 4'h3 : _GEN_11186; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11188 = 10'h37 == _T_244[9:0] ? 4'h1 : _GEN_11187; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11189 = 10'h38 == _T_244[9:0] ? 4'h1 : _GEN_11188; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11190 = 10'h39 == _T_244[9:0] ? 4'h3 : _GEN_11189; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11191 = 10'h3a == _T_244[9:0] ? 4'h3 : _GEN_11190; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11192 = 10'h3b == _T_244[9:0] ? 4'h5 : _GEN_11191; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11193 = 10'h3c == _T_244[9:0] ? 4'h3 : _GEN_11192; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11194 = 10'h3d == _T_244[9:0] ? 4'ha : _GEN_11193; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11195 = 10'h3e == _T_244[9:0] ? 4'h3 : _GEN_11194; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11196 = 10'h3f == _T_244[9:0] ? 4'h0 : _GEN_11195; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11197 = 10'h40 == _T_244[9:0] ? 4'h3 : _GEN_11196; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11198 = 10'h41 == _T_244[9:0] ? 4'h3 : _GEN_11197; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11199 = 10'h42 == _T_244[9:0] ? 4'h3 : _GEN_11198; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11200 = 10'h43 == _T_244[9:0] ? 4'h7 : _GEN_11199; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11201 = 10'h44 == _T_244[9:0] ? 4'ha : _GEN_11200; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11202 = 10'h45 == _T_244[9:0] ? 4'h0 : _GEN_11201; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11203 = 10'h46 == _T_244[9:0] ? 4'h0 : _GEN_11202; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11204 = 10'h47 == _T_244[9:0] ? 4'h0 : _GEN_11203; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11205 = 10'h48 == _T_244[9:0] ? 4'h0 : _GEN_11204; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11206 = 10'h49 == _T_244[9:0] ? 4'h3 : _GEN_11205; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11207 = 10'h4a == _T_244[9:0] ? 4'h3 : _GEN_11206; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11208 = 10'h4b == _T_244[9:0] ? 4'h3 : _GEN_11207; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11209 = 10'h4c == _T_244[9:0] ? 4'h3 : _GEN_11208; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11210 = 10'h4d == _T_244[9:0] ? 4'h5 : _GEN_11209; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11211 = 10'h4e == _T_244[9:0] ? 4'h3 : _GEN_11210; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11212 = 10'h4f == _T_244[9:0] ? 4'h3 : _GEN_11211; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11213 = 10'h50 == _T_244[9:0] ? 4'h3 : _GEN_11212; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11214 = 10'h51 == _T_244[9:0] ? 4'h3 : _GEN_11213; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11215 = 10'h52 == _T_244[9:0] ? 4'h3 : _GEN_11214; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11216 = 10'h53 == _T_244[9:0] ? 4'h3 : _GEN_11215; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11217 = 10'h54 == _T_244[9:0] ? 4'h1 : _GEN_11216; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11218 = 10'h55 == _T_244[9:0] ? 4'h1 : _GEN_11217; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11219 = 10'h56 == _T_244[9:0] ? 4'h1 : _GEN_11218; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11220 = 10'h57 == _T_244[9:0] ? 4'h0 : _GEN_11219; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11221 = 10'h58 == _T_244[9:0] ? 4'h3 : _GEN_11220; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11222 = 10'h59 == _T_244[9:0] ? 4'h0 : _GEN_11221; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11223 = 10'h5a == _T_244[9:0] ? 4'h3 : _GEN_11222; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11224 = 10'h5b == _T_244[9:0] ? 4'h3 : _GEN_11223; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11225 = 10'h5c == _T_244[9:0] ? 4'h3 : _GEN_11224; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11226 = 10'h5d == _T_244[9:0] ? 4'ha : _GEN_11225; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11227 = 10'h5e == _T_244[9:0] ? 4'h3 : _GEN_11226; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11228 = 10'h5f == _T_244[9:0] ? 4'h0 : _GEN_11227; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11229 = 10'h60 == _T_244[9:0] ? 4'h3 : _GEN_11228; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11230 = 10'h61 == _T_244[9:0] ? 4'h3 : _GEN_11229; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11231 = 10'h62 == _T_244[9:0] ? 4'h3 : _GEN_11230; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11232 = 10'h63 == _T_244[9:0] ? 4'h3 : _GEN_11231; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11233 = 10'h64 == _T_244[9:0] ? 4'ha : _GEN_11232; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11234 = 10'h65 == _T_244[9:0] ? 4'h0 : _GEN_11233; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11235 = 10'h66 == _T_244[9:0] ? 4'h3 : _GEN_11234; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11236 = 10'h67 == _T_244[9:0] ? 4'h3 : _GEN_11235; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11237 = 10'h68 == _T_244[9:0] ? 4'h3 : _GEN_11236; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11238 = 10'h69 == _T_244[9:0] ? 4'h0 : _GEN_11237; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11239 = 10'h6a == _T_244[9:0] ? 4'h1 : _GEN_11238; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11240 = 10'h6b == _T_244[9:0] ? 4'h1 : _GEN_11239; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11241 = 10'h6c == _T_244[9:0] ? 4'h3 : _GEN_11240; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11242 = 10'h6d == _T_244[9:0] ? 4'h3 : _GEN_11241; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11243 = 10'h6e == _T_244[9:0] ? 4'h3 : _GEN_11242; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11244 = 10'h6f == _T_244[9:0] ? 4'h3 : _GEN_11243; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11245 = 10'h70 == _T_244[9:0] ? 4'h3 : _GEN_11244; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11246 = 10'h71 == _T_244[9:0] ? 4'h3 : _GEN_11245; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11247 = 10'h72 == _T_244[9:0] ? 4'h3 : _GEN_11246; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11248 = 10'h73 == _T_244[9:0] ? 4'h1 : _GEN_11247; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11249 = 10'h74 == _T_244[9:0] ? 4'h0 : _GEN_11248; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11250 = 10'h75 == _T_244[9:0] ? 4'h0 : _GEN_11249; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11251 = 10'h76 == _T_244[9:0] ? 4'h0 : _GEN_11250; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11252 = 10'h77 == _T_244[9:0] ? 4'h3 : _GEN_11251; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11253 = 10'h78 == _T_244[9:0] ? 4'h3 : _GEN_11252; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11254 = 10'h79 == _T_244[9:0] ? 4'h3 : _GEN_11253; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11255 = 10'h7a == _T_244[9:0] ? 4'h0 : _GEN_11254; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11256 = 10'h7b == _T_244[9:0] ? 4'h3 : _GEN_11255; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11257 = 10'h7c == _T_244[9:0] ? 4'h3 : _GEN_11256; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11258 = 10'h7d == _T_244[9:0] ? 4'h7 : _GEN_11257; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11259 = 10'h7e == _T_244[9:0] ? 4'ha : _GEN_11258; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11260 = 10'h7f == _T_244[9:0] ? 4'h0 : _GEN_11259; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11261 = 10'h80 == _T_244[9:0] ? 4'h3 : _GEN_11260; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11262 = 10'h81 == _T_244[9:0] ? 4'h3 : _GEN_11261; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11263 = 10'h82 == _T_244[9:0] ? 4'h1 : _GEN_11262; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11264 = 10'h83 == _T_244[9:0] ? 4'h0 : _GEN_11263; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11265 = 10'h84 == _T_244[9:0] ? 4'h7 : _GEN_11264; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11266 = 10'h85 == _T_244[9:0] ? 4'h1 : _GEN_11265; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11267 = 10'h86 == _T_244[9:0] ? 4'h1 : _GEN_11266; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11268 = 10'h87 == _T_244[9:0] ? 4'h3 : _GEN_11267; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11269 = 10'h88 == _T_244[9:0] ? 4'h3 : _GEN_11268; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11270 = 10'h89 == _T_244[9:0] ? 4'h0 : _GEN_11269; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11271 = 10'h8a == _T_244[9:0] ? 4'h0 : _GEN_11270; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11272 = 10'h8b == _T_244[9:0] ? 4'h1 : _GEN_11271; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11273 = 10'h8c == _T_244[9:0] ? 4'h1 : _GEN_11272; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11274 = 10'h8d == _T_244[9:0] ? 4'h1 : _GEN_11273; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11275 = 10'h8e == _T_244[9:0] ? 4'h1 : _GEN_11274; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11276 = 10'h8f == _T_244[9:0] ? 4'h1 : _GEN_11275; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11277 = 10'h90 == _T_244[9:0] ? 4'h1 : _GEN_11276; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11278 = 10'h91 == _T_244[9:0] ? 4'h1 : _GEN_11277; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11279 = 10'h92 == _T_244[9:0] ? 4'h1 : _GEN_11278; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11280 = 10'h93 == _T_244[9:0] ? 4'h0 : _GEN_11279; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11281 = 10'h94 == _T_244[9:0] ? 4'h0 : _GEN_11280; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11282 = 10'h95 == _T_244[9:0] ? 4'h3 : _GEN_11281; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11283 = 10'h96 == _T_244[9:0] ? 4'h3 : _GEN_11282; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11284 = 10'h97 == _T_244[9:0] ? 4'h3 : _GEN_11283; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11285 = 10'h98 == _T_244[9:0] ? 4'h1 : _GEN_11284; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11286 = 10'h99 == _T_244[9:0] ? 4'h0 : _GEN_11285; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11287 = 10'h9a == _T_244[9:0] ? 4'h1 : _GEN_11286; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11288 = 10'h9b == _T_244[9:0] ? 4'h1 : _GEN_11287; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11289 = 10'h9c == _T_244[9:0] ? 4'h3 : _GEN_11288; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11290 = 10'h9d == _T_244[9:0] ? 4'h3 : _GEN_11289; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11291 = 10'h9e == _T_244[9:0] ? 4'ha : _GEN_11290; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11292 = 10'h9f == _T_244[9:0] ? 4'h0 : _GEN_11291; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11293 = 10'ha0 == _T_244[9:0] ? 4'h3 : _GEN_11292; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11294 = 10'ha1 == _T_244[9:0] ? 4'h1 : _GEN_11293; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11295 = 10'ha2 == _T_244[9:0] ? 4'h0 : _GEN_11294; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11296 = 10'ha3 == _T_244[9:0] ? 4'ha : _GEN_11295; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11297 = 10'ha4 == _T_244[9:0] ? 4'h3 : _GEN_11296; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11298 = 10'ha5 == _T_244[9:0] ? 4'h3 : _GEN_11297; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11299 = 10'ha6 == _T_244[9:0] ? 4'h3 : _GEN_11298; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11300 = 10'ha7 == _T_244[9:0] ? 4'h0 : _GEN_11299; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11301 = 10'ha8 == _T_244[9:0] ? 4'h3 : _GEN_11300; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11302 = 10'ha9 == _T_244[9:0] ? 4'h1 : _GEN_11301; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11303 = 10'haa == _T_244[9:0] ? 4'h0 : _GEN_11302; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11304 = 10'hab == _T_244[9:0] ? 4'h0 : _GEN_11303; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11305 = 10'hac == _T_244[9:0] ? 4'h0 : _GEN_11304; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11306 = 10'had == _T_244[9:0] ? 4'h0 : _GEN_11305; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11307 = 10'hae == _T_244[9:0] ? 4'h0 : _GEN_11306; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11308 = 10'haf == _T_244[9:0] ? 4'h0 : _GEN_11307; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11309 = 10'hb0 == _T_244[9:0] ? 4'h0 : _GEN_11308; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11310 = 10'hb1 == _T_244[9:0] ? 4'h0 : _GEN_11309; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11311 = 10'hb2 == _T_244[9:0] ? 4'h0 : _GEN_11310; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11312 = 10'hb3 == _T_244[9:0] ? 4'h0 : _GEN_11311; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11313 = 10'hb4 == _T_244[9:0] ? 4'h1 : _GEN_11312; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11314 = 10'hb5 == _T_244[9:0] ? 4'h1 : _GEN_11313; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11315 = 10'hb6 == _T_244[9:0] ? 4'h3 : _GEN_11314; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11316 = 10'hb7 == _T_244[9:0] ? 4'h0 : _GEN_11315; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11317 = 10'hb8 == _T_244[9:0] ? 4'h3 : _GEN_11316; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11318 = 10'hb9 == _T_244[9:0] ? 4'h3 : _GEN_11317; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11319 = 10'hba == _T_244[9:0] ? 4'h3 : _GEN_11318; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11320 = 10'hbb == _T_244[9:0] ? 4'h0 : _GEN_11319; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11321 = 10'hbc == _T_244[9:0] ? 4'h3 : _GEN_11320; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11322 = 10'hbd == _T_244[9:0] ? 4'h3 : _GEN_11321; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11323 = 10'hbe == _T_244[9:0] ? 4'ha : _GEN_11322; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11324 = 10'hbf == _T_244[9:0] ? 4'h0 : _GEN_11323; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11325 = 10'hc0 == _T_244[9:0] ? 4'h3 : _GEN_11324; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11326 = 10'hc1 == _T_244[9:0] ? 4'h3 : _GEN_11325; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11327 = 10'hc2 == _T_244[9:0] ? 4'ha : _GEN_11326; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11328 = 10'hc3 == _T_244[9:0] ? 4'h7 : _GEN_11327; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11329 = 10'hc4 == _T_244[9:0] ? 4'h0 : _GEN_11328; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11330 = 10'hc5 == _T_244[9:0] ? 4'h0 : _GEN_11329; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11331 = 10'hc6 == _T_244[9:0] ? 4'h0 : _GEN_11330; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11332 = 10'hc7 == _T_244[9:0] ? 4'h3 : _GEN_11331; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11333 = 10'hc8 == _T_244[9:0] ? 4'h1 : _GEN_11332; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11334 = 10'hc9 == _T_244[9:0] ? 4'h0 : _GEN_11333; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11335 = 10'hca == _T_244[9:0] ? 4'h0 : _GEN_11334; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11336 = 10'hcb == _T_244[9:0] ? 4'h0 : _GEN_11335; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11337 = 10'hcc == _T_244[9:0] ? 4'h0 : _GEN_11336; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11338 = 10'hcd == _T_244[9:0] ? 4'h0 : _GEN_11337; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11339 = 10'hce == _T_244[9:0] ? 4'h0 : _GEN_11338; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11340 = 10'hcf == _T_244[9:0] ? 4'h0 : _GEN_11339; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11341 = 10'hd0 == _T_244[9:0] ? 4'h0 : _GEN_11340; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11342 = 10'hd1 == _T_244[9:0] ? 4'h0 : _GEN_11341; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11343 = 10'hd2 == _T_244[9:0] ? 4'h0 : _GEN_11342; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11344 = 10'hd3 == _T_244[9:0] ? 4'h0 : _GEN_11343; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11345 = 10'hd4 == _T_244[9:0] ? 4'h0 : _GEN_11344; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11346 = 10'hd5 == _T_244[9:0] ? 4'h0 : _GEN_11345; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11347 = 10'hd6 == _T_244[9:0] ? 4'h1 : _GEN_11346; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11348 = 10'hd7 == _T_244[9:0] ? 4'h3 : _GEN_11347; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11349 = 10'hd8 == _T_244[9:0] ? 4'h0 : _GEN_11348; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11350 = 10'hd9 == _T_244[9:0] ? 4'h3 : _GEN_11349; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11351 = 10'hda == _T_244[9:0] ? 4'h3 : _GEN_11350; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11352 = 10'hdb == _T_244[9:0] ? 4'h3 : _GEN_11351; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11353 = 10'hdc == _T_244[9:0] ? 4'h3 : _GEN_11352; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11354 = 10'hdd == _T_244[9:0] ? 4'ha : _GEN_11353; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11355 = 10'hde == _T_244[9:0] ? 4'h7 : _GEN_11354; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11356 = 10'hdf == _T_244[9:0] ? 4'h0 : _GEN_11355; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11357 = 10'he0 == _T_244[9:0] ? 4'h3 : _GEN_11356; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11358 = 10'he1 == _T_244[9:0] ? 4'h3 : _GEN_11357; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11359 = 10'he2 == _T_244[9:0] ? 4'ha : _GEN_11358; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11360 = 10'he3 == _T_244[9:0] ? 4'h3 : _GEN_11359; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11361 = 10'he4 == _T_244[9:0] ? 4'h3 : _GEN_11360; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11362 = 10'he5 == _T_244[9:0] ? 4'h3 : _GEN_11361; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11363 = 10'he6 == _T_244[9:0] ? 4'h3 : _GEN_11362; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11364 = 10'he7 == _T_244[9:0] ? 4'h1 : _GEN_11363; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11365 = 10'he8 == _T_244[9:0] ? 4'h1 : _GEN_11364; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11366 = 10'he9 == _T_244[9:0] ? 4'h1 : _GEN_11365; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11367 = 10'hea == _T_244[9:0] ? 4'h0 : _GEN_11366; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11368 = 10'heb == _T_244[9:0] ? 4'h0 : _GEN_11367; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11369 = 10'hec == _T_244[9:0] ? 4'h0 : _GEN_11368; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11370 = 10'hed == _T_244[9:0] ? 4'h0 : _GEN_11369; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11371 = 10'hee == _T_244[9:0] ? 4'h0 : _GEN_11370; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11372 = 10'hef == _T_244[9:0] ? 4'h0 : _GEN_11371; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11373 = 10'hf0 == _T_244[9:0] ? 4'h0 : _GEN_11372; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11374 = 10'hf1 == _T_244[9:0] ? 4'h0 : _GEN_11373; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11375 = 10'hf2 == _T_244[9:0] ? 4'h0 : _GEN_11374; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11376 = 10'hf3 == _T_244[9:0] ? 4'h0 : _GEN_11375; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11377 = 10'hf4 == _T_244[9:0] ? 4'h0 : _GEN_11376; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11378 = 10'hf5 == _T_244[9:0] ? 4'h1 : _GEN_11377; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11379 = 10'hf6 == _T_244[9:0] ? 4'h0 : _GEN_11378; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11380 = 10'hf7 == _T_244[9:0] ? 4'h0 : _GEN_11379; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11381 = 10'hf8 == _T_244[9:0] ? 4'h1 : _GEN_11380; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11382 = 10'hf9 == _T_244[9:0] ? 4'h0 : _GEN_11381; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11383 = 10'hfa == _T_244[9:0] ? 4'h3 : _GEN_11382; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11384 = 10'hfb == _T_244[9:0] ? 4'h3 : _GEN_11383; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11385 = 10'hfc == _T_244[9:0] ? 4'h3 : _GEN_11384; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11386 = 10'hfd == _T_244[9:0] ? 4'ha : _GEN_11385; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11387 = 10'hfe == _T_244[9:0] ? 4'h3 : _GEN_11386; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11388 = 10'hff == _T_244[9:0] ? 4'h0 : _GEN_11387; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11389 = 10'h100 == _T_244[9:0] ? 4'h3 : _GEN_11388; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11390 = 10'h101 == _T_244[9:0] ? 4'h0 : _GEN_11389; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11391 = 10'h102 == _T_244[9:0] ? 4'ha : _GEN_11390; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11392 = 10'h103 == _T_244[9:0] ? 4'h3 : _GEN_11391; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11393 = 10'h104 == _T_244[9:0] ? 4'h3 : _GEN_11392; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11394 = 10'h105 == _T_244[9:0] ? 4'h3 : _GEN_11393; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11395 = 10'h106 == _T_244[9:0] ? 4'h3 : _GEN_11394; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11396 = 10'h107 == _T_244[9:0] ? 4'h3 : _GEN_11395; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11397 = 10'h108 == _T_244[9:0] ? 4'h1 : _GEN_11396; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11398 = 10'h109 == _T_244[9:0] ? 4'h0 : _GEN_11397; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11399 = 10'h10a == _T_244[9:0] ? 4'h0 : _GEN_11398; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11400 = 10'h10b == _T_244[9:0] ? 4'h0 : _GEN_11399; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11401 = 10'h10c == _T_244[9:0] ? 4'h0 : _GEN_11400; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11402 = 10'h10d == _T_244[9:0] ? 4'h0 : _GEN_11401; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11403 = 10'h10e == _T_244[9:0] ? 4'h0 : _GEN_11402; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11404 = 10'h10f == _T_244[9:0] ? 4'h0 : _GEN_11403; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11405 = 10'h110 == _T_244[9:0] ? 4'h0 : _GEN_11404; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11406 = 10'h111 == _T_244[9:0] ? 4'h0 : _GEN_11405; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11407 = 10'h112 == _T_244[9:0] ? 4'h0 : _GEN_11406; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11408 = 10'h113 == _T_244[9:0] ? 4'h0 : _GEN_11407; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11409 = 10'h114 == _T_244[9:0] ? 4'h0 : _GEN_11408; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11410 = 10'h115 == _T_244[9:0] ? 4'h0 : _GEN_11409; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11411 = 10'h116 == _T_244[9:0] ? 4'h1 : _GEN_11410; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11412 = 10'h117 == _T_244[9:0] ? 4'h3 : _GEN_11411; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11413 = 10'h118 == _T_244[9:0] ? 4'h3 : _GEN_11412; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11414 = 10'h119 == _T_244[9:0] ? 4'h3 : _GEN_11413; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11415 = 10'h11a == _T_244[9:0] ? 4'h0 : _GEN_11414; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11416 = 10'h11b == _T_244[9:0] ? 4'h3 : _GEN_11415; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11417 = 10'h11c == _T_244[9:0] ? 4'h3 : _GEN_11416; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11418 = 10'h11d == _T_244[9:0] ? 4'h7 : _GEN_11417; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11419 = 10'h11e == _T_244[9:0] ? 4'ha : _GEN_11418; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11420 = 10'h11f == _T_244[9:0] ? 4'h0 : _GEN_11419; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11421 = 10'h120 == _T_244[9:0] ? 4'h3 : _GEN_11420; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11422 = 10'h121 == _T_244[9:0] ? 4'h3 : _GEN_11421; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11423 = 10'h122 == _T_244[9:0] ? 4'ha : _GEN_11422; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11424 = 10'h123 == _T_244[9:0] ? 4'h3 : _GEN_11423; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11425 = 10'h124 == _T_244[9:0] ? 4'h3 : _GEN_11424; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11426 = 10'h125 == _T_244[9:0] ? 4'h3 : _GEN_11425; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11427 = 10'h126 == _T_244[9:0] ? 4'h3 : _GEN_11426; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11428 = 10'h127 == _T_244[9:0] ? 4'h1 : _GEN_11427; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11429 = 10'h128 == _T_244[9:0] ? 4'h0 : _GEN_11428; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11430 = 10'h129 == _T_244[9:0] ? 4'h3 : _GEN_11429; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11431 = 10'h12a == _T_244[9:0] ? 4'h3 : _GEN_11430; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11432 = 10'h12b == _T_244[9:0] ? 4'h0 : _GEN_11431; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11433 = 10'h12c == _T_244[9:0] ? 4'h0 : _GEN_11432; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11434 = 10'h12d == _T_244[9:0] ? 4'h0 : _GEN_11433; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11435 = 10'h12e == _T_244[9:0] ? 4'h0 : _GEN_11434; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11436 = 10'h12f == _T_244[9:0] ? 4'h0 : _GEN_11435; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11437 = 10'h130 == _T_244[9:0] ? 4'h0 : _GEN_11436; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11438 = 10'h131 == _T_244[9:0] ? 4'h0 : _GEN_11437; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11439 = 10'h132 == _T_244[9:0] ? 4'h0 : _GEN_11438; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11440 = 10'h133 == _T_244[9:0] ? 4'h0 : _GEN_11439; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11441 = 10'h134 == _T_244[9:0] ? 4'h3 : _GEN_11440; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11442 = 10'h135 == _T_244[9:0] ? 4'h3 : _GEN_11441; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11443 = 10'h136 == _T_244[9:0] ? 4'h0 : _GEN_11442; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11444 = 10'h137 == _T_244[9:0] ? 4'h1 : _GEN_11443; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11445 = 10'h138 == _T_244[9:0] ? 4'h3 : _GEN_11444; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11446 = 10'h139 == _T_244[9:0] ? 4'h3 : _GEN_11445; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11447 = 10'h13a == _T_244[9:0] ? 4'h3 : _GEN_11446; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11448 = 10'h13b == _T_244[9:0] ? 4'h3 : _GEN_11447; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11449 = 10'h13c == _T_244[9:0] ? 4'h3 : _GEN_11448; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11450 = 10'h13d == _T_244[9:0] ? 4'h3 : _GEN_11449; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11451 = 10'h13e == _T_244[9:0] ? 4'ha : _GEN_11450; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11452 = 10'h13f == _T_244[9:0] ? 4'h0 : _GEN_11451; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11453 = 10'h140 == _T_244[9:0] ? 4'h5 : _GEN_11452; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11454 = 10'h141 == _T_244[9:0] ? 4'h3 : _GEN_11453; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11455 = 10'h142 == _T_244[9:0] ? 4'h7 : _GEN_11454; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11456 = 10'h143 == _T_244[9:0] ? 4'ha : _GEN_11455; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11457 = 10'h144 == _T_244[9:0] ? 4'h3 : _GEN_11456; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11458 = 10'h145 == _T_244[9:0] ? 4'h3 : _GEN_11457; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11459 = 10'h146 == _T_244[9:0] ? 4'h1 : _GEN_11458; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11460 = 10'h147 == _T_244[9:0] ? 4'h0 : _GEN_11459; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11461 = 10'h148 == _T_244[9:0] ? 4'h3 : _GEN_11460; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11462 = 10'h149 == _T_244[9:0] ? 4'h3 : _GEN_11461; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11463 = 10'h14a == _T_244[9:0] ? 4'h3 : _GEN_11462; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11464 = 10'h14b == _T_244[9:0] ? 4'h3 : _GEN_11463; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11465 = 10'h14c == _T_244[9:0] ? 4'h3 : _GEN_11464; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11466 = 10'h14d == _T_244[9:0] ? 4'h3 : _GEN_11465; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11467 = 10'h14e == _T_244[9:0] ? 4'h3 : _GEN_11466; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11468 = 10'h14f == _T_244[9:0] ? 4'h3 : _GEN_11467; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11469 = 10'h150 == _T_244[9:0] ? 4'h3 : _GEN_11468; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11470 = 10'h151 == _T_244[9:0] ? 4'h3 : _GEN_11469; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11471 = 10'h152 == _T_244[9:0] ? 4'h3 : _GEN_11470; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11472 = 10'h153 == _T_244[9:0] ? 4'h3 : _GEN_11471; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11473 = 10'h154 == _T_244[9:0] ? 4'h3 : _GEN_11472; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11474 = 10'h155 == _T_244[9:0] ? 4'h3 : _GEN_11473; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11475 = 10'h156 == _T_244[9:0] ? 4'h3 : _GEN_11474; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11476 = 10'h157 == _T_244[9:0] ? 4'h0 : _GEN_11475; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11477 = 10'h158 == _T_244[9:0] ? 4'h3 : _GEN_11476; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11478 = 10'h159 == _T_244[9:0] ? 4'h3 : _GEN_11477; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11479 = 10'h15a == _T_244[9:0] ? 4'h3 : _GEN_11478; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11480 = 10'h15b == _T_244[9:0] ? 4'h3 : _GEN_11479; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11481 = 10'h15c == _T_244[9:0] ? 4'h3 : _GEN_11480; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11482 = 10'h15d == _T_244[9:0] ? 4'ha : _GEN_11481; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11483 = 10'h15e == _T_244[9:0] ? 4'h7 : _GEN_11482; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11484 = 10'h15f == _T_244[9:0] ? 4'h0 : _GEN_11483; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11485 = 10'h160 == _T_244[9:0] ? 4'h3 : _GEN_11484; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11486 = 10'h161 == _T_244[9:0] ? 4'h3 : _GEN_11485; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11487 = 10'h162 == _T_244[9:0] ? 4'h3 : _GEN_11486; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11488 = 10'h163 == _T_244[9:0] ? 4'h7 : _GEN_11487; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11489 = 10'h164 == _T_244[9:0] ? 4'ha : _GEN_11488; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11490 = 10'h165 == _T_244[9:0] ? 4'h1 : _GEN_11489; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11491 = 10'h166 == _T_244[9:0] ? 4'h0 : _GEN_11490; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11492 = 10'h167 == _T_244[9:0] ? 4'h0 : _GEN_11491; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11493 = 10'h168 == _T_244[9:0] ? 4'hc : _GEN_11492; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11494 = 10'h169 == _T_244[9:0] ? 4'h9 : _GEN_11493; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11495 = 10'h16a == _T_244[9:0] ? 4'hc : _GEN_11494; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11496 = 10'h16b == _T_244[9:0] ? 4'hc : _GEN_11495; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11497 = 10'h16c == _T_244[9:0] ? 4'h3 : _GEN_11496; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11498 = 10'h16d == _T_244[9:0] ? 4'h3 : _GEN_11497; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11499 = 10'h16e == _T_244[9:0] ? 4'h3 : _GEN_11498; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11500 = 10'h16f == _T_244[9:0] ? 4'h3 : _GEN_11499; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11501 = 10'h170 == _T_244[9:0] ? 4'h5 : _GEN_11500; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11502 = 10'h171 == _T_244[9:0] ? 4'h3 : _GEN_11501; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11503 = 10'h172 == _T_244[9:0] ? 4'h3 : _GEN_11502; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11504 = 10'h173 == _T_244[9:0] ? 4'h3 : _GEN_11503; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11505 = 10'h174 == _T_244[9:0] ? 4'h3 : _GEN_11504; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11506 = 10'h175 == _T_244[9:0] ? 4'h3 : _GEN_11505; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11507 = 10'h176 == _T_244[9:0] ? 4'h0 : _GEN_11506; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11508 = 10'h177 == _T_244[9:0] ? 4'h0 : _GEN_11507; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11509 = 10'h178 == _T_244[9:0] ? 4'h1 : _GEN_11508; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11510 = 10'h179 == _T_244[9:0] ? 4'h3 : _GEN_11509; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11511 = 10'h17a == _T_244[9:0] ? 4'h5 : _GEN_11510; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11512 = 10'h17b == _T_244[9:0] ? 4'h3 : _GEN_11511; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11513 = 10'h17c == _T_244[9:0] ? 4'ha : _GEN_11512; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11514 = 10'h17d == _T_244[9:0] ? 4'h7 : _GEN_11513; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11515 = 10'h17e == _T_244[9:0] ? 4'h3 : _GEN_11514; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11516 = 10'h17f == _T_244[9:0] ? 4'h0 : _GEN_11515; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11517 = 10'h180 == _T_244[9:0] ? 4'hc : _GEN_11516; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11518 = 10'h181 == _T_244[9:0] ? 4'hc : _GEN_11517; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11519 = 10'h182 == _T_244[9:0] ? 4'hc : _GEN_11518; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11520 = 10'h183 == _T_244[9:0] ? 4'hc : _GEN_11519; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11521 = 10'h184 == _T_244[9:0] ? 4'ha : _GEN_11520; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11522 = 10'h185 == _T_244[9:0] ? 4'h1 : _GEN_11521; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11523 = 10'h186 == _T_244[9:0] ? 4'hc : _GEN_11522; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11524 = 10'h187 == _T_244[9:0] ? 4'h0 : _GEN_11523; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11525 = 10'h188 == _T_244[9:0] ? 4'hc : _GEN_11524; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11526 = 10'h189 == _T_244[9:0] ? 4'hc : _GEN_11525; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11527 = 10'h18a == _T_244[9:0] ? 4'hc : _GEN_11526; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11528 = 10'h18b == _T_244[9:0] ? 4'hc : _GEN_11527; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11529 = 10'h18c == _T_244[9:0] ? 4'hc : _GEN_11528; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11530 = 10'h18d == _T_244[9:0] ? 4'hc : _GEN_11529; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11531 = 10'h18e == _T_244[9:0] ? 4'hc : _GEN_11530; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11532 = 10'h18f == _T_244[9:0] ? 4'hc : _GEN_11531; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11533 = 10'h190 == _T_244[9:0] ? 4'hc : _GEN_11532; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11534 = 10'h191 == _T_244[9:0] ? 4'hc : _GEN_11533; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11535 = 10'h192 == _T_244[9:0] ? 4'h9 : _GEN_11534; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11536 = 10'h193 == _T_244[9:0] ? 4'hc : _GEN_11535; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11537 = 10'h194 == _T_244[9:0] ? 4'hc : _GEN_11536; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11538 = 10'h195 == _T_244[9:0] ? 4'hc : _GEN_11537; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11539 = 10'h196 == _T_244[9:0] ? 4'h0 : _GEN_11538; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11540 = 10'h197 == _T_244[9:0] ? 4'h3 : _GEN_11539; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11541 = 10'h198 == _T_244[9:0] ? 4'h1 : _GEN_11540; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11542 = 10'h199 == _T_244[9:0] ? 4'h3 : _GEN_11541; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11543 = 10'h19a == _T_244[9:0] ? 4'h3 : _GEN_11542; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11544 = 10'h19b == _T_244[9:0] ? 4'h3 : _GEN_11543; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11545 = 10'h19c == _T_244[9:0] ? 4'ha : _GEN_11544; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11546 = 10'h19d == _T_244[9:0] ? 4'h3 : _GEN_11545; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11547 = 10'h19e == _T_244[9:0] ? 4'h3 : _GEN_11546; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11548 = 10'h19f == _T_244[9:0] ? 4'h0 : _GEN_11547; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11549 = 10'h1a0 == _T_244[9:0] ? 4'hc : _GEN_11548; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11550 = 10'h1a1 == _T_244[9:0] ? 4'hc : _GEN_11549; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11551 = 10'h1a2 == _T_244[9:0] ? 4'h9 : _GEN_11550; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11552 = 10'h1a3 == _T_244[9:0] ? 4'hc : _GEN_11551; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11553 = 10'h1a4 == _T_244[9:0] ? 4'ha : _GEN_11552; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11554 = 10'h1a5 == _T_244[9:0] ? 4'h0 : _GEN_11553; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11555 = 10'h1a6 == _T_244[9:0] ? 4'hc : _GEN_11554; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11556 = 10'h1a7 == _T_244[9:0] ? 4'h0 : _GEN_11555; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11557 = 10'h1a8 == _T_244[9:0] ? 4'hc : _GEN_11556; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11558 = 10'h1a9 == _T_244[9:0] ? 4'hc : _GEN_11557; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11559 = 10'h1aa == _T_244[9:0] ? 4'hc : _GEN_11558; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11560 = 10'h1ab == _T_244[9:0] ? 4'h9 : _GEN_11559; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11561 = 10'h1ac == _T_244[9:0] ? 4'hc : _GEN_11560; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11562 = 10'h1ad == _T_244[9:0] ? 4'hc : _GEN_11561; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11563 = 10'h1ae == _T_244[9:0] ? 4'hc : _GEN_11562; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11564 = 10'h1af == _T_244[9:0] ? 4'hc : _GEN_11563; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11565 = 10'h1b0 == _T_244[9:0] ? 4'hc : _GEN_11564; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11566 = 10'h1b1 == _T_244[9:0] ? 4'hc : _GEN_11565; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11567 = 10'h1b2 == _T_244[9:0] ? 4'hc : _GEN_11566; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11568 = 10'h1b3 == _T_244[9:0] ? 4'hc : _GEN_11567; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11569 = 10'h1b4 == _T_244[9:0] ? 4'hc : _GEN_11568; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11570 = 10'h1b5 == _T_244[9:0] ? 4'hc : _GEN_11569; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11571 = 10'h1b6 == _T_244[9:0] ? 4'h0 : _GEN_11570; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11572 = 10'h1b7 == _T_244[9:0] ? 4'hc : _GEN_11571; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11573 = 10'h1b8 == _T_244[9:0] ? 4'h0 : _GEN_11572; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11574 = 10'h1b9 == _T_244[9:0] ? 4'hc : _GEN_11573; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11575 = 10'h1ba == _T_244[9:0] ? 4'hc : _GEN_11574; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11576 = 10'h1bb == _T_244[9:0] ? 4'hc : _GEN_11575; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11577 = 10'h1bc == _T_244[9:0] ? 4'h7 : _GEN_11576; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11578 = 10'h1bd == _T_244[9:0] ? 4'ha : _GEN_11577; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11579 = 10'h1be == _T_244[9:0] ? 4'hc : _GEN_11578; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11580 = 10'h1bf == _T_244[9:0] ? 4'h0 : _GEN_11579; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11581 = 10'h1c0 == _T_244[9:0] ? 4'hc : _GEN_11580; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11582 = 10'h1c1 == _T_244[9:0] ? 4'hc : _GEN_11581; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11583 = 10'h1c2 == _T_244[9:0] ? 4'hc : _GEN_11582; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11584 = 10'h1c3 == _T_244[9:0] ? 4'h7 : _GEN_11583; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11585 = 10'h1c4 == _T_244[9:0] ? 4'h7 : _GEN_11584; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11586 = 10'h1c5 == _T_244[9:0] ? 4'hc : _GEN_11585; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11587 = 10'h1c6 == _T_244[9:0] ? 4'hc : _GEN_11586; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11588 = 10'h1c7 == _T_244[9:0] ? 4'hc : _GEN_11587; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11589 = 10'h1c8 == _T_244[9:0] ? 4'hc : _GEN_11588; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11590 = 10'h1c9 == _T_244[9:0] ? 4'hc : _GEN_11589; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11591 = 10'h1ca == _T_244[9:0] ? 4'hc : _GEN_11590; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11592 = 10'h1cb == _T_244[9:0] ? 4'hc : _GEN_11591; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11593 = 10'h1cc == _T_244[9:0] ? 4'hc : _GEN_11592; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11594 = 10'h1cd == _T_244[9:0] ? 4'hc : _GEN_11593; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11595 = 10'h1ce == _T_244[9:0] ? 4'hc : _GEN_11594; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11596 = 10'h1cf == _T_244[9:0] ? 4'hc : _GEN_11595; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11597 = 10'h1d0 == _T_244[9:0] ? 4'hc : _GEN_11596; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11598 = 10'h1d1 == _T_244[9:0] ? 4'hc : _GEN_11597; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11599 = 10'h1d2 == _T_244[9:0] ? 4'hc : _GEN_11598; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11600 = 10'h1d3 == _T_244[9:0] ? 4'hc : _GEN_11599; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11601 = 10'h1d4 == _T_244[9:0] ? 4'hc : _GEN_11600; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11602 = 10'h1d5 == _T_244[9:0] ? 4'hc : _GEN_11601; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11603 = 10'h1d6 == _T_244[9:0] ? 4'hc : _GEN_11602; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11604 = 10'h1d7 == _T_244[9:0] ? 4'hc : _GEN_11603; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11605 = 10'h1d8 == _T_244[9:0] ? 4'hc : _GEN_11604; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11606 = 10'h1d9 == _T_244[9:0] ? 4'hc : _GEN_11605; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11607 = 10'h1da == _T_244[9:0] ? 4'hc : _GEN_11606; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11608 = 10'h1db == _T_244[9:0] ? 4'hc : _GEN_11607; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11609 = 10'h1dc == _T_244[9:0] ? 4'hc : _GEN_11608; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11610 = 10'h1dd == _T_244[9:0] ? 4'ha : _GEN_11609; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11611 = 10'h1de == _T_244[9:0] ? 4'hc : _GEN_11610; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11612 = 10'h1df == _T_244[9:0] ? 4'h0 : _GEN_11611; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11613 = 10'h1e0 == _T_244[9:0] ? 4'h9 : _GEN_11612; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11614 = 10'h1e1 == _T_244[9:0] ? 4'hc : _GEN_11613; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11615 = 10'h1e2 == _T_244[9:0] ? 4'h7 : _GEN_11614; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11616 = 10'h1e3 == _T_244[9:0] ? 4'h7 : _GEN_11615; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11617 = 10'h1e4 == _T_244[9:0] ? 4'hc : _GEN_11616; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11618 = 10'h1e5 == _T_244[9:0] ? 4'hc : _GEN_11617; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11619 = 10'h1e6 == _T_244[9:0] ? 4'hc : _GEN_11618; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11620 = 10'h1e7 == _T_244[9:0] ? 4'hc : _GEN_11619; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11621 = 10'h1e8 == _T_244[9:0] ? 4'hc : _GEN_11620; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11622 = 10'h1e9 == _T_244[9:0] ? 4'hc : _GEN_11621; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11623 = 10'h1ea == _T_244[9:0] ? 4'hc : _GEN_11622; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11624 = 10'h1eb == _T_244[9:0] ? 4'hc : _GEN_11623; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11625 = 10'h1ec == _T_244[9:0] ? 4'hc : _GEN_11624; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11626 = 10'h1ed == _T_244[9:0] ? 4'hc : _GEN_11625; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11627 = 10'h1ee == _T_244[9:0] ? 4'hc : _GEN_11626; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11628 = 10'h1ef == _T_244[9:0] ? 4'hc : _GEN_11627; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11629 = 10'h1f0 == _T_244[9:0] ? 4'hc : _GEN_11628; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11630 = 10'h1f1 == _T_244[9:0] ? 4'hc : _GEN_11629; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11631 = 10'h1f2 == _T_244[9:0] ? 4'hc : _GEN_11630; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11632 = 10'h1f3 == _T_244[9:0] ? 4'hc : _GEN_11631; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11633 = 10'h1f4 == _T_244[9:0] ? 4'hc : _GEN_11632; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11634 = 10'h1f5 == _T_244[9:0] ? 4'hc : _GEN_11633; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11635 = 10'h1f6 == _T_244[9:0] ? 4'hc : _GEN_11634; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11636 = 10'h1f7 == _T_244[9:0] ? 4'hc : _GEN_11635; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11637 = 10'h1f8 == _T_244[9:0] ? 4'hc : _GEN_11636; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11638 = 10'h1f9 == _T_244[9:0] ? 4'hc : _GEN_11637; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11639 = 10'h1fa == _T_244[9:0] ? 4'h9 : _GEN_11638; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11640 = 10'h1fb == _T_244[9:0] ? 4'hc : _GEN_11639; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11641 = 10'h1fc == _T_244[9:0] ? 4'hc : _GEN_11640; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11642 = 10'h1fd == _T_244[9:0] ? 4'h7 : _GEN_11641; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11643 = 10'h1fe == _T_244[9:0] ? 4'hc : _GEN_11642; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11644 = 10'h1ff == _T_244[9:0] ? 4'h0 : _GEN_11643; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11645 = 10'h200 == _T_244[9:0] ? 4'hc : _GEN_11644; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11646 = 10'h201 == _T_244[9:0] ? 4'hc : _GEN_11645; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11647 = 10'h202 == _T_244[9:0] ? 4'ha : _GEN_11646; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11648 = 10'h203 == _T_244[9:0] ? 4'hc : _GEN_11647; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11649 = 10'h204 == _T_244[9:0] ? 4'hc : _GEN_11648; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11650 = 10'h205 == _T_244[9:0] ? 4'hc : _GEN_11649; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11651 = 10'h206 == _T_244[9:0] ? 4'hc : _GEN_11650; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11652 = 10'h207 == _T_244[9:0] ? 4'hc : _GEN_11651; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11653 = 10'h208 == _T_244[9:0] ? 4'hc : _GEN_11652; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11654 = 10'h209 == _T_244[9:0] ? 4'hc : _GEN_11653; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11655 = 10'h20a == _T_244[9:0] ? 4'hc : _GEN_11654; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11656 = 10'h20b == _T_244[9:0] ? 4'hc : _GEN_11655; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11657 = 10'h20c == _T_244[9:0] ? 4'hc : _GEN_11656; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11658 = 10'h20d == _T_244[9:0] ? 4'hc : _GEN_11657; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11659 = 10'h20e == _T_244[9:0] ? 4'hc : _GEN_11658; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11660 = 10'h20f == _T_244[9:0] ? 4'hc : _GEN_11659; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11661 = 10'h210 == _T_244[9:0] ? 4'hc : _GEN_11660; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11662 = 10'h211 == _T_244[9:0] ? 4'hc : _GEN_11661; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11663 = 10'h212 == _T_244[9:0] ? 4'hc : _GEN_11662; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11664 = 10'h213 == _T_244[9:0] ? 4'hc : _GEN_11663; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11665 = 10'h214 == _T_244[9:0] ? 4'hc : _GEN_11664; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11666 = 10'h215 == _T_244[9:0] ? 4'hc : _GEN_11665; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11667 = 10'h216 == _T_244[9:0] ? 4'hc : _GEN_11666; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11668 = 10'h217 == _T_244[9:0] ? 4'hc : _GEN_11667; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11669 = 10'h218 == _T_244[9:0] ? 4'hc : _GEN_11668; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11670 = 10'h219 == _T_244[9:0] ? 4'hc : _GEN_11669; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11671 = 10'h21a == _T_244[9:0] ? 4'hc : _GEN_11670; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11672 = 10'h21b == _T_244[9:0] ? 4'hc : _GEN_11671; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11673 = 10'h21c == _T_244[9:0] ? 4'ha : _GEN_11672; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11674 = 10'h21d == _T_244[9:0] ? 4'h7 : _GEN_11673; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11675 = 10'h21e == _T_244[9:0] ? 4'hc : _GEN_11674; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11676 = 10'h21f == _T_244[9:0] ? 4'h0 : _GEN_11675; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11677 = 10'h220 == _T_244[9:0] ? 4'h0 : _GEN_11676; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11678 = 10'h221 == _T_244[9:0] ? 4'h0 : _GEN_11677; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11679 = 10'h222 == _T_244[9:0] ? 4'h0 : _GEN_11678; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11680 = 10'h223 == _T_244[9:0] ? 4'h0 : _GEN_11679; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11681 = 10'h224 == _T_244[9:0] ? 4'h0 : _GEN_11680; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11682 = 10'h225 == _T_244[9:0] ? 4'h0 : _GEN_11681; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11683 = 10'h226 == _T_244[9:0] ? 4'h0 : _GEN_11682; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11684 = 10'h227 == _T_244[9:0] ? 4'h0 : _GEN_11683; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11685 = 10'h228 == _T_244[9:0] ? 4'h0 : _GEN_11684; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11686 = 10'h229 == _T_244[9:0] ? 4'h0 : _GEN_11685; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11687 = 10'h22a == _T_244[9:0] ? 4'h0 : _GEN_11686; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11688 = 10'h22b == _T_244[9:0] ? 4'h0 : _GEN_11687; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11689 = 10'h22c == _T_244[9:0] ? 4'h0 : _GEN_11688; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11690 = 10'h22d == _T_244[9:0] ? 4'h0 : _GEN_11689; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11691 = 10'h22e == _T_244[9:0] ? 4'h0 : _GEN_11690; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11692 = 10'h22f == _T_244[9:0] ? 4'h0 : _GEN_11691; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11693 = 10'h230 == _T_244[9:0] ? 4'h0 : _GEN_11692; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11694 = 10'h231 == _T_244[9:0] ? 4'h0 : _GEN_11693; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11695 = 10'h232 == _T_244[9:0] ? 4'h0 : _GEN_11694; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11696 = 10'h233 == _T_244[9:0] ? 4'h0 : _GEN_11695; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11697 = 10'h234 == _T_244[9:0] ? 4'h0 : _GEN_11696; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11698 = 10'h235 == _T_244[9:0] ? 4'h0 : _GEN_11697; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11699 = 10'h236 == _T_244[9:0] ? 4'h0 : _GEN_11698; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11700 = 10'h237 == _T_244[9:0] ? 4'h0 : _GEN_11699; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11701 = 10'h238 == _T_244[9:0] ? 4'h0 : _GEN_11700; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11702 = 10'h239 == _T_244[9:0] ? 4'h0 : _GEN_11701; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11703 = 10'h23a == _T_244[9:0] ? 4'h0 : _GEN_11702; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11704 = 10'h23b == _T_244[9:0] ? 4'h0 : _GEN_11703; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11705 = 10'h23c == _T_244[9:0] ? 4'h0 : _GEN_11704; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11706 = 10'h23d == _T_244[9:0] ? 4'h0 : _GEN_11705; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11707 = 10'h23e == _T_244[9:0] ? 4'h0 : _GEN_11706; // @[Filter.scala 191:102]
  wire [3:0] _GEN_11708 = 10'h23f == _T_244[9:0] ? 4'h0 : _GEN_11707; // @[Filter.scala 191:102]
  wire [6:0] _GEN_28336 = {{3'd0}, _GEN_11708}; // @[Filter.scala 191:102]
  wire [10:0] _T_251 = _GEN_28336 * 7'h46; // @[Filter.scala 191:102]
  wire [10:0] _GEN_28337 = {{2'd0}, _T_246}; // @[Filter.scala 191:69]
  wire [10:0] _T_253 = _GEN_28337 + _T_251; // @[Filter.scala 191:69]
  wire [3:0] _GEN_11740 = 10'h1f == _T_244[9:0] ? 4'h0 : 4'h3; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11741 = 10'h20 == _T_244[9:0] ? 4'h3 : _GEN_11740; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11742 = 10'h21 == _T_244[9:0] ? 4'h3 : _GEN_11741; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11743 = 10'h22 == _T_244[9:0] ? 4'h3 : _GEN_11742; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11744 = 10'h23 == _T_244[9:0] ? 4'h3 : _GEN_11743; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11745 = 10'h24 == _T_244[9:0] ? 4'h3 : _GEN_11744; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11746 = 10'h25 == _T_244[9:0] ? 4'h3 : _GEN_11745; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11747 = 10'h26 == _T_244[9:0] ? 4'h3 : _GEN_11746; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11748 = 10'h27 == _T_244[9:0] ? 4'h9 : _GEN_11747; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11749 = 10'h28 == _T_244[9:0] ? 4'h9 : _GEN_11748; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11750 = 10'h29 == _T_244[9:0] ? 4'h3 : _GEN_11749; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11751 = 10'h2a == _T_244[9:0] ? 4'h3 : _GEN_11750; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11752 = 10'h2b == _T_244[9:0] ? 4'h3 : _GEN_11751; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11753 = 10'h2c == _T_244[9:0] ? 4'h3 : _GEN_11752; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11754 = 10'h2d == _T_244[9:0] ? 4'h3 : _GEN_11753; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11755 = 10'h2e == _T_244[9:0] ? 4'h3 : _GEN_11754; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11756 = 10'h2f == _T_244[9:0] ? 4'h3 : _GEN_11755; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11757 = 10'h30 == _T_244[9:0] ? 4'h3 : _GEN_11756; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11758 = 10'h31 == _T_244[9:0] ? 4'h3 : _GEN_11757; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11759 = 10'h32 == _T_244[9:0] ? 4'h3 : _GEN_11758; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11760 = 10'h33 == _T_244[9:0] ? 4'h3 : _GEN_11759; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11761 = 10'h34 == _T_244[9:0] ? 4'h3 : _GEN_11760; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11762 = 10'h35 == _T_244[9:0] ? 4'h3 : _GEN_11761; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11763 = 10'h36 == _T_244[9:0] ? 4'h3 : _GEN_11762; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11764 = 10'h37 == _T_244[9:0] ? 4'h9 : _GEN_11763; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11765 = 10'h38 == _T_244[9:0] ? 4'h9 : _GEN_11764; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11766 = 10'h39 == _T_244[9:0] ? 4'h3 : _GEN_11765; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11767 = 10'h3a == _T_244[9:0] ? 4'h3 : _GEN_11766; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11768 = 10'h3b == _T_244[9:0] ? 4'h3 : _GEN_11767; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11769 = 10'h3c == _T_244[9:0] ? 4'h3 : _GEN_11768; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11770 = 10'h3d == _T_244[9:0] ? 4'h3 : _GEN_11769; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11771 = 10'h3e == _T_244[9:0] ? 4'h3 : _GEN_11770; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11772 = 10'h3f == _T_244[9:0] ? 4'h0 : _GEN_11771; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11773 = 10'h40 == _T_244[9:0] ? 4'h3 : _GEN_11772; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11774 = 10'h41 == _T_244[9:0] ? 4'h3 : _GEN_11773; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11775 = 10'h42 == _T_244[9:0] ? 4'h3 : _GEN_11774; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11776 = 10'h43 == _T_244[9:0] ? 4'h2 : _GEN_11775; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11777 = 10'h44 == _T_244[9:0] ? 4'h3 : _GEN_11776; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11778 = 10'h45 == _T_244[9:0] ? 4'hf : _GEN_11777; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11779 = 10'h46 == _T_244[9:0] ? 4'hf : _GEN_11778; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11780 = 10'h47 == _T_244[9:0] ? 4'hf : _GEN_11779; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11781 = 10'h48 == _T_244[9:0] ? 4'hf : _GEN_11780; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11782 = 10'h49 == _T_244[9:0] ? 4'h3 : _GEN_11781; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11783 = 10'h4a == _T_244[9:0] ? 4'h3 : _GEN_11782; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11784 = 10'h4b == _T_244[9:0] ? 4'h3 : _GEN_11783; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11785 = 10'h4c == _T_244[9:0] ? 4'h3 : _GEN_11784; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11786 = 10'h4d == _T_244[9:0] ? 4'h3 : _GEN_11785; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11787 = 10'h4e == _T_244[9:0] ? 4'h3 : _GEN_11786; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11788 = 10'h4f == _T_244[9:0] ? 4'h3 : _GEN_11787; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11789 = 10'h50 == _T_244[9:0] ? 4'h3 : _GEN_11788; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11790 = 10'h51 == _T_244[9:0] ? 4'h3 : _GEN_11789; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11791 = 10'h52 == _T_244[9:0] ? 4'h3 : _GEN_11790; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11792 = 10'h53 == _T_244[9:0] ? 4'h3 : _GEN_11791; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11793 = 10'h54 == _T_244[9:0] ? 4'h9 : _GEN_11792; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11794 = 10'h55 == _T_244[9:0] ? 4'h9 : _GEN_11793; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11795 = 10'h56 == _T_244[9:0] ? 4'h9 : _GEN_11794; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11796 = 10'h57 == _T_244[9:0] ? 4'hf : _GEN_11795; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11797 = 10'h58 == _T_244[9:0] ? 4'h3 : _GEN_11796; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11798 = 10'h59 == _T_244[9:0] ? 4'hf : _GEN_11797; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11799 = 10'h5a == _T_244[9:0] ? 4'h3 : _GEN_11798; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11800 = 10'h5b == _T_244[9:0] ? 4'h3 : _GEN_11799; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11801 = 10'h5c == _T_244[9:0] ? 4'h3 : _GEN_11800; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11802 = 10'h5d == _T_244[9:0] ? 4'h3 : _GEN_11801; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11803 = 10'h5e == _T_244[9:0] ? 4'h3 : _GEN_11802; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11804 = 10'h5f == _T_244[9:0] ? 4'h0 : _GEN_11803; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11805 = 10'h60 == _T_244[9:0] ? 4'h3 : _GEN_11804; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11806 = 10'h61 == _T_244[9:0] ? 4'h3 : _GEN_11805; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11807 = 10'h62 == _T_244[9:0] ? 4'h3 : _GEN_11806; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11808 = 10'h63 == _T_244[9:0] ? 4'h3 : _GEN_11807; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11809 = 10'h64 == _T_244[9:0] ? 4'h3 : _GEN_11808; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11810 = 10'h65 == _T_244[9:0] ? 4'hf : _GEN_11809; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11811 = 10'h66 == _T_244[9:0] ? 4'h3 : _GEN_11810; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11812 = 10'h67 == _T_244[9:0] ? 4'h3 : _GEN_11811; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11813 = 10'h68 == _T_244[9:0] ? 4'h3 : _GEN_11812; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11814 = 10'h69 == _T_244[9:0] ? 4'hf : _GEN_11813; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11815 = 10'h6a == _T_244[9:0] ? 4'h9 : _GEN_11814; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11816 = 10'h6b == _T_244[9:0] ? 4'h9 : _GEN_11815; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11817 = 10'h6c == _T_244[9:0] ? 4'h3 : _GEN_11816; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11818 = 10'h6d == _T_244[9:0] ? 4'h3 : _GEN_11817; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11819 = 10'h6e == _T_244[9:0] ? 4'h3 : _GEN_11818; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11820 = 10'h6f == _T_244[9:0] ? 4'h3 : _GEN_11819; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11821 = 10'h70 == _T_244[9:0] ? 4'h3 : _GEN_11820; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11822 = 10'h71 == _T_244[9:0] ? 4'h3 : _GEN_11821; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11823 = 10'h72 == _T_244[9:0] ? 4'h3 : _GEN_11822; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11824 = 10'h73 == _T_244[9:0] ? 4'h9 : _GEN_11823; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11825 = 10'h74 == _T_244[9:0] ? 4'hf : _GEN_11824; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11826 = 10'h75 == _T_244[9:0] ? 4'hf : _GEN_11825; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11827 = 10'h76 == _T_244[9:0] ? 4'hf : _GEN_11826; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11828 = 10'h77 == _T_244[9:0] ? 4'h3 : _GEN_11827; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11829 = 10'h78 == _T_244[9:0] ? 4'h3 : _GEN_11828; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11830 = 10'h79 == _T_244[9:0] ? 4'h3 : _GEN_11829; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11831 = 10'h7a == _T_244[9:0] ? 4'hf : _GEN_11830; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11832 = 10'h7b == _T_244[9:0] ? 4'h3 : _GEN_11831; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11833 = 10'h7c == _T_244[9:0] ? 4'h3 : _GEN_11832; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11834 = 10'h7d == _T_244[9:0] ? 4'h2 : _GEN_11833; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11835 = 10'h7e == _T_244[9:0] ? 4'h3 : _GEN_11834; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11836 = 10'h7f == _T_244[9:0] ? 4'h0 : _GEN_11835; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11837 = 10'h80 == _T_244[9:0] ? 4'h3 : _GEN_11836; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11838 = 10'h81 == _T_244[9:0] ? 4'h3 : _GEN_11837; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11839 = 10'h82 == _T_244[9:0] ? 4'h9 : _GEN_11838; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11840 = 10'h83 == _T_244[9:0] ? 4'hf : _GEN_11839; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11841 = 10'h84 == _T_244[9:0] ? 4'h2 : _GEN_11840; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11842 = 10'h85 == _T_244[9:0] ? 4'h9 : _GEN_11841; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11843 = 10'h86 == _T_244[9:0] ? 4'h9 : _GEN_11842; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11844 = 10'h87 == _T_244[9:0] ? 4'h3 : _GEN_11843; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11845 = 10'h88 == _T_244[9:0] ? 4'h3 : _GEN_11844; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11846 = 10'h89 == _T_244[9:0] ? 4'hf : _GEN_11845; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11847 = 10'h8a == _T_244[9:0] ? 4'hf : _GEN_11846; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11848 = 10'h8b == _T_244[9:0] ? 4'h9 : _GEN_11847; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11849 = 10'h8c == _T_244[9:0] ? 4'h9 : _GEN_11848; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11850 = 10'h8d == _T_244[9:0] ? 4'h9 : _GEN_11849; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11851 = 10'h8e == _T_244[9:0] ? 4'h9 : _GEN_11850; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11852 = 10'h8f == _T_244[9:0] ? 4'h9 : _GEN_11851; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11853 = 10'h90 == _T_244[9:0] ? 4'h9 : _GEN_11852; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11854 = 10'h91 == _T_244[9:0] ? 4'h9 : _GEN_11853; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11855 = 10'h92 == _T_244[9:0] ? 4'h9 : _GEN_11854; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11856 = 10'h93 == _T_244[9:0] ? 4'hf : _GEN_11855; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11857 = 10'h94 == _T_244[9:0] ? 4'hf : _GEN_11856; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11858 = 10'h95 == _T_244[9:0] ? 4'h3 : _GEN_11857; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11859 = 10'h96 == _T_244[9:0] ? 4'h3 : _GEN_11858; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11860 = 10'h97 == _T_244[9:0] ? 4'h3 : _GEN_11859; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11861 = 10'h98 == _T_244[9:0] ? 4'h9 : _GEN_11860; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11862 = 10'h99 == _T_244[9:0] ? 4'hf : _GEN_11861; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11863 = 10'h9a == _T_244[9:0] ? 4'h9 : _GEN_11862; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11864 = 10'h9b == _T_244[9:0] ? 4'h9 : _GEN_11863; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11865 = 10'h9c == _T_244[9:0] ? 4'h3 : _GEN_11864; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11866 = 10'h9d == _T_244[9:0] ? 4'h3 : _GEN_11865; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11867 = 10'h9e == _T_244[9:0] ? 4'h3 : _GEN_11866; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11868 = 10'h9f == _T_244[9:0] ? 4'h0 : _GEN_11867; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11869 = 10'ha0 == _T_244[9:0] ? 4'h3 : _GEN_11868; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11870 = 10'ha1 == _T_244[9:0] ? 4'h9 : _GEN_11869; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11871 = 10'ha2 == _T_244[9:0] ? 4'hf : _GEN_11870; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11872 = 10'ha3 == _T_244[9:0] ? 4'h3 : _GEN_11871; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11873 = 10'ha4 == _T_244[9:0] ? 4'h3 : _GEN_11872; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11874 = 10'ha5 == _T_244[9:0] ? 4'h3 : _GEN_11873; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11875 = 10'ha6 == _T_244[9:0] ? 4'h3 : _GEN_11874; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11876 = 10'ha7 == _T_244[9:0] ? 4'hf : _GEN_11875; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11877 = 10'ha8 == _T_244[9:0] ? 4'h3 : _GEN_11876; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11878 = 10'ha9 == _T_244[9:0] ? 4'h9 : _GEN_11877; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11879 = 10'haa == _T_244[9:0] ? 4'hf : _GEN_11878; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11880 = 10'hab == _T_244[9:0] ? 4'hf : _GEN_11879; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11881 = 10'hac == _T_244[9:0] ? 4'hf : _GEN_11880; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11882 = 10'had == _T_244[9:0] ? 4'hf : _GEN_11881; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11883 = 10'hae == _T_244[9:0] ? 4'hf : _GEN_11882; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11884 = 10'haf == _T_244[9:0] ? 4'hf : _GEN_11883; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11885 = 10'hb0 == _T_244[9:0] ? 4'hf : _GEN_11884; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11886 = 10'hb1 == _T_244[9:0] ? 4'hf : _GEN_11885; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11887 = 10'hb2 == _T_244[9:0] ? 4'hf : _GEN_11886; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11888 = 10'hb3 == _T_244[9:0] ? 4'hf : _GEN_11887; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11889 = 10'hb4 == _T_244[9:0] ? 4'h9 : _GEN_11888; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11890 = 10'hb5 == _T_244[9:0] ? 4'h9 : _GEN_11889; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11891 = 10'hb6 == _T_244[9:0] ? 4'h3 : _GEN_11890; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11892 = 10'hb7 == _T_244[9:0] ? 4'hf : _GEN_11891; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11893 = 10'hb8 == _T_244[9:0] ? 4'h3 : _GEN_11892; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11894 = 10'hb9 == _T_244[9:0] ? 4'h3 : _GEN_11893; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11895 = 10'hba == _T_244[9:0] ? 4'h3 : _GEN_11894; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11896 = 10'hbb == _T_244[9:0] ? 4'hf : _GEN_11895; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11897 = 10'hbc == _T_244[9:0] ? 4'h3 : _GEN_11896; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11898 = 10'hbd == _T_244[9:0] ? 4'h3 : _GEN_11897; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11899 = 10'hbe == _T_244[9:0] ? 4'h3 : _GEN_11898; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11900 = 10'hbf == _T_244[9:0] ? 4'h0 : _GEN_11899; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11901 = 10'hc0 == _T_244[9:0] ? 4'h3 : _GEN_11900; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11902 = 10'hc1 == _T_244[9:0] ? 4'h3 : _GEN_11901; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11903 = 10'hc2 == _T_244[9:0] ? 4'h3 : _GEN_11902; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11904 = 10'hc3 == _T_244[9:0] ? 4'h2 : _GEN_11903; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11905 = 10'hc4 == _T_244[9:0] ? 4'hf : _GEN_11904; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11906 = 10'hc5 == _T_244[9:0] ? 4'hf : _GEN_11905; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11907 = 10'hc6 == _T_244[9:0] ? 4'hf : _GEN_11906; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11908 = 10'hc7 == _T_244[9:0] ? 4'h3 : _GEN_11907; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11909 = 10'hc8 == _T_244[9:0] ? 4'h9 : _GEN_11908; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11910 = 10'hc9 == _T_244[9:0] ? 4'hf : _GEN_11909; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11911 = 10'hca == _T_244[9:0] ? 4'hf : _GEN_11910; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11912 = 10'hcb == _T_244[9:0] ? 4'hf : _GEN_11911; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11913 = 10'hcc == _T_244[9:0] ? 4'hf : _GEN_11912; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11914 = 10'hcd == _T_244[9:0] ? 4'hf : _GEN_11913; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11915 = 10'hce == _T_244[9:0] ? 4'hf : _GEN_11914; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11916 = 10'hcf == _T_244[9:0] ? 4'hf : _GEN_11915; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11917 = 10'hd0 == _T_244[9:0] ? 4'hf : _GEN_11916; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11918 = 10'hd1 == _T_244[9:0] ? 4'hf : _GEN_11917; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11919 = 10'hd2 == _T_244[9:0] ? 4'hf : _GEN_11918; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11920 = 10'hd3 == _T_244[9:0] ? 4'hf : _GEN_11919; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11921 = 10'hd4 == _T_244[9:0] ? 4'hf : _GEN_11920; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11922 = 10'hd5 == _T_244[9:0] ? 4'hf : _GEN_11921; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11923 = 10'hd6 == _T_244[9:0] ? 4'h9 : _GEN_11922; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11924 = 10'hd7 == _T_244[9:0] ? 4'h3 : _GEN_11923; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11925 = 10'hd8 == _T_244[9:0] ? 4'hf : _GEN_11924; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11926 = 10'hd9 == _T_244[9:0] ? 4'h3 : _GEN_11925; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11927 = 10'hda == _T_244[9:0] ? 4'h3 : _GEN_11926; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11928 = 10'hdb == _T_244[9:0] ? 4'h3 : _GEN_11927; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11929 = 10'hdc == _T_244[9:0] ? 4'h3 : _GEN_11928; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11930 = 10'hdd == _T_244[9:0] ? 4'h3 : _GEN_11929; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11931 = 10'hde == _T_244[9:0] ? 4'h2 : _GEN_11930; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11932 = 10'hdf == _T_244[9:0] ? 4'h0 : _GEN_11931; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11933 = 10'he0 == _T_244[9:0] ? 4'h3 : _GEN_11932; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11934 = 10'he1 == _T_244[9:0] ? 4'h3 : _GEN_11933; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11935 = 10'he2 == _T_244[9:0] ? 4'h3 : _GEN_11934; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11936 = 10'he3 == _T_244[9:0] ? 4'h3 : _GEN_11935; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11937 = 10'he4 == _T_244[9:0] ? 4'h3 : _GEN_11936; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11938 = 10'he5 == _T_244[9:0] ? 4'h3 : _GEN_11937; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11939 = 10'he6 == _T_244[9:0] ? 4'h3 : _GEN_11938; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11940 = 10'he7 == _T_244[9:0] ? 4'h9 : _GEN_11939; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11941 = 10'he8 == _T_244[9:0] ? 4'h9 : _GEN_11940; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11942 = 10'he9 == _T_244[9:0] ? 4'h9 : _GEN_11941; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11943 = 10'hea == _T_244[9:0] ? 4'hf : _GEN_11942; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11944 = 10'heb == _T_244[9:0] ? 4'hf : _GEN_11943; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11945 = 10'hec == _T_244[9:0] ? 4'hf : _GEN_11944; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11946 = 10'hed == _T_244[9:0] ? 4'hf : _GEN_11945; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11947 = 10'hee == _T_244[9:0] ? 4'hf : _GEN_11946; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11948 = 10'hef == _T_244[9:0] ? 4'hf : _GEN_11947; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11949 = 10'hf0 == _T_244[9:0] ? 4'hf : _GEN_11948; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11950 = 10'hf1 == _T_244[9:0] ? 4'hf : _GEN_11949; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11951 = 10'hf2 == _T_244[9:0] ? 4'hf : _GEN_11950; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11952 = 10'hf3 == _T_244[9:0] ? 4'hf : _GEN_11951; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11953 = 10'hf4 == _T_244[9:0] ? 4'hf : _GEN_11952; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11954 = 10'hf5 == _T_244[9:0] ? 4'h9 : _GEN_11953; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11955 = 10'hf6 == _T_244[9:0] ? 4'hf : _GEN_11954; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11956 = 10'hf7 == _T_244[9:0] ? 4'hf : _GEN_11955; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11957 = 10'hf8 == _T_244[9:0] ? 4'h9 : _GEN_11956; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11958 = 10'hf9 == _T_244[9:0] ? 4'hf : _GEN_11957; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11959 = 10'hfa == _T_244[9:0] ? 4'h3 : _GEN_11958; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11960 = 10'hfb == _T_244[9:0] ? 4'h3 : _GEN_11959; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11961 = 10'hfc == _T_244[9:0] ? 4'h3 : _GEN_11960; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11962 = 10'hfd == _T_244[9:0] ? 4'h3 : _GEN_11961; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11963 = 10'hfe == _T_244[9:0] ? 4'h3 : _GEN_11962; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11964 = 10'hff == _T_244[9:0] ? 4'h0 : _GEN_11963; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11965 = 10'h100 == _T_244[9:0] ? 4'h3 : _GEN_11964; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11966 = 10'h101 == _T_244[9:0] ? 4'hf : _GEN_11965; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11967 = 10'h102 == _T_244[9:0] ? 4'h3 : _GEN_11966; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11968 = 10'h103 == _T_244[9:0] ? 4'h3 : _GEN_11967; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11969 = 10'h104 == _T_244[9:0] ? 4'h3 : _GEN_11968; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11970 = 10'h105 == _T_244[9:0] ? 4'h3 : _GEN_11969; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11971 = 10'h106 == _T_244[9:0] ? 4'h3 : _GEN_11970; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11972 = 10'h107 == _T_244[9:0] ? 4'h3 : _GEN_11971; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11973 = 10'h108 == _T_244[9:0] ? 4'h9 : _GEN_11972; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11974 = 10'h109 == _T_244[9:0] ? 4'hf : _GEN_11973; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11975 = 10'h10a == _T_244[9:0] ? 4'hf : _GEN_11974; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11976 = 10'h10b == _T_244[9:0] ? 4'hf : _GEN_11975; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11977 = 10'h10c == _T_244[9:0] ? 4'hf : _GEN_11976; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11978 = 10'h10d == _T_244[9:0] ? 4'h0 : _GEN_11977; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11979 = 10'h10e == _T_244[9:0] ? 4'hf : _GEN_11978; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11980 = 10'h10f == _T_244[9:0] ? 4'hf : _GEN_11979; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11981 = 10'h110 == _T_244[9:0] ? 4'hf : _GEN_11980; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11982 = 10'h111 == _T_244[9:0] ? 4'h0 : _GEN_11981; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11983 = 10'h112 == _T_244[9:0] ? 4'hf : _GEN_11982; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11984 = 10'h113 == _T_244[9:0] ? 4'hf : _GEN_11983; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11985 = 10'h114 == _T_244[9:0] ? 4'hf : _GEN_11984; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11986 = 10'h115 == _T_244[9:0] ? 4'hf : _GEN_11985; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11987 = 10'h116 == _T_244[9:0] ? 4'h9 : _GEN_11986; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11988 = 10'h117 == _T_244[9:0] ? 4'h3 : _GEN_11987; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11989 = 10'h118 == _T_244[9:0] ? 4'h3 : _GEN_11988; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11990 = 10'h119 == _T_244[9:0] ? 4'h3 : _GEN_11989; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11991 = 10'h11a == _T_244[9:0] ? 4'hf : _GEN_11990; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11992 = 10'h11b == _T_244[9:0] ? 4'h3 : _GEN_11991; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11993 = 10'h11c == _T_244[9:0] ? 4'h3 : _GEN_11992; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11994 = 10'h11d == _T_244[9:0] ? 4'h2 : _GEN_11993; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11995 = 10'h11e == _T_244[9:0] ? 4'h3 : _GEN_11994; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11996 = 10'h11f == _T_244[9:0] ? 4'h0 : _GEN_11995; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11997 = 10'h120 == _T_244[9:0] ? 4'h3 : _GEN_11996; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11998 = 10'h121 == _T_244[9:0] ? 4'h3 : _GEN_11997; // @[Filter.scala 191:142]
  wire [3:0] _GEN_11999 = 10'h122 == _T_244[9:0] ? 4'h3 : _GEN_11998; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12000 = 10'h123 == _T_244[9:0] ? 4'h3 : _GEN_11999; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12001 = 10'h124 == _T_244[9:0] ? 4'h3 : _GEN_12000; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12002 = 10'h125 == _T_244[9:0] ? 4'h3 : _GEN_12001; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12003 = 10'h126 == _T_244[9:0] ? 4'h3 : _GEN_12002; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12004 = 10'h127 == _T_244[9:0] ? 4'h9 : _GEN_12003; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12005 = 10'h128 == _T_244[9:0] ? 4'hf : _GEN_12004; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12006 = 10'h129 == _T_244[9:0] ? 4'h3 : _GEN_12005; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12007 = 10'h12a == _T_244[9:0] ? 4'h3 : _GEN_12006; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12008 = 10'h12b == _T_244[9:0] ? 4'hf : _GEN_12007; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12009 = 10'h12c == _T_244[9:0] ? 4'hf : _GEN_12008; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12010 = 10'h12d == _T_244[9:0] ? 4'hf : _GEN_12009; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12011 = 10'h12e == _T_244[9:0] ? 4'hf : _GEN_12010; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12012 = 10'h12f == _T_244[9:0] ? 4'hf : _GEN_12011; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12013 = 10'h130 == _T_244[9:0] ? 4'hf : _GEN_12012; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12014 = 10'h131 == _T_244[9:0] ? 4'hf : _GEN_12013; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12015 = 10'h132 == _T_244[9:0] ? 4'hf : _GEN_12014; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12016 = 10'h133 == _T_244[9:0] ? 4'hf : _GEN_12015; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12017 = 10'h134 == _T_244[9:0] ? 4'h3 : _GEN_12016; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12018 = 10'h135 == _T_244[9:0] ? 4'h3 : _GEN_12017; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12019 = 10'h136 == _T_244[9:0] ? 4'hf : _GEN_12018; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12020 = 10'h137 == _T_244[9:0] ? 4'h9 : _GEN_12019; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12021 = 10'h138 == _T_244[9:0] ? 4'h3 : _GEN_12020; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12022 = 10'h139 == _T_244[9:0] ? 4'h3 : _GEN_12021; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12023 = 10'h13a == _T_244[9:0] ? 4'h3 : _GEN_12022; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12024 = 10'h13b == _T_244[9:0] ? 4'h3 : _GEN_12023; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12025 = 10'h13c == _T_244[9:0] ? 4'h3 : _GEN_12024; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12026 = 10'h13d == _T_244[9:0] ? 4'h3 : _GEN_12025; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12027 = 10'h13e == _T_244[9:0] ? 4'h3 : _GEN_12026; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12028 = 10'h13f == _T_244[9:0] ? 4'h0 : _GEN_12027; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12029 = 10'h140 == _T_244[9:0] ? 4'h3 : _GEN_12028; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12030 = 10'h141 == _T_244[9:0] ? 4'h3 : _GEN_12029; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12031 = 10'h142 == _T_244[9:0] ? 4'h2 : _GEN_12030; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12032 = 10'h143 == _T_244[9:0] ? 4'h3 : _GEN_12031; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12033 = 10'h144 == _T_244[9:0] ? 4'h3 : _GEN_12032; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12034 = 10'h145 == _T_244[9:0] ? 4'h3 : _GEN_12033; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12035 = 10'h146 == _T_244[9:0] ? 4'h9 : _GEN_12034; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12036 = 10'h147 == _T_244[9:0] ? 4'hf : _GEN_12035; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12037 = 10'h148 == _T_244[9:0] ? 4'h3 : _GEN_12036; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12038 = 10'h149 == _T_244[9:0] ? 4'h3 : _GEN_12037; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12039 = 10'h14a == _T_244[9:0] ? 4'h3 : _GEN_12038; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12040 = 10'h14b == _T_244[9:0] ? 4'h3 : _GEN_12039; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12041 = 10'h14c == _T_244[9:0] ? 4'h3 : _GEN_12040; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12042 = 10'h14d == _T_244[9:0] ? 4'h3 : _GEN_12041; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12043 = 10'h14e == _T_244[9:0] ? 4'h3 : _GEN_12042; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12044 = 10'h14f == _T_244[9:0] ? 4'h3 : _GEN_12043; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12045 = 10'h150 == _T_244[9:0] ? 4'h3 : _GEN_12044; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12046 = 10'h151 == _T_244[9:0] ? 4'h3 : _GEN_12045; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12047 = 10'h152 == _T_244[9:0] ? 4'h3 : _GEN_12046; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12048 = 10'h153 == _T_244[9:0] ? 4'h3 : _GEN_12047; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12049 = 10'h154 == _T_244[9:0] ? 4'h3 : _GEN_12048; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12050 = 10'h155 == _T_244[9:0] ? 4'h3 : _GEN_12049; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12051 = 10'h156 == _T_244[9:0] ? 4'h3 : _GEN_12050; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12052 = 10'h157 == _T_244[9:0] ? 4'hf : _GEN_12051; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12053 = 10'h158 == _T_244[9:0] ? 4'h3 : _GEN_12052; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12054 = 10'h159 == _T_244[9:0] ? 4'h3 : _GEN_12053; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12055 = 10'h15a == _T_244[9:0] ? 4'h3 : _GEN_12054; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12056 = 10'h15b == _T_244[9:0] ? 4'h3 : _GEN_12055; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12057 = 10'h15c == _T_244[9:0] ? 4'h3 : _GEN_12056; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12058 = 10'h15d == _T_244[9:0] ? 4'h3 : _GEN_12057; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12059 = 10'h15e == _T_244[9:0] ? 4'h2 : _GEN_12058; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12060 = 10'h15f == _T_244[9:0] ? 4'h0 : _GEN_12059; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12061 = 10'h160 == _T_244[9:0] ? 4'h3 : _GEN_12060; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12062 = 10'h161 == _T_244[9:0] ? 4'h3 : _GEN_12061; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12063 = 10'h162 == _T_244[9:0] ? 4'h3 : _GEN_12062; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12064 = 10'h163 == _T_244[9:0] ? 4'h2 : _GEN_12063; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12065 = 10'h164 == _T_244[9:0] ? 4'h3 : _GEN_12064; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12066 = 10'h165 == _T_244[9:0] ? 4'h9 : _GEN_12065; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12067 = 10'h166 == _T_244[9:0] ? 4'hf : _GEN_12066; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12068 = 10'h167 == _T_244[9:0] ? 4'hf : _GEN_12067; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12069 = 10'h168 == _T_244[9:0] ? 4'hd : _GEN_12068; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12070 = 10'h169 == _T_244[9:0] ? 4'h9 : _GEN_12069; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12071 = 10'h16a == _T_244[9:0] ? 4'hd : _GEN_12070; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12072 = 10'h16b == _T_244[9:0] ? 4'hd : _GEN_12071; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12073 = 10'h16c == _T_244[9:0] ? 4'h3 : _GEN_12072; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12074 = 10'h16d == _T_244[9:0] ? 4'h3 : _GEN_12073; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12075 = 10'h16e == _T_244[9:0] ? 4'h3 : _GEN_12074; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12076 = 10'h16f == _T_244[9:0] ? 4'h3 : _GEN_12075; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12077 = 10'h170 == _T_244[9:0] ? 4'h3 : _GEN_12076; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12078 = 10'h171 == _T_244[9:0] ? 4'h3 : _GEN_12077; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12079 = 10'h172 == _T_244[9:0] ? 4'h3 : _GEN_12078; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12080 = 10'h173 == _T_244[9:0] ? 4'h3 : _GEN_12079; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12081 = 10'h174 == _T_244[9:0] ? 4'h3 : _GEN_12080; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12082 = 10'h175 == _T_244[9:0] ? 4'h3 : _GEN_12081; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12083 = 10'h176 == _T_244[9:0] ? 4'hf : _GEN_12082; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12084 = 10'h177 == _T_244[9:0] ? 4'hf : _GEN_12083; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12085 = 10'h178 == _T_244[9:0] ? 4'h9 : _GEN_12084; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12086 = 10'h179 == _T_244[9:0] ? 4'h3 : _GEN_12085; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12087 = 10'h17a == _T_244[9:0] ? 4'h3 : _GEN_12086; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12088 = 10'h17b == _T_244[9:0] ? 4'h3 : _GEN_12087; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12089 = 10'h17c == _T_244[9:0] ? 4'h3 : _GEN_12088; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12090 = 10'h17d == _T_244[9:0] ? 4'h2 : _GEN_12089; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12091 = 10'h17e == _T_244[9:0] ? 4'h3 : _GEN_12090; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12092 = 10'h17f == _T_244[9:0] ? 4'h0 : _GEN_12091; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12093 = 10'h180 == _T_244[9:0] ? 4'hd : _GEN_12092; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12094 = 10'h181 == _T_244[9:0] ? 4'hd : _GEN_12093; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12095 = 10'h182 == _T_244[9:0] ? 4'hd : _GEN_12094; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12096 = 10'h183 == _T_244[9:0] ? 4'hd : _GEN_12095; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12097 = 10'h184 == _T_244[9:0] ? 4'h3 : _GEN_12096; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12098 = 10'h185 == _T_244[9:0] ? 4'h9 : _GEN_12097; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12099 = 10'h186 == _T_244[9:0] ? 4'hb : _GEN_12098; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12100 = 10'h187 == _T_244[9:0] ? 4'hf : _GEN_12099; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12101 = 10'h188 == _T_244[9:0] ? 4'hd : _GEN_12100; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12102 = 10'h189 == _T_244[9:0] ? 4'hd : _GEN_12101; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12103 = 10'h18a == _T_244[9:0] ? 4'hd : _GEN_12102; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12104 = 10'h18b == _T_244[9:0] ? 4'hd : _GEN_12103; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12105 = 10'h18c == _T_244[9:0] ? 4'hd : _GEN_12104; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12106 = 10'h18d == _T_244[9:0] ? 4'hd : _GEN_12105; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12107 = 10'h18e == _T_244[9:0] ? 4'hd : _GEN_12106; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12108 = 10'h18f == _T_244[9:0] ? 4'hd : _GEN_12107; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12109 = 10'h190 == _T_244[9:0] ? 4'hd : _GEN_12108; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12110 = 10'h191 == _T_244[9:0] ? 4'hd : _GEN_12109; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12111 = 10'h192 == _T_244[9:0] ? 4'h9 : _GEN_12110; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12112 = 10'h193 == _T_244[9:0] ? 4'hd : _GEN_12111; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12113 = 10'h194 == _T_244[9:0] ? 4'hd : _GEN_12112; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12114 = 10'h195 == _T_244[9:0] ? 4'hd : _GEN_12113; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12115 = 10'h196 == _T_244[9:0] ? 4'hf : _GEN_12114; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12116 = 10'h197 == _T_244[9:0] ? 4'h3 : _GEN_12115; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12117 = 10'h198 == _T_244[9:0] ? 4'h9 : _GEN_12116; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12118 = 10'h199 == _T_244[9:0] ? 4'h3 : _GEN_12117; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12119 = 10'h19a == _T_244[9:0] ? 4'h3 : _GEN_12118; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12120 = 10'h19b == _T_244[9:0] ? 4'h3 : _GEN_12119; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12121 = 10'h19c == _T_244[9:0] ? 4'h3 : _GEN_12120; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12122 = 10'h19d == _T_244[9:0] ? 4'h3 : _GEN_12121; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12123 = 10'h19e == _T_244[9:0] ? 4'h3 : _GEN_12122; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12124 = 10'h19f == _T_244[9:0] ? 4'h0 : _GEN_12123; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12125 = 10'h1a0 == _T_244[9:0] ? 4'hd : _GEN_12124; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12126 = 10'h1a1 == _T_244[9:0] ? 4'hd : _GEN_12125; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12127 = 10'h1a2 == _T_244[9:0] ? 4'h9 : _GEN_12126; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12128 = 10'h1a3 == _T_244[9:0] ? 4'hd : _GEN_12127; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12129 = 10'h1a4 == _T_244[9:0] ? 4'h3 : _GEN_12128; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12130 = 10'h1a5 == _T_244[9:0] ? 4'hf : _GEN_12129; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12131 = 10'h1a6 == _T_244[9:0] ? 4'hd : _GEN_12130; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12132 = 10'h1a7 == _T_244[9:0] ? 4'hf : _GEN_12131; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12133 = 10'h1a8 == _T_244[9:0] ? 4'hb : _GEN_12132; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12134 = 10'h1a9 == _T_244[9:0] ? 4'hd : _GEN_12133; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12135 = 10'h1aa == _T_244[9:0] ? 4'hd : _GEN_12134; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12136 = 10'h1ab == _T_244[9:0] ? 4'h9 : _GEN_12135; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12137 = 10'h1ac == _T_244[9:0] ? 4'hd : _GEN_12136; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12138 = 10'h1ad == _T_244[9:0] ? 4'hd : _GEN_12137; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12139 = 10'h1ae == _T_244[9:0] ? 4'hd : _GEN_12138; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12140 = 10'h1af == _T_244[9:0] ? 4'hd : _GEN_12139; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12141 = 10'h1b0 == _T_244[9:0] ? 4'hd : _GEN_12140; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12142 = 10'h1b1 == _T_244[9:0] ? 4'hd : _GEN_12141; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12143 = 10'h1b2 == _T_244[9:0] ? 4'hd : _GEN_12142; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12144 = 10'h1b3 == _T_244[9:0] ? 4'hd : _GEN_12143; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12145 = 10'h1b4 == _T_244[9:0] ? 4'hd : _GEN_12144; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12146 = 10'h1b5 == _T_244[9:0] ? 4'hd : _GEN_12145; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12147 = 10'h1b6 == _T_244[9:0] ? 4'hf : _GEN_12146; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12148 = 10'h1b7 == _T_244[9:0] ? 4'hd : _GEN_12147; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12149 = 10'h1b8 == _T_244[9:0] ? 4'hf : _GEN_12148; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12150 = 10'h1b9 == _T_244[9:0] ? 4'hd : _GEN_12149; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12151 = 10'h1ba == _T_244[9:0] ? 4'hd : _GEN_12150; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12152 = 10'h1bb == _T_244[9:0] ? 4'hd : _GEN_12151; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12153 = 10'h1bc == _T_244[9:0] ? 4'h2 : _GEN_12152; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12154 = 10'h1bd == _T_244[9:0] ? 4'h3 : _GEN_12153; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12155 = 10'h1be == _T_244[9:0] ? 4'hd : _GEN_12154; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12156 = 10'h1bf == _T_244[9:0] ? 4'h0 : _GEN_12155; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12157 = 10'h1c0 == _T_244[9:0] ? 4'hd : _GEN_12156; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12158 = 10'h1c1 == _T_244[9:0] ? 4'hd : _GEN_12157; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12159 = 10'h1c2 == _T_244[9:0] ? 4'hd : _GEN_12158; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12160 = 10'h1c3 == _T_244[9:0] ? 4'h2 : _GEN_12159; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12161 = 10'h1c4 == _T_244[9:0] ? 4'h2 : _GEN_12160; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12162 = 10'h1c5 == _T_244[9:0] ? 4'hd : _GEN_12161; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12163 = 10'h1c6 == _T_244[9:0] ? 4'hd : _GEN_12162; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12164 = 10'h1c7 == _T_244[9:0] ? 4'hd : _GEN_12163; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12165 = 10'h1c8 == _T_244[9:0] ? 4'hd : _GEN_12164; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12166 = 10'h1c9 == _T_244[9:0] ? 4'hb : _GEN_12165; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12167 = 10'h1ca == _T_244[9:0] ? 4'hb : _GEN_12166; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12168 = 10'h1cb == _T_244[9:0] ? 4'hb : _GEN_12167; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12169 = 10'h1cc == _T_244[9:0] ? 4'hb : _GEN_12168; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12170 = 10'h1cd == _T_244[9:0] ? 4'hb : _GEN_12169; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12171 = 10'h1ce == _T_244[9:0] ? 4'hb : _GEN_12170; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12172 = 10'h1cf == _T_244[9:0] ? 4'hb : _GEN_12171; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12173 = 10'h1d0 == _T_244[9:0] ? 4'hb : _GEN_12172; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12174 = 10'h1d1 == _T_244[9:0] ? 4'hb : _GEN_12173; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12175 = 10'h1d2 == _T_244[9:0] ? 4'hb : _GEN_12174; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12176 = 10'h1d3 == _T_244[9:0] ? 4'hb : _GEN_12175; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12177 = 10'h1d4 == _T_244[9:0] ? 4'hb : _GEN_12176; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12178 = 10'h1d5 == _T_244[9:0] ? 4'hb : _GEN_12177; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12179 = 10'h1d6 == _T_244[9:0] ? 4'hd : _GEN_12178; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12180 = 10'h1d7 == _T_244[9:0] ? 4'hd : _GEN_12179; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12181 = 10'h1d8 == _T_244[9:0] ? 4'hd : _GEN_12180; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12182 = 10'h1d9 == _T_244[9:0] ? 4'hd : _GEN_12181; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12183 = 10'h1da == _T_244[9:0] ? 4'hd : _GEN_12182; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12184 = 10'h1db == _T_244[9:0] ? 4'hd : _GEN_12183; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12185 = 10'h1dc == _T_244[9:0] ? 4'hd : _GEN_12184; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12186 = 10'h1dd == _T_244[9:0] ? 4'h3 : _GEN_12185; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12187 = 10'h1de == _T_244[9:0] ? 4'hd : _GEN_12186; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12188 = 10'h1df == _T_244[9:0] ? 4'h0 : _GEN_12187; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12189 = 10'h1e0 == _T_244[9:0] ? 4'h9 : _GEN_12188; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12190 = 10'h1e1 == _T_244[9:0] ? 4'hd : _GEN_12189; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12191 = 10'h1e2 == _T_244[9:0] ? 4'h2 : _GEN_12190; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12192 = 10'h1e3 == _T_244[9:0] ? 4'h2 : _GEN_12191; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12193 = 10'h1e4 == _T_244[9:0] ? 4'hd : _GEN_12192; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12194 = 10'h1e5 == _T_244[9:0] ? 4'hd : _GEN_12193; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12195 = 10'h1e6 == _T_244[9:0] ? 4'hd : _GEN_12194; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12196 = 10'h1e7 == _T_244[9:0] ? 4'hd : _GEN_12195; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12197 = 10'h1e8 == _T_244[9:0] ? 4'hb : _GEN_12196; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12198 = 10'h1e9 == _T_244[9:0] ? 4'hd : _GEN_12197; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12199 = 10'h1ea == _T_244[9:0] ? 4'hd : _GEN_12198; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12200 = 10'h1eb == _T_244[9:0] ? 4'hb : _GEN_12199; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12201 = 10'h1ec == _T_244[9:0] ? 4'hd : _GEN_12200; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12202 = 10'h1ed == _T_244[9:0] ? 4'hb : _GEN_12201; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12203 = 10'h1ee == _T_244[9:0] ? 4'hd : _GEN_12202; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12204 = 10'h1ef == _T_244[9:0] ? 4'hb : _GEN_12203; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12205 = 10'h1f0 == _T_244[9:0] ? 4'hd : _GEN_12204; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12206 = 10'h1f1 == _T_244[9:0] ? 4'hb : _GEN_12205; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12207 = 10'h1f2 == _T_244[9:0] ? 4'hb : _GEN_12206; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12208 = 10'h1f3 == _T_244[9:0] ? 4'hd : _GEN_12207; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12209 = 10'h1f4 == _T_244[9:0] ? 4'hb : _GEN_12208; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12210 = 10'h1f5 == _T_244[9:0] ? 4'hb : _GEN_12209; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12211 = 10'h1f6 == _T_244[9:0] ? 4'hd : _GEN_12210; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12212 = 10'h1f7 == _T_244[9:0] ? 4'hd : _GEN_12211; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12213 = 10'h1f8 == _T_244[9:0] ? 4'hd : _GEN_12212; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12214 = 10'h1f9 == _T_244[9:0] ? 4'hd : _GEN_12213; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12215 = 10'h1fa == _T_244[9:0] ? 4'h9 : _GEN_12214; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12216 = 10'h1fb == _T_244[9:0] ? 4'hd : _GEN_12215; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12217 = 10'h1fc == _T_244[9:0] ? 4'hd : _GEN_12216; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12218 = 10'h1fd == _T_244[9:0] ? 4'h2 : _GEN_12217; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12219 = 10'h1fe == _T_244[9:0] ? 4'hd : _GEN_12218; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12220 = 10'h1ff == _T_244[9:0] ? 4'h0 : _GEN_12219; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12221 = 10'h200 == _T_244[9:0] ? 4'hd : _GEN_12220; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12222 = 10'h201 == _T_244[9:0] ? 4'hd : _GEN_12221; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12223 = 10'h202 == _T_244[9:0] ? 4'h3 : _GEN_12222; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12224 = 10'h203 == _T_244[9:0] ? 4'hd : _GEN_12223; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12225 = 10'h204 == _T_244[9:0] ? 4'hd : _GEN_12224; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12226 = 10'h205 == _T_244[9:0] ? 4'hd : _GEN_12225; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12227 = 10'h206 == _T_244[9:0] ? 4'hb : _GEN_12226; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12228 = 10'h207 == _T_244[9:0] ? 4'hb : _GEN_12227; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12229 = 10'h208 == _T_244[9:0] ? 4'hd : _GEN_12228; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12230 = 10'h209 == _T_244[9:0] ? 4'hd : _GEN_12229; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12231 = 10'h20a == _T_244[9:0] ? 4'hd : _GEN_12230; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12232 = 10'h20b == _T_244[9:0] ? 4'hb : _GEN_12231; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12233 = 10'h20c == _T_244[9:0] ? 4'hd : _GEN_12232; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12234 = 10'h20d == _T_244[9:0] ? 4'hb : _GEN_12233; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12235 = 10'h20e == _T_244[9:0] ? 4'hd : _GEN_12234; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12236 = 10'h20f == _T_244[9:0] ? 4'hb : _GEN_12235; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12237 = 10'h210 == _T_244[9:0] ? 4'hd : _GEN_12236; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12238 = 10'h211 == _T_244[9:0] ? 4'hd : _GEN_12237; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12239 = 10'h212 == _T_244[9:0] ? 4'hb : _GEN_12238; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12240 = 10'h213 == _T_244[9:0] ? 4'hb : _GEN_12239; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12241 = 10'h214 == _T_244[9:0] ? 4'hb : _GEN_12240; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12242 = 10'h215 == _T_244[9:0] ? 4'hd : _GEN_12241; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12243 = 10'h216 == _T_244[9:0] ? 4'hd : _GEN_12242; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12244 = 10'h217 == _T_244[9:0] ? 4'hd : _GEN_12243; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12245 = 10'h218 == _T_244[9:0] ? 4'hd : _GEN_12244; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12246 = 10'h219 == _T_244[9:0] ? 4'hd : _GEN_12245; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12247 = 10'h21a == _T_244[9:0] ? 4'hd : _GEN_12246; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12248 = 10'h21b == _T_244[9:0] ? 4'hd : _GEN_12247; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12249 = 10'h21c == _T_244[9:0] ? 4'h3 : _GEN_12248; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12250 = 10'h21d == _T_244[9:0] ? 4'h2 : _GEN_12249; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12251 = 10'h21e == _T_244[9:0] ? 4'hd : _GEN_12250; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12252 = 10'h21f == _T_244[9:0] ? 4'h0 : _GEN_12251; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12253 = 10'h220 == _T_244[9:0] ? 4'h0 : _GEN_12252; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12254 = 10'h221 == _T_244[9:0] ? 4'h0 : _GEN_12253; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12255 = 10'h222 == _T_244[9:0] ? 4'h0 : _GEN_12254; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12256 = 10'h223 == _T_244[9:0] ? 4'h0 : _GEN_12255; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12257 = 10'h224 == _T_244[9:0] ? 4'h0 : _GEN_12256; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12258 = 10'h225 == _T_244[9:0] ? 4'h0 : _GEN_12257; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12259 = 10'h226 == _T_244[9:0] ? 4'h0 : _GEN_12258; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12260 = 10'h227 == _T_244[9:0] ? 4'h0 : _GEN_12259; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12261 = 10'h228 == _T_244[9:0] ? 4'h0 : _GEN_12260; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12262 = 10'h229 == _T_244[9:0] ? 4'h0 : _GEN_12261; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12263 = 10'h22a == _T_244[9:0] ? 4'h0 : _GEN_12262; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12264 = 10'h22b == _T_244[9:0] ? 4'h0 : _GEN_12263; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12265 = 10'h22c == _T_244[9:0] ? 4'h0 : _GEN_12264; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12266 = 10'h22d == _T_244[9:0] ? 4'h0 : _GEN_12265; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12267 = 10'h22e == _T_244[9:0] ? 4'h0 : _GEN_12266; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12268 = 10'h22f == _T_244[9:0] ? 4'h0 : _GEN_12267; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12269 = 10'h230 == _T_244[9:0] ? 4'h0 : _GEN_12268; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12270 = 10'h231 == _T_244[9:0] ? 4'h0 : _GEN_12269; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12271 = 10'h232 == _T_244[9:0] ? 4'h0 : _GEN_12270; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12272 = 10'h233 == _T_244[9:0] ? 4'h0 : _GEN_12271; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12273 = 10'h234 == _T_244[9:0] ? 4'h0 : _GEN_12272; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12274 = 10'h235 == _T_244[9:0] ? 4'h0 : _GEN_12273; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12275 = 10'h236 == _T_244[9:0] ? 4'h0 : _GEN_12274; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12276 = 10'h237 == _T_244[9:0] ? 4'h0 : _GEN_12275; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12277 = 10'h238 == _T_244[9:0] ? 4'h0 : _GEN_12276; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12278 = 10'h239 == _T_244[9:0] ? 4'h0 : _GEN_12277; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12279 = 10'h23a == _T_244[9:0] ? 4'h0 : _GEN_12278; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12280 = 10'h23b == _T_244[9:0] ? 4'h0 : _GEN_12279; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12281 = 10'h23c == _T_244[9:0] ? 4'h0 : _GEN_12280; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12282 = 10'h23d == _T_244[9:0] ? 4'h0 : _GEN_12281; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12283 = 10'h23e == _T_244[9:0] ? 4'h0 : _GEN_12282; // @[Filter.scala 191:142]
  wire [3:0] _GEN_12284 = 10'h23f == _T_244[9:0] ? 4'h0 : _GEN_12283; // @[Filter.scala 191:142]
  wire [7:0] _T_258 = _GEN_12284 * 4'ha; // @[Filter.scala 191:142]
  wire [10:0] _GEN_28339 = {{3'd0}, _T_258}; // @[Filter.scala 191:109]
  wire [10:0] _T_260 = _T_253 + _GEN_28339; // @[Filter.scala 191:109]
  wire [10:0] _T_261 = _T_260 / 11'h64; // @[Filter.scala 191:150]
  wire  _T_263 = _T_234 >= 6'h20; // @[Filter.scala 194:31]
  wire  _T_267 = _T_241 >= 32'h12; // @[Filter.scala 194:63]
  wire  _T_268 = _T_263 | _T_267; // @[Filter.scala 194:58]
  wire [10:0] _GEN_12861 = io_SPI_distort ? _T_261 : {{7'd0}, _GEN_11132}; // @[Filter.scala 196:35]
  wire [10:0] _GEN_12862 = _T_268 ? 11'h0 : _GEN_12861; // @[Filter.scala 194:80]
  wire [10:0] _GEN_13439 = io_SPI_distort ? _T_261 : {{7'd0}, _GEN_11708}; // @[Filter.scala 196:35]
  wire [10:0] _GEN_13440 = _T_268 ? 11'h0 : _GEN_13439; // @[Filter.scala 194:80]
  wire [10:0] _GEN_14017 = io_SPI_distort ? _T_261 : {{7'd0}, _GEN_12284}; // @[Filter.scala 196:35]
  wire [10:0] _GEN_14018 = _T_268 ? 11'h0 : _GEN_14017; // @[Filter.scala 194:80]
  wire [31:0] _T_296 = pixelIndex + 32'h4; // @[Filter.scala 189:31]
  wire [31:0] _GEN_4 = _T_296 % 32'h20; // @[Filter.scala 189:38]
  wire [5:0] _T_297 = _GEN_4[5:0]; // @[Filter.scala 189:38]
  wire [5:0] _T_299 = _T_297 + _GEN_28295; // @[Filter.scala 189:53]
  wire [5:0] _T_301 = _T_299 - 6'h1; // @[Filter.scala 189:69]
  wire [31:0] _T_304 = _T_296 / 32'h20; // @[Filter.scala 190:38]
  wire [31:0] _T_306 = _T_304 + _GEN_28296; // @[Filter.scala 190:53]
  wire [31:0] _T_308 = _T_306 - 32'h1; // @[Filter.scala 190:69]
  wire [37:0] _T_309 = _T_308 * 32'h20; // @[Filter.scala 191:42]
  wire [37:0] _GEN_28345 = {{32'd0}, _T_301}; // @[Filter.scala 191:57]
  wire [37:0] _T_311 = _T_309 + _GEN_28345; // @[Filter.scala 191:57]
  wire [3:0] _GEN_14022 = 10'h3 == _T_311[9:0] ? 4'h3 : 4'ha; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14023 = 10'h4 == _T_311[9:0] ? 4'ha : _GEN_14022; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14024 = 10'h5 == _T_311[9:0] ? 4'ha : _GEN_14023; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14025 = 10'h6 == _T_311[9:0] ? 4'ha : _GEN_14024; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14026 = 10'h7 == _T_311[9:0] ? 4'ha : _GEN_14025; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14027 = 10'h8 == _T_311[9:0] ? 4'ha : _GEN_14026; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14028 = 10'h9 == _T_311[9:0] ? 4'ha : _GEN_14027; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14029 = 10'ha == _T_311[9:0] ? 4'ha : _GEN_14028; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14030 = 10'hb == _T_311[9:0] ? 4'ha : _GEN_14029; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14031 = 10'hc == _T_311[9:0] ? 4'ha : _GEN_14030; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14032 = 10'hd == _T_311[9:0] ? 4'ha : _GEN_14031; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14033 = 10'he == _T_311[9:0] ? 4'ha : _GEN_14032; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14034 = 10'hf == _T_311[9:0] ? 4'ha : _GEN_14033; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14035 = 10'h10 == _T_311[9:0] ? 4'ha : _GEN_14034; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14036 = 10'h11 == _T_311[9:0] ? 4'ha : _GEN_14035; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14037 = 10'h12 == _T_311[9:0] ? 4'ha : _GEN_14036; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14038 = 10'h13 == _T_311[9:0] ? 4'ha : _GEN_14037; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14039 = 10'h14 == _T_311[9:0] ? 4'ha : _GEN_14038; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14040 = 10'h15 == _T_311[9:0] ? 4'ha : _GEN_14039; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14041 = 10'h16 == _T_311[9:0] ? 4'ha : _GEN_14040; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14042 = 10'h17 == _T_311[9:0] ? 4'ha : _GEN_14041; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14043 = 10'h18 == _T_311[9:0] ? 4'ha : _GEN_14042; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14044 = 10'h19 == _T_311[9:0] ? 4'ha : _GEN_14043; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14045 = 10'h1a == _T_311[9:0] ? 4'ha : _GEN_14044; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14046 = 10'h1b == _T_311[9:0] ? 4'ha : _GEN_14045; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14047 = 10'h1c == _T_311[9:0] ? 4'ha : _GEN_14046; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14048 = 10'h1d == _T_311[9:0] ? 4'ha : _GEN_14047; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14049 = 10'h1e == _T_311[9:0] ? 4'ha : _GEN_14048; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14050 = 10'h1f == _T_311[9:0] ? 4'h0 : _GEN_14049; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14051 = 10'h20 == _T_311[9:0] ? 4'ha : _GEN_14050; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14052 = 10'h21 == _T_311[9:0] ? 4'ha : _GEN_14051; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14053 = 10'h22 == _T_311[9:0] ? 4'ha : _GEN_14052; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14054 = 10'h23 == _T_311[9:0] ? 4'h3 : _GEN_14053; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14055 = 10'h24 == _T_311[9:0] ? 4'ha : _GEN_14054; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14056 = 10'h25 == _T_311[9:0] ? 4'ha : _GEN_14055; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14057 = 10'h26 == _T_311[9:0] ? 4'ha : _GEN_14056; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14058 = 10'h27 == _T_311[9:0] ? 4'h1 : _GEN_14057; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14059 = 10'h28 == _T_311[9:0] ? 4'h1 : _GEN_14058; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14060 = 10'h29 == _T_311[9:0] ? 4'ha : _GEN_14059; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14061 = 10'h2a == _T_311[9:0] ? 4'ha : _GEN_14060; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14062 = 10'h2b == _T_311[9:0] ? 4'ha : _GEN_14061; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14063 = 10'h2c == _T_311[9:0] ? 4'ha : _GEN_14062; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14064 = 10'h2d == _T_311[9:0] ? 4'ha : _GEN_14063; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14065 = 10'h2e == _T_311[9:0] ? 4'ha : _GEN_14064; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14066 = 10'h2f == _T_311[9:0] ? 4'ha : _GEN_14065; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14067 = 10'h30 == _T_311[9:0] ? 4'ha : _GEN_14066; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14068 = 10'h31 == _T_311[9:0] ? 4'ha : _GEN_14067; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14069 = 10'h32 == _T_311[9:0] ? 4'ha : _GEN_14068; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14070 = 10'h33 == _T_311[9:0] ? 4'ha : _GEN_14069; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14071 = 10'h34 == _T_311[9:0] ? 4'ha : _GEN_14070; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14072 = 10'h35 == _T_311[9:0] ? 4'ha : _GEN_14071; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14073 = 10'h36 == _T_311[9:0] ? 4'ha : _GEN_14072; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14074 = 10'h37 == _T_311[9:0] ? 4'h1 : _GEN_14073; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14075 = 10'h38 == _T_311[9:0] ? 4'h1 : _GEN_14074; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14076 = 10'h39 == _T_311[9:0] ? 4'ha : _GEN_14075; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14077 = 10'h3a == _T_311[9:0] ? 4'ha : _GEN_14076; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14078 = 10'h3b == _T_311[9:0] ? 4'ha : _GEN_14077; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14079 = 10'h3c == _T_311[9:0] ? 4'ha : _GEN_14078; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14080 = 10'h3d == _T_311[9:0] ? 4'h3 : _GEN_14079; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14081 = 10'h3e == _T_311[9:0] ? 4'ha : _GEN_14080; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14082 = 10'h3f == _T_311[9:0] ? 4'h0 : _GEN_14081; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14083 = 10'h40 == _T_311[9:0] ? 4'ha : _GEN_14082; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14084 = 10'h41 == _T_311[9:0] ? 4'ha : _GEN_14083; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14085 = 10'h42 == _T_311[9:0] ? 4'ha : _GEN_14084; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14086 = 10'h43 == _T_311[9:0] ? 4'h2 : _GEN_14085; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14087 = 10'h44 == _T_311[9:0] ? 4'h3 : _GEN_14086; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14088 = 10'h45 == _T_311[9:0] ? 4'h0 : _GEN_14087; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14089 = 10'h46 == _T_311[9:0] ? 4'h0 : _GEN_14088; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14090 = 10'h47 == _T_311[9:0] ? 4'h0 : _GEN_14089; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14091 = 10'h48 == _T_311[9:0] ? 4'h0 : _GEN_14090; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14092 = 10'h49 == _T_311[9:0] ? 4'ha : _GEN_14091; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14093 = 10'h4a == _T_311[9:0] ? 4'ha : _GEN_14092; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14094 = 10'h4b == _T_311[9:0] ? 4'ha : _GEN_14093; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14095 = 10'h4c == _T_311[9:0] ? 4'ha : _GEN_14094; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14096 = 10'h4d == _T_311[9:0] ? 4'ha : _GEN_14095; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14097 = 10'h4e == _T_311[9:0] ? 4'ha : _GEN_14096; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14098 = 10'h4f == _T_311[9:0] ? 4'ha : _GEN_14097; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14099 = 10'h50 == _T_311[9:0] ? 4'ha : _GEN_14098; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14100 = 10'h51 == _T_311[9:0] ? 4'ha : _GEN_14099; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14101 = 10'h52 == _T_311[9:0] ? 4'ha : _GEN_14100; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14102 = 10'h53 == _T_311[9:0] ? 4'ha : _GEN_14101; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14103 = 10'h54 == _T_311[9:0] ? 4'h1 : _GEN_14102; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14104 = 10'h55 == _T_311[9:0] ? 4'h1 : _GEN_14103; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14105 = 10'h56 == _T_311[9:0] ? 4'h1 : _GEN_14104; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14106 = 10'h57 == _T_311[9:0] ? 4'h0 : _GEN_14105; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14107 = 10'h58 == _T_311[9:0] ? 4'ha : _GEN_14106; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14108 = 10'h59 == _T_311[9:0] ? 4'h0 : _GEN_14107; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14109 = 10'h5a == _T_311[9:0] ? 4'ha : _GEN_14108; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14110 = 10'h5b == _T_311[9:0] ? 4'ha : _GEN_14109; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14111 = 10'h5c == _T_311[9:0] ? 4'ha : _GEN_14110; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14112 = 10'h5d == _T_311[9:0] ? 4'h3 : _GEN_14111; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14113 = 10'h5e == _T_311[9:0] ? 4'ha : _GEN_14112; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14114 = 10'h5f == _T_311[9:0] ? 4'h0 : _GEN_14113; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14115 = 10'h60 == _T_311[9:0] ? 4'ha : _GEN_14114; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14116 = 10'h61 == _T_311[9:0] ? 4'ha : _GEN_14115; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14117 = 10'h62 == _T_311[9:0] ? 4'ha : _GEN_14116; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14118 = 10'h63 == _T_311[9:0] ? 4'ha : _GEN_14117; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14119 = 10'h64 == _T_311[9:0] ? 4'h3 : _GEN_14118; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14120 = 10'h65 == _T_311[9:0] ? 4'h0 : _GEN_14119; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14121 = 10'h66 == _T_311[9:0] ? 4'ha : _GEN_14120; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14122 = 10'h67 == _T_311[9:0] ? 4'ha : _GEN_14121; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14123 = 10'h68 == _T_311[9:0] ? 4'ha : _GEN_14122; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14124 = 10'h69 == _T_311[9:0] ? 4'h0 : _GEN_14123; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14125 = 10'h6a == _T_311[9:0] ? 4'h1 : _GEN_14124; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14126 = 10'h6b == _T_311[9:0] ? 4'h1 : _GEN_14125; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14127 = 10'h6c == _T_311[9:0] ? 4'ha : _GEN_14126; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14128 = 10'h6d == _T_311[9:0] ? 4'ha : _GEN_14127; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14129 = 10'h6e == _T_311[9:0] ? 4'ha : _GEN_14128; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14130 = 10'h6f == _T_311[9:0] ? 4'ha : _GEN_14129; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14131 = 10'h70 == _T_311[9:0] ? 4'ha : _GEN_14130; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14132 = 10'h71 == _T_311[9:0] ? 4'ha : _GEN_14131; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14133 = 10'h72 == _T_311[9:0] ? 4'ha : _GEN_14132; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14134 = 10'h73 == _T_311[9:0] ? 4'h1 : _GEN_14133; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14135 = 10'h74 == _T_311[9:0] ? 4'h0 : _GEN_14134; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14136 = 10'h75 == _T_311[9:0] ? 4'h0 : _GEN_14135; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14137 = 10'h76 == _T_311[9:0] ? 4'h0 : _GEN_14136; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14138 = 10'h77 == _T_311[9:0] ? 4'ha : _GEN_14137; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14139 = 10'h78 == _T_311[9:0] ? 4'ha : _GEN_14138; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14140 = 10'h79 == _T_311[9:0] ? 4'ha : _GEN_14139; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14141 = 10'h7a == _T_311[9:0] ? 4'h0 : _GEN_14140; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14142 = 10'h7b == _T_311[9:0] ? 4'ha : _GEN_14141; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14143 = 10'h7c == _T_311[9:0] ? 4'ha : _GEN_14142; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14144 = 10'h7d == _T_311[9:0] ? 4'h2 : _GEN_14143; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14145 = 10'h7e == _T_311[9:0] ? 4'h3 : _GEN_14144; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14146 = 10'h7f == _T_311[9:0] ? 4'h0 : _GEN_14145; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14147 = 10'h80 == _T_311[9:0] ? 4'ha : _GEN_14146; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14148 = 10'h81 == _T_311[9:0] ? 4'ha : _GEN_14147; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14149 = 10'h82 == _T_311[9:0] ? 4'h1 : _GEN_14148; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14150 = 10'h83 == _T_311[9:0] ? 4'h0 : _GEN_14149; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14151 = 10'h84 == _T_311[9:0] ? 4'h2 : _GEN_14150; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14152 = 10'h85 == _T_311[9:0] ? 4'h1 : _GEN_14151; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14153 = 10'h86 == _T_311[9:0] ? 4'h1 : _GEN_14152; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14154 = 10'h87 == _T_311[9:0] ? 4'ha : _GEN_14153; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14155 = 10'h88 == _T_311[9:0] ? 4'ha : _GEN_14154; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14156 = 10'h89 == _T_311[9:0] ? 4'h0 : _GEN_14155; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14157 = 10'h8a == _T_311[9:0] ? 4'h0 : _GEN_14156; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14158 = 10'h8b == _T_311[9:0] ? 4'h1 : _GEN_14157; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14159 = 10'h8c == _T_311[9:0] ? 4'h1 : _GEN_14158; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14160 = 10'h8d == _T_311[9:0] ? 4'h1 : _GEN_14159; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14161 = 10'h8e == _T_311[9:0] ? 4'h1 : _GEN_14160; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14162 = 10'h8f == _T_311[9:0] ? 4'h1 : _GEN_14161; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14163 = 10'h90 == _T_311[9:0] ? 4'h1 : _GEN_14162; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14164 = 10'h91 == _T_311[9:0] ? 4'h1 : _GEN_14163; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14165 = 10'h92 == _T_311[9:0] ? 4'h1 : _GEN_14164; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14166 = 10'h93 == _T_311[9:0] ? 4'h0 : _GEN_14165; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14167 = 10'h94 == _T_311[9:0] ? 4'h0 : _GEN_14166; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14168 = 10'h95 == _T_311[9:0] ? 4'ha : _GEN_14167; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14169 = 10'h96 == _T_311[9:0] ? 4'ha : _GEN_14168; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14170 = 10'h97 == _T_311[9:0] ? 4'ha : _GEN_14169; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14171 = 10'h98 == _T_311[9:0] ? 4'h1 : _GEN_14170; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14172 = 10'h99 == _T_311[9:0] ? 4'h0 : _GEN_14171; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14173 = 10'h9a == _T_311[9:0] ? 4'h1 : _GEN_14172; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14174 = 10'h9b == _T_311[9:0] ? 4'h1 : _GEN_14173; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14175 = 10'h9c == _T_311[9:0] ? 4'ha : _GEN_14174; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14176 = 10'h9d == _T_311[9:0] ? 4'ha : _GEN_14175; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14177 = 10'h9e == _T_311[9:0] ? 4'h3 : _GEN_14176; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14178 = 10'h9f == _T_311[9:0] ? 4'h0 : _GEN_14177; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14179 = 10'ha0 == _T_311[9:0] ? 4'ha : _GEN_14178; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14180 = 10'ha1 == _T_311[9:0] ? 4'h1 : _GEN_14179; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14181 = 10'ha2 == _T_311[9:0] ? 4'h0 : _GEN_14180; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14182 = 10'ha3 == _T_311[9:0] ? 4'h3 : _GEN_14181; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14183 = 10'ha4 == _T_311[9:0] ? 4'ha : _GEN_14182; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14184 = 10'ha5 == _T_311[9:0] ? 4'ha : _GEN_14183; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14185 = 10'ha6 == _T_311[9:0] ? 4'ha : _GEN_14184; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14186 = 10'ha7 == _T_311[9:0] ? 4'h0 : _GEN_14185; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14187 = 10'ha8 == _T_311[9:0] ? 4'ha : _GEN_14186; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14188 = 10'ha9 == _T_311[9:0] ? 4'h1 : _GEN_14187; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14189 = 10'haa == _T_311[9:0] ? 4'h0 : _GEN_14188; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14190 = 10'hab == _T_311[9:0] ? 4'h0 : _GEN_14189; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14191 = 10'hac == _T_311[9:0] ? 4'h0 : _GEN_14190; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14192 = 10'had == _T_311[9:0] ? 4'h0 : _GEN_14191; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14193 = 10'hae == _T_311[9:0] ? 4'h0 : _GEN_14192; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14194 = 10'haf == _T_311[9:0] ? 4'h0 : _GEN_14193; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14195 = 10'hb0 == _T_311[9:0] ? 4'h0 : _GEN_14194; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14196 = 10'hb1 == _T_311[9:0] ? 4'h0 : _GEN_14195; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14197 = 10'hb2 == _T_311[9:0] ? 4'h0 : _GEN_14196; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14198 = 10'hb3 == _T_311[9:0] ? 4'h0 : _GEN_14197; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14199 = 10'hb4 == _T_311[9:0] ? 4'h1 : _GEN_14198; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14200 = 10'hb5 == _T_311[9:0] ? 4'h1 : _GEN_14199; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14201 = 10'hb6 == _T_311[9:0] ? 4'ha : _GEN_14200; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14202 = 10'hb7 == _T_311[9:0] ? 4'h0 : _GEN_14201; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14203 = 10'hb8 == _T_311[9:0] ? 4'ha : _GEN_14202; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14204 = 10'hb9 == _T_311[9:0] ? 4'ha : _GEN_14203; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14205 = 10'hba == _T_311[9:0] ? 4'ha : _GEN_14204; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14206 = 10'hbb == _T_311[9:0] ? 4'h0 : _GEN_14205; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14207 = 10'hbc == _T_311[9:0] ? 4'ha : _GEN_14206; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14208 = 10'hbd == _T_311[9:0] ? 4'ha : _GEN_14207; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14209 = 10'hbe == _T_311[9:0] ? 4'h3 : _GEN_14208; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14210 = 10'hbf == _T_311[9:0] ? 4'h0 : _GEN_14209; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14211 = 10'hc0 == _T_311[9:0] ? 4'ha : _GEN_14210; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14212 = 10'hc1 == _T_311[9:0] ? 4'ha : _GEN_14211; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14213 = 10'hc2 == _T_311[9:0] ? 4'h3 : _GEN_14212; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14214 = 10'hc3 == _T_311[9:0] ? 4'h2 : _GEN_14213; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14215 = 10'hc4 == _T_311[9:0] ? 4'h0 : _GEN_14214; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14216 = 10'hc5 == _T_311[9:0] ? 4'h0 : _GEN_14215; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14217 = 10'hc6 == _T_311[9:0] ? 4'h0 : _GEN_14216; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14218 = 10'hc7 == _T_311[9:0] ? 4'ha : _GEN_14217; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14219 = 10'hc8 == _T_311[9:0] ? 4'h1 : _GEN_14218; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14220 = 10'hc9 == _T_311[9:0] ? 4'h0 : _GEN_14219; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14221 = 10'hca == _T_311[9:0] ? 4'h0 : _GEN_14220; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14222 = 10'hcb == _T_311[9:0] ? 4'h0 : _GEN_14221; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14223 = 10'hcc == _T_311[9:0] ? 4'h0 : _GEN_14222; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14224 = 10'hcd == _T_311[9:0] ? 4'h0 : _GEN_14223; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14225 = 10'hce == _T_311[9:0] ? 4'h0 : _GEN_14224; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14226 = 10'hcf == _T_311[9:0] ? 4'h0 : _GEN_14225; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14227 = 10'hd0 == _T_311[9:0] ? 4'h0 : _GEN_14226; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14228 = 10'hd1 == _T_311[9:0] ? 4'h0 : _GEN_14227; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14229 = 10'hd2 == _T_311[9:0] ? 4'h0 : _GEN_14228; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14230 = 10'hd3 == _T_311[9:0] ? 4'h0 : _GEN_14229; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14231 = 10'hd4 == _T_311[9:0] ? 4'h0 : _GEN_14230; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14232 = 10'hd5 == _T_311[9:0] ? 4'h0 : _GEN_14231; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14233 = 10'hd6 == _T_311[9:0] ? 4'h1 : _GEN_14232; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14234 = 10'hd7 == _T_311[9:0] ? 4'ha : _GEN_14233; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14235 = 10'hd8 == _T_311[9:0] ? 4'h0 : _GEN_14234; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14236 = 10'hd9 == _T_311[9:0] ? 4'ha : _GEN_14235; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14237 = 10'hda == _T_311[9:0] ? 4'ha : _GEN_14236; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14238 = 10'hdb == _T_311[9:0] ? 4'ha : _GEN_14237; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14239 = 10'hdc == _T_311[9:0] ? 4'ha : _GEN_14238; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14240 = 10'hdd == _T_311[9:0] ? 4'h3 : _GEN_14239; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14241 = 10'hde == _T_311[9:0] ? 4'h2 : _GEN_14240; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14242 = 10'hdf == _T_311[9:0] ? 4'h0 : _GEN_14241; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14243 = 10'he0 == _T_311[9:0] ? 4'ha : _GEN_14242; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14244 = 10'he1 == _T_311[9:0] ? 4'ha : _GEN_14243; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14245 = 10'he2 == _T_311[9:0] ? 4'h3 : _GEN_14244; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14246 = 10'he3 == _T_311[9:0] ? 4'ha : _GEN_14245; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14247 = 10'he4 == _T_311[9:0] ? 4'ha : _GEN_14246; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14248 = 10'he5 == _T_311[9:0] ? 4'ha : _GEN_14247; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14249 = 10'he6 == _T_311[9:0] ? 4'ha : _GEN_14248; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14250 = 10'he7 == _T_311[9:0] ? 4'h1 : _GEN_14249; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14251 = 10'he8 == _T_311[9:0] ? 4'h1 : _GEN_14250; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14252 = 10'he9 == _T_311[9:0] ? 4'h1 : _GEN_14251; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14253 = 10'hea == _T_311[9:0] ? 4'h0 : _GEN_14252; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14254 = 10'heb == _T_311[9:0] ? 4'h0 : _GEN_14253; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14255 = 10'hec == _T_311[9:0] ? 4'h0 : _GEN_14254; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14256 = 10'hed == _T_311[9:0] ? 4'h0 : _GEN_14255; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14257 = 10'hee == _T_311[9:0] ? 4'h0 : _GEN_14256; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14258 = 10'hef == _T_311[9:0] ? 4'h0 : _GEN_14257; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14259 = 10'hf0 == _T_311[9:0] ? 4'h0 : _GEN_14258; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14260 = 10'hf1 == _T_311[9:0] ? 4'h0 : _GEN_14259; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14261 = 10'hf2 == _T_311[9:0] ? 4'h0 : _GEN_14260; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14262 = 10'hf3 == _T_311[9:0] ? 4'h0 : _GEN_14261; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14263 = 10'hf4 == _T_311[9:0] ? 4'h0 : _GEN_14262; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14264 = 10'hf5 == _T_311[9:0] ? 4'h1 : _GEN_14263; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14265 = 10'hf6 == _T_311[9:0] ? 4'h0 : _GEN_14264; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14266 = 10'hf7 == _T_311[9:0] ? 4'h0 : _GEN_14265; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14267 = 10'hf8 == _T_311[9:0] ? 4'h1 : _GEN_14266; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14268 = 10'hf9 == _T_311[9:0] ? 4'h0 : _GEN_14267; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14269 = 10'hfa == _T_311[9:0] ? 4'ha : _GEN_14268; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14270 = 10'hfb == _T_311[9:0] ? 4'ha : _GEN_14269; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14271 = 10'hfc == _T_311[9:0] ? 4'ha : _GEN_14270; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14272 = 10'hfd == _T_311[9:0] ? 4'h3 : _GEN_14271; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14273 = 10'hfe == _T_311[9:0] ? 4'ha : _GEN_14272; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14274 = 10'hff == _T_311[9:0] ? 4'h0 : _GEN_14273; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14275 = 10'h100 == _T_311[9:0] ? 4'ha : _GEN_14274; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14276 = 10'h101 == _T_311[9:0] ? 4'h0 : _GEN_14275; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14277 = 10'h102 == _T_311[9:0] ? 4'h3 : _GEN_14276; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14278 = 10'h103 == _T_311[9:0] ? 4'ha : _GEN_14277; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14279 = 10'h104 == _T_311[9:0] ? 4'ha : _GEN_14278; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14280 = 10'h105 == _T_311[9:0] ? 4'ha : _GEN_14279; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14281 = 10'h106 == _T_311[9:0] ? 4'ha : _GEN_14280; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14282 = 10'h107 == _T_311[9:0] ? 4'ha : _GEN_14281; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14283 = 10'h108 == _T_311[9:0] ? 4'h1 : _GEN_14282; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14284 = 10'h109 == _T_311[9:0] ? 4'h0 : _GEN_14283; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14285 = 10'h10a == _T_311[9:0] ? 4'h0 : _GEN_14284; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14286 = 10'h10b == _T_311[9:0] ? 4'h0 : _GEN_14285; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14287 = 10'h10c == _T_311[9:0] ? 4'h0 : _GEN_14286; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14288 = 10'h10d == _T_311[9:0] ? 4'h0 : _GEN_14287; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14289 = 10'h10e == _T_311[9:0] ? 4'h0 : _GEN_14288; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14290 = 10'h10f == _T_311[9:0] ? 4'h0 : _GEN_14289; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14291 = 10'h110 == _T_311[9:0] ? 4'h0 : _GEN_14290; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14292 = 10'h111 == _T_311[9:0] ? 4'h0 : _GEN_14291; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14293 = 10'h112 == _T_311[9:0] ? 4'h0 : _GEN_14292; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14294 = 10'h113 == _T_311[9:0] ? 4'h0 : _GEN_14293; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14295 = 10'h114 == _T_311[9:0] ? 4'h0 : _GEN_14294; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14296 = 10'h115 == _T_311[9:0] ? 4'h0 : _GEN_14295; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14297 = 10'h116 == _T_311[9:0] ? 4'h1 : _GEN_14296; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14298 = 10'h117 == _T_311[9:0] ? 4'ha : _GEN_14297; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14299 = 10'h118 == _T_311[9:0] ? 4'ha : _GEN_14298; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14300 = 10'h119 == _T_311[9:0] ? 4'ha : _GEN_14299; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14301 = 10'h11a == _T_311[9:0] ? 4'h0 : _GEN_14300; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14302 = 10'h11b == _T_311[9:0] ? 4'ha : _GEN_14301; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14303 = 10'h11c == _T_311[9:0] ? 4'ha : _GEN_14302; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14304 = 10'h11d == _T_311[9:0] ? 4'h2 : _GEN_14303; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14305 = 10'h11e == _T_311[9:0] ? 4'h3 : _GEN_14304; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14306 = 10'h11f == _T_311[9:0] ? 4'h0 : _GEN_14305; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14307 = 10'h120 == _T_311[9:0] ? 4'ha : _GEN_14306; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14308 = 10'h121 == _T_311[9:0] ? 4'ha : _GEN_14307; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14309 = 10'h122 == _T_311[9:0] ? 4'h3 : _GEN_14308; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14310 = 10'h123 == _T_311[9:0] ? 4'ha : _GEN_14309; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14311 = 10'h124 == _T_311[9:0] ? 4'ha : _GEN_14310; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14312 = 10'h125 == _T_311[9:0] ? 4'ha : _GEN_14311; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14313 = 10'h126 == _T_311[9:0] ? 4'ha : _GEN_14312; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14314 = 10'h127 == _T_311[9:0] ? 4'h1 : _GEN_14313; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14315 = 10'h128 == _T_311[9:0] ? 4'h0 : _GEN_14314; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14316 = 10'h129 == _T_311[9:0] ? 4'ha : _GEN_14315; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14317 = 10'h12a == _T_311[9:0] ? 4'ha : _GEN_14316; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14318 = 10'h12b == _T_311[9:0] ? 4'h0 : _GEN_14317; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14319 = 10'h12c == _T_311[9:0] ? 4'h0 : _GEN_14318; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14320 = 10'h12d == _T_311[9:0] ? 4'h0 : _GEN_14319; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14321 = 10'h12e == _T_311[9:0] ? 4'h0 : _GEN_14320; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14322 = 10'h12f == _T_311[9:0] ? 4'h0 : _GEN_14321; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14323 = 10'h130 == _T_311[9:0] ? 4'h0 : _GEN_14322; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14324 = 10'h131 == _T_311[9:0] ? 4'h0 : _GEN_14323; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14325 = 10'h132 == _T_311[9:0] ? 4'h0 : _GEN_14324; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14326 = 10'h133 == _T_311[9:0] ? 4'h0 : _GEN_14325; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14327 = 10'h134 == _T_311[9:0] ? 4'ha : _GEN_14326; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14328 = 10'h135 == _T_311[9:0] ? 4'ha : _GEN_14327; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14329 = 10'h136 == _T_311[9:0] ? 4'h0 : _GEN_14328; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14330 = 10'h137 == _T_311[9:0] ? 4'h1 : _GEN_14329; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14331 = 10'h138 == _T_311[9:0] ? 4'ha : _GEN_14330; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14332 = 10'h139 == _T_311[9:0] ? 4'ha : _GEN_14331; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14333 = 10'h13a == _T_311[9:0] ? 4'ha : _GEN_14332; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14334 = 10'h13b == _T_311[9:0] ? 4'ha : _GEN_14333; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14335 = 10'h13c == _T_311[9:0] ? 4'ha : _GEN_14334; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14336 = 10'h13d == _T_311[9:0] ? 4'ha : _GEN_14335; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14337 = 10'h13e == _T_311[9:0] ? 4'h3 : _GEN_14336; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14338 = 10'h13f == _T_311[9:0] ? 4'h0 : _GEN_14337; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14339 = 10'h140 == _T_311[9:0] ? 4'ha : _GEN_14338; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14340 = 10'h141 == _T_311[9:0] ? 4'ha : _GEN_14339; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14341 = 10'h142 == _T_311[9:0] ? 4'h2 : _GEN_14340; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14342 = 10'h143 == _T_311[9:0] ? 4'h3 : _GEN_14341; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14343 = 10'h144 == _T_311[9:0] ? 4'ha : _GEN_14342; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14344 = 10'h145 == _T_311[9:0] ? 4'ha : _GEN_14343; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14345 = 10'h146 == _T_311[9:0] ? 4'h1 : _GEN_14344; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14346 = 10'h147 == _T_311[9:0] ? 4'h0 : _GEN_14345; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14347 = 10'h148 == _T_311[9:0] ? 4'ha : _GEN_14346; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14348 = 10'h149 == _T_311[9:0] ? 4'ha : _GEN_14347; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14349 = 10'h14a == _T_311[9:0] ? 4'ha : _GEN_14348; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14350 = 10'h14b == _T_311[9:0] ? 4'ha : _GEN_14349; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14351 = 10'h14c == _T_311[9:0] ? 4'ha : _GEN_14350; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14352 = 10'h14d == _T_311[9:0] ? 4'ha : _GEN_14351; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14353 = 10'h14e == _T_311[9:0] ? 4'ha : _GEN_14352; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14354 = 10'h14f == _T_311[9:0] ? 4'ha : _GEN_14353; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14355 = 10'h150 == _T_311[9:0] ? 4'ha : _GEN_14354; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14356 = 10'h151 == _T_311[9:0] ? 4'ha : _GEN_14355; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14357 = 10'h152 == _T_311[9:0] ? 4'ha : _GEN_14356; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14358 = 10'h153 == _T_311[9:0] ? 4'ha : _GEN_14357; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14359 = 10'h154 == _T_311[9:0] ? 4'ha : _GEN_14358; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14360 = 10'h155 == _T_311[9:0] ? 4'ha : _GEN_14359; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14361 = 10'h156 == _T_311[9:0] ? 4'ha : _GEN_14360; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14362 = 10'h157 == _T_311[9:0] ? 4'h0 : _GEN_14361; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14363 = 10'h158 == _T_311[9:0] ? 4'ha : _GEN_14362; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14364 = 10'h159 == _T_311[9:0] ? 4'ha : _GEN_14363; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14365 = 10'h15a == _T_311[9:0] ? 4'ha : _GEN_14364; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14366 = 10'h15b == _T_311[9:0] ? 4'ha : _GEN_14365; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14367 = 10'h15c == _T_311[9:0] ? 4'ha : _GEN_14366; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14368 = 10'h15d == _T_311[9:0] ? 4'h3 : _GEN_14367; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14369 = 10'h15e == _T_311[9:0] ? 4'h2 : _GEN_14368; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14370 = 10'h15f == _T_311[9:0] ? 4'h0 : _GEN_14369; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14371 = 10'h160 == _T_311[9:0] ? 4'ha : _GEN_14370; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14372 = 10'h161 == _T_311[9:0] ? 4'ha : _GEN_14371; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14373 = 10'h162 == _T_311[9:0] ? 4'ha : _GEN_14372; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14374 = 10'h163 == _T_311[9:0] ? 4'h2 : _GEN_14373; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14375 = 10'h164 == _T_311[9:0] ? 4'h3 : _GEN_14374; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14376 = 10'h165 == _T_311[9:0] ? 4'h1 : _GEN_14375; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14377 = 10'h166 == _T_311[9:0] ? 4'h0 : _GEN_14376; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14378 = 10'h167 == _T_311[9:0] ? 4'h0 : _GEN_14377; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14379 = 10'h168 == _T_311[9:0] ? 4'h5 : _GEN_14378; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14380 = 10'h169 == _T_311[9:0] ? 4'h3 : _GEN_14379; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14381 = 10'h16a == _T_311[9:0] ? 4'h5 : _GEN_14380; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14382 = 10'h16b == _T_311[9:0] ? 4'h5 : _GEN_14381; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14383 = 10'h16c == _T_311[9:0] ? 4'ha : _GEN_14382; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14384 = 10'h16d == _T_311[9:0] ? 4'ha : _GEN_14383; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14385 = 10'h16e == _T_311[9:0] ? 4'ha : _GEN_14384; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14386 = 10'h16f == _T_311[9:0] ? 4'ha : _GEN_14385; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14387 = 10'h170 == _T_311[9:0] ? 4'ha : _GEN_14386; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14388 = 10'h171 == _T_311[9:0] ? 4'ha : _GEN_14387; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14389 = 10'h172 == _T_311[9:0] ? 4'ha : _GEN_14388; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14390 = 10'h173 == _T_311[9:0] ? 4'ha : _GEN_14389; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14391 = 10'h174 == _T_311[9:0] ? 4'ha : _GEN_14390; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14392 = 10'h175 == _T_311[9:0] ? 4'ha : _GEN_14391; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14393 = 10'h176 == _T_311[9:0] ? 4'h0 : _GEN_14392; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14394 = 10'h177 == _T_311[9:0] ? 4'h0 : _GEN_14393; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14395 = 10'h178 == _T_311[9:0] ? 4'h1 : _GEN_14394; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14396 = 10'h179 == _T_311[9:0] ? 4'ha : _GEN_14395; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14397 = 10'h17a == _T_311[9:0] ? 4'ha : _GEN_14396; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14398 = 10'h17b == _T_311[9:0] ? 4'ha : _GEN_14397; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14399 = 10'h17c == _T_311[9:0] ? 4'h3 : _GEN_14398; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14400 = 10'h17d == _T_311[9:0] ? 4'h2 : _GEN_14399; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14401 = 10'h17e == _T_311[9:0] ? 4'ha : _GEN_14400; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14402 = 10'h17f == _T_311[9:0] ? 4'h0 : _GEN_14401; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14403 = 10'h180 == _T_311[9:0] ? 4'h5 : _GEN_14402; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14404 = 10'h181 == _T_311[9:0] ? 4'h5 : _GEN_14403; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14405 = 10'h182 == _T_311[9:0] ? 4'h5 : _GEN_14404; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14406 = 10'h183 == _T_311[9:0] ? 4'h5 : _GEN_14405; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14407 = 10'h184 == _T_311[9:0] ? 4'h3 : _GEN_14406; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14408 = 10'h185 == _T_311[9:0] ? 4'h1 : _GEN_14407; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14409 = 10'h186 == _T_311[9:0] ? 4'hb : _GEN_14408; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14410 = 10'h187 == _T_311[9:0] ? 4'h0 : _GEN_14409; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14411 = 10'h188 == _T_311[9:0] ? 4'h5 : _GEN_14410; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14412 = 10'h189 == _T_311[9:0] ? 4'h5 : _GEN_14411; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14413 = 10'h18a == _T_311[9:0] ? 4'h5 : _GEN_14412; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14414 = 10'h18b == _T_311[9:0] ? 4'h5 : _GEN_14413; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14415 = 10'h18c == _T_311[9:0] ? 4'h5 : _GEN_14414; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14416 = 10'h18d == _T_311[9:0] ? 4'h5 : _GEN_14415; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14417 = 10'h18e == _T_311[9:0] ? 4'h5 : _GEN_14416; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14418 = 10'h18f == _T_311[9:0] ? 4'h5 : _GEN_14417; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14419 = 10'h190 == _T_311[9:0] ? 4'h5 : _GEN_14418; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14420 = 10'h191 == _T_311[9:0] ? 4'h5 : _GEN_14419; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14421 = 10'h192 == _T_311[9:0] ? 4'h3 : _GEN_14420; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14422 = 10'h193 == _T_311[9:0] ? 4'h5 : _GEN_14421; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14423 = 10'h194 == _T_311[9:0] ? 4'h5 : _GEN_14422; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14424 = 10'h195 == _T_311[9:0] ? 4'h5 : _GEN_14423; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14425 = 10'h196 == _T_311[9:0] ? 4'h0 : _GEN_14424; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14426 = 10'h197 == _T_311[9:0] ? 4'ha : _GEN_14425; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14427 = 10'h198 == _T_311[9:0] ? 4'h1 : _GEN_14426; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14428 = 10'h199 == _T_311[9:0] ? 4'ha : _GEN_14427; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14429 = 10'h19a == _T_311[9:0] ? 4'ha : _GEN_14428; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14430 = 10'h19b == _T_311[9:0] ? 4'ha : _GEN_14429; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14431 = 10'h19c == _T_311[9:0] ? 4'h3 : _GEN_14430; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14432 = 10'h19d == _T_311[9:0] ? 4'ha : _GEN_14431; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14433 = 10'h19e == _T_311[9:0] ? 4'ha : _GEN_14432; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14434 = 10'h19f == _T_311[9:0] ? 4'h0 : _GEN_14433; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14435 = 10'h1a0 == _T_311[9:0] ? 4'h5 : _GEN_14434; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14436 = 10'h1a1 == _T_311[9:0] ? 4'h5 : _GEN_14435; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14437 = 10'h1a2 == _T_311[9:0] ? 4'h3 : _GEN_14436; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14438 = 10'h1a3 == _T_311[9:0] ? 4'h5 : _GEN_14437; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14439 = 10'h1a4 == _T_311[9:0] ? 4'h3 : _GEN_14438; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14440 = 10'h1a5 == _T_311[9:0] ? 4'h0 : _GEN_14439; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14441 = 10'h1a6 == _T_311[9:0] ? 4'h5 : _GEN_14440; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14442 = 10'h1a7 == _T_311[9:0] ? 4'h0 : _GEN_14441; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14443 = 10'h1a8 == _T_311[9:0] ? 4'hb : _GEN_14442; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14444 = 10'h1a9 == _T_311[9:0] ? 4'h5 : _GEN_14443; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14445 = 10'h1aa == _T_311[9:0] ? 4'h5 : _GEN_14444; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14446 = 10'h1ab == _T_311[9:0] ? 4'h3 : _GEN_14445; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14447 = 10'h1ac == _T_311[9:0] ? 4'h5 : _GEN_14446; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14448 = 10'h1ad == _T_311[9:0] ? 4'h5 : _GEN_14447; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14449 = 10'h1ae == _T_311[9:0] ? 4'h5 : _GEN_14448; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14450 = 10'h1af == _T_311[9:0] ? 4'h5 : _GEN_14449; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14451 = 10'h1b0 == _T_311[9:0] ? 4'h5 : _GEN_14450; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14452 = 10'h1b1 == _T_311[9:0] ? 4'h5 : _GEN_14451; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14453 = 10'h1b2 == _T_311[9:0] ? 4'h5 : _GEN_14452; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14454 = 10'h1b3 == _T_311[9:0] ? 4'h5 : _GEN_14453; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14455 = 10'h1b4 == _T_311[9:0] ? 4'h5 : _GEN_14454; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14456 = 10'h1b5 == _T_311[9:0] ? 4'h5 : _GEN_14455; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14457 = 10'h1b6 == _T_311[9:0] ? 4'h0 : _GEN_14456; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14458 = 10'h1b7 == _T_311[9:0] ? 4'h5 : _GEN_14457; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14459 = 10'h1b8 == _T_311[9:0] ? 4'h0 : _GEN_14458; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14460 = 10'h1b9 == _T_311[9:0] ? 4'h5 : _GEN_14459; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14461 = 10'h1ba == _T_311[9:0] ? 4'h5 : _GEN_14460; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14462 = 10'h1bb == _T_311[9:0] ? 4'h5 : _GEN_14461; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14463 = 10'h1bc == _T_311[9:0] ? 4'h2 : _GEN_14462; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14464 = 10'h1bd == _T_311[9:0] ? 4'h3 : _GEN_14463; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14465 = 10'h1be == _T_311[9:0] ? 4'h5 : _GEN_14464; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14466 = 10'h1bf == _T_311[9:0] ? 4'h0 : _GEN_14465; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14467 = 10'h1c0 == _T_311[9:0] ? 4'h5 : _GEN_14466; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14468 = 10'h1c1 == _T_311[9:0] ? 4'h5 : _GEN_14467; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14469 = 10'h1c2 == _T_311[9:0] ? 4'h5 : _GEN_14468; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14470 = 10'h1c3 == _T_311[9:0] ? 4'h2 : _GEN_14469; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14471 = 10'h1c4 == _T_311[9:0] ? 4'h2 : _GEN_14470; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14472 = 10'h1c5 == _T_311[9:0] ? 4'h5 : _GEN_14471; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14473 = 10'h1c6 == _T_311[9:0] ? 4'h5 : _GEN_14472; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14474 = 10'h1c7 == _T_311[9:0] ? 4'h5 : _GEN_14473; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14475 = 10'h1c8 == _T_311[9:0] ? 4'h5 : _GEN_14474; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14476 = 10'h1c9 == _T_311[9:0] ? 4'hb : _GEN_14475; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14477 = 10'h1ca == _T_311[9:0] ? 4'hb : _GEN_14476; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14478 = 10'h1cb == _T_311[9:0] ? 4'hb : _GEN_14477; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14479 = 10'h1cc == _T_311[9:0] ? 4'hb : _GEN_14478; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14480 = 10'h1cd == _T_311[9:0] ? 4'hb : _GEN_14479; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14481 = 10'h1ce == _T_311[9:0] ? 4'hb : _GEN_14480; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14482 = 10'h1cf == _T_311[9:0] ? 4'hb : _GEN_14481; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14483 = 10'h1d0 == _T_311[9:0] ? 4'hb : _GEN_14482; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14484 = 10'h1d1 == _T_311[9:0] ? 4'hb : _GEN_14483; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14485 = 10'h1d2 == _T_311[9:0] ? 4'hb : _GEN_14484; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14486 = 10'h1d3 == _T_311[9:0] ? 4'hb : _GEN_14485; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14487 = 10'h1d4 == _T_311[9:0] ? 4'hb : _GEN_14486; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14488 = 10'h1d5 == _T_311[9:0] ? 4'hb : _GEN_14487; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14489 = 10'h1d6 == _T_311[9:0] ? 4'h5 : _GEN_14488; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14490 = 10'h1d7 == _T_311[9:0] ? 4'h5 : _GEN_14489; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14491 = 10'h1d8 == _T_311[9:0] ? 4'h5 : _GEN_14490; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14492 = 10'h1d9 == _T_311[9:0] ? 4'h5 : _GEN_14491; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14493 = 10'h1da == _T_311[9:0] ? 4'h5 : _GEN_14492; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14494 = 10'h1db == _T_311[9:0] ? 4'h5 : _GEN_14493; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14495 = 10'h1dc == _T_311[9:0] ? 4'h5 : _GEN_14494; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14496 = 10'h1dd == _T_311[9:0] ? 4'h3 : _GEN_14495; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14497 = 10'h1de == _T_311[9:0] ? 4'h5 : _GEN_14496; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14498 = 10'h1df == _T_311[9:0] ? 4'h0 : _GEN_14497; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14499 = 10'h1e0 == _T_311[9:0] ? 4'h3 : _GEN_14498; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14500 = 10'h1e1 == _T_311[9:0] ? 4'h5 : _GEN_14499; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14501 = 10'h1e2 == _T_311[9:0] ? 4'h2 : _GEN_14500; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14502 = 10'h1e3 == _T_311[9:0] ? 4'h2 : _GEN_14501; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14503 = 10'h1e4 == _T_311[9:0] ? 4'h5 : _GEN_14502; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14504 = 10'h1e5 == _T_311[9:0] ? 4'h5 : _GEN_14503; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14505 = 10'h1e6 == _T_311[9:0] ? 4'h5 : _GEN_14504; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14506 = 10'h1e7 == _T_311[9:0] ? 4'h5 : _GEN_14505; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14507 = 10'h1e8 == _T_311[9:0] ? 4'hb : _GEN_14506; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14508 = 10'h1e9 == _T_311[9:0] ? 4'h5 : _GEN_14507; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14509 = 10'h1ea == _T_311[9:0] ? 4'h5 : _GEN_14508; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14510 = 10'h1eb == _T_311[9:0] ? 4'hb : _GEN_14509; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14511 = 10'h1ec == _T_311[9:0] ? 4'h5 : _GEN_14510; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14512 = 10'h1ed == _T_311[9:0] ? 4'hb : _GEN_14511; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14513 = 10'h1ee == _T_311[9:0] ? 4'h5 : _GEN_14512; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14514 = 10'h1ef == _T_311[9:0] ? 4'hb : _GEN_14513; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14515 = 10'h1f0 == _T_311[9:0] ? 4'h5 : _GEN_14514; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14516 = 10'h1f1 == _T_311[9:0] ? 4'hb : _GEN_14515; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14517 = 10'h1f2 == _T_311[9:0] ? 4'hb : _GEN_14516; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14518 = 10'h1f3 == _T_311[9:0] ? 4'h5 : _GEN_14517; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14519 = 10'h1f4 == _T_311[9:0] ? 4'hb : _GEN_14518; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14520 = 10'h1f5 == _T_311[9:0] ? 4'hb : _GEN_14519; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14521 = 10'h1f6 == _T_311[9:0] ? 4'h5 : _GEN_14520; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14522 = 10'h1f7 == _T_311[9:0] ? 4'h5 : _GEN_14521; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14523 = 10'h1f8 == _T_311[9:0] ? 4'h5 : _GEN_14522; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14524 = 10'h1f9 == _T_311[9:0] ? 4'h5 : _GEN_14523; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14525 = 10'h1fa == _T_311[9:0] ? 4'h3 : _GEN_14524; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14526 = 10'h1fb == _T_311[9:0] ? 4'h5 : _GEN_14525; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14527 = 10'h1fc == _T_311[9:0] ? 4'h5 : _GEN_14526; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14528 = 10'h1fd == _T_311[9:0] ? 4'h2 : _GEN_14527; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14529 = 10'h1fe == _T_311[9:0] ? 4'h5 : _GEN_14528; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14530 = 10'h1ff == _T_311[9:0] ? 4'h0 : _GEN_14529; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14531 = 10'h200 == _T_311[9:0] ? 4'h5 : _GEN_14530; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14532 = 10'h201 == _T_311[9:0] ? 4'h5 : _GEN_14531; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14533 = 10'h202 == _T_311[9:0] ? 4'h3 : _GEN_14532; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14534 = 10'h203 == _T_311[9:0] ? 4'h5 : _GEN_14533; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14535 = 10'h204 == _T_311[9:0] ? 4'h5 : _GEN_14534; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14536 = 10'h205 == _T_311[9:0] ? 4'h5 : _GEN_14535; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14537 = 10'h206 == _T_311[9:0] ? 4'hb : _GEN_14536; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14538 = 10'h207 == _T_311[9:0] ? 4'hb : _GEN_14537; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14539 = 10'h208 == _T_311[9:0] ? 4'h5 : _GEN_14538; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14540 = 10'h209 == _T_311[9:0] ? 4'h5 : _GEN_14539; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14541 = 10'h20a == _T_311[9:0] ? 4'h5 : _GEN_14540; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14542 = 10'h20b == _T_311[9:0] ? 4'hb : _GEN_14541; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14543 = 10'h20c == _T_311[9:0] ? 4'h5 : _GEN_14542; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14544 = 10'h20d == _T_311[9:0] ? 4'hb : _GEN_14543; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14545 = 10'h20e == _T_311[9:0] ? 4'h5 : _GEN_14544; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14546 = 10'h20f == _T_311[9:0] ? 4'hb : _GEN_14545; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14547 = 10'h210 == _T_311[9:0] ? 4'h5 : _GEN_14546; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14548 = 10'h211 == _T_311[9:0] ? 4'h5 : _GEN_14547; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14549 = 10'h212 == _T_311[9:0] ? 4'hb : _GEN_14548; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14550 = 10'h213 == _T_311[9:0] ? 4'hb : _GEN_14549; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14551 = 10'h214 == _T_311[9:0] ? 4'hb : _GEN_14550; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14552 = 10'h215 == _T_311[9:0] ? 4'h5 : _GEN_14551; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14553 = 10'h216 == _T_311[9:0] ? 4'h5 : _GEN_14552; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14554 = 10'h217 == _T_311[9:0] ? 4'h5 : _GEN_14553; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14555 = 10'h218 == _T_311[9:0] ? 4'h5 : _GEN_14554; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14556 = 10'h219 == _T_311[9:0] ? 4'h5 : _GEN_14555; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14557 = 10'h21a == _T_311[9:0] ? 4'h5 : _GEN_14556; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14558 = 10'h21b == _T_311[9:0] ? 4'h5 : _GEN_14557; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14559 = 10'h21c == _T_311[9:0] ? 4'h3 : _GEN_14558; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14560 = 10'h21d == _T_311[9:0] ? 4'h2 : _GEN_14559; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14561 = 10'h21e == _T_311[9:0] ? 4'h5 : _GEN_14560; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14562 = 10'h21f == _T_311[9:0] ? 4'h0 : _GEN_14561; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14563 = 10'h220 == _T_311[9:0] ? 4'h0 : _GEN_14562; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14564 = 10'h221 == _T_311[9:0] ? 4'h0 : _GEN_14563; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14565 = 10'h222 == _T_311[9:0] ? 4'h0 : _GEN_14564; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14566 = 10'h223 == _T_311[9:0] ? 4'h0 : _GEN_14565; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14567 = 10'h224 == _T_311[9:0] ? 4'h0 : _GEN_14566; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14568 = 10'h225 == _T_311[9:0] ? 4'h0 : _GEN_14567; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14569 = 10'h226 == _T_311[9:0] ? 4'h0 : _GEN_14568; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14570 = 10'h227 == _T_311[9:0] ? 4'h0 : _GEN_14569; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14571 = 10'h228 == _T_311[9:0] ? 4'h0 : _GEN_14570; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14572 = 10'h229 == _T_311[9:0] ? 4'h0 : _GEN_14571; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14573 = 10'h22a == _T_311[9:0] ? 4'h0 : _GEN_14572; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14574 = 10'h22b == _T_311[9:0] ? 4'h0 : _GEN_14573; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14575 = 10'h22c == _T_311[9:0] ? 4'h0 : _GEN_14574; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14576 = 10'h22d == _T_311[9:0] ? 4'h0 : _GEN_14575; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14577 = 10'h22e == _T_311[9:0] ? 4'h0 : _GEN_14576; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14578 = 10'h22f == _T_311[9:0] ? 4'h0 : _GEN_14577; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14579 = 10'h230 == _T_311[9:0] ? 4'h0 : _GEN_14578; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14580 = 10'h231 == _T_311[9:0] ? 4'h0 : _GEN_14579; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14581 = 10'h232 == _T_311[9:0] ? 4'h0 : _GEN_14580; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14582 = 10'h233 == _T_311[9:0] ? 4'h0 : _GEN_14581; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14583 = 10'h234 == _T_311[9:0] ? 4'h0 : _GEN_14582; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14584 = 10'h235 == _T_311[9:0] ? 4'h0 : _GEN_14583; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14585 = 10'h236 == _T_311[9:0] ? 4'h0 : _GEN_14584; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14586 = 10'h237 == _T_311[9:0] ? 4'h0 : _GEN_14585; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14587 = 10'h238 == _T_311[9:0] ? 4'h0 : _GEN_14586; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14588 = 10'h239 == _T_311[9:0] ? 4'h0 : _GEN_14587; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14589 = 10'h23a == _T_311[9:0] ? 4'h0 : _GEN_14588; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14590 = 10'h23b == _T_311[9:0] ? 4'h0 : _GEN_14589; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14591 = 10'h23c == _T_311[9:0] ? 4'h0 : _GEN_14590; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14592 = 10'h23d == _T_311[9:0] ? 4'h0 : _GEN_14591; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14593 = 10'h23e == _T_311[9:0] ? 4'h0 : _GEN_14592; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14594 = 10'h23f == _T_311[9:0] ? 4'h0 : _GEN_14593; // @[Filter.scala 191:62]
  wire [4:0] _GEN_28346 = {{1'd0}, _GEN_14594}; // @[Filter.scala 191:62]
  wire [8:0] _T_313 = _GEN_28346 * 5'h14; // @[Filter.scala 191:62]
  wire [3:0] _GEN_14598 = 10'h3 == _T_311[9:0] ? 4'ha : 4'h3; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14599 = 10'h4 == _T_311[9:0] ? 4'h3 : _GEN_14598; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14600 = 10'h5 == _T_311[9:0] ? 4'h3 : _GEN_14599; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14601 = 10'h6 == _T_311[9:0] ? 4'h3 : _GEN_14600; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14602 = 10'h7 == _T_311[9:0] ? 4'h3 : _GEN_14601; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14603 = 10'h8 == _T_311[9:0] ? 4'h3 : _GEN_14602; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14604 = 10'h9 == _T_311[9:0] ? 4'h3 : _GEN_14603; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14605 = 10'ha == _T_311[9:0] ? 4'h3 : _GEN_14604; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14606 = 10'hb == _T_311[9:0] ? 4'h3 : _GEN_14605; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14607 = 10'hc == _T_311[9:0] ? 4'h5 : _GEN_14606; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14608 = 10'hd == _T_311[9:0] ? 4'h3 : _GEN_14607; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14609 = 10'he == _T_311[9:0] ? 4'h3 : _GEN_14608; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14610 = 10'hf == _T_311[9:0] ? 4'h3 : _GEN_14609; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14611 = 10'h10 == _T_311[9:0] ? 4'h3 : _GEN_14610; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14612 = 10'h11 == _T_311[9:0] ? 4'h3 : _GEN_14611; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14613 = 10'h12 == _T_311[9:0] ? 4'h3 : _GEN_14612; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14614 = 10'h13 == _T_311[9:0] ? 4'h3 : _GEN_14613; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14615 = 10'h14 == _T_311[9:0] ? 4'h3 : _GEN_14614; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14616 = 10'h15 == _T_311[9:0] ? 4'h3 : _GEN_14615; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14617 = 10'h16 == _T_311[9:0] ? 4'h3 : _GEN_14616; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14618 = 10'h17 == _T_311[9:0] ? 4'h3 : _GEN_14617; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14619 = 10'h18 == _T_311[9:0] ? 4'h3 : _GEN_14618; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14620 = 10'h19 == _T_311[9:0] ? 4'h3 : _GEN_14619; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14621 = 10'h1a == _T_311[9:0] ? 4'h3 : _GEN_14620; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14622 = 10'h1b == _T_311[9:0] ? 4'h3 : _GEN_14621; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14623 = 10'h1c == _T_311[9:0] ? 4'h3 : _GEN_14622; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14624 = 10'h1d == _T_311[9:0] ? 4'h3 : _GEN_14623; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14625 = 10'h1e == _T_311[9:0] ? 4'h3 : _GEN_14624; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14626 = 10'h1f == _T_311[9:0] ? 4'h0 : _GEN_14625; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14627 = 10'h20 == _T_311[9:0] ? 4'h3 : _GEN_14626; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14628 = 10'h21 == _T_311[9:0] ? 4'h5 : _GEN_14627; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14629 = 10'h22 == _T_311[9:0] ? 4'h3 : _GEN_14628; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14630 = 10'h23 == _T_311[9:0] ? 4'ha : _GEN_14629; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14631 = 10'h24 == _T_311[9:0] ? 4'h3 : _GEN_14630; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14632 = 10'h25 == _T_311[9:0] ? 4'h3 : _GEN_14631; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14633 = 10'h26 == _T_311[9:0] ? 4'h3 : _GEN_14632; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14634 = 10'h27 == _T_311[9:0] ? 4'h1 : _GEN_14633; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14635 = 10'h28 == _T_311[9:0] ? 4'h1 : _GEN_14634; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14636 = 10'h29 == _T_311[9:0] ? 4'h3 : _GEN_14635; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14637 = 10'h2a == _T_311[9:0] ? 4'h3 : _GEN_14636; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14638 = 10'h2b == _T_311[9:0] ? 4'h3 : _GEN_14637; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14639 = 10'h2c == _T_311[9:0] ? 4'h3 : _GEN_14638; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14640 = 10'h2d == _T_311[9:0] ? 4'h3 : _GEN_14639; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14641 = 10'h2e == _T_311[9:0] ? 4'h3 : _GEN_14640; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14642 = 10'h2f == _T_311[9:0] ? 4'h3 : _GEN_14641; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14643 = 10'h30 == _T_311[9:0] ? 4'h3 : _GEN_14642; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14644 = 10'h31 == _T_311[9:0] ? 4'h5 : _GEN_14643; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14645 = 10'h32 == _T_311[9:0] ? 4'h3 : _GEN_14644; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14646 = 10'h33 == _T_311[9:0] ? 4'h3 : _GEN_14645; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14647 = 10'h34 == _T_311[9:0] ? 4'h3 : _GEN_14646; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14648 = 10'h35 == _T_311[9:0] ? 4'h3 : _GEN_14647; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14649 = 10'h36 == _T_311[9:0] ? 4'h3 : _GEN_14648; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14650 = 10'h37 == _T_311[9:0] ? 4'h1 : _GEN_14649; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14651 = 10'h38 == _T_311[9:0] ? 4'h1 : _GEN_14650; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14652 = 10'h39 == _T_311[9:0] ? 4'h3 : _GEN_14651; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14653 = 10'h3a == _T_311[9:0] ? 4'h3 : _GEN_14652; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14654 = 10'h3b == _T_311[9:0] ? 4'h5 : _GEN_14653; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14655 = 10'h3c == _T_311[9:0] ? 4'h3 : _GEN_14654; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14656 = 10'h3d == _T_311[9:0] ? 4'ha : _GEN_14655; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14657 = 10'h3e == _T_311[9:0] ? 4'h3 : _GEN_14656; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14658 = 10'h3f == _T_311[9:0] ? 4'h0 : _GEN_14657; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14659 = 10'h40 == _T_311[9:0] ? 4'h3 : _GEN_14658; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14660 = 10'h41 == _T_311[9:0] ? 4'h3 : _GEN_14659; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14661 = 10'h42 == _T_311[9:0] ? 4'h3 : _GEN_14660; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14662 = 10'h43 == _T_311[9:0] ? 4'h7 : _GEN_14661; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14663 = 10'h44 == _T_311[9:0] ? 4'ha : _GEN_14662; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14664 = 10'h45 == _T_311[9:0] ? 4'h0 : _GEN_14663; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14665 = 10'h46 == _T_311[9:0] ? 4'h0 : _GEN_14664; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14666 = 10'h47 == _T_311[9:0] ? 4'h0 : _GEN_14665; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14667 = 10'h48 == _T_311[9:0] ? 4'h0 : _GEN_14666; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14668 = 10'h49 == _T_311[9:0] ? 4'h3 : _GEN_14667; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14669 = 10'h4a == _T_311[9:0] ? 4'h3 : _GEN_14668; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14670 = 10'h4b == _T_311[9:0] ? 4'h3 : _GEN_14669; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14671 = 10'h4c == _T_311[9:0] ? 4'h3 : _GEN_14670; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14672 = 10'h4d == _T_311[9:0] ? 4'h5 : _GEN_14671; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14673 = 10'h4e == _T_311[9:0] ? 4'h3 : _GEN_14672; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14674 = 10'h4f == _T_311[9:0] ? 4'h3 : _GEN_14673; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14675 = 10'h50 == _T_311[9:0] ? 4'h3 : _GEN_14674; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14676 = 10'h51 == _T_311[9:0] ? 4'h3 : _GEN_14675; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14677 = 10'h52 == _T_311[9:0] ? 4'h3 : _GEN_14676; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14678 = 10'h53 == _T_311[9:0] ? 4'h3 : _GEN_14677; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14679 = 10'h54 == _T_311[9:0] ? 4'h1 : _GEN_14678; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14680 = 10'h55 == _T_311[9:0] ? 4'h1 : _GEN_14679; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14681 = 10'h56 == _T_311[9:0] ? 4'h1 : _GEN_14680; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14682 = 10'h57 == _T_311[9:0] ? 4'h0 : _GEN_14681; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14683 = 10'h58 == _T_311[9:0] ? 4'h3 : _GEN_14682; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14684 = 10'h59 == _T_311[9:0] ? 4'h0 : _GEN_14683; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14685 = 10'h5a == _T_311[9:0] ? 4'h3 : _GEN_14684; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14686 = 10'h5b == _T_311[9:0] ? 4'h3 : _GEN_14685; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14687 = 10'h5c == _T_311[9:0] ? 4'h3 : _GEN_14686; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14688 = 10'h5d == _T_311[9:0] ? 4'ha : _GEN_14687; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14689 = 10'h5e == _T_311[9:0] ? 4'h3 : _GEN_14688; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14690 = 10'h5f == _T_311[9:0] ? 4'h0 : _GEN_14689; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14691 = 10'h60 == _T_311[9:0] ? 4'h3 : _GEN_14690; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14692 = 10'h61 == _T_311[9:0] ? 4'h3 : _GEN_14691; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14693 = 10'h62 == _T_311[9:0] ? 4'h3 : _GEN_14692; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14694 = 10'h63 == _T_311[9:0] ? 4'h3 : _GEN_14693; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14695 = 10'h64 == _T_311[9:0] ? 4'ha : _GEN_14694; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14696 = 10'h65 == _T_311[9:0] ? 4'h0 : _GEN_14695; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14697 = 10'h66 == _T_311[9:0] ? 4'h3 : _GEN_14696; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14698 = 10'h67 == _T_311[9:0] ? 4'h3 : _GEN_14697; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14699 = 10'h68 == _T_311[9:0] ? 4'h3 : _GEN_14698; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14700 = 10'h69 == _T_311[9:0] ? 4'h0 : _GEN_14699; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14701 = 10'h6a == _T_311[9:0] ? 4'h1 : _GEN_14700; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14702 = 10'h6b == _T_311[9:0] ? 4'h1 : _GEN_14701; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14703 = 10'h6c == _T_311[9:0] ? 4'h3 : _GEN_14702; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14704 = 10'h6d == _T_311[9:0] ? 4'h3 : _GEN_14703; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14705 = 10'h6e == _T_311[9:0] ? 4'h3 : _GEN_14704; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14706 = 10'h6f == _T_311[9:0] ? 4'h3 : _GEN_14705; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14707 = 10'h70 == _T_311[9:0] ? 4'h3 : _GEN_14706; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14708 = 10'h71 == _T_311[9:0] ? 4'h3 : _GEN_14707; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14709 = 10'h72 == _T_311[9:0] ? 4'h3 : _GEN_14708; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14710 = 10'h73 == _T_311[9:0] ? 4'h1 : _GEN_14709; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14711 = 10'h74 == _T_311[9:0] ? 4'h0 : _GEN_14710; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14712 = 10'h75 == _T_311[9:0] ? 4'h0 : _GEN_14711; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14713 = 10'h76 == _T_311[9:0] ? 4'h0 : _GEN_14712; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14714 = 10'h77 == _T_311[9:0] ? 4'h3 : _GEN_14713; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14715 = 10'h78 == _T_311[9:0] ? 4'h3 : _GEN_14714; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14716 = 10'h79 == _T_311[9:0] ? 4'h3 : _GEN_14715; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14717 = 10'h7a == _T_311[9:0] ? 4'h0 : _GEN_14716; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14718 = 10'h7b == _T_311[9:0] ? 4'h3 : _GEN_14717; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14719 = 10'h7c == _T_311[9:0] ? 4'h3 : _GEN_14718; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14720 = 10'h7d == _T_311[9:0] ? 4'h7 : _GEN_14719; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14721 = 10'h7e == _T_311[9:0] ? 4'ha : _GEN_14720; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14722 = 10'h7f == _T_311[9:0] ? 4'h0 : _GEN_14721; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14723 = 10'h80 == _T_311[9:0] ? 4'h3 : _GEN_14722; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14724 = 10'h81 == _T_311[9:0] ? 4'h3 : _GEN_14723; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14725 = 10'h82 == _T_311[9:0] ? 4'h1 : _GEN_14724; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14726 = 10'h83 == _T_311[9:0] ? 4'h0 : _GEN_14725; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14727 = 10'h84 == _T_311[9:0] ? 4'h7 : _GEN_14726; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14728 = 10'h85 == _T_311[9:0] ? 4'h1 : _GEN_14727; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14729 = 10'h86 == _T_311[9:0] ? 4'h1 : _GEN_14728; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14730 = 10'h87 == _T_311[9:0] ? 4'h3 : _GEN_14729; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14731 = 10'h88 == _T_311[9:0] ? 4'h3 : _GEN_14730; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14732 = 10'h89 == _T_311[9:0] ? 4'h0 : _GEN_14731; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14733 = 10'h8a == _T_311[9:0] ? 4'h0 : _GEN_14732; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14734 = 10'h8b == _T_311[9:0] ? 4'h1 : _GEN_14733; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14735 = 10'h8c == _T_311[9:0] ? 4'h1 : _GEN_14734; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14736 = 10'h8d == _T_311[9:0] ? 4'h1 : _GEN_14735; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14737 = 10'h8e == _T_311[9:0] ? 4'h1 : _GEN_14736; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14738 = 10'h8f == _T_311[9:0] ? 4'h1 : _GEN_14737; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14739 = 10'h90 == _T_311[9:0] ? 4'h1 : _GEN_14738; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14740 = 10'h91 == _T_311[9:0] ? 4'h1 : _GEN_14739; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14741 = 10'h92 == _T_311[9:0] ? 4'h1 : _GEN_14740; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14742 = 10'h93 == _T_311[9:0] ? 4'h0 : _GEN_14741; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14743 = 10'h94 == _T_311[9:0] ? 4'h0 : _GEN_14742; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14744 = 10'h95 == _T_311[9:0] ? 4'h3 : _GEN_14743; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14745 = 10'h96 == _T_311[9:0] ? 4'h3 : _GEN_14744; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14746 = 10'h97 == _T_311[9:0] ? 4'h3 : _GEN_14745; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14747 = 10'h98 == _T_311[9:0] ? 4'h1 : _GEN_14746; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14748 = 10'h99 == _T_311[9:0] ? 4'h0 : _GEN_14747; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14749 = 10'h9a == _T_311[9:0] ? 4'h1 : _GEN_14748; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14750 = 10'h9b == _T_311[9:0] ? 4'h1 : _GEN_14749; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14751 = 10'h9c == _T_311[9:0] ? 4'h3 : _GEN_14750; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14752 = 10'h9d == _T_311[9:0] ? 4'h3 : _GEN_14751; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14753 = 10'h9e == _T_311[9:0] ? 4'ha : _GEN_14752; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14754 = 10'h9f == _T_311[9:0] ? 4'h0 : _GEN_14753; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14755 = 10'ha0 == _T_311[9:0] ? 4'h3 : _GEN_14754; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14756 = 10'ha1 == _T_311[9:0] ? 4'h1 : _GEN_14755; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14757 = 10'ha2 == _T_311[9:0] ? 4'h0 : _GEN_14756; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14758 = 10'ha3 == _T_311[9:0] ? 4'ha : _GEN_14757; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14759 = 10'ha4 == _T_311[9:0] ? 4'h3 : _GEN_14758; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14760 = 10'ha5 == _T_311[9:0] ? 4'h3 : _GEN_14759; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14761 = 10'ha6 == _T_311[9:0] ? 4'h3 : _GEN_14760; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14762 = 10'ha7 == _T_311[9:0] ? 4'h0 : _GEN_14761; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14763 = 10'ha8 == _T_311[9:0] ? 4'h3 : _GEN_14762; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14764 = 10'ha9 == _T_311[9:0] ? 4'h1 : _GEN_14763; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14765 = 10'haa == _T_311[9:0] ? 4'h0 : _GEN_14764; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14766 = 10'hab == _T_311[9:0] ? 4'h0 : _GEN_14765; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14767 = 10'hac == _T_311[9:0] ? 4'h0 : _GEN_14766; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14768 = 10'had == _T_311[9:0] ? 4'h0 : _GEN_14767; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14769 = 10'hae == _T_311[9:0] ? 4'h0 : _GEN_14768; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14770 = 10'haf == _T_311[9:0] ? 4'h0 : _GEN_14769; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14771 = 10'hb0 == _T_311[9:0] ? 4'h0 : _GEN_14770; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14772 = 10'hb1 == _T_311[9:0] ? 4'h0 : _GEN_14771; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14773 = 10'hb2 == _T_311[9:0] ? 4'h0 : _GEN_14772; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14774 = 10'hb3 == _T_311[9:0] ? 4'h0 : _GEN_14773; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14775 = 10'hb4 == _T_311[9:0] ? 4'h1 : _GEN_14774; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14776 = 10'hb5 == _T_311[9:0] ? 4'h1 : _GEN_14775; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14777 = 10'hb6 == _T_311[9:0] ? 4'h3 : _GEN_14776; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14778 = 10'hb7 == _T_311[9:0] ? 4'h0 : _GEN_14777; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14779 = 10'hb8 == _T_311[9:0] ? 4'h3 : _GEN_14778; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14780 = 10'hb9 == _T_311[9:0] ? 4'h3 : _GEN_14779; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14781 = 10'hba == _T_311[9:0] ? 4'h3 : _GEN_14780; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14782 = 10'hbb == _T_311[9:0] ? 4'h0 : _GEN_14781; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14783 = 10'hbc == _T_311[9:0] ? 4'h3 : _GEN_14782; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14784 = 10'hbd == _T_311[9:0] ? 4'h3 : _GEN_14783; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14785 = 10'hbe == _T_311[9:0] ? 4'ha : _GEN_14784; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14786 = 10'hbf == _T_311[9:0] ? 4'h0 : _GEN_14785; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14787 = 10'hc0 == _T_311[9:0] ? 4'h3 : _GEN_14786; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14788 = 10'hc1 == _T_311[9:0] ? 4'h3 : _GEN_14787; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14789 = 10'hc2 == _T_311[9:0] ? 4'ha : _GEN_14788; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14790 = 10'hc3 == _T_311[9:0] ? 4'h7 : _GEN_14789; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14791 = 10'hc4 == _T_311[9:0] ? 4'h0 : _GEN_14790; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14792 = 10'hc5 == _T_311[9:0] ? 4'h0 : _GEN_14791; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14793 = 10'hc6 == _T_311[9:0] ? 4'h0 : _GEN_14792; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14794 = 10'hc7 == _T_311[9:0] ? 4'h3 : _GEN_14793; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14795 = 10'hc8 == _T_311[9:0] ? 4'h1 : _GEN_14794; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14796 = 10'hc9 == _T_311[9:0] ? 4'h0 : _GEN_14795; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14797 = 10'hca == _T_311[9:0] ? 4'h0 : _GEN_14796; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14798 = 10'hcb == _T_311[9:0] ? 4'h0 : _GEN_14797; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14799 = 10'hcc == _T_311[9:0] ? 4'h0 : _GEN_14798; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14800 = 10'hcd == _T_311[9:0] ? 4'h0 : _GEN_14799; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14801 = 10'hce == _T_311[9:0] ? 4'h0 : _GEN_14800; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14802 = 10'hcf == _T_311[9:0] ? 4'h0 : _GEN_14801; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14803 = 10'hd0 == _T_311[9:0] ? 4'h0 : _GEN_14802; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14804 = 10'hd1 == _T_311[9:0] ? 4'h0 : _GEN_14803; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14805 = 10'hd2 == _T_311[9:0] ? 4'h0 : _GEN_14804; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14806 = 10'hd3 == _T_311[9:0] ? 4'h0 : _GEN_14805; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14807 = 10'hd4 == _T_311[9:0] ? 4'h0 : _GEN_14806; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14808 = 10'hd5 == _T_311[9:0] ? 4'h0 : _GEN_14807; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14809 = 10'hd6 == _T_311[9:0] ? 4'h1 : _GEN_14808; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14810 = 10'hd7 == _T_311[9:0] ? 4'h3 : _GEN_14809; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14811 = 10'hd8 == _T_311[9:0] ? 4'h0 : _GEN_14810; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14812 = 10'hd9 == _T_311[9:0] ? 4'h3 : _GEN_14811; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14813 = 10'hda == _T_311[9:0] ? 4'h3 : _GEN_14812; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14814 = 10'hdb == _T_311[9:0] ? 4'h3 : _GEN_14813; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14815 = 10'hdc == _T_311[9:0] ? 4'h3 : _GEN_14814; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14816 = 10'hdd == _T_311[9:0] ? 4'ha : _GEN_14815; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14817 = 10'hde == _T_311[9:0] ? 4'h7 : _GEN_14816; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14818 = 10'hdf == _T_311[9:0] ? 4'h0 : _GEN_14817; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14819 = 10'he0 == _T_311[9:0] ? 4'h3 : _GEN_14818; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14820 = 10'he1 == _T_311[9:0] ? 4'h3 : _GEN_14819; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14821 = 10'he2 == _T_311[9:0] ? 4'ha : _GEN_14820; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14822 = 10'he3 == _T_311[9:0] ? 4'h3 : _GEN_14821; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14823 = 10'he4 == _T_311[9:0] ? 4'h3 : _GEN_14822; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14824 = 10'he5 == _T_311[9:0] ? 4'h3 : _GEN_14823; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14825 = 10'he6 == _T_311[9:0] ? 4'h3 : _GEN_14824; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14826 = 10'he7 == _T_311[9:0] ? 4'h1 : _GEN_14825; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14827 = 10'he8 == _T_311[9:0] ? 4'h1 : _GEN_14826; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14828 = 10'he9 == _T_311[9:0] ? 4'h1 : _GEN_14827; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14829 = 10'hea == _T_311[9:0] ? 4'h0 : _GEN_14828; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14830 = 10'heb == _T_311[9:0] ? 4'h0 : _GEN_14829; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14831 = 10'hec == _T_311[9:0] ? 4'h0 : _GEN_14830; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14832 = 10'hed == _T_311[9:0] ? 4'h0 : _GEN_14831; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14833 = 10'hee == _T_311[9:0] ? 4'h0 : _GEN_14832; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14834 = 10'hef == _T_311[9:0] ? 4'h0 : _GEN_14833; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14835 = 10'hf0 == _T_311[9:0] ? 4'h0 : _GEN_14834; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14836 = 10'hf1 == _T_311[9:0] ? 4'h0 : _GEN_14835; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14837 = 10'hf2 == _T_311[9:0] ? 4'h0 : _GEN_14836; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14838 = 10'hf3 == _T_311[9:0] ? 4'h0 : _GEN_14837; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14839 = 10'hf4 == _T_311[9:0] ? 4'h0 : _GEN_14838; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14840 = 10'hf5 == _T_311[9:0] ? 4'h1 : _GEN_14839; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14841 = 10'hf6 == _T_311[9:0] ? 4'h0 : _GEN_14840; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14842 = 10'hf7 == _T_311[9:0] ? 4'h0 : _GEN_14841; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14843 = 10'hf8 == _T_311[9:0] ? 4'h1 : _GEN_14842; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14844 = 10'hf9 == _T_311[9:0] ? 4'h0 : _GEN_14843; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14845 = 10'hfa == _T_311[9:0] ? 4'h3 : _GEN_14844; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14846 = 10'hfb == _T_311[9:0] ? 4'h3 : _GEN_14845; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14847 = 10'hfc == _T_311[9:0] ? 4'h3 : _GEN_14846; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14848 = 10'hfd == _T_311[9:0] ? 4'ha : _GEN_14847; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14849 = 10'hfe == _T_311[9:0] ? 4'h3 : _GEN_14848; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14850 = 10'hff == _T_311[9:0] ? 4'h0 : _GEN_14849; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14851 = 10'h100 == _T_311[9:0] ? 4'h3 : _GEN_14850; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14852 = 10'h101 == _T_311[9:0] ? 4'h0 : _GEN_14851; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14853 = 10'h102 == _T_311[9:0] ? 4'ha : _GEN_14852; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14854 = 10'h103 == _T_311[9:0] ? 4'h3 : _GEN_14853; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14855 = 10'h104 == _T_311[9:0] ? 4'h3 : _GEN_14854; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14856 = 10'h105 == _T_311[9:0] ? 4'h3 : _GEN_14855; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14857 = 10'h106 == _T_311[9:0] ? 4'h3 : _GEN_14856; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14858 = 10'h107 == _T_311[9:0] ? 4'h3 : _GEN_14857; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14859 = 10'h108 == _T_311[9:0] ? 4'h1 : _GEN_14858; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14860 = 10'h109 == _T_311[9:0] ? 4'h0 : _GEN_14859; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14861 = 10'h10a == _T_311[9:0] ? 4'h0 : _GEN_14860; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14862 = 10'h10b == _T_311[9:0] ? 4'h0 : _GEN_14861; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14863 = 10'h10c == _T_311[9:0] ? 4'h0 : _GEN_14862; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14864 = 10'h10d == _T_311[9:0] ? 4'h0 : _GEN_14863; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14865 = 10'h10e == _T_311[9:0] ? 4'h0 : _GEN_14864; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14866 = 10'h10f == _T_311[9:0] ? 4'h0 : _GEN_14865; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14867 = 10'h110 == _T_311[9:0] ? 4'h0 : _GEN_14866; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14868 = 10'h111 == _T_311[9:0] ? 4'h0 : _GEN_14867; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14869 = 10'h112 == _T_311[9:0] ? 4'h0 : _GEN_14868; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14870 = 10'h113 == _T_311[9:0] ? 4'h0 : _GEN_14869; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14871 = 10'h114 == _T_311[9:0] ? 4'h0 : _GEN_14870; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14872 = 10'h115 == _T_311[9:0] ? 4'h0 : _GEN_14871; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14873 = 10'h116 == _T_311[9:0] ? 4'h1 : _GEN_14872; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14874 = 10'h117 == _T_311[9:0] ? 4'h3 : _GEN_14873; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14875 = 10'h118 == _T_311[9:0] ? 4'h3 : _GEN_14874; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14876 = 10'h119 == _T_311[9:0] ? 4'h3 : _GEN_14875; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14877 = 10'h11a == _T_311[9:0] ? 4'h0 : _GEN_14876; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14878 = 10'h11b == _T_311[9:0] ? 4'h3 : _GEN_14877; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14879 = 10'h11c == _T_311[9:0] ? 4'h3 : _GEN_14878; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14880 = 10'h11d == _T_311[9:0] ? 4'h7 : _GEN_14879; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14881 = 10'h11e == _T_311[9:0] ? 4'ha : _GEN_14880; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14882 = 10'h11f == _T_311[9:0] ? 4'h0 : _GEN_14881; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14883 = 10'h120 == _T_311[9:0] ? 4'h3 : _GEN_14882; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14884 = 10'h121 == _T_311[9:0] ? 4'h3 : _GEN_14883; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14885 = 10'h122 == _T_311[9:0] ? 4'ha : _GEN_14884; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14886 = 10'h123 == _T_311[9:0] ? 4'h3 : _GEN_14885; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14887 = 10'h124 == _T_311[9:0] ? 4'h3 : _GEN_14886; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14888 = 10'h125 == _T_311[9:0] ? 4'h3 : _GEN_14887; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14889 = 10'h126 == _T_311[9:0] ? 4'h3 : _GEN_14888; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14890 = 10'h127 == _T_311[9:0] ? 4'h1 : _GEN_14889; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14891 = 10'h128 == _T_311[9:0] ? 4'h0 : _GEN_14890; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14892 = 10'h129 == _T_311[9:0] ? 4'h3 : _GEN_14891; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14893 = 10'h12a == _T_311[9:0] ? 4'h3 : _GEN_14892; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14894 = 10'h12b == _T_311[9:0] ? 4'h0 : _GEN_14893; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14895 = 10'h12c == _T_311[9:0] ? 4'h0 : _GEN_14894; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14896 = 10'h12d == _T_311[9:0] ? 4'h0 : _GEN_14895; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14897 = 10'h12e == _T_311[9:0] ? 4'h0 : _GEN_14896; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14898 = 10'h12f == _T_311[9:0] ? 4'h0 : _GEN_14897; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14899 = 10'h130 == _T_311[9:0] ? 4'h0 : _GEN_14898; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14900 = 10'h131 == _T_311[9:0] ? 4'h0 : _GEN_14899; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14901 = 10'h132 == _T_311[9:0] ? 4'h0 : _GEN_14900; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14902 = 10'h133 == _T_311[9:0] ? 4'h0 : _GEN_14901; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14903 = 10'h134 == _T_311[9:0] ? 4'h3 : _GEN_14902; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14904 = 10'h135 == _T_311[9:0] ? 4'h3 : _GEN_14903; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14905 = 10'h136 == _T_311[9:0] ? 4'h0 : _GEN_14904; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14906 = 10'h137 == _T_311[9:0] ? 4'h1 : _GEN_14905; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14907 = 10'h138 == _T_311[9:0] ? 4'h3 : _GEN_14906; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14908 = 10'h139 == _T_311[9:0] ? 4'h3 : _GEN_14907; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14909 = 10'h13a == _T_311[9:0] ? 4'h3 : _GEN_14908; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14910 = 10'h13b == _T_311[9:0] ? 4'h3 : _GEN_14909; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14911 = 10'h13c == _T_311[9:0] ? 4'h3 : _GEN_14910; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14912 = 10'h13d == _T_311[9:0] ? 4'h3 : _GEN_14911; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14913 = 10'h13e == _T_311[9:0] ? 4'ha : _GEN_14912; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14914 = 10'h13f == _T_311[9:0] ? 4'h0 : _GEN_14913; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14915 = 10'h140 == _T_311[9:0] ? 4'h5 : _GEN_14914; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14916 = 10'h141 == _T_311[9:0] ? 4'h3 : _GEN_14915; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14917 = 10'h142 == _T_311[9:0] ? 4'h7 : _GEN_14916; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14918 = 10'h143 == _T_311[9:0] ? 4'ha : _GEN_14917; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14919 = 10'h144 == _T_311[9:0] ? 4'h3 : _GEN_14918; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14920 = 10'h145 == _T_311[9:0] ? 4'h3 : _GEN_14919; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14921 = 10'h146 == _T_311[9:0] ? 4'h1 : _GEN_14920; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14922 = 10'h147 == _T_311[9:0] ? 4'h0 : _GEN_14921; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14923 = 10'h148 == _T_311[9:0] ? 4'h3 : _GEN_14922; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14924 = 10'h149 == _T_311[9:0] ? 4'h3 : _GEN_14923; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14925 = 10'h14a == _T_311[9:0] ? 4'h3 : _GEN_14924; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14926 = 10'h14b == _T_311[9:0] ? 4'h3 : _GEN_14925; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14927 = 10'h14c == _T_311[9:0] ? 4'h3 : _GEN_14926; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14928 = 10'h14d == _T_311[9:0] ? 4'h3 : _GEN_14927; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14929 = 10'h14e == _T_311[9:0] ? 4'h3 : _GEN_14928; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14930 = 10'h14f == _T_311[9:0] ? 4'h3 : _GEN_14929; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14931 = 10'h150 == _T_311[9:0] ? 4'h3 : _GEN_14930; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14932 = 10'h151 == _T_311[9:0] ? 4'h3 : _GEN_14931; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14933 = 10'h152 == _T_311[9:0] ? 4'h3 : _GEN_14932; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14934 = 10'h153 == _T_311[9:0] ? 4'h3 : _GEN_14933; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14935 = 10'h154 == _T_311[9:0] ? 4'h3 : _GEN_14934; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14936 = 10'h155 == _T_311[9:0] ? 4'h3 : _GEN_14935; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14937 = 10'h156 == _T_311[9:0] ? 4'h3 : _GEN_14936; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14938 = 10'h157 == _T_311[9:0] ? 4'h0 : _GEN_14937; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14939 = 10'h158 == _T_311[9:0] ? 4'h3 : _GEN_14938; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14940 = 10'h159 == _T_311[9:0] ? 4'h3 : _GEN_14939; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14941 = 10'h15a == _T_311[9:0] ? 4'h3 : _GEN_14940; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14942 = 10'h15b == _T_311[9:0] ? 4'h3 : _GEN_14941; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14943 = 10'h15c == _T_311[9:0] ? 4'h3 : _GEN_14942; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14944 = 10'h15d == _T_311[9:0] ? 4'ha : _GEN_14943; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14945 = 10'h15e == _T_311[9:0] ? 4'h7 : _GEN_14944; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14946 = 10'h15f == _T_311[9:0] ? 4'h0 : _GEN_14945; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14947 = 10'h160 == _T_311[9:0] ? 4'h3 : _GEN_14946; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14948 = 10'h161 == _T_311[9:0] ? 4'h3 : _GEN_14947; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14949 = 10'h162 == _T_311[9:0] ? 4'h3 : _GEN_14948; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14950 = 10'h163 == _T_311[9:0] ? 4'h7 : _GEN_14949; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14951 = 10'h164 == _T_311[9:0] ? 4'ha : _GEN_14950; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14952 = 10'h165 == _T_311[9:0] ? 4'h1 : _GEN_14951; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14953 = 10'h166 == _T_311[9:0] ? 4'h0 : _GEN_14952; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14954 = 10'h167 == _T_311[9:0] ? 4'h0 : _GEN_14953; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14955 = 10'h168 == _T_311[9:0] ? 4'hc : _GEN_14954; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14956 = 10'h169 == _T_311[9:0] ? 4'h9 : _GEN_14955; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14957 = 10'h16a == _T_311[9:0] ? 4'hc : _GEN_14956; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14958 = 10'h16b == _T_311[9:0] ? 4'hc : _GEN_14957; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14959 = 10'h16c == _T_311[9:0] ? 4'h3 : _GEN_14958; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14960 = 10'h16d == _T_311[9:0] ? 4'h3 : _GEN_14959; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14961 = 10'h16e == _T_311[9:0] ? 4'h3 : _GEN_14960; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14962 = 10'h16f == _T_311[9:0] ? 4'h3 : _GEN_14961; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14963 = 10'h170 == _T_311[9:0] ? 4'h5 : _GEN_14962; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14964 = 10'h171 == _T_311[9:0] ? 4'h3 : _GEN_14963; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14965 = 10'h172 == _T_311[9:0] ? 4'h3 : _GEN_14964; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14966 = 10'h173 == _T_311[9:0] ? 4'h3 : _GEN_14965; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14967 = 10'h174 == _T_311[9:0] ? 4'h3 : _GEN_14966; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14968 = 10'h175 == _T_311[9:0] ? 4'h3 : _GEN_14967; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14969 = 10'h176 == _T_311[9:0] ? 4'h0 : _GEN_14968; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14970 = 10'h177 == _T_311[9:0] ? 4'h0 : _GEN_14969; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14971 = 10'h178 == _T_311[9:0] ? 4'h1 : _GEN_14970; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14972 = 10'h179 == _T_311[9:0] ? 4'h3 : _GEN_14971; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14973 = 10'h17a == _T_311[9:0] ? 4'h5 : _GEN_14972; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14974 = 10'h17b == _T_311[9:0] ? 4'h3 : _GEN_14973; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14975 = 10'h17c == _T_311[9:0] ? 4'ha : _GEN_14974; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14976 = 10'h17d == _T_311[9:0] ? 4'h7 : _GEN_14975; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14977 = 10'h17e == _T_311[9:0] ? 4'h3 : _GEN_14976; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14978 = 10'h17f == _T_311[9:0] ? 4'h0 : _GEN_14977; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14979 = 10'h180 == _T_311[9:0] ? 4'hc : _GEN_14978; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14980 = 10'h181 == _T_311[9:0] ? 4'hc : _GEN_14979; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14981 = 10'h182 == _T_311[9:0] ? 4'hc : _GEN_14980; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14982 = 10'h183 == _T_311[9:0] ? 4'hc : _GEN_14981; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14983 = 10'h184 == _T_311[9:0] ? 4'ha : _GEN_14982; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14984 = 10'h185 == _T_311[9:0] ? 4'h1 : _GEN_14983; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14985 = 10'h186 == _T_311[9:0] ? 4'hc : _GEN_14984; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14986 = 10'h187 == _T_311[9:0] ? 4'h0 : _GEN_14985; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14987 = 10'h188 == _T_311[9:0] ? 4'hc : _GEN_14986; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14988 = 10'h189 == _T_311[9:0] ? 4'hc : _GEN_14987; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14989 = 10'h18a == _T_311[9:0] ? 4'hc : _GEN_14988; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14990 = 10'h18b == _T_311[9:0] ? 4'hc : _GEN_14989; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14991 = 10'h18c == _T_311[9:0] ? 4'hc : _GEN_14990; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14992 = 10'h18d == _T_311[9:0] ? 4'hc : _GEN_14991; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14993 = 10'h18e == _T_311[9:0] ? 4'hc : _GEN_14992; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14994 = 10'h18f == _T_311[9:0] ? 4'hc : _GEN_14993; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14995 = 10'h190 == _T_311[9:0] ? 4'hc : _GEN_14994; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14996 = 10'h191 == _T_311[9:0] ? 4'hc : _GEN_14995; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14997 = 10'h192 == _T_311[9:0] ? 4'h9 : _GEN_14996; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14998 = 10'h193 == _T_311[9:0] ? 4'hc : _GEN_14997; // @[Filter.scala 191:102]
  wire [3:0] _GEN_14999 = 10'h194 == _T_311[9:0] ? 4'hc : _GEN_14998; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15000 = 10'h195 == _T_311[9:0] ? 4'hc : _GEN_14999; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15001 = 10'h196 == _T_311[9:0] ? 4'h0 : _GEN_15000; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15002 = 10'h197 == _T_311[9:0] ? 4'h3 : _GEN_15001; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15003 = 10'h198 == _T_311[9:0] ? 4'h1 : _GEN_15002; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15004 = 10'h199 == _T_311[9:0] ? 4'h3 : _GEN_15003; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15005 = 10'h19a == _T_311[9:0] ? 4'h3 : _GEN_15004; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15006 = 10'h19b == _T_311[9:0] ? 4'h3 : _GEN_15005; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15007 = 10'h19c == _T_311[9:0] ? 4'ha : _GEN_15006; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15008 = 10'h19d == _T_311[9:0] ? 4'h3 : _GEN_15007; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15009 = 10'h19e == _T_311[9:0] ? 4'h3 : _GEN_15008; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15010 = 10'h19f == _T_311[9:0] ? 4'h0 : _GEN_15009; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15011 = 10'h1a0 == _T_311[9:0] ? 4'hc : _GEN_15010; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15012 = 10'h1a1 == _T_311[9:0] ? 4'hc : _GEN_15011; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15013 = 10'h1a2 == _T_311[9:0] ? 4'h9 : _GEN_15012; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15014 = 10'h1a3 == _T_311[9:0] ? 4'hc : _GEN_15013; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15015 = 10'h1a4 == _T_311[9:0] ? 4'ha : _GEN_15014; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15016 = 10'h1a5 == _T_311[9:0] ? 4'h0 : _GEN_15015; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15017 = 10'h1a6 == _T_311[9:0] ? 4'hc : _GEN_15016; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15018 = 10'h1a7 == _T_311[9:0] ? 4'h0 : _GEN_15017; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15019 = 10'h1a8 == _T_311[9:0] ? 4'hc : _GEN_15018; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15020 = 10'h1a9 == _T_311[9:0] ? 4'hc : _GEN_15019; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15021 = 10'h1aa == _T_311[9:0] ? 4'hc : _GEN_15020; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15022 = 10'h1ab == _T_311[9:0] ? 4'h9 : _GEN_15021; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15023 = 10'h1ac == _T_311[9:0] ? 4'hc : _GEN_15022; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15024 = 10'h1ad == _T_311[9:0] ? 4'hc : _GEN_15023; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15025 = 10'h1ae == _T_311[9:0] ? 4'hc : _GEN_15024; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15026 = 10'h1af == _T_311[9:0] ? 4'hc : _GEN_15025; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15027 = 10'h1b0 == _T_311[9:0] ? 4'hc : _GEN_15026; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15028 = 10'h1b1 == _T_311[9:0] ? 4'hc : _GEN_15027; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15029 = 10'h1b2 == _T_311[9:0] ? 4'hc : _GEN_15028; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15030 = 10'h1b3 == _T_311[9:0] ? 4'hc : _GEN_15029; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15031 = 10'h1b4 == _T_311[9:0] ? 4'hc : _GEN_15030; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15032 = 10'h1b5 == _T_311[9:0] ? 4'hc : _GEN_15031; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15033 = 10'h1b6 == _T_311[9:0] ? 4'h0 : _GEN_15032; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15034 = 10'h1b7 == _T_311[9:0] ? 4'hc : _GEN_15033; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15035 = 10'h1b8 == _T_311[9:0] ? 4'h0 : _GEN_15034; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15036 = 10'h1b9 == _T_311[9:0] ? 4'hc : _GEN_15035; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15037 = 10'h1ba == _T_311[9:0] ? 4'hc : _GEN_15036; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15038 = 10'h1bb == _T_311[9:0] ? 4'hc : _GEN_15037; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15039 = 10'h1bc == _T_311[9:0] ? 4'h7 : _GEN_15038; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15040 = 10'h1bd == _T_311[9:0] ? 4'ha : _GEN_15039; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15041 = 10'h1be == _T_311[9:0] ? 4'hc : _GEN_15040; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15042 = 10'h1bf == _T_311[9:0] ? 4'h0 : _GEN_15041; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15043 = 10'h1c0 == _T_311[9:0] ? 4'hc : _GEN_15042; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15044 = 10'h1c1 == _T_311[9:0] ? 4'hc : _GEN_15043; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15045 = 10'h1c2 == _T_311[9:0] ? 4'hc : _GEN_15044; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15046 = 10'h1c3 == _T_311[9:0] ? 4'h7 : _GEN_15045; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15047 = 10'h1c4 == _T_311[9:0] ? 4'h7 : _GEN_15046; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15048 = 10'h1c5 == _T_311[9:0] ? 4'hc : _GEN_15047; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15049 = 10'h1c6 == _T_311[9:0] ? 4'hc : _GEN_15048; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15050 = 10'h1c7 == _T_311[9:0] ? 4'hc : _GEN_15049; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15051 = 10'h1c8 == _T_311[9:0] ? 4'hc : _GEN_15050; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15052 = 10'h1c9 == _T_311[9:0] ? 4'hc : _GEN_15051; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15053 = 10'h1ca == _T_311[9:0] ? 4'hc : _GEN_15052; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15054 = 10'h1cb == _T_311[9:0] ? 4'hc : _GEN_15053; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15055 = 10'h1cc == _T_311[9:0] ? 4'hc : _GEN_15054; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15056 = 10'h1cd == _T_311[9:0] ? 4'hc : _GEN_15055; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15057 = 10'h1ce == _T_311[9:0] ? 4'hc : _GEN_15056; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15058 = 10'h1cf == _T_311[9:0] ? 4'hc : _GEN_15057; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15059 = 10'h1d0 == _T_311[9:0] ? 4'hc : _GEN_15058; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15060 = 10'h1d1 == _T_311[9:0] ? 4'hc : _GEN_15059; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15061 = 10'h1d2 == _T_311[9:0] ? 4'hc : _GEN_15060; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15062 = 10'h1d3 == _T_311[9:0] ? 4'hc : _GEN_15061; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15063 = 10'h1d4 == _T_311[9:0] ? 4'hc : _GEN_15062; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15064 = 10'h1d5 == _T_311[9:0] ? 4'hc : _GEN_15063; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15065 = 10'h1d6 == _T_311[9:0] ? 4'hc : _GEN_15064; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15066 = 10'h1d7 == _T_311[9:0] ? 4'hc : _GEN_15065; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15067 = 10'h1d8 == _T_311[9:0] ? 4'hc : _GEN_15066; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15068 = 10'h1d9 == _T_311[9:0] ? 4'hc : _GEN_15067; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15069 = 10'h1da == _T_311[9:0] ? 4'hc : _GEN_15068; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15070 = 10'h1db == _T_311[9:0] ? 4'hc : _GEN_15069; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15071 = 10'h1dc == _T_311[9:0] ? 4'hc : _GEN_15070; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15072 = 10'h1dd == _T_311[9:0] ? 4'ha : _GEN_15071; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15073 = 10'h1de == _T_311[9:0] ? 4'hc : _GEN_15072; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15074 = 10'h1df == _T_311[9:0] ? 4'h0 : _GEN_15073; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15075 = 10'h1e0 == _T_311[9:0] ? 4'h9 : _GEN_15074; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15076 = 10'h1e1 == _T_311[9:0] ? 4'hc : _GEN_15075; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15077 = 10'h1e2 == _T_311[9:0] ? 4'h7 : _GEN_15076; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15078 = 10'h1e3 == _T_311[9:0] ? 4'h7 : _GEN_15077; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15079 = 10'h1e4 == _T_311[9:0] ? 4'hc : _GEN_15078; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15080 = 10'h1e5 == _T_311[9:0] ? 4'hc : _GEN_15079; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15081 = 10'h1e6 == _T_311[9:0] ? 4'hc : _GEN_15080; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15082 = 10'h1e7 == _T_311[9:0] ? 4'hc : _GEN_15081; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15083 = 10'h1e8 == _T_311[9:0] ? 4'hc : _GEN_15082; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15084 = 10'h1e9 == _T_311[9:0] ? 4'hc : _GEN_15083; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15085 = 10'h1ea == _T_311[9:0] ? 4'hc : _GEN_15084; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15086 = 10'h1eb == _T_311[9:0] ? 4'hc : _GEN_15085; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15087 = 10'h1ec == _T_311[9:0] ? 4'hc : _GEN_15086; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15088 = 10'h1ed == _T_311[9:0] ? 4'hc : _GEN_15087; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15089 = 10'h1ee == _T_311[9:0] ? 4'hc : _GEN_15088; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15090 = 10'h1ef == _T_311[9:0] ? 4'hc : _GEN_15089; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15091 = 10'h1f0 == _T_311[9:0] ? 4'hc : _GEN_15090; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15092 = 10'h1f1 == _T_311[9:0] ? 4'hc : _GEN_15091; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15093 = 10'h1f2 == _T_311[9:0] ? 4'hc : _GEN_15092; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15094 = 10'h1f3 == _T_311[9:0] ? 4'hc : _GEN_15093; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15095 = 10'h1f4 == _T_311[9:0] ? 4'hc : _GEN_15094; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15096 = 10'h1f5 == _T_311[9:0] ? 4'hc : _GEN_15095; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15097 = 10'h1f6 == _T_311[9:0] ? 4'hc : _GEN_15096; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15098 = 10'h1f7 == _T_311[9:0] ? 4'hc : _GEN_15097; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15099 = 10'h1f8 == _T_311[9:0] ? 4'hc : _GEN_15098; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15100 = 10'h1f9 == _T_311[9:0] ? 4'hc : _GEN_15099; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15101 = 10'h1fa == _T_311[9:0] ? 4'h9 : _GEN_15100; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15102 = 10'h1fb == _T_311[9:0] ? 4'hc : _GEN_15101; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15103 = 10'h1fc == _T_311[9:0] ? 4'hc : _GEN_15102; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15104 = 10'h1fd == _T_311[9:0] ? 4'h7 : _GEN_15103; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15105 = 10'h1fe == _T_311[9:0] ? 4'hc : _GEN_15104; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15106 = 10'h1ff == _T_311[9:0] ? 4'h0 : _GEN_15105; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15107 = 10'h200 == _T_311[9:0] ? 4'hc : _GEN_15106; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15108 = 10'h201 == _T_311[9:0] ? 4'hc : _GEN_15107; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15109 = 10'h202 == _T_311[9:0] ? 4'ha : _GEN_15108; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15110 = 10'h203 == _T_311[9:0] ? 4'hc : _GEN_15109; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15111 = 10'h204 == _T_311[9:0] ? 4'hc : _GEN_15110; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15112 = 10'h205 == _T_311[9:0] ? 4'hc : _GEN_15111; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15113 = 10'h206 == _T_311[9:0] ? 4'hc : _GEN_15112; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15114 = 10'h207 == _T_311[9:0] ? 4'hc : _GEN_15113; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15115 = 10'h208 == _T_311[9:0] ? 4'hc : _GEN_15114; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15116 = 10'h209 == _T_311[9:0] ? 4'hc : _GEN_15115; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15117 = 10'h20a == _T_311[9:0] ? 4'hc : _GEN_15116; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15118 = 10'h20b == _T_311[9:0] ? 4'hc : _GEN_15117; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15119 = 10'h20c == _T_311[9:0] ? 4'hc : _GEN_15118; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15120 = 10'h20d == _T_311[9:0] ? 4'hc : _GEN_15119; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15121 = 10'h20e == _T_311[9:0] ? 4'hc : _GEN_15120; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15122 = 10'h20f == _T_311[9:0] ? 4'hc : _GEN_15121; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15123 = 10'h210 == _T_311[9:0] ? 4'hc : _GEN_15122; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15124 = 10'h211 == _T_311[9:0] ? 4'hc : _GEN_15123; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15125 = 10'h212 == _T_311[9:0] ? 4'hc : _GEN_15124; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15126 = 10'h213 == _T_311[9:0] ? 4'hc : _GEN_15125; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15127 = 10'h214 == _T_311[9:0] ? 4'hc : _GEN_15126; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15128 = 10'h215 == _T_311[9:0] ? 4'hc : _GEN_15127; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15129 = 10'h216 == _T_311[9:0] ? 4'hc : _GEN_15128; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15130 = 10'h217 == _T_311[9:0] ? 4'hc : _GEN_15129; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15131 = 10'h218 == _T_311[9:0] ? 4'hc : _GEN_15130; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15132 = 10'h219 == _T_311[9:0] ? 4'hc : _GEN_15131; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15133 = 10'h21a == _T_311[9:0] ? 4'hc : _GEN_15132; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15134 = 10'h21b == _T_311[9:0] ? 4'hc : _GEN_15133; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15135 = 10'h21c == _T_311[9:0] ? 4'ha : _GEN_15134; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15136 = 10'h21d == _T_311[9:0] ? 4'h7 : _GEN_15135; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15137 = 10'h21e == _T_311[9:0] ? 4'hc : _GEN_15136; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15138 = 10'h21f == _T_311[9:0] ? 4'h0 : _GEN_15137; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15139 = 10'h220 == _T_311[9:0] ? 4'h0 : _GEN_15138; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15140 = 10'h221 == _T_311[9:0] ? 4'h0 : _GEN_15139; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15141 = 10'h222 == _T_311[9:0] ? 4'h0 : _GEN_15140; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15142 = 10'h223 == _T_311[9:0] ? 4'h0 : _GEN_15141; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15143 = 10'h224 == _T_311[9:0] ? 4'h0 : _GEN_15142; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15144 = 10'h225 == _T_311[9:0] ? 4'h0 : _GEN_15143; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15145 = 10'h226 == _T_311[9:0] ? 4'h0 : _GEN_15144; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15146 = 10'h227 == _T_311[9:0] ? 4'h0 : _GEN_15145; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15147 = 10'h228 == _T_311[9:0] ? 4'h0 : _GEN_15146; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15148 = 10'h229 == _T_311[9:0] ? 4'h0 : _GEN_15147; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15149 = 10'h22a == _T_311[9:0] ? 4'h0 : _GEN_15148; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15150 = 10'h22b == _T_311[9:0] ? 4'h0 : _GEN_15149; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15151 = 10'h22c == _T_311[9:0] ? 4'h0 : _GEN_15150; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15152 = 10'h22d == _T_311[9:0] ? 4'h0 : _GEN_15151; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15153 = 10'h22e == _T_311[9:0] ? 4'h0 : _GEN_15152; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15154 = 10'h22f == _T_311[9:0] ? 4'h0 : _GEN_15153; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15155 = 10'h230 == _T_311[9:0] ? 4'h0 : _GEN_15154; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15156 = 10'h231 == _T_311[9:0] ? 4'h0 : _GEN_15155; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15157 = 10'h232 == _T_311[9:0] ? 4'h0 : _GEN_15156; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15158 = 10'h233 == _T_311[9:0] ? 4'h0 : _GEN_15157; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15159 = 10'h234 == _T_311[9:0] ? 4'h0 : _GEN_15158; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15160 = 10'h235 == _T_311[9:0] ? 4'h0 : _GEN_15159; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15161 = 10'h236 == _T_311[9:0] ? 4'h0 : _GEN_15160; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15162 = 10'h237 == _T_311[9:0] ? 4'h0 : _GEN_15161; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15163 = 10'h238 == _T_311[9:0] ? 4'h0 : _GEN_15162; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15164 = 10'h239 == _T_311[9:0] ? 4'h0 : _GEN_15163; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15165 = 10'h23a == _T_311[9:0] ? 4'h0 : _GEN_15164; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15166 = 10'h23b == _T_311[9:0] ? 4'h0 : _GEN_15165; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15167 = 10'h23c == _T_311[9:0] ? 4'h0 : _GEN_15166; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15168 = 10'h23d == _T_311[9:0] ? 4'h0 : _GEN_15167; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15169 = 10'h23e == _T_311[9:0] ? 4'h0 : _GEN_15168; // @[Filter.scala 191:102]
  wire [3:0] _GEN_15170 = 10'h23f == _T_311[9:0] ? 4'h0 : _GEN_15169; // @[Filter.scala 191:102]
  wire [6:0] _GEN_28348 = {{3'd0}, _GEN_15170}; // @[Filter.scala 191:102]
  wire [10:0] _T_318 = _GEN_28348 * 7'h46; // @[Filter.scala 191:102]
  wire [10:0] _GEN_28349 = {{2'd0}, _T_313}; // @[Filter.scala 191:69]
  wire [10:0] _T_320 = _GEN_28349 + _T_318; // @[Filter.scala 191:69]
  wire [3:0] _GEN_15202 = 10'h1f == _T_311[9:0] ? 4'h0 : 4'h3; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15203 = 10'h20 == _T_311[9:0] ? 4'h3 : _GEN_15202; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15204 = 10'h21 == _T_311[9:0] ? 4'h3 : _GEN_15203; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15205 = 10'h22 == _T_311[9:0] ? 4'h3 : _GEN_15204; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15206 = 10'h23 == _T_311[9:0] ? 4'h3 : _GEN_15205; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15207 = 10'h24 == _T_311[9:0] ? 4'h3 : _GEN_15206; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15208 = 10'h25 == _T_311[9:0] ? 4'h3 : _GEN_15207; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15209 = 10'h26 == _T_311[9:0] ? 4'h3 : _GEN_15208; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15210 = 10'h27 == _T_311[9:0] ? 4'h9 : _GEN_15209; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15211 = 10'h28 == _T_311[9:0] ? 4'h9 : _GEN_15210; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15212 = 10'h29 == _T_311[9:0] ? 4'h3 : _GEN_15211; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15213 = 10'h2a == _T_311[9:0] ? 4'h3 : _GEN_15212; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15214 = 10'h2b == _T_311[9:0] ? 4'h3 : _GEN_15213; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15215 = 10'h2c == _T_311[9:0] ? 4'h3 : _GEN_15214; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15216 = 10'h2d == _T_311[9:0] ? 4'h3 : _GEN_15215; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15217 = 10'h2e == _T_311[9:0] ? 4'h3 : _GEN_15216; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15218 = 10'h2f == _T_311[9:0] ? 4'h3 : _GEN_15217; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15219 = 10'h30 == _T_311[9:0] ? 4'h3 : _GEN_15218; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15220 = 10'h31 == _T_311[9:0] ? 4'h3 : _GEN_15219; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15221 = 10'h32 == _T_311[9:0] ? 4'h3 : _GEN_15220; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15222 = 10'h33 == _T_311[9:0] ? 4'h3 : _GEN_15221; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15223 = 10'h34 == _T_311[9:0] ? 4'h3 : _GEN_15222; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15224 = 10'h35 == _T_311[9:0] ? 4'h3 : _GEN_15223; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15225 = 10'h36 == _T_311[9:0] ? 4'h3 : _GEN_15224; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15226 = 10'h37 == _T_311[9:0] ? 4'h9 : _GEN_15225; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15227 = 10'h38 == _T_311[9:0] ? 4'h9 : _GEN_15226; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15228 = 10'h39 == _T_311[9:0] ? 4'h3 : _GEN_15227; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15229 = 10'h3a == _T_311[9:0] ? 4'h3 : _GEN_15228; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15230 = 10'h3b == _T_311[9:0] ? 4'h3 : _GEN_15229; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15231 = 10'h3c == _T_311[9:0] ? 4'h3 : _GEN_15230; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15232 = 10'h3d == _T_311[9:0] ? 4'h3 : _GEN_15231; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15233 = 10'h3e == _T_311[9:0] ? 4'h3 : _GEN_15232; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15234 = 10'h3f == _T_311[9:0] ? 4'h0 : _GEN_15233; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15235 = 10'h40 == _T_311[9:0] ? 4'h3 : _GEN_15234; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15236 = 10'h41 == _T_311[9:0] ? 4'h3 : _GEN_15235; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15237 = 10'h42 == _T_311[9:0] ? 4'h3 : _GEN_15236; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15238 = 10'h43 == _T_311[9:0] ? 4'h2 : _GEN_15237; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15239 = 10'h44 == _T_311[9:0] ? 4'h3 : _GEN_15238; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15240 = 10'h45 == _T_311[9:0] ? 4'hf : _GEN_15239; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15241 = 10'h46 == _T_311[9:0] ? 4'hf : _GEN_15240; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15242 = 10'h47 == _T_311[9:0] ? 4'hf : _GEN_15241; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15243 = 10'h48 == _T_311[9:0] ? 4'hf : _GEN_15242; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15244 = 10'h49 == _T_311[9:0] ? 4'h3 : _GEN_15243; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15245 = 10'h4a == _T_311[9:0] ? 4'h3 : _GEN_15244; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15246 = 10'h4b == _T_311[9:0] ? 4'h3 : _GEN_15245; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15247 = 10'h4c == _T_311[9:0] ? 4'h3 : _GEN_15246; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15248 = 10'h4d == _T_311[9:0] ? 4'h3 : _GEN_15247; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15249 = 10'h4e == _T_311[9:0] ? 4'h3 : _GEN_15248; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15250 = 10'h4f == _T_311[9:0] ? 4'h3 : _GEN_15249; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15251 = 10'h50 == _T_311[9:0] ? 4'h3 : _GEN_15250; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15252 = 10'h51 == _T_311[9:0] ? 4'h3 : _GEN_15251; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15253 = 10'h52 == _T_311[9:0] ? 4'h3 : _GEN_15252; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15254 = 10'h53 == _T_311[9:0] ? 4'h3 : _GEN_15253; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15255 = 10'h54 == _T_311[9:0] ? 4'h9 : _GEN_15254; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15256 = 10'h55 == _T_311[9:0] ? 4'h9 : _GEN_15255; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15257 = 10'h56 == _T_311[9:0] ? 4'h9 : _GEN_15256; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15258 = 10'h57 == _T_311[9:0] ? 4'hf : _GEN_15257; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15259 = 10'h58 == _T_311[9:0] ? 4'h3 : _GEN_15258; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15260 = 10'h59 == _T_311[9:0] ? 4'hf : _GEN_15259; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15261 = 10'h5a == _T_311[9:0] ? 4'h3 : _GEN_15260; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15262 = 10'h5b == _T_311[9:0] ? 4'h3 : _GEN_15261; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15263 = 10'h5c == _T_311[9:0] ? 4'h3 : _GEN_15262; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15264 = 10'h5d == _T_311[9:0] ? 4'h3 : _GEN_15263; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15265 = 10'h5e == _T_311[9:0] ? 4'h3 : _GEN_15264; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15266 = 10'h5f == _T_311[9:0] ? 4'h0 : _GEN_15265; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15267 = 10'h60 == _T_311[9:0] ? 4'h3 : _GEN_15266; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15268 = 10'h61 == _T_311[9:0] ? 4'h3 : _GEN_15267; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15269 = 10'h62 == _T_311[9:0] ? 4'h3 : _GEN_15268; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15270 = 10'h63 == _T_311[9:0] ? 4'h3 : _GEN_15269; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15271 = 10'h64 == _T_311[9:0] ? 4'h3 : _GEN_15270; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15272 = 10'h65 == _T_311[9:0] ? 4'hf : _GEN_15271; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15273 = 10'h66 == _T_311[9:0] ? 4'h3 : _GEN_15272; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15274 = 10'h67 == _T_311[9:0] ? 4'h3 : _GEN_15273; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15275 = 10'h68 == _T_311[9:0] ? 4'h3 : _GEN_15274; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15276 = 10'h69 == _T_311[9:0] ? 4'hf : _GEN_15275; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15277 = 10'h6a == _T_311[9:0] ? 4'h9 : _GEN_15276; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15278 = 10'h6b == _T_311[9:0] ? 4'h9 : _GEN_15277; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15279 = 10'h6c == _T_311[9:0] ? 4'h3 : _GEN_15278; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15280 = 10'h6d == _T_311[9:0] ? 4'h3 : _GEN_15279; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15281 = 10'h6e == _T_311[9:0] ? 4'h3 : _GEN_15280; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15282 = 10'h6f == _T_311[9:0] ? 4'h3 : _GEN_15281; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15283 = 10'h70 == _T_311[9:0] ? 4'h3 : _GEN_15282; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15284 = 10'h71 == _T_311[9:0] ? 4'h3 : _GEN_15283; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15285 = 10'h72 == _T_311[9:0] ? 4'h3 : _GEN_15284; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15286 = 10'h73 == _T_311[9:0] ? 4'h9 : _GEN_15285; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15287 = 10'h74 == _T_311[9:0] ? 4'hf : _GEN_15286; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15288 = 10'h75 == _T_311[9:0] ? 4'hf : _GEN_15287; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15289 = 10'h76 == _T_311[9:0] ? 4'hf : _GEN_15288; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15290 = 10'h77 == _T_311[9:0] ? 4'h3 : _GEN_15289; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15291 = 10'h78 == _T_311[9:0] ? 4'h3 : _GEN_15290; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15292 = 10'h79 == _T_311[9:0] ? 4'h3 : _GEN_15291; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15293 = 10'h7a == _T_311[9:0] ? 4'hf : _GEN_15292; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15294 = 10'h7b == _T_311[9:0] ? 4'h3 : _GEN_15293; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15295 = 10'h7c == _T_311[9:0] ? 4'h3 : _GEN_15294; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15296 = 10'h7d == _T_311[9:0] ? 4'h2 : _GEN_15295; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15297 = 10'h7e == _T_311[9:0] ? 4'h3 : _GEN_15296; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15298 = 10'h7f == _T_311[9:0] ? 4'h0 : _GEN_15297; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15299 = 10'h80 == _T_311[9:0] ? 4'h3 : _GEN_15298; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15300 = 10'h81 == _T_311[9:0] ? 4'h3 : _GEN_15299; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15301 = 10'h82 == _T_311[9:0] ? 4'h9 : _GEN_15300; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15302 = 10'h83 == _T_311[9:0] ? 4'hf : _GEN_15301; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15303 = 10'h84 == _T_311[9:0] ? 4'h2 : _GEN_15302; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15304 = 10'h85 == _T_311[9:0] ? 4'h9 : _GEN_15303; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15305 = 10'h86 == _T_311[9:0] ? 4'h9 : _GEN_15304; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15306 = 10'h87 == _T_311[9:0] ? 4'h3 : _GEN_15305; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15307 = 10'h88 == _T_311[9:0] ? 4'h3 : _GEN_15306; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15308 = 10'h89 == _T_311[9:0] ? 4'hf : _GEN_15307; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15309 = 10'h8a == _T_311[9:0] ? 4'hf : _GEN_15308; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15310 = 10'h8b == _T_311[9:0] ? 4'h9 : _GEN_15309; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15311 = 10'h8c == _T_311[9:0] ? 4'h9 : _GEN_15310; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15312 = 10'h8d == _T_311[9:0] ? 4'h9 : _GEN_15311; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15313 = 10'h8e == _T_311[9:0] ? 4'h9 : _GEN_15312; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15314 = 10'h8f == _T_311[9:0] ? 4'h9 : _GEN_15313; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15315 = 10'h90 == _T_311[9:0] ? 4'h9 : _GEN_15314; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15316 = 10'h91 == _T_311[9:0] ? 4'h9 : _GEN_15315; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15317 = 10'h92 == _T_311[9:0] ? 4'h9 : _GEN_15316; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15318 = 10'h93 == _T_311[9:0] ? 4'hf : _GEN_15317; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15319 = 10'h94 == _T_311[9:0] ? 4'hf : _GEN_15318; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15320 = 10'h95 == _T_311[9:0] ? 4'h3 : _GEN_15319; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15321 = 10'h96 == _T_311[9:0] ? 4'h3 : _GEN_15320; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15322 = 10'h97 == _T_311[9:0] ? 4'h3 : _GEN_15321; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15323 = 10'h98 == _T_311[9:0] ? 4'h9 : _GEN_15322; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15324 = 10'h99 == _T_311[9:0] ? 4'hf : _GEN_15323; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15325 = 10'h9a == _T_311[9:0] ? 4'h9 : _GEN_15324; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15326 = 10'h9b == _T_311[9:0] ? 4'h9 : _GEN_15325; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15327 = 10'h9c == _T_311[9:0] ? 4'h3 : _GEN_15326; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15328 = 10'h9d == _T_311[9:0] ? 4'h3 : _GEN_15327; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15329 = 10'h9e == _T_311[9:0] ? 4'h3 : _GEN_15328; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15330 = 10'h9f == _T_311[9:0] ? 4'h0 : _GEN_15329; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15331 = 10'ha0 == _T_311[9:0] ? 4'h3 : _GEN_15330; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15332 = 10'ha1 == _T_311[9:0] ? 4'h9 : _GEN_15331; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15333 = 10'ha2 == _T_311[9:0] ? 4'hf : _GEN_15332; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15334 = 10'ha3 == _T_311[9:0] ? 4'h3 : _GEN_15333; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15335 = 10'ha4 == _T_311[9:0] ? 4'h3 : _GEN_15334; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15336 = 10'ha5 == _T_311[9:0] ? 4'h3 : _GEN_15335; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15337 = 10'ha6 == _T_311[9:0] ? 4'h3 : _GEN_15336; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15338 = 10'ha7 == _T_311[9:0] ? 4'hf : _GEN_15337; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15339 = 10'ha8 == _T_311[9:0] ? 4'h3 : _GEN_15338; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15340 = 10'ha9 == _T_311[9:0] ? 4'h9 : _GEN_15339; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15341 = 10'haa == _T_311[9:0] ? 4'hf : _GEN_15340; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15342 = 10'hab == _T_311[9:0] ? 4'hf : _GEN_15341; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15343 = 10'hac == _T_311[9:0] ? 4'hf : _GEN_15342; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15344 = 10'had == _T_311[9:0] ? 4'hf : _GEN_15343; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15345 = 10'hae == _T_311[9:0] ? 4'hf : _GEN_15344; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15346 = 10'haf == _T_311[9:0] ? 4'hf : _GEN_15345; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15347 = 10'hb0 == _T_311[9:0] ? 4'hf : _GEN_15346; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15348 = 10'hb1 == _T_311[9:0] ? 4'hf : _GEN_15347; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15349 = 10'hb2 == _T_311[9:0] ? 4'hf : _GEN_15348; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15350 = 10'hb3 == _T_311[9:0] ? 4'hf : _GEN_15349; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15351 = 10'hb4 == _T_311[9:0] ? 4'h9 : _GEN_15350; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15352 = 10'hb5 == _T_311[9:0] ? 4'h9 : _GEN_15351; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15353 = 10'hb6 == _T_311[9:0] ? 4'h3 : _GEN_15352; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15354 = 10'hb7 == _T_311[9:0] ? 4'hf : _GEN_15353; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15355 = 10'hb8 == _T_311[9:0] ? 4'h3 : _GEN_15354; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15356 = 10'hb9 == _T_311[9:0] ? 4'h3 : _GEN_15355; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15357 = 10'hba == _T_311[9:0] ? 4'h3 : _GEN_15356; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15358 = 10'hbb == _T_311[9:0] ? 4'hf : _GEN_15357; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15359 = 10'hbc == _T_311[9:0] ? 4'h3 : _GEN_15358; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15360 = 10'hbd == _T_311[9:0] ? 4'h3 : _GEN_15359; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15361 = 10'hbe == _T_311[9:0] ? 4'h3 : _GEN_15360; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15362 = 10'hbf == _T_311[9:0] ? 4'h0 : _GEN_15361; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15363 = 10'hc0 == _T_311[9:0] ? 4'h3 : _GEN_15362; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15364 = 10'hc1 == _T_311[9:0] ? 4'h3 : _GEN_15363; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15365 = 10'hc2 == _T_311[9:0] ? 4'h3 : _GEN_15364; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15366 = 10'hc3 == _T_311[9:0] ? 4'h2 : _GEN_15365; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15367 = 10'hc4 == _T_311[9:0] ? 4'hf : _GEN_15366; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15368 = 10'hc5 == _T_311[9:0] ? 4'hf : _GEN_15367; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15369 = 10'hc6 == _T_311[9:0] ? 4'hf : _GEN_15368; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15370 = 10'hc7 == _T_311[9:0] ? 4'h3 : _GEN_15369; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15371 = 10'hc8 == _T_311[9:0] ? 4'h9 : _GEN_15370; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15372 = 10'hc9 == _T_311[9:0] ? 4'hf : _GEN_15371; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15373 = 10'hca == _T_311[9:0] ? 4'hf : _GEN_15372; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15374 = 10'hcb == _T_311[9:0] ? 4'hf : _GEN_15373; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15375 = 10'hcc == _T_311[9:0] ? 4'hf : _GEN_15374; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15376 = 10'hcd == _T_311[9:0] ? 4'hf : _GEN_15375; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15377 = 10'hce == _T_311[9:0] ? 4'hf : _GEN_15376; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15378 = 10'hcf == _T_311[9:0] ? 4'hf : _GEN_15377; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15379 = 10'hd0 == _T_311[9:0] ? 4'hf : _GEN_15378; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15380 = 10'hd1 == _T_311[9:0] ? 4'hf : _GEN_15379; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15381 = 10'hd2 == _T_311[9:0] ? 4'hf : _GEN_15380; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15382 = 10'hd3 == _T_311[9:0] ? 4'hf : _GEN_15381; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15383 = 10'hd4 == _T_311[9:0] ? 4'hf : _GEN_15382; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15384 = 10'hd5 == _T_311[9:0] ? 4'hf : _GEN_15383; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15385 = 10'hd6 == _T_311[9:0] ? 4'h9 : _GEN_15384; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15386 = 10'hd7 == _T_311[9:0] ? 4'h3 : _GEN_15385; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15387 = 10'hd8 == _T_311[9:0] ? 4'hf : _GEN_15386; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15388 = 10'hd9 == _T_311[9:0] ? 4'h3 : _GEN_15387; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15389 = 10'hda == _T_311[9:0] ? 4'h3 : _GEN_15388; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15390 = 10'hdb == _T_311[9:0] ? 4'h3 : _GEN_15389; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15391 = 10'hdc == _T_311[9:0] ? 4'h3 : _GEN_15390; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15392 = 10'hdd == _T_311[9:0] ? 4'h3 : _GEN_15391; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15393 = 10'hde == _T_311[9:0] ? 4'h2 : _GEN_15392; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15394 = 10'hdf == _T_311[9:0] ? 4'h0 : _GEN_15393; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15395 = 10'he0 == _T_311[9:0] ? 4'h3 : _GEN_15394; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15396 = 10'he1 == _T_311[9:0] ? 4'h3 : _GEN_15395; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15397 = 10'he2 == _T_311[9:0] ? 4'h3 : _GEN_15396; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15398 = 10'he3 == _T_311[9:0] ? 4'h3 : _GEN_15397; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15399 = 10'he4 == _T_311[9:0] ? 4'h3 : _GEN_15398; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15400 = 10'he5 == _T_311[9:0] ? 4'h3 : _GEN_15399; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15401 = 10'he6 == _T_311[9:0] ? 4'h3 : _GEN_15400; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15402 = 10'he7 == _T_311[9:0] ? 4'h9 : _GEN_15401; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15403 = 10'he8 == _T_311[9:0] ? 4'h9 : _GEN_15402; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15404 = 10'he9 == _T_311[9:0] ? 4'h9 : _GEN_15403; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15405 = 10'hea == _T_311[9:0] ? 4'hf : _GEN_15404; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15406 = 10'heb == _T_311[9:0] ? 4'hf : _GEN_15405; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15407 = 10'hec == _T_311[9:0] ? 4'hf : _GEN_15406; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15408 = 10'hed == _T_311[9:0] ? 4'hf : _GEN_15407; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15409 = 10'hee == _T_311[9:0] ? 4'hf : _GEN_15408; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15410 = 10'hef == _T_311[9:0] ? 4'hf : _GEN_15409; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15411 = 10'hf0 == _T_311[9:0] ? 4'hf : _GEN_15410; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15412 = 10'hf1 == _T_311[9:0] ? 4'hf : _GEN_15411; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15413 = 10'hf2 == _T_311[9:0] ? 4'hf : _GEN_15412; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15414 = 10'hf3 == _T_311[9:0] ? 4'hf : _GEN_15413; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15415 = 10'hf4 == _T_311[9:0] ? 4'hf : _GEN_15414; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15416 = 10'hf5 == _T_311[9:0] ? 4'h9 : _GEN_15415; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15417 = 10'hf6 == _T_311[9:0] ? 4'hf : _GEN_15416; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15418 = 10'hf7 == _T_311[9:0] ? 4'hf : _GEN_15417; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15419 = 10'hf8 == _T_311[9:0] ? 4'h9 : _GEN_15418; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15420 = 10'hf9 == _T_311[9:0] ? 4'hf : _GEN_15419; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15421 = 10'hfa == _T_311[9:0] ? 4'h3 : _GEN_15420; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15422 = 10'hfb == _T_311[9:0] ? 4'h3 : _GEN_15421; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15423 = 10'hfc == _T_311[9:0] ? 4'h3 : _GEN_15422; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15424 = 10'hfd == _T_311[9:0] ? 4'h3 : _GEN_15423; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15425 = 10'hfe == _T_311[9:0] ? 4'h3 : _GEN_15424; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15426 = 10'hff == _T_311[9:0] ? 4'h0 : _GEN_15425; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15427 = 10'h100 == _T_311[9:0] ? 4'h3 : _GEN_15426; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15428 = 10'h101 == _T_311[9:0] ? 4'hf : _GEN_15427; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15429 = 10'h102 == _T_311[9:0] ? 4'h3 : _GEN_15428; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15430 = 10'h103 == _T_311[9:0] ? 4'h3 : _GEN_15429; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15431 = 10'h104 == _T_311[9:0] ? 4'h3 : _GEN_15430; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15432 = 10'h105 == _T_311[9:0] ? 4'h3 : _GEN_15431; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15433 = 10'h106 == _T_311[9:0] ? 4'h3 : _GEN_15432; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15434 = 10'h107 == _T_311[9:0] ? 4'h3 : _GEN_15433; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15435 = 10'h108 == _T_311[9:0] ? 4'h9 : _GEN_15434; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15436 = 10'h109 == _T_311[9:0] ? 4'hf : _GEN_15435; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15437 = 10'h10a == _T_311[9:0] ? 4'hf : _GEN_15436; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15438 = 10'h10b == _T_311[9:0] ? 4'hf : _GEN_15437; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15439 = 10'h10c == _T_311[9:0] ? 4'hf : _GEN_15438; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15440 = 10'h10d == _T_311[9:0] ? 4'h0 : _GEN_15439; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15441 = 10'h10e == _T_311[9:0] ? 4'hf : _GEN_15440; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15442 = 10'h10f == _T_311[9:0] ? 4'hf : _GEN_15441; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15443 = 10'h110 == _T_311[9:0] ? 4'hf : _GEN_15442; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15444 = 10'h111 == _T_311[9:0] ? 4'h0 : _GEN_15443; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15445 = 10'h112 == _T_311[9:0] ? 4'hf : _GEN_15444; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15446 = 10'h113 == _T_311[9:0] ? 4'hf : _GEN_15445; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15447 = 10'h114 == _T_311[9:0] ? 4'hf : _GEN_15446; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15448 = 10'h115 == _T_311[9:0] ? 4'hf : _GEN_15447; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15449 = 10'h116 == _T_311[9:0] ? 4'h9 : _GEN_15448; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15450 = 10'h117 == _T_311[9:0] ? 4'h3 : _GEN_15449; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15451 = 10'h118 == _T_311[9:0] ? 4'h3 : _GEN_15450; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15452 = 10'h119 == _T_311[9:0] ? 4'h3 : _GEN_15451; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15453 = 10'h11a == _T_311[9:0] ? 4'hf : _GEN_15452; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15454 = 10'h11b == _T_311[9:0] ? 4'h3 : _GEN_15453; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15455 = 10'h11c == _T_311[9:0] ? 4'h3 : _GEN_15454; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15456 = 10'h11d == _T_311[9:0] ? 4'h2 : _GEN_15455; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15457 = 10'h11e == _T_311[9:0] ? 4'h3 : _GEN_15456; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15458 = 10'h11f == _T_311[9:0] ? 4'h0 : _GEN_15457; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15459 = 10'h120 == _T_311[9:0] ? 4'h3 : _GEN_15458; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15460 = 10'h121 == _T_311[9:0] ? 4'h3 : _GEN_15459; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15461 = 10'h122 == _T_311[9:0] ? 4'h3 : _GEN_15460; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15462 = 10'h123 == _T_311[9:0] ? 4'h3 : _GEN_15461; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15463 = 10'h124 == _T_311[9:0] ? 4'h3 : _GEN_15462; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15464 = 10'h125 == _T_311[9:0] ? 4'h3 : _GEN_15463; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15465 = 10'h126 == _T_311[9:0] ? 4'h3 : _GEN_15464; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15466 = 10'h127 == _T_311[9:0] ? 4'h9 : _GEN_15465; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15467 = 10'h128 == _T_311[9:0] ? 4'hf : _GEN_15466; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15468 = 10'h129 == _T_311[9:0] ? 4'h3 : _GEN_15467; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15469 = 10'h12a == _T_311[9:0] ? 4'h3 : _GEN_15468; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15470 = 10'h12b == _T_311[9:0] ? 4'hf : _GEN_15469; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15471 = 10'h12c == _T_311[9:0] ? 4'hf : _GEN_15470; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15472 = 10'h12d == _T_311[9:0] ? 4'hf : _GEN_15471; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15473 = 10'h12e == _T_311[9:0] ? 4'hf : _GEN_15472; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15474 = 10'h12f == _T_311[9:0] ? 4'hf : _GEN_15473; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15475 = 10'h130 == _T_311[9:0] ? 4'hf : _GEN_15474; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15476 = 10'h131 == _T_311[9:0] ? 4'hf : _GEN_15475; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15477 = 10'h132 == _T_311[9:0] ? 4'hf : _GEN_15476; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15478 = 10'h133 == _T_311[9:0] ? 4'hf : _GEN_15477; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15479 = 10'h134 == _T_311[9:0] ? 4'h3 : _GEN_15478; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15480 = 10'h135 == _T_311[9:0] ? 4'h3 : _GEN_15479; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15481 = 10'h136 == _T_311[9:0] ? 4'hf : _GEN_15480; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15482 = 10'h137 == _T_311[9:0] ? 4'h9 : _GEN_15481; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15483 = 10'h138 == _T_311[9:0] ? 4'h3 : _GEN_15482; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15484 = 10'h139 == _T_311[9:0] ? 4'h3 : _GEN_15483; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15485 = 10'h13a == _T_311[9:0] ? 4'h3 : _GEN_15484; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15486 = 10'h13b == _T_311[9:0] ? 4'h3 : _GEN_15485; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15487 = 10'h13c == _T_311[9:0] ? 4'h3 : _GEN_15486; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15488 = 10'h13d == _T_311[9:0] ? 4'h3 : _GEN_15487; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15489 = 10'h13e == _T_311[9:0] ? 4'h3 : _GEN_15488; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15490 = 10'h13f == _T_311[9:0] ? 4'h0 : _GEN_15489; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15491 = 10'h140 == _T_311[9:0] ? 4'h3 : _GEN_15490; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15492 = 10'h141 == _T_311[9:0] ? 4'h3 : _GEN_15491; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15493 = 10'h142 == _T_311[9:0] ? 4'h2 : _GEN_15492; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15494 = 10'h143 == _T_311[9:0] ? 4'h3 : _GEN_15493; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15495 = 10'h144 == _T_311[9:0] ? 4'h3 : _GEN_15494; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15496 = 10'h145 == _T_311[9:0] ? 4'h3 : _GEN_15495; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15497 = 10'h146 == _T_311[9:0] ? 4'h9 : _GEN_15496; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15498 = 10'h147 == _T_311[9:0] ? 4'hf : _GEN_15497; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15499 = 10'h148 == _T_311[9:0] ? 4'h3 : _GEN_15498; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15500 = 10'h149 == _T_311[9:0] ? 4'h3 : _GEN_15499; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15501 = 10'h14a == _T_311[9:0] ? 4'h3 : _GEN_15500; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15502 = 10'h14b == _T_311[9:0] ? 4'h3 : _GEN_15501; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15503 = 10'h14c == _T_311[9:0] ? 4'h3 : _GEN_15502; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15504 = 10'h14d == _T_311[9:0] ? 4'h3 : _GEN_15503; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15505 = 10'h14e == _T_311[9:0] ? 4'h3 : _GEN_15504; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15506 = 10'h14f == _T_311[9:0] ? 4'h3 : _GEN_15505; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15507 = 10'h150 == _T_311[9:0] ? 4'h3 : _GEN_15506; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15508 = 10'h151 == _T_311[9:0] ? 4'h3 : _GEN_15507; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15509 = 10'h152 == _T_311[9:0] ? 4'h3 : _GEN_15508; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15510 = 10'h153 == _T_311[9:0] ? 4'h3 : _GEN_15509; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15511 = 10'h154 == _T_311[9:0] ? 4'h3 : _GEN_15510; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15512 = 10'h155 == _T_311[9:0] ? 4'h3 : _GEN_15511; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15513 = 10'h156 == _T_311[9:0] ? 4'h3 : _GEN_15512; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15514 = 10'h157 == _T_311[9:0] ? 4'hf : _GEN_15513; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15515 = 10'h158 == _T_311[9:0] ? 4'h3 : _GEN_15514; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15516 = 10'h159 == _T_311[9:0] ? 4'h3 : _GEN_15515; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15517 = 10'h15a == _T_311[9:0] ? 4'h3 : _GEN_15516; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15518 = 10'h15b == _T_311[9:0] ? 4'h3 : _GEN_15517; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15519 = 10'h15c == _T_311[9:0] ? 4'h3 : _GEN_15518; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15520 = 10'h15d == _T_311[9:0] ? 4'h3 : _GEN_15519; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15521 = 10'h15e == _T_311[9:0] ? 4'h2 : _GEN_15520; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15522 = 10'h15f == _T_311[9:0] ? 4'h0 : _GEN_15521; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15523 = 10'h160 == _T_311[9:0] ? 4'h3 : _GEN_15522; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15524 = 10'h161 == _T_311[9:0] ? 4'h3 : _GEN_15523; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15525 = 10'h162 == _T_311[9:0] ? 4'h3 : _GEN_15524; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15526 = 10'h163 == _T_311[9:0] ? 4'h2 : _GEN_15525; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15527 = 10'h164 == _T_311[9:0] ? 4'h3 : _GEN_15526; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15528 = 10'h165 == _T_311[9:0] ? 4'h9 : _GEN_15527; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15529 = 10'h166 == _T_311[9:0] ? 4'hf : _GEN_15528; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15530 = 10'h167 == _T_311[9:0] ? 4'hf : _GEN_15529; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15531 = 10'h168 == _T_311[9:0] ? 4'hd : _GEN_15530; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15532 = 10'h169 == _T_311[9:0] ? 4'h9 : _GEN_15531; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15533 = 10'h16a == _T_311[9:0] ? 4'hd : _GEN_15532; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15534 = 10'h16b == _T_311[9:0] ? 4'hd : _GEN_15533; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15535 = 10'h16c == _T_311[9:0] ? 4'h3 : _GEN_15534; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15536 = 10'h16d == _T_311[9:0] ? 4'h3 : _GEN_15535; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15537 = 10'h16e == _T_311[9:0] ? 4'h3 : _GEN_15536; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15538 = 10'h16f == _T_311[9:0] ? 4'h3 : _GEN_15537; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15539 = 10'h170 == _T_311[9:0] ? 4'h3 : _GEN_15538; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15540 = 10'h171 == _T_311[9:0] ? 4'h3 : _GEN_15539; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15541 = 10'h172 == _T_311[9:0] ? 4'h3 : _GEN_15540; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15542 = 10'h173 == _T_311[9:0] ? 4'h3 : _GEN_15541; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15543 = 10'h174 == _T_311[9:0] ? 4'h3 : _GEN_15542; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15544 = 10'h175 == _T_311[9:0] ? 4'h3 : _GEN_15543; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15545 = 10'h176 == _T_311[9:0] ? 4'hf : _GEN_15544; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15546 = 10'h177 == _T_311[9:0] ? 4'hf : _GEN_15545; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15547 = 10'h178 == _T_311[9:0] ? 4'h9 : _GEN_15546; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15548 = 10'h179 == _T_311[9:0] ? 4'h3 : _GEN_15547; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15549 = 10'h17a == _T_311[9:0] ? 4'h3 : _GEN_15548; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15550 = 10'h17b == _T_311[9:0] ? 4'h3 : _GEN_15549; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15551 = 10'h17c == _T_311[9:0] ? 4'h3 : _GEN_15550; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15552 = 10'h17d == _T_311[9:0] ? 4'h2 : _GEN_15551; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15553 = 10'h17e == _T_311[9:0] ? 4'h3 : _GEN_15552; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15554 = 10'h17f == _T_311[9:0] ? 4'h0 : _GEN_15553; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15555 = 10'h180 == _T_311[9:0] ? 4'hd : _GEN_15554; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15556 = 10'h181 == _T_311[9:0] ? 4'hd : _GEN_15555; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15557 = 10'h182 == _T_311[9:0] ? 4'hd : _GEN_15556; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15558 = 10'h183 == _T_311[9:0] ? 4'hd : _GEN_15557; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15559 = 10'h184 == _T_311[9:0] ? 4'h3 : _GEN_15558; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15560 = 10'h185 == _T_311[9:0] ? 4'h9 : _GEN_15559; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15561 = 10'h186 == _T_311[9:0] ? 4'hb : _GEN_15560; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15562 = 10'h187 == _T_311[9:0] ? 4'hf : _GEN_15561; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15563 = 10'h188 == _T_311[9:0] ? 4'hd : _GEN_15562; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15564 = 10'h189 == _T_311[9:0] ? 4'hd : _GEN_15563; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15565 = 10'h18a == _T_311[9:0] ? 4'hd : _GEN_15564; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15566 = 10'h18b == _T_311[9:0] ? 4'hd : _GEN_15565; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15567 = 10'h18c == _T_311[9:0] ? 4'hd : _GEN_15566; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15568 = 10'h18d == _T_311[9:0] ? 4'hd : _GEN_15567; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15569 = 10'h18e == _T_311[9:0] ? 4'hd : _GEN_15568; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15570 = 10'h18f == _T_311[9:0] ? 4'hd : _GEN_15569; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15571 = 10'h190 == _T_311[9:0] ? 4'hd : _GEN_15570; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15572 = 10'h191 == _T_311[9:0] ? 4'hd : _GEN_15571; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15573 = 10'h192 == _T_311[9:0] ? 4'h9 : _GEN_15572; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15574 = 10'h193 == _T_311[9:0] ? 4'hd : _GEN_15573; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15575 = 10'h194 == _T_311[9:0] ? 4'hd : _GEN_15574; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15576 = 10'h195 == _T_311[9:0] ? 4'hd : _GEN_15575; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15577 = 10'h196 == _T_311[9:0] ? 4'hf : _GEN_15576; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15578 = 10'h197 == _T_311[9:0] ? 4'h3 : _GEN_15577; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15579 = 10'h198 == _T_311[9:0] ? 4'h9 : _GEN_15578; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15580 = 10'h199 == _T_311[9:0] ? 4'h3 : _GEN_15579; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15581 = 10'h19a == _T_311[9:0] ? 4'h3 : _GEN_15580; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15582 = 10'h19b == _T_311[9:0] ? 4'h3 : _GEN_15581; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15583 = 10'h19c == _T_311[9:0] ? 4'h3 : _GEN_15582; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15584 = 10'h19d == _T_311[9:0] ? 4'h3 : _GEN_15583; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15585 = 10'h19e == _T_311[9:0] ? 4'h3 : _GEN_15584; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15586 = 10'h19f == _T_311[9:0] ? 4'h0 : _GEN_15585; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15587 = 10'h1a0 == _T_311[9:0] ? 4'hd : _GEN_15586; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15588 = 10'h1a1 == _T_311[9:0] ? 4'hd : _GEN_15587; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15589 = 10'h1a2 == _T_311[9:0] ? 4'h9 : _GEN_15588; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15590 = 10'h1a3 == _T_311[9:0] ? 4'hd : _GEN_15589; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15591 = 10'h1a4 == _T_311[9:0] ? 4'h3 : _GEN_15590; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15592 = 10'h1a5 == _T_311[9:0] ? 4'hf : _GEN_15591; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15593 = 10'h1a6 == _T_311[9:0] ? 4'hd : _GEN_15592; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15594 = 10'h1a7 == _T_311[9:0] ? 4'hf : _GEN_15593; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15595 = 10'h1a8 == _T_311[9:0] ? 4'hb : _GEN_15594; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15596 = 10'h1a9 == _T_311[9:0] ? 4'hd : _GEN_15595; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15597 = 10'h1aa == _T_311[9:0] ? 4'hd : _GEN_15596; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15598 = 10'h1ab == _T_311[9:0] ? 4'h9 : _GEN_15597; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15599 = 10'h1ac == _T_311[9:0] ? 4'hd : _GEN_15598; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15600 = 10'h1ad == _T_311[9:0] ? 4'hd : _GEN_15599; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15601 = 10'h1ae == _T_311[9:0] ? 4'hd : _GEN_15600; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15602 = 10'h1af == _T_311[9:0] ? 4'hd : _GEN_15601; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15603 = 10'h1b0 == _T_311[9:0] ? 4'hd : _GEN_15602; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15604 = 10'h1b1 == _T_311[9:0] ? 4'hd : _GEN_15603; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15605 = 10'h1b2 == _T_311[9:0] ? 4'hd : _GEN_15604; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15606 = 10'h1b3 == _T_311[9:0] ? 4'hd : _GEN_15605; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15607 = 10'h1b4 == _T_311[9:0] ? 4'hd : _GEN_15606; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15608 = 10'h1b5 == _T_311[9:0] ? 4'hd : _GEN_15607; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15609 = 10'h1b6 == _T_311[9:0] ? 4'hf : _GEN_15608; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15610 = 10'h1b7 == _T_311[9:0] ? 4'hd : _GEN_15609; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15611 = 10'h1b8 == _T_311[9:0] ? 4'hf : _GEN_15610; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15612 = 10'h1b9 == _T_311[9:0] ? 4'hd : _GEN_15611; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15613 = 10'h1ba == _T_311[9:0] ? 4'hd : _GEN_15612; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15614 = 10'h1bb == _T_311[9:0] ? 4'hd : _GEN_15613; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15615 = 10'h1bc == _T_311[9:0] ? 4'h2 : _GEN_15614; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15616 = 10'h1bd == _T_311[9:0] ? 4'h3 : _GEN_15615; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15617 = 10'h1be == _T_311[9:0] ? 4'hd : _GEN_15616; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15618 = 10'h1bf == _T_311[9:0] ? 4'h0 : _GEN_15617; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15619 = 10'h1c0 == _T_311[9:0] ? 4'hd : _GEN_15618; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15620 = 10'h1c1 == _T_311[9:0] ? 4'hd : _GEN_15619; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15621 = 10'h1c2 == _T_311[9:0] ? 4'hd : _GEN_15620; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15622 = 10'h1c3 == _T_311[9:0] ? 4'h2 : _GEN_15621; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15623 = 10'h1c4 == _T_311[9:0] ? 4'h2 : _GEN_15622; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15624 = 10'h1c5 == _T_311[9:0] ? 4'hd : _GEN_15623; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15625 = 10'h1c6 == _T_311[9:0] ? 4'hd : _GEN_15624; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15626 = 10'h1c7 == _T_311[9:0] ? 4'hd : _GEN_15625; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15627 = 10'h1c8 == _T_311[9:0] ? 4'hd : _GEN_15626; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15628 = 10'h1c9 == _T_311[9:0] ? 4'hb : _GEN_15627; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15629 = 10'h1ca == _T_311[9:0] ? 4'hb : _GEN_15628; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15630 = 10'h1cb == _T_311[9:0] ? 4'hb : _GEN_15629; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15631 = 10'h1cc == _T_311[9:0] ? 4'hb : _GEN_15630; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15632 = 10'h1cd == _T_311[9:0] ? 4'hb : _GEN_15631; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15633 = 10'h1ce == _T_311[9:0] ? 4'hb : _GEN_15632; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15634 = 10'h1cf == _T_311[9:0] ? 4'hb : _GEN_15633; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15635 = 10'h1d0 == _T_311[9:0] ? 4'hb : _GEN_15634; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15636 = 10'h1d1 == _T_311[9:0] ? 4'hb : _GEN_15635; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15637 = 10'h1d2 == _T_311[9:0] ? 4'hb : _GEN_15636; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15638 = 10'h1d3 == _T_311[9:0] ? 4'hb : _GEN_15637; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15639 = 10'h1d4 == _T_311[9:0] ? 4'hb : _GEN_15638; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15640 = 10'h1d5 == _T_311[9:0] ? 4'hb : _GEN_15639; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15641 = 10'h1d6 == _T_311[9:0] ? 4'hd : _GEN_15640; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15642 = 10'h1d7 == _T_311[9:0] ? 4'hd : _GEN_15641; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15643 = 10'h1d8 == _T_311[9:0] ? 4'hd : _GEN_15642; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15644 = 10'h1d9 == _T_311[9:0] ? 4'hd : _GEN_15643; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15645 = 10'h1da == _T_311[9:0] ? 4'hd : _GEN_15644; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15646 = 10'h1db == _T_311[9:0] ? 4'hd : _GEN_15645; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15647 = 10'h1dc == _T_311[9:0] ? 4'hd : _GEN_15646; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15648 = 10'h1dd == _T_311[9:0] ? 4'h3 : _GEN_15647; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15649 = 10'h1de == _T_311[9:0] ? 4'hd : _GEN_15648; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15650 = 10'h1df == _T_311[9:0] ? 4'h0 : _GEN_15649; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15651 = 10'h1e0 == _T_311[9:0] ? 4'h9 : _GEN_15650; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15652 = 10'h1e1 == _T_311[9:0] ? 4'hd : _GEN_15651; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15653 = 10'h1e2 == _T_311[9:0] ? 4'h2 : _GEN_15652; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15654 = 10'h1e3 == _T_311[9:0] ? 4'h2 : _GEN_15653; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15655 = 10'h1e4 == _T_311[9:0] ? 4'hd : _GEN_15654; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15656 = 10'h1e5 == _T_311[9:0] ? 4'hd : _GEN_15655; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15657 = 10'h1e6 == _T_311[9:0] ? 4'hd : _GEN_15656; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15658 = 10'h1e7 == _T_311[9:0] ? 4'hd : _GEN_15657; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15659 = 10'h1e8 == _T_311[9:0] ? 4'hb : _GEN_15658; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15660 = 10'h1e9 == _T_311[9:0] ? 4'hd : _GEN_15659; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15661 = 10'h1ea == _T_311[9:0] ? 4'hd : _GEN_15660; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15662 = 10'h1eb == _T_311[9:0] ? 4'hb : _GEN_15661; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15663 = 10'h1ec == _T_311[9:0] ? 4'hd : _GEN_15662; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15664 = 10'h1ed == _T_311[9:0] ? 4'hb : _GEN_15663; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15665 = 10'h1ee == _T_311[9:0] ? 4'hd : _GEN_15664; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15666 = 10'h1ef == _T_311[9:0] ? 4'hb : _GEN_15665; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15667 = 10'h1f0 == _T_311[9:0] ? 4'hd : _GEN_15666; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15668 = 10'h1f1 == _T_311[9:0] ? 4'hb : _GEN_15667; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15669 = 10'h1f2 == _T_311[9:0] ? 4'hb : _GEN_15668; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15670 = 10'h1f3 == _T_311[9:0] ? 4'hd : _GEN_15669; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15671 = 10'h1f4 == _T_311[9:0] ? 4'hb : _GEN_15670; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15672 = 10'h1f5 == _T_311[9:0] ? 4'hb : _GEN_15671; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15673 = 10'h1f6 == _T_311[9:0] ? 4'hd : _GEN_15672; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15674 = 10'h1f7 == _T_311[9:0] ? 4'hd : _GEN_15673; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15675 = 10'h1f8 == _T_311[9:0] ? 4'hd : _GEN_15674; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15676 = 10'h1f9 == _T_311[9:0] ? 4'hd : _GEN_15675; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15677 = 10'h1fa == _T_311[9:0] ? 4'h9 : _GEN_15676; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15678 = 10'h1fb == _T_311[9:0] ? 4'hd : _GEN_15677; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15679 = 10'h1fc == _T_311[9:0] ? 4'hd : _GEN_15678; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15680 = 10'h1fd == _T_311[9:0] ? 4'h2 : _GEN_15679; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15681 = 10'h1fe == _T_311[9:0] ? 4'hd : _GEN_15680; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15682 = 10'h1ff == _T_311[9:0] ? 4'h0 : _GEN_15681; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15683 = 10'h200 == _T_311[9:0] ? 4'hd : _GEN_15682; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15684 = 10'h201 == _T_311[9:0] ? 4'hd : _GEN_15683; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15685 = 10'h202 == _T_311[9:0] ? 4'h3 : _GEN_15684; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15686 = 10'h203 == _T_311[9:0] ? 4'hd : _GEN_15685; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15687 = 10'h204 == _T_311[9:0] ? 4'hd : _GEN_15686; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15688 = 10'h205 == _T_311[9:0] ? 4'hd : _GEN_15687; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15689 = 10'h206 == _T_311[9:0] ? 4'hb : _GEN_15688; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15690 = 10'h207 == _T_311[9:0] ? 4'hb : _GEN_15689; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15691 = 10'h208 == _T_311[9:0] ? 4'hd : _GEN_15690; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15692 = 10'h209 == _T_311[9:0] ? 4'hd : _GEN_15691; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15693 = 10'h20a == _T_311[9:0] ? 4'hd : _GEN_15692; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15694 = 10'h20b == _T_311[9:0] ? 4'hb : _GEN_15693; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15695 = 10'h20c == _T_311[9:0] ? 4'hd : _GEN_15694; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15696 = 10'h20d == _T_311[9:0] ? 4'hb : _GEN_15695; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15697 = 10'h20e == _T_311[9:0] ? 4'hd : _GEN_15696; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15698 = 10'h20f == _T_311[9:0] ? 4'hb : _GEN_15697; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15699 = 10'h210 == _T_311[9:0] ? 4'hd : _GEN_15698; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15700 = 10'h211 == _T_311[9:0] ? 4'hd : _GEN_15699; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15701 = 10'h212 == _T_311[9:0] ? 4'hb : _GEN_15700; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15702 = 10'h213 == _T_311[9:0] ? 4'hb : _GEN_15701; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15703 = 10'h214 == _T_311[9:0] ? 4'hb : _GEN_15702; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15704 = 10'h215 == _T_311[9:0] ? 4'hd : _GEN_15703; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15705 = 10'h216 == _T_311[9:0] ? 4'hd : _GEN_15704; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15706 = 10'h217 == _T_311[9:0] ? 4'hd : _GEN_15705; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15707 = 10'h218 == _T_311[9:0] ? 4'hd : _GEN_15706; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15708 = 10'h219 == _T_311[9:0] ? 4'hd : _GEN_15707; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15709 = 10'h21a == _T_311[9:0] ? 4'hd : _GEN_15708; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15710 = 10'h21b == _T_311[9:0] ? 4'hd : _GEN_15709; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15711 = 10'h21c == _T_311[9:0] ? 4'h3 : _GEN_15710; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15712 = 10'h21d == _T_311[9:0] ? 4'h2 : _GEN_15711; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15713 = 10'h21e == _T_311[9:0] ? 4'hd : _GEN_15712; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15714 = 10'h21f == _T_311[9:0] ? 4'h0 : _GEN_15713; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15715 = 10'h220 == _T_311[9:0] ? 4'h0 : _GEN_15714; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15716 = 10'h221 == _T_311[9:0] ? 4'h0 : _GEN_15715; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15717 = 10'h222 == _T_311[9:0] ? 4'h0 : _GEN_15716; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15718 = 10'h223 == _T_311[9:0] ? 4'h0 : _GEN_15717; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15719 = 10'h224 == _T_311[9:0] ? 4'h0 : _GEN_15718; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15720 = 10'h225 == _T_311[9:0] ? 4'h0 : _GEN_15719; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15721 = 10'h226 == _T_311[9:0] ? 4'h0 : _GEN_15720; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15722 = 10'h227 == _T_311[9:0] ? 4'h0 : _GEN_15721; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15723 = 10'h228 == _T_311[9:0] ? 4'h0 : _GEN_15722; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15724 = 10'h229 == _T_311[9:0] ? 4'h0 : _GEN_15723; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15725 = 10'h22a == _T_311[9:0] ? 4'h0 : _GEN_15724; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15726 = 10'h22b == _T_311[9:0] ? 4'h0 : _GEN_15725; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15727 = 10'h22c == _T_311[9:0] ? 4'h0 : _GEN_15726; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15728 = 10'h22d == _T_311[9:0] ? 4'h0 : _GEN_15727; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15729 = 10'h22e == _T_311[9:0] ? 4'h0 : _GEN_15728; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15730 = 10'h22f == _T_311[9:0] ? 4'h0 : _GEN_15729; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15731 = 10'h230 == _T_311[9:0] ? 4'h0 : _GEN_15730; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15732 = 10'h231 == _T_311[9:0] ? 4'h0 : _GEN_15731; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15733 = 10'h232 == _T_311[9:0] ? 4'h0 : _GEN_15732; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15734 = 10'h233 == _T_311[9:0] ? 4'h0 : _GEN_15733; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15735 = 10'h234 == _T_311[9:0] ? 4'h0 : _GEN_15734; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15736 = 10'h235 == _T_311[9:0] ? 4'h0 : _GEN_15735; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15737 = 10'h236 == _T_311[9:0] ? 4'h0 : _GEN_15736; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15738 = 10'h237 == _T_311[9:0] ? 4'h0 : _GEN_15737; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15739 = 10'h238 == _T_311[9:0] ? 4'h0 : _GEN_15738; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15740 = 10'h239 == _T_311[9:0] ? 4'h0 : _GEN_15739; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15741 = 10'h23a == _T_311[9:0] ? 4'h0 : _GEN_15740; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15742 = 10'h23b == _T_311[9:0] ? 4'h0 : _GEN_15741; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15743 = 10'h23c == _T_311[9:0] ? 4'h0 : _GEN_15742; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15744 = 10'h23d == _T_311[9:0] ? 4'h0 : _GEN_15743; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15745 = 10'h23e == _T_311[9:0] ? 4'h0 : _GEN_15744; // @[Filter.scala 191:142]
  wire [3:0] _GEN_15746 = 10'h23f == _T_311[9:0] ? 4'h0 : _GEN_15745; // @[Filter.scala 191:142]
  wire [7:0] _T_325 = _GEN_15746 * 4'ha; // @[Filter.scala 191:142]
  wire [10:0] _GEN_28351 = {{3'd0}, _T_325}; // @[Filter.scala 191:109]
  wire [10:0] _T_327 = _T_320 + _GEN_28351; // @[Filter.scala 191:109]
  wire [10:0] _T_328 = _T_327 / 11'h64; // @[Filter.scala 191:150]
  wire  _T_330 = _T_301 >= 6'h20; // @[Filter.scala 194:31]
  wire  _T_334 = _T_308 >= 32'h12; // @[Filter.scala 194:63]
  wire  _T_335 = _T_330 | _T_334; // @[Filter.scala 194:58]
  wire [10:0] _GEN_16323 = io_SPI_distort ? _T_328 : {{7'd0}, _GEN_14594}; // @[Filter.scala 196:35]
  wire [10:0] _GEN_16324 = _T_335 ? 11'h0 : _GEN_16323; // @[Filter.scala 194:80]
  wire [10:0] _GEN_16901 = io_SPI_distort ? _T_328 : {{7'd0}, _GEN_15170}; // @[Filter.scala 196:35]
  wire [10:0] _GEN_16902 = _T_335 ? 11'h0 : _GEN_16901; // @[Filter.scala 194:80]
  wire [10:0] _GEN_17479 = io_SPI_distort ? _T_328 : {{7'd0}, _GEN_15746}; // @[Filter.scala 196:35]
  wire [10:0] _GEN_17480 = _T_335 ? 11'h0 : _GEN_17479; // @[Filter.scala 194:80]
  wire [31:0] _T_363 = pixelIndex + 32'h5; // @[Filter.scala 189:31]
  wire [31:0] _GEN_5 = _T_363 % 32'h20; // @[Filter.scala 189:38]
  wire [5:0] _T_364 = _GEN_5[5:0]; // @[Filter.scala 189:38]
  wire [5:0] _T_366 = _T_364 + _GEN_28295; // @[Filter.scala 189:53]
  wire [5:0] _T_368 = _T_366 - 6'h1; // @[Filter.scala 189:69]
  wire [31:0] _T_371 = _T_363 / 32'h20; // @[Filter.scala 190:38]
  wire [31:0] _T_373 = _T_371 + _GEN_28296; // @[Filter.scala 190:53]
  wire [31:0] _T_375 = _T_373 - 32'h1; // @[Filter.scala 190:69]
  wire [37:0] _T_376 = _T_375 * 32'h20; // @[Filter.scala 191:42]
  wire [37:0] _GEN_28357 = {{32'd0}, _T_368}; // @[Filter.scala 191:57]
  wire [37:0] _T_378 = _T_376 + _GEN_28357; // @[Filter.scala 191:57]
  wire [3:0] _GEN_17484 = 10'h3 == _T_378[9:0] ? 4'h3 : 4'ha; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17485 = 10'h4 == _T_378[9:0] ? 4'ha : _GEN_17484; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17486 = 10'h5 == _T_378[9:0] ? 4'ha : _GEN_17485; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17487 = 10'h6 == _T_378[9:0] ? 4'ha : _GEN_17486; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17488 = 10'h7 == _T_378[9:0] ? 4'ha : _GEN_17487; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17489 = 10'h8 == _T_378[9:0] ? 4'ha : _GEN_17488; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17490 = 10'h9 == _T_378[9:0] ? 4'ha : _GEN_17489; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17491 = 10'ha == _T_378[9:0] ? 4'ha : _GEN_17490; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17492 = 10'hb == _T_378[9:0] ? 4'ha : _GEN_17491; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17493 = 10'hc == _T_378[9:0] ? 4'ha : _GEN_17492; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17494 = 10'hd == _T_378[9:0] ? 4'ha : _GEN_17493; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17495 = 10'he == _T_378[9:0] ? 4'ha : _GEN_17494; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17496 = 10'hf == _T_378[9:0] ? 4'ha : _GEN_17495; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17497 = 10'h10 == _T_378[9:0] ? 4'ha : _GEN_17496; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17498 = 10'h11 == _T_378[9:0] ? 4'ha : _GEN_17497; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17499 = 10'h12 == _T_378[9:0] ? 4'ha : _GEN_17498; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17500 = 10'h13 == _T_378[9:0] ? 4'ha : _GEN_17499; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17501 = 10'h14 == _T_378[9:0] ? 4'ha : _GEN_17500; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17502 = 10'h15 == _T_378[9:0] ? 4'ha : _GEN_17501; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17503 = 10'h16 == _T_378[9:0] ? 4'ha : _GEN_17502; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17504 = 10'h17 == _T_378[9:0] ? 4'ha : _GEN_17503; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17505 = 10'h18 == _T_378[9:0] ? 4'ha : _GEN_17504; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17506 = 10'h19 == _T_378[9:0] ? 4'ha : _GEN_17505; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17507 = 10'h1a == _T_378[9:0] ? 4'ha : _GEN_17506; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17508 = 10'h1b == _T_378[9:0] ? 4'ha : _GEN_17507; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17509 = 10'h1c == _T_378[9:0] ? 4'ha : _GEN_17508; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17510 = 10'h1d == _T_378[9:0] ? 4'ha : _GEN_17509; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17511 = 10'h1e == _T_378[9:0] ? 4'ha : _GEN_17510; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17512 = 10'h1f == _T_378[9:0] ? 4'h0 : _GEN_17511; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17513 = 10'h20 == _T_378[9:0] ? 4'ha : _GEN_17512; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17514 = 10'h21 == _T_378[9:0] ? 4'ha : _GEN_17513; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17515 = 10'h22 == _T_378[9:0] ? 4'ha : _GEN_17514; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17516 = 10'h23 == _T_378[9:0] ? 4'h3 : _GEN_17515; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17517 = 10'h24 == _T_378[9:0] ? 4'ha : _GEN_17516; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17518 = 10'h25 == _T_378[9:0] ? 4'ha : _GEN_17517; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17519 = 10'h26 == _T_378[9:0] ? 4'ha : _GEN_17518; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17520 = 10'h27 == _T_378[9:0] ? 4'h1 : _GEN_17519; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17521 = 10'h28 == _T_378[9:0] ? 4'h1 : _GEN_17520; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17522 = 10'h29 == _T_378[9:0] ? 4'ha : _GEN_17521; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17523 = 10'h2a == _T_378[9:0] ? 4'ha : _GEN_17522; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17524 = 10'h2b == _T_378[9:0] ? 4'ha : _GEN_17523; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17525 = 10'h2c == _T_378[9:0] ? 4'ha : _GEN_17524; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17526 = 10'h2d == _T_378[9:0] ? 4'ha : _GEN_17525; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17527 = 10'h2e == _T_378[9:0] ? 4'ha : _GEN_17526; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17528 = 10'h2f == _T_378[9:0] ? 4'ha : _GEN_17527; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17529 = 10'h30 == _T_378[9:0] ? 4'ha : _GEN_17528; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17530 = 10'h31 == _T_378[9:0] ? 4'ha : _GEN_17529; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17531 = 10'h32 == _T_378[9:0] ? 4'ha : _GEN_17530; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17532 = 10'h33 == _T_378[9:0] ? 4'ha : _GEN_17531; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17533 = 10'h34 == _T_378[9:0] ? 4'ha : _GEN_17532; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17534 = 10'h35 == _T_378[9:0] ? 4'ha : _GEN_17533; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17535 = 10'h36 == _T_378[9:0] ? 4'ha : _GEN_17534; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17536 = 10'h37 == _T_378[9:0] ? 4'h1 : _GEN_17535; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17537 = 10'h38 == _T_378[9:0] ? 4'h1 : _GEN_17536; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17538 = 10'h39 == _T_378[9:0] ? 4'ha : _GEN_17537; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17539 = 10'h3a == _T_378[9:0] ? 4'ha : _GEN_17538; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17540 = 10'h3b == _T_378[9:0] ? 4'ha : _GEN_17539; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17541 = 10'h3c == _T_378[9:0] ? 4'ha : _GEN_17540; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17542 = 10'h3d == _T_378[9:0] ? 4'h3 : _GEN_17541; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17543 = 10'h3e == _T_378[9:0] ? 4'ha : _GEN_17542; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17544 = 10'h3f == _T_378[9:0] ? 4'h0 : _GEN_17543; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17545 = 10'h40 == _T_378[9:0] ? 4'ha : _GEN_17544; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17546 = 10'h41 == _T_378[9:0] ? 4'ha : _GEN_17545; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17547 = 10'h42 == _T_378[9:0] ? 4'ha : _GEN_17546; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17548 = 10'h43 == _T_378[9:0] ? 4'h2 : _GEN_17547; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17549 = 10'h44 == _T_378[9:0] ? 4'h3 : _GEN_17548; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17550 = 10'h45 == _T_378[9:0] ? 4'h0 : _GEN_17549; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17551 = 10'h46 == _T_378[9:0] ? 4'h0 : _GEN_17550; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17552 = 10'h47 == _T_378[9:0] ? 4'h0 : _GEN_17551; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17553 = 10'h48 == _T_378[9:0] ? 4'h0 : _GEN_17552; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17554 = 10'h49 == _T_378[9:0] ? 4'ha : _GEN_17553; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17555 = 10'h4a == _T_378[9:0] ? 4'ha : _GEN_17554; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17556 = 10'h4b == _T_378[9:0] ? 4'ha : _GEN_17555; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17557 = 10'h4c == _T_378[9:0] ? 4'ha : _GEN_17556; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17558 = 10'h4d == _T_378[9:0] ? 4'ha : _GEN_17557; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17559 = 10'h4e == _T_378[9:0] ? 4'ha : _GEN_17558; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17560 = 10'h4f == _T_378[9:0] ? 4'ha : _GEN_17559; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17561 = 10'h50 == _T_378[9:0] ? 4'ha : _GEN_17560; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17562 = 10'h51 == _T_378[9:0] ? 4'ha : _GEN_17561; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17563 = 10'h52 == _T_378[9:0] ? 4'ha : _GEN_17562; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17564 = 10'h53 == _T_378[9:0] ? 4'ha : _GEN_17563; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17565 = 10'h54 == _T_378[9:0] ? 4'h1 : _GEN_17564; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17566 = 10'h55 == _T_378[9:0] ? 4'h1 : _GEN_17565; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17567 = 10'h56 == _T_378[9:0] ? 4'h1 : _GEN_17566; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17568 = 10'h57 == _T_378[9:0] ? 4'h0 : _GEN_17567; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17569 = 10'h58 == _T_378[9:0] ? 4'ha : _GEN_17568; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17570 = 10'h59 == _T_378[9:0] ? 4'h0 : _GEN_17569; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17571 = 10'h5a == _T_378[9:0] ? 4'ha : _GEN_17570; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17572 = 10'h5b == _T_378[9:0] ? 4'ha : _GEN_17571; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17573 = 10'h5c == _T_378[9:0] ? 4'ha : _GEN_17572; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17574 = 10'h5d == _T_378[9:0] ? 4'h3 : _GEN_17573; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17575 = 10'h5e == _T_378[9:0] ? 4'ha : _GEN_17574; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17576 = 10'h5f == _T_378[9:0] ? 4'h0 : _GEN_17575; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17577 = 10'h60 == _T_378[9:0] ? 4'ha : _GEN_17576; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17578 = 10'h61 == _T_378[9:0] ? 4'ha : _GEN_17577; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17579 = 10'h62 == _T_378[9:0] ? 4'ha : _GEN_17578; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17580 = 10'h63 == _T_378[9:0] ? 4'ha : _GEN_17579; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17581 = 10'h64 == _T_378[9:0] ? 4'h3 : _GEN_17580; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17582 = 10'h65 == _T_378[9:0] ? 4'h0 : _GEN_17581; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17583 = 10'h66 == _T_378[9:0] ? 4'ha : _GEN_17582; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17584 = 10'h67 == _T_378[9:0] ? 4'ha : _GEN_17583; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17585 = 10'h68 == _T_378[9:0] ? 4'ha : _GEN_17584; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17586 = 10'h69 == _T_378[9:0] ? 4'h0 : _GEN_17585; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17587 = 10'h6a == _T_378[9:0] ? 4'h1 : _GEN_17586; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17588 = 10'h6b == _T_378[9:0] ? 4'h1 : _GEN_17587; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17589 = 10'h6c == _T_378[9:0] ? 4'ha : _GEN_17588; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17590 = 10'h6d == _T_378[9:0] ? 4'ha : _GEN_17589; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17591 = 10'h6e == _T_378[9:0] ? 4'ha : _GEN_17590; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17592 = 10'h6f == _T_378[9:0] ? 4'ha : _GEN_17591; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17593 = 10'h70 == _T_378[9:0] ? 4'ha : _GEN_17592; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17594 = 10'h71 == _T_378[9:0] ? 4'ha : _GEN_17593; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17595 = 10'h72 == _T_378[9:0] ? 4'ha : _GEN_17594; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17596 = 10'h73 == _T_378[9:0] ? 4'h1 : _GEN_17595; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17597 = 10'h74 == _T_378[9:0] ? 4'h0 : _GEN_17596; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17598 = 10'h75 == _T_378[9:0] ? 4'h0 : _GEN_17597; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17599 = 10'h76 == _T_378[9:0] ? 4'h0 : _GEN_17598; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17600 = 10'h77 == _T_378[9:0] ? 4'ha : _GEN_17599; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17601 = 10'h78 == _T_378[9:0] ? 4'ha : _GEN_17600; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17602 = 10'h79 == _T_378[9:0] ? 4'ha : _GEN_17601; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17603 = 10'h7a == _T_378[9:0] ? 4'h0 : _GEN_17602; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17604 = 10'h7b == _T_378[9:0] ? 4'ha : _GEN_17603; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17605 = 10'h7c == _T_378[9:0] ? 4'ha : _GEN_17604; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17606 = 10'h7d == _T_378[9:0] ? 4'h2 : _GEN_17605; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17607 = 10'h7e == _T_378[9:0] ? 4'h3 : _GEN_17606; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17608 = 10'h7f == _T_378[9:0] ? 4'h0 : _GEN_17607; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17609 = 10'h80 == _T_378[9:0] ? 4'ha : _GEN_17608; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17610 = 10'h81 == _T_378[9:0] ? 4'ha : _GEN_17609; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17611 = 10'h82 == _T_378[9:0] ? 4'h1 : _GEN_17610; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17612 = 10'h83 == _T_378[9:0] ? 4'h0 : _GEN_17611; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17613 = 10'h84 == _T_378[9:0] ? 4'h2 : _GEN_17612; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17614 = 10'h85 == _T_378[9:0] ? 4'h1 : _GEN_17613; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17615 = 10'h86 == _T_378[9:0] ? 4'h1 : _GEN_17614; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17616 = 10'h87 == _T_378[9:0] ? 4'ha : _GEN_17615; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17617 = 10'h88 == _T_378[9:0] ? 4'ha : _GEN_17616; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17618 = 10'h89 == _T_378[9:0] ? 4'h0 : _GEN_17617; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17619 = 10'h8a == _T_378[9:0] ? 4'h0 : _GEN_17618; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17620 = 10'h8b == _T_378[9:0] ? 4'h1 : _GEN_17619; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17621 = 10'h8c == _T_378[9:0] ? 4'h1 : _GEN_17620; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17622 = 10'h8d == _T_378[9:0] ? 4'h1 : _GEN_17621; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17623 = 10'h8e == _T_378[9:0] ? 4'h1 : _GEN_17622; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17624 = 10'h8f == _T_378[9:0] ? 4'h1 : _GEN_17623; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17625 = 10'h90 == _T_378[9:0] ? 4'h1 : _GEN_17624; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17626 = 10'h91 == _T_378[9:0] ? 4'h1 : _GEN_17625; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17627 = 10'h92 == _T_378[9:0] ? 4'h1 : _GEN_17626; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17628 = 10'h93 == _T_378[9:0] ? 4'h0 : _GEN_17627; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17629 = 10'h94 == _T_378[9:0] ? 4'h0 : _GEN_17628; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17630 = 10'h95 == _T_378[9:0] ? 4'ha : _GEN_17629; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17631 = 10'h96 == _T_378[9:0] ? 4'ha : _GEN_17630; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17632 = 10'h97 == _T_378[9:0] ? 4'ha : _GEN_17631; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17633 = 10'h98 == _T_378[9:0] ? 4'h1 : _GEN_17632; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17634 = 10'h99 == _T_378[9:0] ? 4'h0 : _GEN_17633; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17635 = 10'h9a == _T_378[9:0] ? 4'h1 : _GEN_17634; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17636 = 10'h9b == _T_378[9:0] ? 4'h1 : _GEN_17635; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17637 = 10'h9c == _T_378[9:0] ? 4'ha : _GEN_17636; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17638 = 10'h9d == _T_378[9:0] ? 4'ha : _GEN_17637; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17639 = 10'h9e == _T_378[9:0] ? 4'h3 : _GEN_17638; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17640 = 10'h9f == _T_378[9:0] ? 4'h0 : _GEN_17639; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17641 = 10'ha0 == _T_378[9:0] ? 4'ha : _GEN_17640; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17642 = 10'ha1 == _T_378[9:0] ? 4'h1 : _GEN_17641; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17643 = 10'ha2 == _T_378[9:0] ? 4'h0 : _GEN_17642; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17644 = 10'ha3 == _T_378[9:0] ? 4'h3 : _GEN_17643; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17645 = 10'ha4 == _T_378[9:0] ? 4'ha : _GEN_17644; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17646 = 10'ha5 == _T_378[9:0] ? 4'ha : _GEN_17645; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17647 = 10'ha6 == _T_378[9:0] ? 4'ha : _GEN_17646; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17648 = 10'ha7 == _T_378[9:0] ? 4'h0 : _GEN_17647; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17649 = 10'ha8 == _T_378[9:0] ? 4'ha : _GEN_17648; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17650 = 10'ha9 == _T_378[9:0] ? 4'h1 : _GEN_17649; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17651 = 10'haa == _T_378[9:0] ? 4'h0 : _GEN_17650; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17652 = 10'hab == _T_378[9:0] ? 4'h0 : _GEN_17651; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17653 = 10'hac == _T_378[9:0] ? 4'h0 : _GEN_17652; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17654 = 10'had == _T_378[9:0] ? 4'h0 : _GEN_17653; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17655 = 10'hae == _T_378[9:0] ? 4'h0 : _GEN_17654; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17656 = 10'haf == _T_378[9:0] ? 4'h0 : _GEN_17655; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17657 = 10'hb0 == _T_378[9:0] ? 4'h0 : _GEN_17656; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17658 = 10'hb1 == _T_378[9:0] ? 4'h0 : _GEN_17657; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17659 = 10'hb2 == _T_378[9:0] ? 4'h0 : _GEN_17658; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17660 = 10'hb3 == _T_378[9:0] ? 4'h0 : _GEN_17659; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17661 = 10'hb4 == _T_378[9:0] ? 4'h1 : _GEN_17660; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17662 = 10'hb5 == _T_378[9:0] ? 4'h1 : _GEN_17661; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17663 = 10'hb6 == _T_378[9:0] ? 4'ha : _GEN_17662; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17664 = 10'hb7 == _T_378[9:0] ? 4'h0 : _GEN_17663; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17665 = 10'hb8 == _T_378[9:0] ? 4'ha : _GEN_17664; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17666 = 10'hb9 == _T_378[9:0] ? 4'ha : _GEN_17665; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17667 = 10'hba == _T_378[9:0] ? 4'ha : _GEN_17666; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17668 = 10'hbb == _T_378[9:0] ? 4'h0 : _GEN_17667; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17669 = 10'hbc == _T_378[9:0] ? 4'ha : _GEN_17668; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17670 = 10'hbd == _T_378[9:0] ? 4'ha : _GEN_17669; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17671 = 10'hbe == _T_378[9:0] ? 4'h3 : _GEN_17670; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17672 = 10'hbf == _T_378[9:0] ? 4'h0 : _GEN_17671; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17673 = 10'hc0 == _T_378[9:0] ? 4'ha : _GEN_17672; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17674 = 10'hc1 == _T_378[9:0] ? 4'ha : _GEN_17673; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17675 = 10'hc2 == _T_378[9:0] ? 4'h3 : _GEN_17674; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17676 = 10'hc3 == _T_378[9:0] ? 4'h2 : _GEN_17675; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17677 = 10'hc4 == _T_378[9:0] ? 4'h0 : _GEN_17676; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17678 = 10'hc5 == _T_378[9:0] ? 4'h0 : _GEN_17677; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17679 = 10'hc6 == _T_378[9:0] ? 4'h0 : _GEN_17678; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17680 = 10'hc7 == _T_378[9:0] ? 4'ha : _GEN_17679; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17681 = 10'hc8 == _T_378[9:0] ? 4'h1 : _GEN_17680; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17682 = 10'hc9 == _T_378[9:0] ? 4'h0 : _GEN_17681; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17683 = 10'hca == _T_378[9:0] ? 4'h0 : _GEN_17682; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17684 = 10'hcb == _T_378[9:0] ? 4'h0 : _GEN_17683; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17685 = 10'hcc == _T_378[9:0] ? 4'h0 : _GEN_17684; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17686 = 10'hcd == _T_378[9:0] ? 4'h0 : _GEN_17685; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17687 = 10'hce == _T_378[9:0] ? 4'h0 : _GEN_17686; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17688 = 10'hcf == _T_378[9:0] ? 4'h0 : _GEN_17687; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17689 = 10'hd0 == _T_378[9:0] ? 4'h0 : _GEN_17688; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17690 = 10'hd1 == _T_378[9:0] ? 4'h0 : _GEN_17689; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17691 = 10'hd2 == _T_378[9:0] ? 4'h0 : _GEN_17690; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17692 = 10'hd3 == _T_378[9:0] ? 4'h0 : _GEN_17691; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17693 = 10'hd4 == _T_378[9:0] ? 4'h0 : _GEN_17692; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17694 = 10'hd5 == _T_378[9:0] ? 4'h0 : _GEN_17693; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17695 = 10'hd6 == _T_378[9:0] ? 4'h1 : _GEN_17694; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17696 = 10'hd7 == _T_378[9:0] ? 4'ha : _GEN_17695; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17697 = 10'hd8 == _T_378[9:0] ? 4'h0 : _GEN_17696; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17698 = 10'hd9 == _T_378[9:0] ? 4'ha : _GEN_17697; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17699 = 10'hda == _T_378[9:0] ? 4'ha : _GEN_17698; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17700 = 10'hdb == _T_378[9:0] ? 4'ha : _GEN_17699; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17701 = 10'hdc == _T_378[9:0] ? 4'ha : _GEN_17700; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17702 = 10'hdd == _T_378[9:0] ? 4'h3 : _GEN_17701; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17703 = 10'hde == _T_378[9:0] ? 4'h2 : _GEN_17702; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17704 = 10'hdf == _T_378[9:0] ? 4'h0 : _GEN_17703; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17705 = 10'he0 == _T_378[9:0] ? 4'ha : _GEN_17704; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17706 = 10'he1 == _T_378[9:0] ? 4'ha : _GEN_17705; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17707 = 10'he2 == _T_378[9:0] ? 4'h3 : _GEN_17706; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17708 = 10'he3 == _T_378[9:0] ? 4'ha : _GEN_17707; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17709 = 10'he4 == _T_378[9:0] ? 4'ha : _GEN_17708; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17710 = 10'he5 == _T_378[9:0] ? 4'ha : _GEN_17709; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17711 = 10'he6 == _T_378[9:0] ? 4'ha : _GEN_17710; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17712 = 10'he7 == _T_378[9:0] ? 4'h1 : _GEN_17711; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17713 = 10'he8 == _T_378[9:0] ? 4'h1 : _GEN_17712; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17714 = 10'he9 == _T_378[9:0] ? 4'h1 : _GEN_17713; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17715 = 10'hea == _T_378[9:0] ? 4'h0 : _GEN_17714; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17716 = 10'heb == _T_378[9:0] ? 4'h0 : _GEN_17715; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17717 = 10'hec == _T_378[9:0] ? 4'h0 : _GEN_17716; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17718 = 10'hed == _T_378[9:0] ? 4'h0 : _GEN_17717; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17719 = 10'hee == _T_378[9:0] ? 4'h0 : _GEN_17718; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17720 = 10'hef == _T_378[9:0] ? 4'h0 : _GEN_17719; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17721 = 10'hf0 == _T_378[9:0] ? 4'h0 : _GEN_17720; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17722 = 10'hf1 == _T_378[9:0] ? 4'h0 : _GEN_17721; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17723 = 10'hf2 == _T_378[9:0] ? 4'h0 : _GEN_17722; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17724 = 10'hf3 == _T_378[9:0] ? 4'h0 : _GEN_17723; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17725 = 10'hf4 == _T_378[9:0] ? 4'h0 : _GEN_17724; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17726 = 10'hf5 == _T_378[9:0] ? 4'h1 : _GEN_17725; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17727 = 10'hf6 == _T_378[9:0] ? 4'h0 : _GEN_17726; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17728 = 10'hf7 == _T_378[9:0] ? 4'h0 : _GEN_17727; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17729 = 10'hf8 == _T_378[9:0] ? 4'h1 : _GEN_17728; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17730 = 10'hf9 == _T_378[9:0] ? 4'h0 : _GEN_17729; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17731 = 10'hfa == _T_378[9:0] ? 4'ha : _GEN_17730; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17732 = 10'hfb == _T_378[9:0] ? 4'ha : _GEN_17731; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17733 = 10'hfc == _T_378[9:0] ? 4'ha : _GEN_17732; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17734 = 10'hfd == _T_378[9:0] ? 4'h3 : _GEN_17733; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17735 = 10'hfe == _T_378[9:0] ? 4'ha : _GEN_17734; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17736 = 10'hff == _T_378[9:0] ? 4'h0 : _GEN_17735; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17737 = 10'h100 == _T_378[9:0] ? 4'ha : _GEN_17736; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17738 = 10'h101 == _T_378[9:0] ? 4'h0 : _GEN_17737; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17739 = 10'h102 == _T_378[9:0] ? 4'h3 : _GEN_17738; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17740 = 10'h103 == _T_378[9:0] ? 4'ha : _GEN_17739; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17741 = 10'h104 == _T_378[9:0] ? 4'ha : _GEN_17740; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17742 = 10'h105 == _T_378[9:0] ? 4'ha : _GEN_17741; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17743 = 10'h106 == _T_378[9:0] ? 4'ha : _GEN_17742; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17744 = 10'h107 == _T_378[9:0] ? 4'ha : _GEN_17743; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17745 = 10'h108 == _T_378[9:0] ? 4'h1 : _GEN_17744; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17746 = 10'h109 == _T_378[9:0] ? 4'h0 : _GEN_17745; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17747 = 10'h10a == _T_378[9:0] ? 4'h0 : _GEN_17746; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17748 = 10'h10b == _T_378[9:0] ? 4'h0 : _GEN_17747; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17749 = 10'h10c == _T_378[9:0] ? 4'h0 : _GEN_17748; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17750 = 10'h10d == _T_378[9:0] ? 4'h0 : _GEN_17749; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17751 = 10'h10e == _T_378[9:0] ? 4'h0 : _GEN_17750; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17752 = 10'h10f == _T_378[9:0] ? 4'h0 : _GEN_17751; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17753 = 10'h110 == _T_378[9:0] ? 4'h0 : _GEN_17752; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17754 = 10'h111 == _T_378[9:0] ? 4'h0 : _GEN_17753; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17755 = 10'h112 == _T_378[9:0] ? 4'h0 : _GEN_17754; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17756 = 10'h113 == _T_378[9:0] ? 4'h0 : _GEN_17755; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17757 = 10'h114 == _T_378[9:0] ? 4'h0 : _GEN_17756; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17758 = 10'h115 == _T_378[9:0] ? 4'h0 : _GEN_17757; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17759 = 10'h116 == _T_378[9:0] ? 4'h1 : _GEN_17758; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17760 = 10'h117 == _T_378[9:0] ? 4'ha : _GEN_17759; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17761 = 10'h118 == _T_378[9:0] ? 4'ha : _GEN_17760; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17762 = 10'h119 == _T_378[9:0] ? 4'ha : _GEN_17761; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17763 = 10'h11a == _T_378[9:0] ? 4'h0 : _GEN_17762; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17764 = 10'h11b == _T_378[9:0] ? 4'ha : _GEN_17763; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17765 = 10'h11c == _T_378[9:0] ? 4'ha : _GEN_17764; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17766 = 10'h11d == _T_378[9:0] ? 4'h2 : _GEN_17765; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17767 = 10'h11e == _T_378[9:0] ? 4'h3 : _GEN_17766; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17768 = 10'h11f == _T_378[9:0] ? 4'h0 : _GEN_17767; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17769 = 10'h120 == _T_378[9:0] ? 4'ha : _GEN_17768; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17770 = 10'h121 == _T_378[9:0] ? 4'ha : _GEN_17769; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17771 = 10'h122 == _T_378[9:0] ? 4'h3 : _GEN_17770; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17772 = 10'h123 == _T_378[9:0] ? 4'ha : _GEN_17771; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17773 = 10'h124 == _T_378[9:0] ? 4'ha : _GEN_17772; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17774 = 10'h125 == _T_378[9:0] ? 4'ha : _GEN_17773; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17775 = 10'h126 == _T_378[9:0] ? 4'ha : _GEN_17774; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17776 = 10'h127 == _T_378[9:0] ? 4'h1 : _GEN_17775; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17777 = 10'h128 == _T_378[9:0] ? 4'h0 : _GEN_17776; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17778 = 10'h129 == _T_378[9:0] ? 4'ha : _GEN_17777; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17779 = 10'h12a == _T_378[9:0] ? 4'ha : _GEN_17778; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17780 = 10'h12b == _T_378[9:0] ? 4'h0 : _GEN_17779; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17781 = 10'h12c == _T_378[9:0] ? 4'h0 : _GEN_17780; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17782 = 10'h12d == _T_378[9:0] ? 4'h0 : _GEN_17781; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17783 = 10'h12e == _T_378[9:0] ? 4'h0 : _GEN_17782; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17784 = 10'h12f == _T_378[9:0] ? 4'h0 : _GEN_17783; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17785 = 10'h130 == _T_378[9:0] ? 4'h0 : _GEN_17784; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17786 = 10'h131 == _T_378[9:0] ? 4'h0 : _GEN_17785; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17787 = 10'h132 == _T_378[9:0] ? 4'h0 : _GEN_17786; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17788 = 10'h133 == _T_378[9:0] ? 4'h0 : _GEN_17787; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17789 = 10'h134 == _T_378[9:0] ? 4'ha : _GEN_17788; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17790 = 10'h135 == _T_378[9:0] ? 4'ha : _GEN_17789; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17791 = 10'h136 == _T_378[9:0] ? 4'h0 : _GEN_17790; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17792 = 10'h137 == _T_378[9:0] ? 4'h1 : _GEN_17791; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17793 = 10'h138 == _T_378[9:0] ? 4'ha : _GEN_17792; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17794 = 10'h139 == _T_378[9:0] ? 4'ha : _GEN_17793; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17795 = 10'h13a == _T_378[9:0] ? 4'ha : _GEN_17794; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17796 = 10'h13b == _T_378[9:0] ? 4'ha : _GEN_17795; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17797 = 10'h13c == _T_378[9:0] ? 4'ha : _GEN_17796; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17798 = 10'h13d == _T_378[9:0] ? 4'ha : _GEN_17797; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17799 = 10'h13e == _T_378[9:0] ? 4'h3 : _GEN_17798; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17800 = 10'h13f == _T_378[9:0] ? 4'h0 : _GEN_17799; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17801 = 10'h140 == _T_378[9:0] ? 4'ha : _GEN_17800; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17802 = 10'h141 == _T_378[9:0] ? 4'ha : _GEN_17801; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17803 = 10'h142 == _T_378[9:0] ? 4'h2 : _GEN_17802; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17804 = 10'h143 == _T_378[9:0] ? 4'h3 : _GEN_17803; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17805 = 10'h144 == _T_378[9:0] ? 4'ha : _GEN_17804; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17806 = 10'h145 == _T_378[9:0] ? 4'ha : _GEN_17805; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17807 = 10'h146 == _T_378[9:0] ? 4'h1 : _GEN_17806; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17808 = 10'h147 == _T_378[9:0] ? 4'h0 : _GEN_17807; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17809 = 10'h148 == _T_378[9:0] ? 4'ha : _GEN_17808; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17810 = 10'h149 == _T_378[9:0] ? 4'ha : _GEN_17809; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17811 = 10'h14a == _T_378[9:0] ? 4'ha : _GEN_17810; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17812 = 10'h14b == _T_378[9:0] ? 4'ha : _GEN_17811; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17813 = 10'h14c == _T_378[9:0] ? 4'ha : _GEN_17812; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17814 = 10'h14d == _T_378[9:0] ? 4'ha : _GEN_17813; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17815 = 10'h14e == _T_378[9:0] ? 4'ha : _GEN_17814; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17816 = 10'h14f == _T_378[9:0] ? 4'ha : _GEN_17815; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17817 = 10'h150 == _T_378[9:0] ? 4'ha : _GEN_17816; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17818 = 10'h151 == _T_378[9:0] ? 4'ha : _GEN_17817; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17819 = 10'h152 == _T_378[9:0] ? 4'ha : _GEN_17818; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17820 = 10'h153 == _T_378[9:0] ? 4'ha : _GEN_17819; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17821 = 10'h154 == _T_378[9:0] ? 4'ha : _GEN_17820; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17822 = 10'h155 == _T_378[9:0] ? 4'ha : _GEN_17821; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17823 = 10'h156 == _T_378[9:0] ? 4'ha : _GEN_17822; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17824 = 10'h157 == _T_378[9:0] ? 4'h0 : _GEN_17823; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17825 = 10'h158 == _T_378[9:0] ? 4'ha : _GEN_17824; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17826 = 10'h159 == _T_378[9:0] ? 4'ha : _GEN_17825; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17827 = 10'h15a == _T_378[9:0] ? 4'ha : _GEN_17826; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17828 = 10'h15b == _T_378[9:0] ? 4'ha : _GEN_17827; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17829 = 10'h15c == _T_378[9:0] ? 4'ha : _GEN_17828; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17830 = 10'h15d == _T_378[9:0] ? 4'h3 : _GEN_17829; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17831 = 10'h15e == _T_378[9:0] ? 4'h2 : _GEN_17830; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17832 = 10'h15f == _T_378[9:0] ? 4'h0 : _GEN_17831; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17833 = 10'h160 == _T_378[9:0] ? 4'ha : _GEN_17832; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17834 = 10'h161 == _T_378[9:0] ? 4'ha : _GEN_17833; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17835 = 10'h162 == _T_378[9:0] ? 4'ha : _GEN_17834; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17836 = 10'h163 == _T_378[9:0] ? 4'h2 : _GEN_17835; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17837 = 10'h164 == _T_378[9:0] ? 4'h3 : _GEN_17836; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17838 = 10'h165 == _T_378[9:0] ? 4'h1 : _GEN_17837; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17839 = 10'h166 == _T_378[9:0] ? 4'h0 : _GEN_17838; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17840 = 10'h167 == _T_378[9:0] ? 4'h0 : _GEN_17839; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17841 = 10'h168 == _T_378[9:0] ? 4'h5 : _GEN_17840; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17842 = 10'h169 == _T_378[9:0] ? 4'h3 : _GEN_17841; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17843 = 10'h16a == _T_378[9:0] ? 4'h5 : _GEN_17842; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17844 = 10'h16b == _T_378[9:0] ? 4'h5 : _GEN_17843; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17845 = 10'h16c == _T_378[9:0] ? 4'ha : _GEN_17844; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17846 = 10'h16d == _T_378[9:0] ? 4'ha : _GEN_17845; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17847 = 10'h16e == _T_378[9:0] ? 4'ha : _GEN_17846; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17848 = 10'h16f == _T_378[9:0] ? 4'ha : _GEN_17847; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17849 = 10'h170 == _T_378[9:0] ? 4'ha : _GEN_17848; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17850 = 10'h171 == _T_378[9:0] ? 4'ha : _GEN_17849; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17851 = 10'h172 == _T_378[9:0] ? 4'ha : _GEN_17850; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17852 = 10'h173 == _T_378[9:0] ? 4'ha : _GEN_17851; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17853 = 10'h174 == _T_378[9:0] ? 4'ha : _GEN_17852; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17854 = 10'h175 == _T_378[9:0] ? 4'ha : _GEN_17853; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17855 = 10'h176 == _T_378[9:0] ? 4'h0 : _GEN_17854; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17856 = 10'h177 == _T_378[9:0] ? 4'h0 : _GEN_17855; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17857 = 10'h178 == _T_378[9:0] ? 4'h1 : _GEN_17856; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17858 = 10'h179 == _T_378[9:0] ? 4'ha : _GEN_17857; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17859 = 10'h17a == _T_378[9:0] ? 4'ha : _GEN_17858; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17860 = 10'h17b == _T_378[9:0] ? 4'ha : _GEN_17859; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17861 = 10'h17c == _T_378[9:0] ? 4'h3 : _GEN_17860; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17862 = 10'h17d == _T_378[9:0] ? 4'h2 : _GEN_17861; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17863 = 10'h17e == _T_378[9:0] ? 4'ha : _GEN_17862; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17864 = 10'h17f == _T_378[9:0] ? 4'h0 : _GEN_17863; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17865 = 10'h180 == _T_378[9:0] ? 4'h5 : _GEN_17864; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17866 = 10'h181 == _T_378[9:0] ? 4'h5 : _GEN_17865; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17867 = 10'h182 == _T_378[9:0] ? 4'h5 : _GEN_17866; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17868 = 10'h183 == _T_378[9:0] ? 4'h5 : _GEN_17867; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17869 = 10'h184 == _T_378[9:0] ? 4'h3 : _GEN_17868; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17870 = 10'h185 == _T_378[9:0] ? 4'h1 : _GEN_17869; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17871 = 10'h186 == _T_378[9:0] ? 4'hb : _GEN_17870; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17872 = 10'h187 == _T_378[9:0] ? 4'h0 : _GEN_17871; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17873 = 10'h188 == _T_378[9:0] ? 4'h5 : _GEN_17872; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17874 = 10'h189 == _T_378[9:0] ? 4'h5 : _GEN_17873; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17875 = 10'h18a == _T_378[9:0] ? 4'h5 : _GEN_17874; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17876 = 10'h18b == _T_378[9:0] ? 4'h5 : _GEN_17875; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17877 = 10'h18c == _T_378[9:0] ? 4'h5 : _GEN_17876; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17878 = 10'h18d == _T_378[9:0] ? 4'h5 : _GEN_17877; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17879 = 10'h18e == _T_378[9:0] ? 4'h5 : _GEN_17878; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17880 = 10'h18f == _T_378[9:0] ? 4'h5 : _GEN_17879; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17881 = 10'h190 == _T_378[9:0] ? 4'h5 : _GEN_17880; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17882 = 10'h191 == _T_378[9:0] ? 4'h5 : _GEN_17881; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17883 = 10'h192 == _T_378[9:0] ? 4'h3 : _GEN_17882; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17884 = 10'h193 == _T_378[9:0] ? 4'h5 : _GEN_17883; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17885 = 10'h194 == _T_378[9:0] ? 4'h5 : _GEN_17884; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17886 = 10'h195 == _T_378[9:0] ? 4'h5 : _GEN_17885; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17887 = 10'h196 == _T_378[9:0] ? 4'h0 : _GEN_17886; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17888 = 10'h197 == _T_378[9:0] ? 4'ha : _GEN_17887; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17889 = 10'h198 == _T_378[9:0] ? 4'h1 : _GEN_17888; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17890 = 10'h199 == _T_378[9:0] ? 4'ha : _GEN_17889; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17891 = 10'h19a == _T_378[9:0] ? 4'ha : _GEN_17890; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17892 = 10'h19b == _T_378[9:0] ? 4'ha : _GEN_17891; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17893 = 10'h19c == _T_378[9:0] ? 4'h3 : _GEN_17892; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17894 = 10'h19d == _T_378[9:0] ? 4'ha : _GEN_17893; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17895 = 10'h19e == _T_378[9:0] ? 4'ha : _GEN_17894; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17896 = 10'h19f == _T_378[9:0] ? 4'h0 : _GEN_17895; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17897 = 10'h1a0 == _T_378[9:0] ? 4'h5 : _GEN_17896; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17898 = 10'h1a1 == _T_378[9:0] ? 4'h5 : _GEN_17897; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17899 = 10'h1a2 == _T_378[9:0] ? 4'h3 : _GEN_17898; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17900 = 10'h1a3 == _T_378[9:0] ? 4'h5 : _GEN_17899; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17901 = 10'h1a4 == _T_378[9:0] ? 4'h3 : _GEN_17900; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17902 = 10'h1a5 == _T_378[9:0] ? 4'h0 : _GEN_17901; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17903 = 10'h1a6 == _T_378[9:0] ? 4'h5 : _GEN_17902; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17904 = 10'h1a7 == _T_378[9:0] ? 4'h0 : _GEN_17903; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17905 = 10'h1a8 == _T_378[9:0] ? 4'hb : _GEN_17904; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17906 = 10'h1a9 == _T_378[9:0] ? 4'h5 : _GEN_17905; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17907 = 10'h1aa == _T_378[9:0] ? 4'h5 : _GEN_17906; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17908 = 10'h1ab == _T_378[9:0] ? 4'h3 : _GEN_17907; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17909 = 10'h1ac == _T_378[9:0] ? 4'h5 : _GEN_17908; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17910 = 10'h1ad == _T_378[9:0] ? 4'h5 : _GEN_17909; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17911 = 10'h1ae == _T_378[9:0] ? 4'h5 : _GEN_17910; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17912 = 10'h1af == _T_378[9:0] ? 4'h5 : _GEN_17911; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17913 = 10'h1b0 == _T_378[9:0] ? 4'h5 : _GEN_17912; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17914 = 10'h1b1 == _T_378[9:0] ? 4'h5 : _GEN_17913; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17915 = 10'h1b2 == _T_378[9:0] ? 4'h5 : _GEN_17914; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17916 = 10'h1b3 == _T_378[9:0] ? 4'h5 : _GEN_17915; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17917 = 10'h1b4 == _T_378[9:0] ? 4'h5 : _GEN_17916; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17918 = 10'h1b5 == _T_378[9:0] ? 4'h5 : _GEN_17917; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17919 = 10'h1b6 == _T_378[9:0] ? 4'h0 : _GEN_17918; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17920 = 10'h1b7 == _T_378[9:0] ? 4'h5 : _GEN_17919; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17921 = 10'h1b8 == _T_378[9:0] ? 4'h0 : _GEN_17920; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17922 = 10'h1b9 == _T_378[9:0] ? 4'h5 : _GEN_17921; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17923 = 10'h1ba == _T_378[9:0] ? 4'h5 : _GEN_17922; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17924 = 10'h1bb == _T_378[9:0] ? 4'h5 : _GEN_17923; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17925 = 10'h1bc == _T_378[9:0] ? 4'h2 : _GEN_17924; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17926 = 10'h1bd == _T_378[9:0] ? 4'h3 : _GEN_17925; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17927 = 10'h1be == _T_378[9:0] ? 4'h5 : _GEN_17926; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17928 = 10'h1bf == _T_378[9:0] ? 4'h0 : _GEN_17927; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17929 = 10'h1c0 == _T_378[9:0] ? 4'h5 : _GEN_17928; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17930 = 10'h1c1 == _T_378[9:0] ? 4'h5 : _GEN_17929; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17931 = 10'h1c2 == _T_378[9:0] ? 4'h5 : _GEN_17930; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17932 = 10'h1c3 == _T_378[9:0] ? 4'h2 : _GEN_17931; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17933 = 10'h1c4 == _T_378[9:0] ? 4'h2 : _GEN_17932; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17934 = 10'h1c5 == _T_378[9:0] ? 4'h5 : _GEN_17933; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17935 = 10'h1c6 == _T_378[9:0] ? 4'h5 : _GEN_17934; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17936 = 10'h1c7 == _T_378[9:0] ? 4'h5 : _GEN_17935; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17937 = 10'h1c8 == _T_378[9:0] ? 4'h5 : _GEN_17936; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17938 = 10'h1c9 == _T_378[9:0] ? 4'hb : _GEN_17937; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17939 = 10'h1ca == _T_378[9:0] ? 4'hb : _GEN_17938; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17940 = 10'h1cb == _T_378[9:0] ? 4'hb : _GEN_17939; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17941 = 10'h1cc == _T_378[9:0] ? 4'hb : _GEN_17940; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17942 = 10'h1cd == _T_378[9:0] ? 4'hb : _GEN_17941; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17943 = 10'h1ce == _T_378[9:0] ? 4'hb : _GEN_17942; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17944 = 10'h1cf == _T_378[9:0] ? 4'hb : _GEN_17943; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17945 = 10'h1d0 == _T_378[9:0] ? 4'hb : _GEN_17944; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17946 = 10'h1d1 == _T_378[9:0] ? 4'hb : _GEN_17945; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17947 = 10'h1d2 == _T_378[9:0] ? 4'hb : _GEN_17946; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17948 = 10'h1d3 == _T_378[9:0] ? 4'hb : _GEN_17947; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17949 = 10'h1d4 == _T_378[9:0] ? 4'hb : _GEN_17948; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17950 = 10'h1d5 == _T_378[9:0] ? 4'hb : _GEN_17949; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17951 = 10'h1d6 == _T_378[9:0] ? 4'h5 : _GEN_17950; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17952 = 10'h1d7 == _T_378[9:0] ? 4'h5 : _GEN_17951; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17953 = 10'h1d8 == _T_378[9:0] ? 4'h5 : _GEN_17952; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17954 = 10'h1d9 == _T_378[9:0] ? 4'h5 : _GEN_17953; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17955 = 10'h1da == _T_378[9:0] ? 4'h5 : _GEN_17954; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17956 = 10'h1db == _T_378[9:0] ? 4'h5 : _GEN_17955; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17957 = 10'h1dc == _T_378[9:0] ? 4'h5 : _GEN_17956; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17958 = 10'h1dd == _T_378[9:0] ? 4'h3 : _GEN_17957; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17959 = 10'h1de == _T_378[9:0] ? 4'h5 : _GEN_17958; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17960 = 10'h1df == _T_378[9:0] ? 4'h0 : _GEN_17959; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17961 = 10'h1e0 == _T_378[9:0] ? 4'h3 : _GEN_17960; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17962 = 10'h1e1 == _T_378[9:0] ? 4'h5 : _GEN_17961; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17963 = 10'h1e2 == _T_378[9:0] ? 4'h2 : _GEN_17962; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17964 = 10'h1e3 == _T_378[9:0] ? 4'h2 : _GEN_17963; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17965 = 10'h1e4 == _T_378[9:0] ? 4'h5 : _GEN_17964; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17966 = 10'h1e5 == _T_378[9:0] ? 4'h5 : _GEN_17965; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17967 = 10'h1e6 == _T_378[9:0] ? 4'h5 : _GEN_17966; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17968 = 10'h1e7 == _T_378[9:0] ? 4'h5 : _GEN_17967; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17969 = 10'h1e8 == _T_378[9:0] ? 4'hb : _GEN_17968; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17970 = 10'h1e9 == _T_378[9:0] ? 4'h5 : _GEN_17969; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17971 = 10'h1ea == _T_378[9:0] ? 4'h5 : _GEN_17970; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17972 = 10'h1eb == _T_378[9:0] ? 4'hb : _GEN_17971; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17973 = 10'h1ec == _T_378[9:0] ? 4'h5 : _GEN_17972; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17974 = 10'h1ed == _T_378[9:0] ? 4'hb : _GEN_17973; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17975 = 10'h1ee == _T_378[9:0] ? 4'h5 : _GEN_17974; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17976 = 10'h1ef == _T_378[9:0] ? 4'hb : _GEN_17975; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17977 = 10'h1f0 == _T_378[9:0] ? 4'h5 : _GEN_17976; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17978 = 10'h1f1 == _T_378[9:0] ? 4'hb : _GEN_17977; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17979 = 10'h1f2 == _T_378[9:0] ? 4'hb : _GEN_17978; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17980 = 10'h1f3 == _T_378[9:0] ? 4'h5 : _GEN_17979; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17981 = 10'h1f4 == _T_378[9:0] ? 4'hb : _GEN_17980; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17982 = 10'h1f5 == _T_378[9:0] ? 4'hb : _GEN_17981; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17983 = 10'h1f6 == _T_378[9:0] ? 4'h5 : _GEN_17982; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17984 = 10'h1f7 == _T_378[9:0] ? 4'h5 : _GEN_17983; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17985 = 10'h1f8 == _T_378[9:0] ? 4'h5 : _GEN_17984; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17986 = 10'h1f9 == _T_378[9:0] ? 4'h5 : _GEN_17985; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17987 = 10'h1fa == _T_378[9:0] ? 4'h3 : _GEN_17986; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17988 = 10'h1fb == _T_378[9:0] ? 4'h5 : _GEN_17987; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17989 = 10'h1fc == _T_378[9:0] ? 4'h5 : _GEN_17988; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17990 = 10'h1fd == _T_378[9:0] ? 4'h2 : _GEN_17989; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17991 = 10'h1fe == _T_378[9:0] ? 4'h5 : _GEN_17990; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17992 = 10'h1ff == _T_378[9:0] ? 4'h0 : _GEN_17991; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17993 = 10'h200 == _T_378[9:0] ? 4'h5 : _GEN_17992; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17994 = 10'h201 == _T_378[9:0] ? 4'h5 : _GEN_17993; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17995 = 10'h202 == _T_378[9:0] ? 4'h3 : _GEN_17994; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17996 = 10'h203 == _T_378[9:0] ? 4'h5 : _GEN_17995; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17997 = 10'h204 == _T_378[9:0] ? 4'h5 : _GEN_17996; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17998 = 10'h205 == _T_378[9:0] ? 4'h5 : _GEN_17997; // @[Filter.scala 191:62]
  wire [3:0] _GEN_17999 = 10'h206 == _T_378[9:0] ? 4'hb : _GEN_17998; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18000 = 10'h207 == _T_378[9:0] ? 4'hb : _GEN_17999; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18001 = 10'h208 == _T_378[9:0] ? 4'h5 : _GEN_18000; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18002 = 10'h209 == _T_378[9:0] ? 4'h5 : _GEN_18001; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18003 = 10'h20a == _T_378[9:0] ? 4'h5 : _GEN_18002; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18004 = 10'h20b == _T_378[9:0] ? 4'hb : _GEN_18003; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18005 = 10'h20c == _T_378[9:0] ? 4'h5 : _GEN_18004; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18006 = 10'h20d == _T_378[9:0] ? 4'hb : _GEN_18005; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18007 = 10'h20e == _T_378[9:0] ? 4'h5 : _GEN_18006; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18008 = 10'h20f == _T_378[9:0] ? 4'hb : _GEN_18007; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18009 = 10'h210 == _T_378[9:0] ? 4'h5 : _GEN_18008; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18010 = 10'h211 == _T_378[9:0] ? 4'h5 : _GEN_18009; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18011 = 10'h212 == _T_378[9:0] ? 4'hb : _GEN_18010; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18012 = 10'h213 == _T_378[9:0] ? 4'hb : _GEN_18011; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18013 = 10'h214 == _T_378[9:0] ? 4'hb : _GEN_18012; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18014 = 10'h215 == _T_378[9:0] ? 4'h5 : _GEN_18013; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18015 = 10'h216 == _T_378[9:0] ? 4'h5 : _GEN_18014; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18016 = 10'h217 == _T_378[9:0] ? 4'h5 : _GEN_18015; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18017 = 10'h218 == _T_378[9:0] ? 4'h5 : _GEN_18016; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18018 = 10'h219 == _T_378[9:0] ? 4'h5 : _GEN_18017; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18019 = 10'h21a == _T_378[9:0] ? 4'h5 : _GEN_18018; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18020 = 10'h21b == _T_378[9:0] ? 4'h5 : _GEN_18019; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18021 = 10'h21c == _T_378[9:0] ? 4'h3 : _GEN_18020; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18022 = 10'h21d == _T_378[9:0] ? 4'h2 : _GEN_18021; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18023 = 10'h21e == _T_378[9:0] ? 4'h5 : _GEN_18022; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18024 = 10'h21f == _T_378[9:0] ? 4'h0 : _GEN_18023; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18025 = 10'h220 == _T_378[9:0] ? 4'h0 : _GEN_18024; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18026 = 10'h221 == _T_378[9:0] ? 4'h0 : _GEN_18025; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18027 = 10'h222 == _T_378[9:0] ? 4'h0 : _GEN_18026; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18028 = 10'h223 == _T_378[9:0] ? 4'h0 : _GEN_18027; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18029 = 10'h224 == _T_378[9:0] ? 4'h0 : _GEN_18028; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18030 = 10'h225 == _T_378[9:0] ? 4'h0 : _GEN_18029; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18031 = 10'h226 == _T_378[9:0] ? 4'h0 : _GEN_18030; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18032 = 10'h227 == _T_378[9:0] ? 4'h0 : _GEN_18031; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18033 = 10'h228 == _T_378[9:0] ? 4'h0 : _GEN_18032; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18034 = 10'h229 == _T_378[9:0] ? 4'h0 : _GEN_18033; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18035 = 10'h22a == _T_378[9:0] ? 4'h0 : _GEN_18034; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18036 = 10'h22b == _T_378[9:0] ? 4'h0 : _GEN_18035; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18037 = 10'h22c == _T_378[9:0] ? 4'h0 : _GEN_18036; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18038 = 10'h22d == _T_378[9:0] ? 4'h0 : _GEN_18037; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18039 = 10'h22e == _T_378[9:0] ? 4'h0 : _GEN_18038; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18040 = 10'h22f == _T_378[9:0] ? 4'h0 : _GEN_18039; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18041 = 10'h230 == _T_378[9:0] ? 4'h0 : _GEN_18040; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18042 = 10'h231 == _T_378[9:0] ? 4'h0 : _GEN_18041; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18043 = 10'h232 == _T_378[9:0] ? 4'h0 : _GEN_18042; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18044 = 10'h233 == _T_378[9:0] ? 4'h0 : _GEN_18043; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18045 = 10'h234 == _T_378[9:0] ? 4'h0 : _GEN_18044; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18046 = 10'h235 == _T_378[9:0] ? 4'h0 : _GEN_18045; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18047 = 10'h236 == _T_378[9:0] ? 4'h0 : _GEN_18046; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18048 = 10'h237 == _T_378[9:0] ? 4'h0 : _GEN_18047; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18049 = 10'h238 == _T_378[9:0] ? 4'h0 : _GEN_18048; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18050 = 10'h239 == _T_378[9:0] ? 4'h0 : _GEN_18049; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18051 = 10'h23a == _T_378[9:0] ? 4'h0 : _GEN_18050; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18052 = 10'h23b == _T_378[9:0] ? 4'h0 : _GEN_18051; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18053 = 10'h23c == _T_378[9:0] ? 4'h0 : _GEN_18052; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18054 = 10'h23d == _T_378[9:0] ? 4'h0 : _GEN_18053; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18055 = 10'h23e == _T_378[9:0] ? 4'h0 : _GEN_18054; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18056 = 10'h23f == _T_378[9:0] ? 4'h0 : _GEN_18055; // @[Filter.scala 191:62]
  wire [4:0] _GEN_28358 = {{1'd0}, _GEN_18056}; // @[Filter.scala 191:62]
  wire [8:0] _T_380 = _GEN_28358 * 5'h14; // @[Filter.scala 191:62]
  wire [3:0] _GEN_18060 = 10'h3 == _T_378[9:0] ? 4'ha : 4'h3; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18061 = 10'h4 == _T_378[9:0] ? 4'h3 : _GEN_18060; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18062 = 10'h5 == _T_378[9:0] ? 4'h3 : _GEN_18061; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18063 = 10'h6 == _T_378[9:0] ? 4'h3 : _GEN_18062; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18064 = 10'h7 == _T_378[9:0] ? 4'h3 : _GEN_18063; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18065 = 10'h8 == _T_378[9:0] ? 4'h3 : _GEN_18064; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18066 = 10'h9 == _T_378[9:0] ? 4'h3 : _GEN_18065; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18067 = 10'ha == _T_378[9:0] ? 4'h3 : _GEN_18066; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18068 = 10'hb == _T_378[9:0] ? 4'h3 : _GEN_18067; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18069 = 10'hc == _T_378[9:0] ? 4'h5 : _GEN_18068; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18070 = 10'hd == _T_378[9:0] ? 4'h3 : _GEN_18069; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18071 = 10'he == _T_378[9:0] ? 4'h3 : _GEN_18070; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18072 = 10'hf == _T_378[9:0] ? 4'h3 : _GEN_18071; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18073 = 10'h10 == _T_378[9:0] ? 4'h3 : _GEN_18072; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18074 = 10'h11 == _T_378[9:0] ? 4'h3 : _GEN_18073; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18075 = 10'h12 == _T_378[9:0] ? 4'h3 : _GEN_18074; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18076 = 10'h13 == _T_378[9:0] ? 4'h3 : _GEN_18075; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18077 = 10'h14 == _T_378[9:0] ? 4'h3 : _GEN_18076; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18078 = 10'h15 == _T_378[9:0] ? 4'h3 : _GEN_18077; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18079 = 10'h16 == _T_378[9:0] ? 4'h3 : _GEN_18078; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18080 = 10'h17 == _T_378[9:0] ? 4'h3 : _GEN_18079; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18081 = 10'h18 == _T_378[9:0] ? 4'h3 : _GEN_18080; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18082 = 10'h19 == _T_378[9:0] ? 4'h3 : _GEN_18081; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18083 = 10'h1a == _T_378[9:0] ? 4'h3 : _GEN_18082; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18084 = 10'h1b == _T_378[9:0] ? 4'h3 : _GEN_18083; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18085 = 10'h1c == _T_378[9:0] ? 4'h3 : _GEN_18084; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18086 = 10'h1d == _T_378[9:0] ? 4'h3 : _GEN_18085; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18087 = 10'h1e == _T_378[9:0] ? 4'h3 : _GEN_18086; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18088 = 10'h1f == _T_378[9:0] ? 4'h0 : _GEN_18087; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18089 = 10'h20 == _T_378[9:0] ? 4'h3 : _GEN_18088; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18090 = 10'h21 == _T_378[9:0] ? 4'h5 : _GEN_18089; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18091 = 10'h22 == _T_378[9:0] ? 4'h3 : _GEN_18090; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18092 = 10'h23 == _T_378[9:0] ? 4'ha : _GEN_18091; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18093 = 10'h24 == _T_378[9:0] ? 4'h3 : _GEN_18092; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18094 = 10'h25 == _T_378[9:0] ? 4'h3 : _GEN_18093; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18095 = 10'h26 == _T_378[9:0] ? 4'h3 : _GEN_18094; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18096 = 10'h27 == _T_378[9:0] ? 4'h1 : _GEN_18095; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18097 = 10'h28 == _T_378[9:0] ? 4'h1 : _GEN_18096; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18098 = 10'h29 == _T_378[9:0] ? 4'h3 : _GEN_18097; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18099 = 10'h2a == _T_378[9:0] ? 4'h3 : _GEN_18098; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18100 = 10'h2b == _T_378[9:0] ? 4'h3 : _GEN_18099; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18101 = 10'h2c == _T_378[9:0] ? 4'h3 : _GEN_18100; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18102 = 10'h2d == _T_378[9:0] ? 4'h3 : _GEN_18101; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18103 = 10'h2e == _T_378[9:0] ? 4'h3 : _GEN_18102; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18104 = 10'h2f == _T_378[9:0] ? 4'h3 : _GEN_18103; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18105 = 10'h30 == _T_378[9:0] ? 4'h3 : _GEN_18104; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18106 = 10'h31 == _T_378[9:0] ? 4'h5 : _GEN_18105; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18107 = 10'h32 == _T_378[9:0] ? 4'h3 : _GEN_18106; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18108 = 10'h33 == _T_378[9:0] ? 4'h3 : _GEN_18107; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18109 = 10'h34 == _T_378[9:0] ? 4'h3 : _GEN_18108; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18110 = 10'h35 == _T_378[9:0] ? 4'h3 : _GEN_18109; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18111 = 10'h36 == _T_378[9:0] ? 4'h3 : _GEN_18110; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18112 = 10'h37 == _T_378[9:0] ? 4'h1 : _GEN_18111; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18113 = 10'h38 == _T_378[9:0] ? 4'h1 : _GEN_18112; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18114 = 10'h39 == _T_378[9:0] ? 4'h3 : _GEN_18113; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18115 = 10'h3a == _T_378[9:0] ? 4'h3 : _GEN_18114; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18116 = 10'h3b == _T_378[9:0] ? 4'h5 : _GEN_18115; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18117 = 10'h3c == _T_378[9:0] ? 4'h3 : _GEN_18116; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18118 = 10'h3d == _T_378[9:0] ? 4'ha : _GEN_18117; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18119 = 10'h3e == _T_378[9:0] ? 4'h3 : _GEN_18118; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18120 = 10'h3f == _T_378[9:0] ? 4'h0 : _GEN_18119; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18121 = 10'h40 == _T_378[9:0] ? 4'h3 : _GEN_18120; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18122 = 10'h41 == _T_378[9:0] ? 4'h3 : _GEN_18121; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18123 = 10'h42 == _T_378[9:0] ? 4'h3 : _GEN_18122; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18124 = 10'h43 == _T_378[9:0] ? 4'h7 : _GEN_18123; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18125 = 10'h44 == _T_378[9:0] ? 4'ha : _GEN_18124; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18126 = 10'h45 == _T_378[9:0] ? 4'h0 : _GEN_18125; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18127 = 10'h46 == _T_378[9:0] ? 4'h0 : _GEN_18126; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18128 = 10'h47 == _T_378[9:0] ? 4'h0 : _GEN_18127; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18129 = 10'h48 == _T_378[9:0] ? 4'h0 : _GEN_18128; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18130 = 10'h49 == _T_378[9:0] ? 4'h3 : _GEN_18129; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18131 = 10'h4a == _T_378[9:0] ? 4'h3 : _GEN_18130; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18132 = 10'h4b == _T_378[9:0] ? 4'h3 : _GEN_18131; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18133 = 10'h4c == _T_378[9:0] ? 4'h3 : _GEN_18132; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18134 = 10'h4d == _T_378[9:0] ? 4'h5 : _GEN_18133; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18135 = 10'h4e == _T_378[9:0] ? 4'h3 : _GEN_18134; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18136 = 10'h4f == _T_378[9:0] ? 4'h3 : _GEN_18135; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18137 = 10'h50 == _T_378[9:0] ? 4'h3 : _GEN_18136; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18138 = 10'h51 == _T_378[9:0] ? 4'h3 : _GEN_18137; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18139 = 10'h52 == _T_378[9:0] ? 4'h3 : _GEN_18138; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18140 = 10'h53 == _T_378[9:0] ? 4'h3 : _GEN_18139; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18141 = 10'h54 == _T_378[9:0] ? 4'h1 : _GEN_18140; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18142 = 10'h55 == _T_378[9:0] ? 4'h1 : _GEN_18141; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18143 = 10'h56 == _T_378[9:0] ? 4'h1 : _GEN_18142; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18144 = 10'h57 == _T_378[9:0] ? 4'h0 : _GEN_18143; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18145 = 10'h58 == _T_378[9:0] ? 4'h3 : _GEN_18144; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18146 = 10'h59 == _T_378[9:0] ? 4'h0 : _GEN_18145; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18147 = 10'h5a == _T_378[9:0] ? 4'h3 : _GEN_18146; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18148 = 10'h5b == _T_378[9:0] ? 4'h3 : _GEN_18147; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18149 = 10'h5c == _T_378[9:0] ? 4'h3 : _GEN_18148; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18150 = 10'h5d == _T_378[9:0] ? 4'ha : _GEN_18149; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18151 = 10'h5e == _T_378[9:0] ? 4'h3 : _GEN_18150; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18152 = 10'h5f == _T_378[9:0] ? 4'h0 : _GEN_18151; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18153 = 10'h60 == _T_378[9:0] ? 4'h3 : _GEN_18152; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18154 = 10'h61 == _T_378[9:0] ? 4'h3 : _GEN_18153; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18155 = 10'h62 == _T_378[9:0] ? 4'h3 : _GEN_18154; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18156 = 10'h63 == _T_378[9:0] ? 4'h3 : _GEN_18155; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18157 = 10'h64 == _T_378[9:0] ? 4'ha : _GEN_18156; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18158 = 10'h65 == _T_378[9:0] ? 4'h0 : _GEN_18157; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18159 = 10'h66 == _T_378[9:0] ? 4'h3 : _GEN_18158; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18160 = 10'h67 == _T_378[9:0] ? 4'h3 : _GEN_18159; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18161 = 10'h68 == _T_378[9:0] ? 4'h3 : _GEN_18160; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18162 = 10'h69 == _T_378[9:0] ? 4'h0 : _GEN_18161; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18163 = 10'h6a == _T_378[9:0] ? 4'h1 : _GEN_18162; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18164 = 10'h6b == _T_378[9:0] ? 4'h1 : _GEN_18163; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18165 = 10'h6c == _T_378[9:0] ? 4'h3 : _GEN_18164; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18166 = 10'h6d == _T_378[9:0] ? 4'h3 : _GEN_18165; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18167 = 10'h6e == _T_378[9:0] ? 4'h3 : _GEN_18166; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18168 = 10'h6f == _T_378[9:0] ? 4'h3 : _GEN_18167; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18169 = 10'h70 == _T_378[9:0] ? 4'h3 : _GEN_18168; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18170 = 10'h71 == _T_378[9:0] ? 4'h3 : _GEN_18169; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18171 = 10'h72 == _T_378[9:0] ? 4'h3 : _GEN_18170; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18172 = 10'h73 == _T_378[9:0] ? 4'h1 : _GEN_18171; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18173 = 10'h74 == _T_378[9:0] ? 4'h0 : _GEN_18172; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18174 = 10'h75 == _T_378[9:0] ? 4'h0 : _GEN_18173; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18175 = 10'h76 == _T_378[9:0] ? 4'h0 : _GEN_18174; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18176 = 10'h77 == _T_378[9:0] ? 4'h3 : _GEN_18175; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18177 = 10'h78 == _T_378[9:0] ? 4'h3 : _GEN_18176; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18178 = 10'h79 == _T_378[9:0] ? 4'h3 : _GEN_18177; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18179 = 10'h7a == _T_378[9:0] ? 4'h0 : _GEN_18178; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18180 = 10'h7b == _T_378[9:0] ? 4'h3 : _GEN_18179; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18181 = 10'h7c == _T_378[9:0] ? 4'h3 : _GEN_18180; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18182 = 10'h7d == _T_378[9:0] ? 4'h7 : _GEN_18181; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18183 = 10'h7e == _T_378[9:0] ? 4'ha : _GEN_18182; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18184 = 10'h7f == _T_378[9:0] ? 4'h0 : _GEN_18183; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18185 = 10'h80 == _T_378[9:0] ? 4'h3 : _GEN_18184; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18186 = 10'h81 == _T_378[9:0] ? 4'h3 : _GEN_18185; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18187 = 10'h82 == _T_378[9:0] ? 4'h1 : _GEN_18186; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18188 = 10'h83 == _T_378[9:0] ? 4'h0 : _GEN_18187; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18189 = 10'h84 == _T_378[9:0] ? 4'h7 : _GEN_18188; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18190 = 10'h85 == _T_378[9:0] ? 4'h1 : _GEN_18189; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18191 = 10'h86 == _T_378[9:0] ? 4'h1 : _GEN_18190; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18192 = 10'h87 == _T_378[9:0] ? 4'h3 : _GEN_18191; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18193 = 10'h88 == _T_378[9:0] ? 4'h3 : _GEN_18192; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18194 = 10'h89 == _T_378[9:0] ? 4'h0 : _GEN_18193; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18195 = 10'h8a == _T_378[9:0] ? 4'h0 : _GEN_18194; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18196 = 10'h8b == _T_378[9:0] ? 4'h1 : _GEN_18195; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18197 = 10'h8c == _T_378[9:0] ? 4'h1 : _GEN_18196; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18198 = 10'h8d == _T_378[9:0] ? 4'h1 : _GEN_18197; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18199 = 10'h8e == _T_378[9:0] ? 4'h1 : _GEN_18198; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18200 = 10'h8f == _T_378[9:0] ? 4'h1 : _GEN_18199; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18201 = 10'h90 == _T_378[9:0] ? 4'h1 : _GEN_18200; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18202 = 10'h91 == _T_378[9:0] ? 4'h1 : _GEN_18201; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18203 = 10'h92 == _T_378[9:0] ? 4'h1 : _GEN_18202; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18204 = 10'h93 == _T_378[9:0] ? 4'h0 : _GEN_18203; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18205 = 10'h94 == _T_378[9:0] ? 4'h0 : _GEN_18204; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18206 = 10'h95 == _T_378[9:0] ? 4'h3 : _GEN_18205; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18207 = 10'h96 == _T_378[9:0] ? 4'h3 : _GEN_18206; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18208 = 10'h97 == _T_378[9:0] ? 4'h3 : _GEN_18207; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18209 = 10'h98 == _T_378[9:0] ? 4'h1 : _GEN_18208; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18210 = 10'h99 == _T_378[9:0] ? 4'h0 : _GEN_18209; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18211 = 10'h9a == _T_378[9:0] ? 4'h1 : _GEN_18210; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18212 = 10'h9b == _T_378[9:0] ? 4'h1 : _GEN_18211; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18213 = 10'h9c == _T_378[9:0] ? 4'h3 : _GEN_18212; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18214 = 10'h9d == _T_378[9:0] ? 4'h3 : _GEN_18213; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18215 = 10'h9e == _T_378[9:0] ? 4'ha : _GEN_18214; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18216 = 10'h9f == _T_378[9:0] ? 4'h0 : _GEN_18215; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18217 = 10'ha0 == _T_378[9:0] ? 4'h3 : _GEN_18216; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18218 = 10'ha1 == _T_378[9:0] ? 4'h1 : _GEN_18217; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18219 = 10'ha2 == _T_378[9:0] ? 4'h0 : _GEN_18218; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18220 = 10'ha3 == _T_378[9:0] ? 4'ha : _GEN_18219; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18221 = 10'ha4 == _T_378[9:0] ? 4'h3 : _GEN_18220; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18222 = 10'ha5 == _T_378[9:0] ? 4'h3 : _GEN_18221; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18223 = 10'ha6 == _T_378[9:0] ? 4'h3 : _GEN_18222; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18224 = 10'ha7 == _T_378[9:0] ? 4'h0 : _GEN_18223; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18225 = 10'ha8 == _T_378[9:0] ? 4'h3 : _GEN_18224; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18226 = 10'ha9 == _T_378[9:0] ? 4'h1 : _GEN_18225; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18227 = 10'haa == _T_378[9:0] ? 4'h0 : _GEN_18226; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18228 = 10'hab == _T_378[9:0] ? 4'h0 : _GEN_18227; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18229 = 10'hac == _T_378[9:0] ? 4'h0 : _GEN_18228; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18230 = 10'had == _T_378[9:0] ? 4'h0 : _GEN_18229; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18231 = 10'hae == _T_378[9:0] ? 4'h0 : _GEN_18230; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18232 = 10'haf == _T_378[9:0] ? 4'h0 : _GEN_18231; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18233 = 10'hb0 == _T_378[9:0] ? 4'h0 : _GEN_18232; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18234 = 10'hb1 == _T_378[9:0] ? 4'h0 : _GEN_18233; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18235 = 10'hb2 == _T_378[9:0] ? 4'h0 : _GEN_18234; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18236 = 10'hb3 == _T_378[9:0] ? 4'h0 : _GEN_18235; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18237 = 10'hb4 == _T_378[9:0] ? 4'h1 : _GEN_18236; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18238 = 10'hb5 == _T_378[9:0] ? 4'h1 : _GEN_18237; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18239 = 10'hb6 == _T_378[9:0] ? 4'h3 : _GEN_18238; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18240 = 10'hb7 == _T_378[9:0] ? 4'h0 : _GEN_18239; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18241 = 10'hb8 == _T_378[9:0] ? 4'h3 : _GEN_18240; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18242 = 10'hb9 == _T_378[9:0] ? 4'h3 : _GEN_18241; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18243 = 10'hba == _T_378[9:0] ? 4'h3 : _GEN_18242; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18244 = 10'hbb == _T_378[9:0] ? 4'h0 : _GEN_18243; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18245 = 10'hbc == _T_378[9:0] ? 4'h3 : _GEN_18244; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18246 = 10'hbd == _T_378[9:0] ? 4'h3 : _GEN_18245; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18247 = 10'hbe == _T_378[9:0] ? 4'ha : _GEN_18246; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18248 = 10'hbf == _T_378[9:0] ? 4'h0 : _GEN_18247; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18249 = 10'hc0 == _T_378[9:0] ? 4'h3 : _GEN_18248; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18250 = 10'hc1 == _T_378[9:0] ? 4'h3 : _GEN_18249; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18251 = 10'hc2 == _T_378[9:0] ? 4'ha : _GEN_18250; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18252 = 10'hc3 == _T_378[9:0] ? 4'h7 : _GEN_18251; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18253 = 10'hc4 == _T_378[9:0] ? 4'h0 : _GEN_18252; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18254 = 10'hc5 == _T_378[9:0] ? 4'h0 : _GEN_18253; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18255 = 10'hc6 == _T_378[9:0] ? 4'h0 : _GEN_18254; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18256 = 10'hc7 == _T_378[9:0] ? 4'h3 : _GEN_18255; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18257 = 10'hc8 == _T_378[9:0] ? 4'h1 : _GEN_18256; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18258 = 10'hc9 == _T_378[9:0] ? 4'h0 : _GEN_18257; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18259 = 10'hca == _T_378[9:0] ? 4'h0 : _GEN_18258; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18260 = 10'hcb == _T_378[9:0] ? 4'h0 : _GEN_18259; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18261 = 10'hcc == _T_378[9:0] ? 4'h0 : _GEN_18260; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18262 = 10'hcd == _T_378[9:0] ? 4'h0 : _GEN_18261; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18263 = 10'hce == _T_378[9:0] ? 4'h0 : _GEN_18262; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18264 = 10'hcf == _T_378[9:0] ? 4'h0 : _GEN_18263; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18265 = 10'hd0 == _T_378[9:0] ? 4'h0 : _GEN_18264; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18266 = 10'hd1 == _T_378[9:0] ? 4'h0 : _GEN_18265; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18267 = 10'hd2 == _T_378[9:0] ? 4'h0 : _GEN_18266; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18268 = 10'hd3 == _T_378[9:0] ? 4'h0 : _GEN_18267; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18269 = 10'hd4 == _T_378[9:0] ? 4'h0 : _GEN_18268; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18270 = 10'hd5 == _T_378[9:0] ? 4'h0 : _GEN_18269; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18271 = 10'hd6 == _T_378[9:0] ? 4'h1 : _GEN_18270; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18272 = 10'hd7 == _T_378[9:0] ? 4'h3 : _GEN_18271; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18273 = 10'hd8 == _T_378[9:0] ? 4'h0 : _GEN_18272; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18274 = 10'hd9 == _T_378[9:0] ? 4'h3 : _GEN_18273; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18275 = 10'hda == _T_378[9:0] ? 4'h3 : _GEN_18274; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18276 = 10'hdb == _T_378[9:0] ? 4'h3 : _GEN_18275; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18277 = 10'hdc == _T_378[9:0] ? 4'h3 : _GEN_18276; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18278 = 10'hdd == _T_378[9:0] ? 4'ha : _GEN_18277; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18279 = 10'hde == _T_378[9:0] ? 4'h7 : _GEN_18278; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18280 = 10'hdf == _T_378[9:0] ? 4'h0 : _GEN_18279; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18281 = 10'he0 == _T_378[9:0] ? 4'h3 : _GEN_18280; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18282 = 10'he1 == _T_378[9:0] ? 4'h3 : _GEN_18281; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18283 = 10'he2 == _T_378[9:0] ? 4'ha : _GEN_18282; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18284 = 10'he3 == _T_378[9:0] ? 4'h3 : _GEN_18283; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18285 = 10'he4 == _T_378[9:0] ? 4'h3 : _GEN_18284; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18286 = 10'he5 == _T_378[9:0] ? 4'h3 : _GEN_18285; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18287 = 10'he6 == _T_378[9:0] ? 4'h3 : _GEN_18286; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18288 = 10'he7 == _T_378[9:0] ? 4'h1 : _GEN_18287; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18289 = 10'he8 == _T_378[9:0] ? 4'h1 : _GEN_18288; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18290 = 10'he9 == _T_378[9:0] ? 4'h1 : _GEN_18289; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18291 = 10'hea == _T_378[9:0] ? 4'h0 : _GEN_18290; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18292 = 10'heb == _T_378[9:0] ? 4'h0 : _GEN_18291; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18293 = 10'hec == _T_378[9:0] ? 4'h0 : _GEN_18292; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18294 = 10'hed == _T_378[9:0] ? 4'h0 : _GEN_18293; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18295 = 10'hee == _T_378[9:0] ? 4'h0 : _GEN_18294; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18296 = 10'hef == _T_378[9:0] ? 4'h0 : _GEN_18295; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18297 = 10'hf0 == _T_378[9:0] ? 4'h0 : _GEN_18296; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18298 = 10'hf1 == _T_378[9:0] ? 4'h0 : _GEN_18297; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18299 = 10'hf2 == _T_378[9:0] ? 4'h0 : _GEN_18298; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18300 = 10'hf3 == _T_378[9:0] ? 4'h0 : _GEN_18299; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18301 = 10'hf4 == _T_378[9:0] ? 4'h0 : _GEN_18300; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18302 = 10'hf5 == _T_378[9:0] ? 4'h1 : _GEN_18301; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18303 = 10'hf6 == _T_378[9:0] ? 4'h0 : _GEN_18302; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18304 = 10'hf7 == _T_378[9:0] ? 4'h0 : _GEN_18303; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18305 = 10'hf8 == _T_378[9:0] ? 4'h1 : _GEN_18304; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18306 = 10'hf9 == _T_378[9:0] ? 4'h0 : _GEN_18305; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18307 = 10'hfa == _T_378[9:0] ? 4'h3 : _GEN_18306; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18308 = 10'hfb == _T_378[9:0] ? 4'h3 : _GEN_18307; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18309 = 10'hfc == _T_378[9:0] ? 4'h3 : _GEN_18308; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18310 = 10'hfd == _T_378[9:0] ? 4'ha : _GEN_18309; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18311 = 10'hfe == _T_378[9:0] ? 4'h3 : _GEN_18310; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18312 = 10'hff == _T_378[9:0] ? 4'h0 : _GEN_18311; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18313 = 10'h100 == _T_378[9:0] ? 4'h3 : _GEN_18312; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18314 = 10'h101 == _T_378[9:0] ? 4'h0 : _GEN_18313; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18315 = 10'h102 == _T_378[9:0] ? 4'ha : _GEN_18314; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18316 = 10'h103 == _T_378[9:0] ? 4'h3 : _GEN_18315; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18317 = 10'h104 == _T_378[9:0] ? 4'h3 : _GEN_18316; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18318 = 10'h105 == _T_378[9:0] ? 4'h3 : _GEN_18317; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18319 = 10'h106 == _T_378[9:0] ? 4'h3 : _GEN_18318; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18320 = 10'h107 == _T_378[9:0] ? 4'h3 : _GEN_18319; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18321 = 10'h108 == _T_378[9:0] ? 4'h1 : _GEN_18320; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18322 = 10'h109 == _T_378[9:0] ? 4'h0 : _GEN_18321; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18323 = 10'h10a == _T_378[9:0] ? 4'h0 : _GEN_18322; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18324 = 10'h10b == _T_378[9:0] ? 4'h0 : _GEN_18323; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18325 = 10'h10c == _T_378[9:0] ? 4'h0 : _GEN_18324; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18326 = 10'h10d == _T_378[9:0] ? 4'h0 : _GEN_18325; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18327 = 10'h10e == _T_378[9:0] ? 4'h0 : _GEN_18326; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18328 = 10'h10f == _T_378[9:0] ? 4'h0 : _GEN_18327; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18329 = 10'h110 == _T_378[9:0] ? 4'h0 : _GEN_18328; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18330 = 10'h111 == _T_378[9:0] ? 4'h0 : _GEN_18329; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18331 = 10'h112 == _T_378[9:0] ? 4'h0 : _GEN_18330; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18332 = 10'h113 == _T_378[9:0] ? 4'h0 : _GEN_18331; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18333 = 10'h114 == _T_378[9:0] ? 4'h0 : _GEN_18332; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18334 = 10'h115 == _T_378[9:0] ? 4'h0 : _GEN_18333; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18335 = 10'h116 == _T_378[9:0] ? 4'h1 : _GEN_18334; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18336 = 10'h117 == _T_378[9:0] ? 4'h3 : _GEN_18335; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18337 = 10'h118 == _T_378[9:0] ? 4'h3 : _GEN_18336; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18338 = 10'h119 == _T_378[9:0] ? 4'h3 : _GEN_18337; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18339 = 10'h11a == _T_378[9:0] ? 4'h0 : _GEN_18338; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18340 = 10'h11b == _T_378[9:0] ? 4'h3 : _GEN_18339; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18341 = 10'h11c == _T_378[9:0] ? 4'h3 : _GEN_18340; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18342 = 10'h11d == _T_378[9:0] ? 4'h7 : _GEN_18341; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18343 = 10'h11e == _T_378[9:0] ? 4'ha : _GEN_18342; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18344 = 10'h11f == _T_378[9:0] ? 4'h0 : _GEN_18343; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18345 = 10'h120 == _T_378[9:0] ? 4'h3 : _GEN_18344; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18346 = 10'h121 == _T_378[9:0] ? 4'h3 : _GEN_18345; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18347 = 10'h122 == _T_378[9:0] ? 4'ha : _GEN_18346; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18348 = 10'h123 == _T_378[9:0] ? 4'h3 : _GEN_18347; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18349 = 10'h124 == _T_378[9:0] ? 4'h3 : _GEN_18348; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18350 = 10'h125 == _T_378[9:0] ? 4'h3 : _GEN_18349; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18351 = 10'h126 == _T_378[9:0] ? 4'h3 : _GEN_18350; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18352 = 10'h127 == _T_378[9:0] ? 4'h1 : _GEN_18351; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18353 = 10'h128 == _T_378[9:0] ? 4'h0 : _GEN_18352; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18354 = 10'h129 == _T_378[9:0] ? 4'h3 : _GEN_18353; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18355 = 10'h12a == _T_378[9:0] ? 4'h3 : _GEN_18354; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18356 = 10'h12b == _T_378[9:0] ? 4'h0 : _GEN_18355; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18357 = 10'h12c == _T_378[9:0] ? 4'h0 : _GEN_18356; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18358 = 10'h12d == _T_378[9:0] ? 4'h0 : _GEN_18357; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18359 = 10'h12e == _T_378[9:0] ? 4'h0 : _GEN_18358; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18360 = 10'h12f == _T_378[9:0] ? 4'h0 : _GEN_18359; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18361 = 10'h130 == _T_378[9:0] ? 4'h0 : _GEN_18360; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18362 = 10'h131 == _T_378[9:0] ? 4'h0 : _GEN_18361; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18363 = 10'h132 == _T_378[9:0] ? 4'h0 : _GEN_18362; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18364 = 10'h133 == _T_378[9:0] ? 4'h0 : _GEN_18363; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18365 = 10'h134 == _T_378[9:0] ? 4'h3 : _GEN_18364; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18366 = 10'h135 == _T_378[9:0] ? 4'h3 : _GEN_18365; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18367 = 10'h136 == _T_378[9:0] ? 4'h0 : _GEN_18366; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18368 = 10'h137 == _T_378[9:0] ? 4'h1 : _GEN_18367; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18369 = 10'h138 == _T_378[9:0] ? 4'h3 : _GEN_18368; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18370 = 10'h139 == _T_378[9:0] ? 4'h3 : _GEN_18369; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18371 = 10'h13a == _T_378[9:0] ? 4'h3 : _GEN_18370; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18372 = 10'h13b == _T_378[9:0] ? 4'h3 : _GEN_18371; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18373 = 10'h13c == _T_378[9:0] ? 4'h3 : _GEN_18372; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18374 = 10'h13d == _T_378[9:0] ? 4'h3 : _GEN_18373; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18375 = 10'h13e == _T_378[9:0] ? 4'ha : _GEN_18374; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18376 = 10'h13f == _T_378[9:0] ? 4'h0 : _GEN_18375; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18377 = 10'h140 == _T_378[9:0] ? 4'h5 : _GEN_18376; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18378 = 10'h141 == _T_378[9:0] ? 4'h3 : _GEN_18377; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18379 = 10'h142 == _T_378[9:0] ? 4'h7 : _GEN_18378; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18380 = 10'h143 == _T_378[9:0] ? 4'ha : _GEN_18379; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18381 = 10'h144 == _T_378[9:0] ? 4'h3 : _GEN_18380; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18382 = 10'h145 == _T_378[9:0] ? 4'h3 : _GEN_18381; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18383 = 10'h146 == _T_378[9:0] ? 4'h1 : _GEN_18382; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18384 = 10'h147 == _T_378[9:0] ? 4'h0 : _GEN_18383; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18385 = 10'h148 == _T_378[9:0] ? 4'h3 : _GEN_18384; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18386 = 10'h149 == _T_378[9:0] ? 4'h3 : _GEN_18385; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18387 = 10'h14a == _T_378[9:0] ? 4'h3 : _GEN_18386; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18388 = 10'h14b == _T_378[9:0] ? 4'h3 : _GEN_18387; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18389 = 10'h14c == _T_378[9:0] ? 4'h3 : _GEN_18388; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18390 = 10'h14d == _T_378[9:0] ? 4'h3 : _GEN_18389; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18391 = 10'h14e == _T_378[9:0] ? 4'h3 : _GEN_18390; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18392 = 10'h14f == _T_378[9:0] ? 4'h3 : _GEN_18391; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18393 = 10'h150 == _T_378[9:0] ? 4'h3 : _GEN_18392; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18394 = 10'h151 == _T_378[9:0] ? 4'h3 : _GEN_18393; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18395 = 10'h152 == _T_378[9:0] ? 4'h3 : _GEN_18394; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18396 = 10'h153 == _T_378[9:0] ? 4'h3 : _GEN_18395; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18397 = 10'h154 == _T_378[9:0] ? 4'h3 : _GEN_18396; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18398 = 10'h155 == _T_378[9:0] ? 4'h3 : _GEN_18397; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18399 = 10'h156 == _T_378[9:0] ? 4'h3 : _GEN_18398; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18400 = 10'h157 == _T_378[9:0] ? 4'h0 : _GEN_18399; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18401 = 10'h158 == _T_378[9:0] ? 4'h3 : _GEN_18400; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18402 = 10'h159 == _T_378[9:0] ? 4'h3 : _GEN_18401; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18403 = 10'h15a == _T_378[9:0] ? 4'h3 : _GEN_18402; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18404 = 10'h15b == _T_378[9:0] ? 4'h3 : _GEN_18403; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18405 = 10'h15c == _T_378[9:0] ? 4'h3 : _GEN_18404; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18406 = 10'h15d == _T_378[9:0] ? 4'ha : _GEN_18405; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18407 = 10'h15e == _T_378[9:0] ? 4'h7 : _GEN_18406; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18408 = 10'h15f == _T_378[9:0] ? 4'h0 : _GEN_18407; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18409 = 10'h160 == _T_378[9:0] ? 4'h3 : _GEN_18408; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18410 = 10'h161 == _T_378[9:0] ? 4'h3 : _GEN_18409; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18411 = 10'h162 == _T_378[9:0] ? 4'h3 : _GEN_18410; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18412 = 10'h163 == _T_378[9:0] ? 4'h7 : _GEN_18411; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18413 = 10'h164 == _T_378[9:0] ? 4'ha : _GEN_18412; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18414 = 10'h165 == _T_378[9:0] ? 4'h1 : _GEN_18413; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18415 = 10'h166 == _T_378[9:0] ? 4'h0 : _GEN_18414; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18416 = 10'h167 == _T_378[9:0] ? 4'h0 : _GEN_18415; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18417 = 10'h168 == _T_378[9:0] ? 4'hc : _GEN_18416; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18418 = 10'h169 == _T_378[9:0] ? 4'h9 : _GEN_18417; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18419 = 10'h16a == _T_378[9:0] ? 4'hc : _GEN_18418; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18420 = 10'h16b == _T_378[9:0] ? 4'hc : _GEN_18419; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18421 = 10'h16c == _T_378[9:0] ? 4'h3 : _GEN_18420; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18422 = 10'h16d == _T_378[9:0] ? 4'h3 : _GEN_18421; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18423 = 10'h16e == _T_378[9:0] ? 4'h3 : _GEN_18422; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18424 = 10'h16f == _T_378[9:0] ? 4'h3 : _GEN_18423; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18425 = 10'h170 == _T_378[9:0] ? 4'h5 : _GEN_18424; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18426 = 10'h171 == _T_378[9:0] ? 4'h3 : _GEN_18425; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18427 = 10'h172 == _T_378[9:0] ? 4'h3 : _GEN_18426; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18428 = 10'h173 == _T_378[9:0] ? 4'h3 : _GEN_18427; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18429 = 10'h174 == _T_378[9:0] ? 4'h3 : _GEN_18428; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18430 = 10'h175 == _T_378[9:0] ? 4'h3 : _GEN_18429; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18431 = 10'h176 == _T_378[9:0] ? 4'h0 : _GEN_18430; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18432 = 10'h177 == _T_378[9:0] ? 4'h0 : _GEN_18431; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18433 = 10'h178 == _T_378[9:0] ? 4'h1 : _GEN_18432; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18434 = 10'h179 == _T_378[9:0] ? 4'h3 : _GEN_18433; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18435 = 10'h17a == _T_378[9:0] ? 4'h5 : _GEN_18434; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18436 = 10'h17b == _T_378[9:0] ? 4'h3 : _GEN_18435; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18437 = 10'h17c == _T_378[9:0] ? 4'ha : _GEN_18436; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18438 = 10'h17d == _T_378[9:0] ? 4'h7 : _GEN_18437; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18439 = 10'h17e == _T_378[9:0] ? 4'h3 : _GEN_18438; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18440 = 10'h17f == _T_378[9:0] ? 4'h0 : _GEN_18439; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18441 = 10'h180 == _T_378[9:0] ? 4'hc : _GEN_18440; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18442 = 10'h181 == _T_378[9:0] ? 4'hc : _GEN_18441; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18443 = 10'h182 == _T_378[9:0] ? 4'hc : _GEN_18442; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18444 = 10'h183 == _T_378[9:0] ? 4'hc : _GEN_18443; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18445 = 10'h184 == _T_378[9:0] ? 4'ha : _GEN_18444; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18446 = 10'h185 == _T_378[9:0] ? 4'h1 : _GEN_18445; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18447 = 10'h186 == _T_378[9:0] ? 4'hc : _GEN_18446; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18448 = 10'h187 == _T_378[9:0] ? 4'h0 : _GEN_18447; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18449 = 10'h188 == _T_378[9:0] ? 4'hc : _GEN_18448; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18450 = 10'h189 == _T_378[9:0] ? 4'hc : _GEN_18449; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18451 = 10'h18a == _T_378[9:0] ? 4'hc : _GEN_18450; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18452 = 10'h18b == _T_378[9:0] ? 4'hc : _GEN_18451; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18453 = 10'h18c == _T_378[9:0] ? 4'hc : _GEN_18452; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18454 = 10'h18d == _T_378[9:0] ? 4'hc : _GEN_18453; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18455 = 10'h18e == _T_378[9:0] ? 4'hc : _GEN_18454; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18456 = 10'h18f == _T_378[9:0] ? 4'hc : _GEN_18455; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18457 = 10'h190 == _T_378[9:0] ? 4'hc : _GEN_18456; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18458 = 10'h191 == _T_378[9:0] ? 4'hc : _GEN_18457; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18459 = 10'h192 == _T_378[9:0] ? 4'h9 : _GEN_18458; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18460 = 10'h193 == _T_378[9:0] ? 4'hc : _GEN_18459; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18461 = 10'h194 == _T_378[9:0] ? 4'hc : _GEN_18460; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18462 = 10'h195 == _T_378[9:0] ? 4'hc : _GEN_18461; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18463 = 10'h196 == _T_378[9:0] ? 4'h0 : _GEN_18462; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18464 = 10'h197 == _T_378[9:0] ? 4'h3 : _GEN_18463; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18465 = 10'h198 == _T_378[9:0] ? 4'h1 : _GEN_18464; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18466 = 10'h199 == _T_378[9:0] ? 4'h3 : _GEN_18465; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18467 = 10'h19a == _T_378[9:0] ? 4'h3 : _GEN_18466; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18468 = 10'h19b == _T_378[9:0] ? 4'h3 : _GEN_18467; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18469 = 10'h19c == _T_378[9:0] ? 4'ha : _GEN_18468; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18470 = 10'h19d == _T_378[9:0] ? 4'h3 : _GEN_18469; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18471 = 10'h19e == _T_378[9:0] ? 4'h3 : _GEN_18470; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18472 = 10'h19f == _T_378[9:0] ? 4'h0 : _GEN_18471; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18473 = 10'h1a0 == _T_378[9:0] ? 4'hc : _GEN_18472; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18474 = 10'h1a1 == _T_378[9:0] ? 4'hc : _GEN_18473; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18475 = 10'h1a2 == _T_378[9:0] ? 4'h9 : _GEN_18474; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18476 = 10'h1a3 == _T_378[9:0] ? 4'hc : _GEN_18475; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18477 = 10'h1a4 == _T_378[9:0] ? 4'ha : _GEN_18476; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18478 = 10'h1a5 == _T_378[9:0] ? 4'h0 : _GEN_18477; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18479 = 10'h1a6 == _T_378[9:0] ? 4'hc : _GEN_18478; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18480 = 10'h1a7 == _T_378[9:0] ? 4'h0 : _GEN_18479; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18481 = 10'h1a8 == _T_378[9:0] ? 4'hc : _GEN_18480; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18482 = 10'h1a9 == _T_378[9:0] ? 4'hc : _GEN_18481; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18483 = 10'h1aa == _T_378[9:0] ? 4'hc : _GEN_18482; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18484 = 10'h1ab == _T_378[9:0] ? 4'h9 : _GEN_18483; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18485 = 10'h1ac == _T_378[9:0] ? 4'hc : _GEN_18484; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18486 = 10'h1ad == _T_378[9:0] ? 4'hc : _GEN_18485; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18487 = 10'h1ae == _T_378[9:0] ? 4'hc : _GEN_18486; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18488 = 10'h1af == _T_378[9:0] ? 4'hc : _GEN_18487; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18489 = 10'h1b0 == _T_378[9:0] ? 4'hc : _GEN_18488; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18490 = 10'h1b1 == _T_378[9:0] ? 4'hc : _GEN_18489; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18491 = 10'h1b2 == _T_378[9:0] ? 4'hc : _GEN_18490; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18492 = 10'h1b3 == _T_378[9:0] ? 4'hc : _GEN_18491; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18493 = 10'h1b4 == _T_378[9:0] ? 4'hc : _GEN_18492; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18494 = 10'h1b5 == _T_378[9:0] ? 4'hc : _GEN_18493; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18495 = 10'h1b6 == _T_378[9:0] ? 4'h0 : _GEN_18494; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18496 = 10'h1b7 == _T_378[9:0] ? 4'hc : _GEN_18495; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18497 = 10'h1b8 == _T_378[9:0] ? 4'h0 : _GEN_18496; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18498 = 10'h1b9 == _T_378[9:0] ? 4'hc : _GEN_18497; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18499 = 10'h1ba == _T_378[9:0] ? 4'hc : _GEN_18498; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18500 = 10'h1bb == _T_378[9:0] ? 4'hc : _GEN_18499; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18501 = 10'h1bc == _T_378[9:0] ? 4'h7 : _GEN_18500; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18502 = 10'h1bd == _T_378[9:0] ? 4'ha : _GEN_18501; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18503 = 10'h1be == _T_378[9:0] ? 4'hc : _GEN_18502; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18504 = 10'h1bf == _T_378[9:0] ? 4'h0 : _GEN_18503; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18505 = 10'h1c0 == _T_378[9:0] ? 4'hc : _GEN_18504; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18506 = 10'h1c1 == _T_378[9:0] ? 4'hc : _GEN_18505; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18507 = 10'h1c2 == _T_378[9:0] ? 4'hc : _GEN_18506; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18508 = 10'h1c3 == _T_378[9:0] ? 4'h7 : _GEN_18507; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18509 = 10'h1c4 == _T_378[9:0] ? 4'h7 : _GEN_18508; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18510 = 10'h1c5 == _T_378[9:0] ? 4'hc : _GEN_18509; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18511 = 10'h1c6 == _T_378[9:0] ? 4'hc : _GEN_18510; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18512 = 10'h1c7 == _T_378[9:0] ? 4'hc : _GEN_18511; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18513 = 10'h1c8 == _T_378[9:0] ? 4'hc : _GEN_18512; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18514 = 10'h1c9 == _T_378[9:0] ? 4'hc : _GEN_18513; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18515 = 10'h1ca == _T_378[9:0] ? 4'hc : _GEN_18514; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18516 = 10'h1cb == _T_378[9:0] ? 4'hc : _GEN_18515; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18517 = 10'h1cc == _T_378[9:0] ? 4'hc : _GEN_18516; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18518 = 10'h1cd == _T_378[9:0] ? 4'hc : _GEN_18517; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18519 = 10'h1ce == _T_378[9:0] ? 4'hc : _GEN_18518; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18520 = 10'h1cf == _T_378[9:0] ? 4'hc : _GEN_18519; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18521 = 10'h1d0 == _T_378[9:0] ? 4'hc : _GEN_18520; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18522 = 10'h1d1 == _T_378[9:0] ? 4'hc : _GEN_18521; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18523 = 10'h1d2 == _T_378[9:0] ? 4'hc : _GEN_18522; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18524 = 10'h1d3 == _T_378[9:0] ? 4'hc : _GEN_18523; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18525 = 10'h1d4 == _T_378[9:0] ? 4'hc : _GEN_18524; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18526 = 10'h1d5 == _T_378[9:0] ? 4'hc : _GEN_18525; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18527 = 10'h1d6 == _T_378[9:0] ? 4'hc : _GEN_18526; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18528 = 10'h1d7 == _T_378[9:0] ? 4'hc : _GEN_18527; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18529 = 10'h1d8 == _T_378[9:0] ? 4'hc : _GEN_18528; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18530 = 10'h1d9 == _T_378[9:0] ? 4'hc : _GEN_18529; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18531 = 10'h1da == _T_378[9:0] ? 4'hc : _GEN_18530; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18532 = 10'h1db == _T_378[9:0] ? 4'hc : _GEN_18531; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18533 = 10'h1dc == _T_378[9:0] ? 4'hc : _GEN_18532; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18534 = 10'h1dd == _T_378[9:0] ? 4'ha : _GEN_18533; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18535 = 10'h1de == _T_378[9:0] ? 4'hc : _GEN_18534; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18536 = 10'h1df == _T_378[9:0] ? 4'h0 : _GEN_18535; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18537 = 10'h1e0 == _T_378[9:0] ? 4'h9 : _GEN_18536; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18538 = 10'h1e1 == _T_378[9:0] ? 4'hc : _GEN_18537; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18539 = 10'h1e2 == _T_378[9:0] ? 4'h7 : _GEN_18538; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18540 = 10'h1e3 == _T_378[9:0] ? 4'h7 : _GEN_18539; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18541 = 10'h1e4 == _T_378[9:0] ? 4'hc : _GEN_18540; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18542 = 10'h1e5 == _T_378[9:0] ? 4'hc : _GEN_18541; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18543 = 10'h1e6 == _T_378[9:0] ? 4'hc : _GEN_18542; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18544 = 10'h1e7 == _T_378[9:0] ? 4'hc : _GEN_18543; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18545 = 10'h1e8 == _T_378[9:0] ? 4'hc : _GEN_18544; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18546 = 10'h1e9 == _T_378[9:0] ? 4'hc : _GEN_18545; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18547 = 10'h1ea == _T_378[9:0] ? 4'hc : _GEN_18546; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18548 = 10'h1eb == _T_378[9:0] ? 4'hc : _GEN_18547; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18549 = 10'h1ec == _T_378[9:0] ? 4'hc : _GEN_18548; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18550 = 10'h1ed == _T_378[9:0] ? 4'hc : _GEN_18549; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18551 = 10'h1ee == _T_378[9:0] ? 4'hc : _GEN_18550; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18552 = 10'h1ef == _T_378[9:0] ? 4'hc : _GEN_18551; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18553 = 10'h1f0 == _T_378[9:0] ? 4'hc : _GEN_18552; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18554 = 10'h1f1 == _T_378[9:0] ? 4'hc : _GEN_18553; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18555 = 10'h1f2 == _T_378[9:0] ? 4'hc : _GEN_18554; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18556 = 10'h1f3 == _T_378[9:0] ? 4'hc : _GEN_18555; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18557 = 10'h1f4 == _T_378[9:0] ? 4'hc : _GEN_18556; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18558 = 10'h1f5 == _T_378[9:0] ? 4'hc : _GEN_18557; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18559 = 10'h1f6 == _T_378[9:0] ? 4'hc : _GEN_18558; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18560 = 10'h1f7 == _T_378[9:0] ? 4'hc : _GEN_18559; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18561 = 10'h1f8 == _T_378[9:0] ? 4'hc : _GEN_18560; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18562 = 10'h1f9 == _T_378[9:0] ? 4'hc : _GEN_18561; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18563 = 10'h1fa == _T_378[9:0] ? 4'h9 : _GEN_18562; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18564 = 10'h1fb == _T_378[9:0] ? 4'hc : _GEN_18563; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18565 = 10'h1fc == _T_378[9:0] ? 4'hc : _GEN_18564; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18566 = 10'h1fd == _T_378[9:0] ? 4'h7 : _GEN_18565; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18567 = 10'h1fe == _T_378[9:0] ? 4'hc : _GEN_18566; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18568 = 10'h1ff == _T_378[9:0] ? 4'h0 : _GEN_18567; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18569 = 10'h200 == _T_378[9:0] ? 4'hc : _GEN_18568; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18570 = 10'h201 == _T_378[9:0] ? 4'hc : _GEN_18569; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18571 = 10'h202 == _T_378[9:0] ? 4'ha : _GEN_18570; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18572 = 10'h203 == _T_378[9:0] ? 4'hc : _GEN_18571; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18573 = 10'h204 == _T_378[9:0] ? 4'hc : _GEN_18572; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18574 = 10'h205 == _T_378[9:0] ? 4'hc : _GEN_18573; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18575 = 10'h206 == _T_378[9:0] ? 4'hc : _GEN_18574; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18576 = 10'h207 == _T_378[9:0] ? 4'hc : _GEN_18575; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18577 = 10'h208 == _T_378[9:0] ? 4'hc : _GEN_18576; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18578 = 10'h209 == _T_378[9:0] ? 4'hc : _GEN_18577; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18579 = 10'h20a == _T_378[9:0] ? 4'hc : _GEN_18578; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18580 = 10'h20b == _T_378[9:0] ? 4'hc : _GEN_18579; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18581 = 10'h20c == _T_378[9:0] ? 4'hc : _GEN_18580; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18582 = 10'h20d == _T_378[9:0] ? 4'hc : _GEN_18581; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18583 = 10'h20e == _T_378[9:0] ? 4'hc : _GEN_18582; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18584 = 10'h20f == _T_378[9:0] ? 4'hc : _GEN_18583; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18585 = 10'h210 == _T_378[9:0] ? 4'hc : _GEN_18584; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18586 = 10'h211 == _T_378[9:0] ? 4'hc : _GEN_18585; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18587 = 10'h212 == _T_378[9:0] ? 4'hc : _GEN_18586; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18588 = 10'h213 == _T_378[9:0] ? 4'hc : _GEN_18587; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18589 = 10'h214 == _T_378[9:0] ? 4'hc : _GEN_18588; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18590 = 10'h215 == _T_378[9:0] ? 4'hc : _GEN_18589; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18591 = 10'h216 == _T_378[9:0] ? 4'hc : _GEN_18590; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18592 = 10'h217 == _T_378[9:0] ? 4'hc : _GEN_18591; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18593 = 10'h218 == _T_378[9:0] ? 4'hc : _GEN_18592; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18594 = 10'h219 == _T_378[9:0] ? 4'hc : _GEN_18593; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18595 = 10'h21a == _T_378[9:0] ? 4'hc : _GEN_18594; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18596 = 10'h21b == _T_378[9:0] ? 4'hc : _GEN_18595; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18597 = 10'h21c == _T_378[9:0] ? 4'ha : _GEN_18596; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18598 = 10'h21d == _T_378[9:0] ? 4'h7 : _GEN_18597; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18599 = 10'h21e == _T_378[9:0] ? 4'hc : _GEN_18598; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18600 = 10'h21f == _T_378[9:0] ? 4'h0 : _GEN_18599; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18601 = 10'h220 == _T_378[9:0] ? 4'h0 : _GEN_18600; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18602 = 10'h221 == _T_378[9:0] ? 4'h0 : _GEN_18601; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18603 = 10'h222 == _T_378[9:0] ? 4'h0 : _GEN_18602; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18604 = 10'h223 == _T_378[9:0] ? 4'h0 : _GEN_18603; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18605 = 10'h224 == _T_378[9:0] ? 4'h0 : _GEN_18604; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18606 = 10'h225 == _T_378[9:0] ? 4'h0 : _GEN_18605; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18607 = 10'h226 == _T_378[9:0] ? 4'h0 : _GEN_18606; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18608 = 10'h227 == _T_378[9:0] ? 4'h0 : _GEN_18607; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18609 = 10'h228 == _T_378[9:0] ? 4'h0 : _GEN_18608; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18610 = 10'h229 == _T_378[9:0] ? 4'h0 : _GEN_18609; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18611 = 10'h22a == _T_378[9:0] ? 4'h0 : _GEN_18610; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18612 = 10'h22b == _T_378[9:0] ? 4'h0 : _GEN_18611; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18613 = 10'h22c == _T_378[9:0] ? 4'h0 : _GEN_18612; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18614 = 10'h22d == _T_378[9:0] ? 4'h0 : _GEN_18613; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18615 = 10'h22e == _T_378[9:0] ? 4'h0 : _GEN_18614; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18616 = 10'h22f == _T_378[9:0] ? 4'h0 : _GEN_18615; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18617 = 10'h230 == _T_378[9:0] ? 4'h0 : _GEN_18616; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18618 = 10'h231 == _T_378[9:0] ? 4'h0 : _GEN_18617; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18619 = 10'h232 == _T_378[9:0] ? 4'h0 : _GEN_18618; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18620 = 10'h233 == _T_378[9:0] ? 4'h0 : _GEN_18619; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18621 = 10'h234 == _T_378[9:0] ? 4'h0 : _GEN_18620; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18622 = 10'h235 == _T_378[9:0] ? 4'h0 : _GEN_18621; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18623 = 10'h236 == _T_378[9:0] ? 4'h0 : _GEN_18622; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18624 = 10'h237 == _T_378[9:0] ? 4'h0 : _GEN_18623; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18625 = 10'h238 == _T_378[9:0] ? 4'h0 : _GEN_18624; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18626 = 10'h239 == _T_378[9:0] ? 4'h0 : _GEN_18625; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18627 = 10'h23a == _T_378[9:0] ? 4'h0 : _GEN_18626; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18628 = 10'h23b == _T_378[9:0] ? 4'h0 : _GEN_18627; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18629 = 10'h23c == _T_378[9:0] ? 4'h0 : _GEN_18628; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18630 = 10'h23d == _T_378[9:0] ? 4'h0 : _GEN_18629; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18631 = 10'h23e == _T_378[9:0] ? 4'h0 : _GEN_18630; // @[Filter.scala 191:102]
  wire [3:0] _GEN_18632 = 10'h23f == _T_378[9:0] ? 4'h0 : _GEN_18631; // @[Filter.scala 191:102]
  wire [6:0] _GEN_28360 = {{3'd0}, _GEN_18632}; // @[Filter.scala 191:102]
  wire [10:0] _T_385 = _GEN_28360 * 7'h46; // @[Filter.scala 191:102]
  wire [10:0] _GEN_28361 = {{2'd0}, _T_380}; // @[Filter.scala 191:69]
  wire [10:0] _T_387 = _GEN_28361 + _T_385; // @[Filter.scala 191:69]
  wire [3:0] _GEN_18664 = 10'h1f == _T_378[9:0] ? 4'h0 : 4'h3; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18665 = 10'h20 == _T_378[9:0] ? 4'h3 : _GEN_18664; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18666 = 10'h21 == _T_378[9:0] ? 4'h3 : _GEN_18665; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18667 = 10'h22 == _T_378[9:0] ? 4'h3 : _GEN_18666; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18668 = 10'h23 == _T_378[9:0] ? 4'h3 : _GEN_18667; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18669 = 10'h24 == _T_378[9:0] ? 4'h3 : _GEN_18668; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18670 = 10'h25 == _T_378[9:0] ? 4'h3 : _GEN_18669; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18671 = 10'h26 == _T_378[9:0] ? 4'h3 : _GEN_18670; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18672 = 10'h27 == _T_378[9:0] ? 4'h9 : _GEN_18671; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18673 = 10'h28 == _T_378[9:0] ? 4'h9 : _GEN_18672; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18674 = 10'h29 == _T_378[9:0] ? 4'h3 : _GEN_18673; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18675 = 10'h2a == _T_378[9:0] ? 4'h3 : _GEN_18674; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18676 = 10'h2b == _T_378[9:0] ? 4'h3 : _GEN_18675; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18677 = 10'h2c == _T_378[9:0] ? 4'h3 : _GEN_18676; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18678 = 10'h2d == _T_378[9:0] ? 4'h3 : _GEN_18677; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18679 = 10'h2e == _T_378[9:0] ? 4'h3 : _GEN_18678; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18680 = 10'h2f == _T_378[9:0] ? 4'h3 : _GEN_18679; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18681 = 10'h30 == _T_378[9:0] ? 4'h3 : _GEN_18680; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18682 = 10'h31 == _T_378[9:0] ? 4'h3 : _GEN_18681; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18683 = 10'h32 == _T_378[9:0] ? 4'h3 : _GEN_18682; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18684 = 10'h33 == _T_378[9:0] ? 4'h3 : _GEN_18683; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18685 = 10'h34 == _T_378[9:0] ? 4'h3 : _GEN_18684; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18686 = 10'h35 == _T_378[9:0] ? 4'h3 : _GEN_18685; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18687 = 10'h36 == _T_378[9:0] ? 4'h3 : _GEN_18686; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18688 = 10'h37 == _T_378[9:0] ? 4'h9 : _GEN_18687; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18689 = 10'h38 == _T_378[9:0] ? 4'h9 : _GEN_18688; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18690 = 10'h39 == _T_378[9:0] ? 4'h3 : _GEN_18689; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18691 = 10'h3a == _T_378[9:0] ? 4'h3 : _GEN_18690; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18692 = 10'h3b == _T_378[9:0] ? 4'h3 : _GEN_18691; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18693 = 10'h3c == _T_378[9:0] ? 4'h3 : _GEN_18692; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18694 = 10'h3d == _T_378[9:0] ? 4'h3 : _GEN_18693; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18695 = 10'h3e == _T_378[9:0] ? 4'h3 : _GEN_18694; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18696 = 10'h3f == _T_378[9:0] ? 4'h0 : _GEN_18695; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18697 = 10'h40 == _T_378[9:0] ? 4'h3 : _GEN_18696; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18698 = 10'h41 == _T_378[9:0] ? 4'h3 : _GEN_18697; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18699 = 10'h42 == _T_378[9:0] ? 4'h3 : _GEN_18698; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18700 = 10'h43 == _T_378[9:0] ? 4'h2 : _GEN_18699; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18701 = 10'h44 == _T_378[9:0] ? 4'h3 : _GEN_18700; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18702 = 10'h45 == _T_378[9:0] ? 4'hf : _GEN_18701; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18703 = 10'h46 == _T_378[9:0] ? 4'hf : _GEN_18702; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18704 = 10'h47 == _T_378[9:0] ? 4'hf : _GEN_18703; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18705 = 10'h48 == _T_378[9:0] ? 4'hf : _GEN_18704; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18706 = 10'h49 == _T_378[9:0] ? 4'h3 : _GEN_18705; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18707 = 10'h4a == _T_378[9:0] ? 4'h3 : _GEN_18706; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18708 = 10'h4b == _T_378[9:0] ? 4'h3 : _GEN_18707; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18709 = 10'h4c == _T_378[9:0] ? 4'h3 : _GEN_18708; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18710 = 10'h4d == _T_378[9:0] ? 4'h3 : _GEN_18709; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18711 = 10'h4e == _T_378[9:0] ? 4'h3 : _GEN_18710; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18712 = 10'h4f == _T_378[9:0] ? 4'h3 : _GEN_18711; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18713 = 10'h50 == _T_378[9:0] ? 4'h3 : _GEN_18712; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18714 = 10'h51 == _T_378[9:0] ? 4'h3 : _GEN_18713; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18715 = 10'h52 == _T_378[9:0] ? 4'h3 : _GEN_18714; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18716 = 10'h53 == _T_378[9:0] ? 4'h3 : _GEN_18715; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18717 = 10'h54 == _T_378[9:0] ? 4'h9 : _GEN_18716; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18718 = 10'h55 == _T_378[9:0] ? 4'h9 : _GEN_18717; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18719 = 10'h56 == _T_378[9:0] ? 4'h9 : _GEN_18718; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18720 = 10'h57 == _T_378[9:0] ? 4'hf : _GEN_18719; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18721 = 10'h58 == _T_378[9:0] ? 4'h3 : _GEN_18720; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18722 = 10'h59 == _T_378[9:0] ? 4'hf : _GEN_18721; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18723 = 10'h5a == _T_378[9:0] ? 4'h3 : _GEN_18722; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18724 = 10'h5b == _T_378[9:0] ? 4'h3 : _GEN_18723; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18725 = 10'h5c == _T_378[9:0] ? 4'h3 : _GEN_18724; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18726 = 10'h5d == _T_378[9:0] ? 4'h3 : _GEN_18725; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18727 = 10'h5e == _T_378[9:0] ? 4'h3 : _GEN_18726; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18728 = 10'h5f == _T_378[9:0] ? 4'h0 : _GEN_18727; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18729 = 10'h60 == _T_378[9:0] ? 4'h3 : _GEN_18728; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18730 = 10'h61 == _T_378[9:0] ? 4'h3 : _GEN_18729; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18731 = 10'h62 == _T_378[9:0] ? 4'h3 : _GEN_18730; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18732 = 10'h63 == _T_378[9:0] ? 4'h3 : _GEN_18731; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18733 = 10'h64 == _T_378[9:0] ? 4'h3 : _GEN_18732; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18734 = 10'h65 == _T_378[9:0] ? 4'hf : _GEN_18733; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18735 = 10'h66 == _T_378[9:0] ? 4'h3 : _GEN_18734; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18736 = 10'h67 == _T_378[9:0] ? 4'h3 : _GEN_18735; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18737 = 10'h68 == _T_378[9:0] ? 4'h3 : _GEN_18736; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18738 = 10'h69 == _T_378[9:0] ? 4'hf : _GEN_18737; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18739 = 10'h6a == _T_378[9:0] ? 4'h9 : _GEN_18738; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18740 = 10'h6b == _T_378[9:0] ? 4'h9 : _GEN_18739; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18741 = 10'h6c == _T_378[9:0] ? 4'h3 : _GEN_18740; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18742 = 10'h6d == _T_378[9:0] ? 4'h3 : _GEN_18741; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18743 = 10'h6e == _T_378[9:0] ? 4'h3 : _GEN_18742; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18744 = 10'h6f == _T_378[9:0] ? 4'h3 : _GEN_18743; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18745 = 10'h70 == _T_378[9:0] ? 4'h3 : _GEN_18744; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18746 = 10'h71 == _T_378[9:0] ? 4'h3 : _GEN_18745; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18747 = 10'h72 == _T_378[9:0] ? 4'h3 : _GEN_18746; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18748 = 10'h73 == _T_378[9:0] ? 4'h9 : _GEN_18747; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18749 = 10'h74 == _T_378[9:0] ? 4'hf : _GEN_18748; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18750 = 10'h75 == _T_378[9:0] ? 4'hf : _GEN_18749; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18751 = 10'h76 == _T_378[9:0] ? 4'hf : _GEN_18750; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18752 = 10'h77 == _T_378[9:0] ? 4'h3 : _GEN_18751; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18753 = 10'h78 == _T_378[9:0] ? 4'h3 : _GEN_18752; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18754 = 10'h79 == _T_378[9:0] ? 4'h3 : _GEN_18753; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18755 = 10'h7a == _T_378[9:0] ? 4'hf : _GEN_18754; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18756 = 10'h7b == _T_378[9:0] ? 4'h3 : _GEN_18755; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18757 = 10'h7c == _T_378[9:0] ? 4'h3 : _GEN_18756; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18758 = 10'h7d == _T_378[9:0] ? 4'h2 : _GEN_18757; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18759 = 10'h7e == _T_378[9:0] ? 4'h3 : _GEN_18758; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18760 = 10'h7f == _T_378[9:0] ? 4'h0 : _GEN_18759; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18761 = 10'h80 == _T_378[9:0] ? 4'h3 : _GEN_18760; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18762 = 10'h81 == _T_378[9:0] ? 4'h3 : _GEN_18761; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18763 = 10'h82 == _T_378[9:0] ? 4'h9 : _GEN_18762; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18764 = 10'h83 == _T_378[9:0] ? 4'hf : _GEN_18763; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18765 = 10'h84 == _T_378[9:0] ? 4'h2 : _GEN_18764; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18766 = 10'h85 == _T_378[9:0] ? 4'h9 : _GEN_18765; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18767 = 10'h86 == _T_378[9:0] ? 4'h9 : _GEN_18766; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18768 = 10'h87 == _T_378[9:0] ? 4'h3 : _GEN_18767; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18769 = 10'h88 == _T_378[9:0] ? 4'h3 : _GEN_18768; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18770 = 10'h89 == _T_378[9:0] ? 4'hf : _GEN_18769; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18771 = 10'h8a == _T_378[9:0] ? 4'hf : _GEN_18770; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18772 = 10'h8b == _T_378[9:0] ? 4'h9 : _GEN_18771; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18773 = 10'h8c == _T_378[9:0] ? 4'h9 : _GEN_18772; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18774 = 10'h8d == _T_378[9:0] ? 4'h9 : _GEN_18773; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18775 = 10'h8e == _T_378[9:0] ? 4'h9 : _GEN_18774; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18776 = 10'h8f == _T_378[9:0] ? 4'h9 : _GEN_18775; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18777 = 10'h90 == _T_378[9:0] ? 4'h9 : _GEN_18776; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18778 = 10'h91 == _T_378[9:0] ? 4'h9 : _GEN_18777; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18779 = 10'h92 == _T_378[9:0] ? 4'h9 : _GEN_18778; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18780 = 10'h93 == _T_378[9:0] ? 4'hf : _GEN_18779; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18781 = 10'h94 == _T_378[9:0] ? 4'hf : _GEN_18780; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18782 = 10'h95 == _T_378[9:0] ? 4'h3 : _GEN_18781; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18783 = 10'h96 == _T_378[9:0] ? 4'h3 : _GEN_18782; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18784 = 10'h97 == _T_378[9:0] ? 4'h3 : _GEN_18783; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18785 = 10'h98 == _T_378[9:0] ? 4'h9 : _GEN_18784; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18786 = 10'h99 == _T_378[9:0] ? 4'hf : _GEN_18785; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18787 = 10'h9a == _T_378[9:0] ? 4'h9 : _GEN_18786; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18788 = 10'h9b == _T_378[9:0] ? 4'h9 : _GEN_18787; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18789 = 10'h9c == _T_378[9:0] ? 4'h3 : _GEN_18788; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18790 = 10'h9d == _T_378[9:0] ? 4'h3 : _GEN_18789; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18791 = 10'h9e == _T_378[9:0] ? 4'h3 : _GEN_18790; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18792 = 10'h9f == _T_378[9:0] ? 4'h0 : _GEN_18791; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18793 = 10'ha0 == _T_378[9:0] ? 4'h3 : _GEN_18792; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18794 = 10'ha1 == _T_378[9:0] ? 4'h9 : _GEN_18793; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18795 = 10'ha2 == _T_378[9:0] ? 4'hf : _GEN_18794; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18796 = 10'ha3 == _T_378[9:0] ? 4'h3 : _GEN_18795; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18797 = 10'ha4 == _T_378[9:0] ? 4'h3 : _GEN_18796; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18798 = 10'ha5 == _T_378[9:0] ? 4'h3 : _GEN_18797; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18799 = 10'ha6 == _T_378[9:0] ? 4'h3 : _GEN_18798; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18800 = 10'ha7 == _T_378[9:0] ? 4'hf : _GEN_18799; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18801 = 10'ha8 == _T_378[9:0] ? 4'h3 : _GEN_18800; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18802 = 10'ha9 == _T_378[9:0] ? 4'h9 : _GEN_18801; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18803 = 10'haa == _T_378[9:0] ? 4'hf : _GEN_18802; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18804 = 10'hab == _T_378[9:0] ? 4'hf : _GEN_18803; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18805 = 10'hac == _T_378[9:0] ? 4'hf : _GEN_18804; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18806 = 10'had == _T_378[9:0] ? 4'hf : _GEN_18805; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18807 = 10'hae == _T_378[9:0] ? 4'hf : _GEN_18806; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18808 = 10'haf == _T_378[9:0] ? 4'hf : _GEN_18807; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18809 = 10'hb0 == _T_378[9:0] ? 4'hf : _GEN_18808; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18810 = 10'hb1 == _T_378[9:0] ? 4'hf : _GEN_18809; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18811 = 10'hb2 == _T_378[9:0] ? 4'hf : _GEN_18810; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18812 = 10'hb3 == _T_378[9:0] ? 4'hf : _GEN_18811; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18813 = 10'hb4 == _T_378[9:0] ? 4'h9 : _GEN_18812; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18814 = 10'hb5 == _T_378[9:0] ? 4'h9 : _GEN_18813; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18815 = 10'hb6 == _T_378[9:0] ? 4'h3 : _GEN_18814; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18816 = 10'hb7 == _T_378[9:0] ? 4'hf : _GEN_18815; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18817 = 10'hb8 == _T_378[9:0] ? 4'h3 : _GEN_18816; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18818 = 10'hb9 == _T_378[9:0] ? 4'h3 : _GEN_18817; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18819 = 10'hba == _T_378[9:0] ? 4'h3 : _GEN_18818; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18820 = 10'hbb == _T_378[9:0] ? 4'hf : _GEN_18819; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18821 = 10'hbc == _T_378[9:0] ? 4'h3 : _GEN_18820; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18822 = 10'hbd == _T_378[9:0] ? 4'h3 : _GEN_18821; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18823 = 10'hbe == _T_378[9:0] ? 4'h3 : _GEN_18822; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18824 = 10'hbf == _T_378[9:0] ? 4'h0 : _GEN_18823; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18825 = 10'hc0 == _T_378[9:0] ? 4'h3 : _GEN_18824; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18826 = 10'hc1 == _T_378[9:0] ? 4'h3 : _GEN_18825; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18827 = 10'hc2 == _T_378[9:0] ? 4'h3 : _GEN_18826; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18828 = 10'hc3 == _T_378[9:0] ? 4'h2 : _GEN_18827; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18829 = 10'hc4 == _T_378[9:0] ? 4'hf : _GEN_18828; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18830 = 10'hc5 == _T_378[9:0] ? 4'hf : _GEN_18829; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18831 = 10'hc6 == _T_378[9:0] ? 4'hf : _GEN_18830; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18832 = 10'hc7 == _T_378[9:0] ? 4'h3 : _GEN_18831; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18833 = 10'hc8 == _T_378[9:0] ? 4'h9 : _GEN_18832; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18834 = 10'hc9 == _T_378[9:0] ? 4'hf : _GEN_18833; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18835 = 10'hca == _T_378[9:0] ? 4'hf : _GEN_18834; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18836 = 10'hcb == _T_378[9:0] ? 4'hf : _GEN_18835; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18837 = 10'hcc == _T_378[9:0] ? 4'hf : _GEN_18836; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18838 = 10'hcd == _T_378[9:0] ? 4'hf : _GEN_18837; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18839 = 10'hce == _T_378[9:0] ? 4'hf : _GEN_18838; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18840 = 10'hcf == _T_378[9:0] ? 4'hf : _GEN_18839; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18841 = 10'hd0 == _T_378[9:0] ? 4'hf : _GEN_18840; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18842 = 10'hd1 == _T_378[9:0] ? 4'hf : _GEN_18841; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18843 = 10'hd2 == _T_378[9:0] ? 4'hf : _GEN_18842; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18844 = 10'hd3 == _T_378[9:0] ? 4'hf : _GEN_18843; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18845 = 10'hd4 == _T_378[9:0] ? 4'hf : _GEN_18844; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18846 = 10'hd5 == _T_378[9:0] ? 4'hf : _GEN_18845; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18847 = 10'hd6 == _T_378[9:0] ? 4'h9 : _GEN_18846; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18848 = 10'hd7 == _T_378[9:0] ? 4'h3 : _GEN_18847; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18849 = 10'hd8 == _T_378[9:0] ? 4'hf : _GEN_18848; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18850 = 10'hd9 == _T_378[9:0] ? 4'h3 : _GEN_18849; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18851 = 10'hda == _T_378[9:0] ? 4'h3 : _GEN_18850; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18852 = 10'hdb == _T_378[9:0] ? 4'h3 : _GEN_18851; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18853 = 10'hdc == _T_378[9:0] ? 4'h3 : _GEN_18852; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18854 = 10'hdd == _T_378[9:0] ? 4'h3 : _GEN_18853; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18855 = 10'hde == _T_378[9:0] ? 4'h2 : _GEN_18854; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18856 = 10'hdf == _T_378[9:0] ? 4'h0 : _GEN_18855; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18857 = 10'he0 == _T_378[9:0] ? 4'h3 : _GEN_18856; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18858 = 10'he1 == _T_378[9:0] ? 4'h3 : _GEN_18857; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18859 = 10'he2 == _T_378[9:0] ? 4'h3 : _GEN_18858; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18860 = 10'he3 == _T_378[9:0] ? 4'h3 : _GEN_18859; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18861 = 10'he4 == _T_378[9:0] ? 4'h3 : _GEN_18860; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18862 = 10'he5 == _T_378[9:0] ? 4'h3 : _GEN_18861; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18863 = 10'he6 == _T_378[9:0] ? 4'h3 : _GEN_18862; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18864 = 10'he7 == _T_378[9:0] ? 4'h9 : _GEN_18863; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18865 = 10'he8 == _T_378[9:0] ? 4'h9 : _GEN_18864; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18866 = 10'he9 == _T_378[9:0] ? 4'h9 : _GEN_18865; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18867 = 10'hea == _T_378[9:0] ? 4'hf : _GEN_18866; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18868 = 10'heb == _T_378[9:0] ? 4'hf : _GEN_18867; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18869 = 10'hec == _T_378[9:0] ? 4'hf : _GEN_18868; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18870 = 10'hed == _T_378[9:0] ? 4'hf : _GEN_18869; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18871 = 10'hee == _T_378[9:0] ? 4'hf : _GEN_18870; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18872 = 10'hef == _T_378[9:0] ? 4'hf : _GEN_18871; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18873 = 10'hf0 == _T_378[9:0] ? 4'hf : _GEN_18872; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18874 = 10'hf1 == _T_378[9:0] ? 4'hf : _GEN_18873; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18875 = 10'hf2 == _T_378[9:0] ? 4'hf : _GEN_18874; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18876 = 10'hf3 == _T_378[9:0] ? 4'hf : _GEN_18875; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18877 = 10'hf4 == _T_378[9:0] ? 4'hf : _GEN_18876; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18878 = 10'hf5 == _T_378[9:0] ? 4'h9 : _GEN_18877; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18879 = 10'hf6 == _T_378[9:0] ? 4'hf : _GEN_18878; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18880 = 10'hf7 == _T_378[9:0] ? 4'hf : _GEN_18879; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18881 = 10'hf8 == _T_378[9:0] ? 4'h9 : _GEN_18880; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18882 = 10'hf9 == _T_378[9:0] ? 4'hf : _GEN_18881; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18883 = 10'hfa == _T_378[9:0] ? 4'h3 : _GEN_18882; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18884 = 10'hfb == _T_378[9:0] ? 4'h3 : _GEN_18883; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18885 = 10'hfc == _T_378[9:0] ? 4'h3 : _GEN_18884; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18886 = 10'hfd == _T_378[9:0] ? 4'h3 : _GEN_18885; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18887 = 10'hfe == _T_378[9:0] ? 4'h3 : _GEN_18886; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18888 = 10'hff == _T_378[9:0] ? 4'h0 : _GEN_18887; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18889 = 10'h100 == _T_378[9:0] ? 4'h3 : _GEN_18888; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18890 = 10'h101 == _T_378[9:0] ? 4'hf : _GEN_18889; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18891 = 10'h102 == _T_378[9:0] ? 4'h3 : _GEN_18890; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18892 = 10'h103 == _T_378[9:0] ? 4'h3 : _GEN_18891; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18893 = 10'h104 == _T_378[9:0] ? 4'h3 : _GEN_18892; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18894 = 10'h105 == _T_378[9:0] ? 4'h3 : _GEN_18893; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18895 = 10'h106 == _T_378[9:0] ? 4'h3 : _GEN_18894; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18896 = 10'h107 == _T_378[9:0] ? 4'h3 : _GEN_18895; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18897 = 10'h108 == _T_378[9:0] ? 4'h9 : _GEN_18896; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18898 = 10'h109 == _T_378[9:0] ? 4'hf : _GEN_18897; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18899 = 10'h10a == _T_378[9:0] ? 4'hf : _GEN_18898; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18900 = 10'h10b == _T_378[9:0] ? 4'hf : _GEN_18899; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18901 = 10'h10c == _T_378[9:0] ? 4'hf : _GEN_18900; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18902 = 10'h10d == _T_378[9:0] ? 4'h0 : _GEN_18901; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18903 = 10'h10e == _T_378[9:0] ? 4'hf : _GEN_18902; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18904 = 10'h10f == _T_378[9:0] ? 4'hf : _GEN_18903; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18905 = 10'h110 == _T_378[9:0] ? 4'hf : _GEN_18904; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18906 = 10'h111 == _T_378[9:0] ? 4'h0 : _GEN_18905; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18907 = 10'h112 == _T_378[9:0] ? 4'hf : _GEN_18906; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18908 = 10'h113 == _T_378[9:0] ? 4'hf : _GEN_18907; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18909 = 10'h114 == _T_378[9:0] ? 4'hf : _GEN_18908; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18910 = 10'h115 == _T_378[9:0] ? 4'hf : _GEN_18909; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18911 = 10'h116 == _T_378[9:0] ? 4'h9 : _GEN_18910; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18912 = 10'h117 == _T_378[9:0] ? 4'h3 : _GEN_18911; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18913 = 10'h118 == _T_378[9:0] ? 4'h3 : _GEN_18912; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18914 = 10'h119 == _T_378[9:0] ? 4'h3 : _GEN_18913; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18915 = 10'h11a == _T_378[9:0] ? 4'hf : _GEN_18914; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18916 = 10'h11b == _T_378[9:0] ? 4'h3 : _GEN_18915; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18917 = 10'h11c == _T_378[9:0] ? 4'h3 : _GEN_18916; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18918 = 10'h11d == _T_378[9:0] ? 4'h2 : _GEN_18917; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18919 = 10'h11e == _T_378[9:0] ? 4'h3 : _GEN_18918; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18920 = 10'h11f == _T_378[9:0] ? 4'h0 : _GEN_18919; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18921 = 10'h120 == _T_378[9:0] ? 4'h3 : _GEN_18920; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18922 = 10'h121 == _T_378[9:0] ? 4'h3 : _GEN_18921; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18923 = 10'h122 == _T_378[9:0] ? 4'h3 : _GEN_18922; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18924 = 10'h123 == _T_378[9:0] ? 4'h3 : _GEN_18923; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18925 = 10'h124 == _T_378[9:0] ? 4'h3 : _GEN_18924; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18926 = 10'h125 == _T_378[9:0] ? 4'h3 : _GEN_18925; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18927 = 10'h126 == _T_378[9:0] ? 4'h3 : _GEN_18926; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18928 = 10'h127 == _T_378[9:0] ? 4'h9 : _GEN_18927; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18929 = 10'h128 == _T_378[9:0] ? 4'hf : _GEN_18928; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18930 = 10'h129 == _T_378[9:0] ? 4'h3 : _GEN_18929; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18931 = 10'h12a == _T_378[9:0] ? 4'h3 : _GEN_18930; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18932 = 10'h12b == _T_378[9:0] ? 4'hf : _GEN_18931; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18933 = 10'h12c == _T_378[9:0] ? 4'hf : _GEN_18932; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18934 = 10'h12d == _T_378[9:0] ? 4'hf : _GEN_18933; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18935 = 10'h12e == _T_378[9:0] ? 4'hf : _GEN_18934; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18936 = 10'h12f == _T_378[9:0] ? 4'hf : _GEN_18935; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18937 = 10'h130 == _T_378[9:0] ? 4'hf : _GEN_18936; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18938 = 10'h131 == _T_378[9:0] ? 4'hf : _GEN_18937; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18939 = 10'h132 == _T_378[9:0] ? 4'hf : _GEN_18938; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18940 = 10'h133 == _T_378[9:0] ? 4'hf : _GEN_18939; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18941 = 10'h134 == _T_378[9:0] ? 4'h3 : _GEN_18940; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18942 = 10'h135 == _T_378[9:0] ? 4'h3 : _GEN_18941; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18943 = 10'h136 == _T_378[9:0] ? 4'hf : _GEN_18942; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18944 = 10'h137 == _T_378[9:0] ? 4'h9 : _GEN_18943; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18945 = 10'h138 == _T_378[9:0] ? 4'h3 : _GEN_18944; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18946 = 10'h139 == _T_378[9:0] ? 4'h3 : _GEN_18945; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18947 = 10'h13a == _T_378[9:0] ? 4'h3 : _GEN_18946; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18948 = 10'h13b == _T_378[9:0] ? 4'h3 : _GEN_18947; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18949 = 10'h13c == _T_378[9:0] ? 4'h3 : _GEN_18948; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18950 = 10'h13d == _T_378[9:0] ? 4'h3 : _GEN_18949; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18951 = 10'h13e == _T_378[9:0] ? 4'h3 : _GEN_18950; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18952 = 10'h13f == _T_378[9:0] ? 4'h0 : _GEN_18951; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18953 = 10'h140 == _T_378[9:0] ? 4'h3 : _GEN_18952; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18954 = 10'h141 == _T_378[9:0] ? 4'h3 : _GEN_18953; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18955 = 10'h142 == _T_378[9:0] ? 4'h2 : _GEN_18954; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18956 = 10'h143 == _T_378[9:0] ? 4'h3 : _GEN_18955; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18957 = 10'h144 == _T_378[9:0] ? 4'h3 : _GEN_18956; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18958 = 10'h145 == _T_378[9:0] ? 4'h3 : _GEN_18957; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18959 = 10'h146 == _T_378[9:0] ? 4'h9 : _GEN_18958; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18960 = 10'h147 == _T_378[9:0] ? 4'hf : _GEN_18959; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18961 = 10'h148 == _T_378[9:0] ? 4'h3 : _GEN_18960; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18962 = 10'h149 == _T_378[9:0] ? 4'h3 : _GEN_18961; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18963 = 10'h14a == _T_378[9:0] ? 4'h3 : _GEN_18962; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18964 = 10'h14b == _T_378[9:0] ? 4'h3 : _GEN_18963; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18965 = 10'h14c == _T_378[9:0] ? 4'h3 : _GEN_18964; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18966 = 10'h14d == _T_378[9:0] ? 4'h3 : _GEN_18965; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18967 = 10'h14e == _T_378[9:0] ? 4'h3 : _GEN_18966; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18968 = 10'h14f == _T_378[9:0] ? 4'h3 : _GEN_18967; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18969 = 10'h150 == _T_378[9:0] ? 4'h3 : _GEN_18968; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18970 = 10'h151 == _T_378[9:0] ? 4'h3 : _GEN_18969; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18971 = 10'h152 == _T_378[9:0] ? 4'h3 : _GEN_18970; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18972 = 10'h153 == _T_378[9:0] ? 4'h3 : _GEN_18971; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18973 = 10'h154 == _T_378[9:0] ? 4'h3 : _GEN_18972; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18974 = 10'h155 == _T_378[9:0] ? 4'h3 : _GEN_18973; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18975 = 10'h156 == _T_378[9:0] ? 4'h3 : _GEN_18974; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18976 = 10'h157 == _T_378[9:0] ? 4'hf : _GEN_18975; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18977 = 10'h158 == _T_378[9:0] ? 4'h3 : _GEN_18976; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18978 = 10'h159 == _T_378[9:0] ? 4'h3 : _GEN_18977; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18979 = 10'h15a == _T_378[9:0] ? 4'h3 : _GEN_18978; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18980 = 10'h15b == _T_378[9:0] ? 4'h3 : _GEN_18979; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18981 = 10'h15c == _T_378[9:0] ? 4'h3 : _GEN_18980; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18982 = 10'h15d == _T_378[9:0] ? 4'h3 : _GEN_18981; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18983 = 10'h15e == _T_378[9:0] ? 4'h2 : _GEN_18982; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18984 = 10'h15f == _T_378[9:0] ? 4'h0 : _GEN_18983; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18985 = 10'h160 == _T_378[9:0] ? 4'h3 : _GEN_18984; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18986 = 10'h161 == _T_378[9:0] ? 4'h3 : _GEN_18985; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18987 = 10'h162 == _T_378[9:0] ? 4'h3 : _GEN_18986; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18988 = 10'h163 == _T_378[9:0] ? 4'h2 : _GEN_18987; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18989 = 10'h164 == _T_378[9:0] ? 4'h3 : _GEN_18988; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18990 = 10'h165 == _T_378[9:0] ? 4'h9 : _GEN_18989; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18991 = 10'h166 == _T_378[9:0] ? 4'hf : _GEN_18990; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18992 = 10'h167 == _T_378[9:0] ? 4'hf : _GEN_18991; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18993 = 10'h168 == _T_378[9:0] ? 4'hd : _GEN_18992; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18994 = 10'h169 == _T_378[9:0] ? 4'h9 : _GEN_18993; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18995 = 10'h16a == _T_378[9:0] ? 4'hd : _GEN_18994; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18996 = 10'h16b == _T_378[9:0] ? 4'hd : _GEN_18995; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18997 = 10'h16c == _T_378[9:0] ? 4'h3 : _GEN_18996; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18998 = 10'h16d == _T_378[9:0] ? 4'h3 : _GEN_18997; // @[Filter.scala 191:142]
  wire [3:0] _GEN_18999 = 10'h16e == _T_378[9:0] ? 4'h3 : _GEN_18998; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19000 = 10'h16f == _T_378[9:0] ? 4'h3 : _GEN_18999; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19001 = 10'h170 == _T_378[9:0] ? 4'h3 : _GEN_19000; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19002 = 10'h171 == _T_378[9:0] ? 4'h3 : _GEN_19001; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19003 = 10'h172 == _T_378[9:0] ? 4'h3 : _GEN_19002; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19004 = 10'h173 == _T_378[9:0] ? 4'h3 : _GEN_19003; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19005 = 10'h174 == _T_378[9:0] ? 4'h3 : _GEN_19004; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19006 = 10'h175 == _T_378[9:0] ? 4'h3 : _GEN_19005; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19007 = 10'h176 == _T_378[9:0] ? 4'hf : _GEN_19006; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19008 = 10'h177 == _T_378[9:0] ? 4'hf : _GEN_19007; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19009 = 10'h178 == _T_378[9:0] ? 4'h9 : _GEN_19008; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19010 = 10'h179 == _T_378[9:0] ? 4'h3 : _GEN_19009; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19011 = 10'h17a == _T_378[9:0] ? 4'h3 : _GEN_19010; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19012 = 10'h17b == _T_378[9:0] ? 4'h3 : _GEN_19011; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19013 = 10'h17c == _T_378[9:0] ? 4'h3 : _GEN_19012; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19014 = 10'h17d == _T_378[9:0] ? 4'h2 : _GEN_19013; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19015 = 10'h17e == _T_378[9:0] ? 4'h3 : _GEN_19014; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19016 = 10'h17f == _T_378[9:0] ? 4'h0 : _GEN_19015; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19017 = 10'h180 == _T_378[9:0] ? 4'hd : _GEN_19016; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19018 = 10'h181 == _T_378[9:0] ? 4'hd : _GEN_19017; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19019 = 10'h182 == _T_378[9:0] ? 4'hd : _GEN_19018; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19020 = 10'h183 == _T_378[9:0] ? 4'hd : _GEN_19019; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19021 = 10'h184 == _T_378[9:0] ? 4'h3 : _GEN_19020; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19022 = 10'h185 == _T_378[9:0] ? 4'h9 : _GEN_19021; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19023 = 10'h186 == _T_378[9:0] ? 4'hb : _GEN_19022; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19024 = 10'h187 == _T_378[9:0] ? 4'hf : _GEN_19023; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19025 = 10'h188 == _T_378[9:0] ? 4'hd : _GEN_19024; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19026 = 10'h189 == _T_378[9:0] ? 4'hd : _GEN_19025; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19027 = 10'h18a == _T_378[9:0] ? 4'hd : _GEN_19026; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19028 = 10'h18b == _T_378[9:0] ? 4'hd : _GEN_19027; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19029 = 10'h18c == _T_378[9:0] ? 4'hd : _GEN_19028; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19030 = 10'h18d == _T_378[9:0] ? 4'hd : _GEN_19029; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19031 = 10'h18e == _T_378[9:0] ? 4'hd : _GEN_19030; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19032 = 10'h18f == _T_378[9:0] ? 4'hd : _GEN_19031; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19033 = 10'h190 == _T_378[9:0] ? 4'hd : _GEN_19032; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19034 = 10'h191 == _T_378[9:0] ? 4'hd : _GEN_19033; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19035 = 10'h192 == _T_378[9:0] ? 4'h9 : _GEN_19034; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19036 = 10'h193 == _T_378[9:0] ? 4'hd : _GEN_19035; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19037 = 10'h194 == _T_378[9:0] ? 4'hd : _GEN_19036; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19038 = 10'h195 == _T_378[9:0] ? 4'hd : _GEN_19037; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19039 = 10'h196 == _T_378[9:0] ? 4'hf : _GEN_19038; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19040 = 10'h197 == _T_378[9:0] ? 4'h3 : _GEN_19039; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19041 = 10'h198 == _T_378[9:0] ? 4'h9 : _GEN_19040; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19042 = 10'h199 == _T_378[9:0] ? 4'h3 : _GEN_19041; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19043 = 10'h19a == _T_378[9:0] ? 4'h3 : _GEN_19042; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19044 = 10'h19b == _T_378[9:0] ? 4'h3 : _GEN_19043; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19045 = 10'h19c == _T_378[9:0] ? 4'h3 : _GEN_19044; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19046 = 10'h19d == _T_378[9:0] ? 4'h3 : _GEN_19045; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19047 = 10'h19e == _T_378[9:0] ? 4'h3 : _GEN_19046; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19048 = 10'h19f == _T_378[9:0] ? 4'h0 : _GEN_19047; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19049 = 10'h1a0 == _T_378[9:0] ? 4'hd : _GEN_19048; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19050 = 10'h1a1 == _T_378[9:0] ? 4'hd : _GEN_19049; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19051 = 10'h1a2 == _T_378[9:0] ? 4'h9 : _GEN_19050; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19052 = 10'h1a3 == _T_378[9:0] ? 4'hd : _GEN_19051; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19053 = 10'h1a4 == _T_378[9:0] ? 4'h3 : _GEN_19052; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19054 = 10'h1a5 == _T_378[9:0] ? 4'hf : _GEN_19053; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19055 = 10'h1a6 == _T_378[9:0] ? 4'hd : _GEN_19054; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19056 = 10'h1a7 == _T_378[9:0] ? 4'hf : _GEN_19055; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19057 = 10'h1a8 == _T_378[9:0] ? 4'hb : _GEN_19056; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19058 = 10'h1a9 == _T_378[9:0] ? 4'hd : _GEN_19057; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19059 = 10'h1aa == _T_378[9:0] ? 4'hd : _GEN_19058; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19060 = 10'h1ab == _T_378[9:0] ? 4'h9 : _GEN_19059; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19061 = 10'h1ac == _T_378[9:0] ? 4'hd : _GEN_19060; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19062 = 10'h1ad == _T_378[9:0] ? 4'hd : _GEN_19061; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19063 = 10'h1ae == _T_378[9:0] ? 4'hd : _GEN_19062; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19064 = 10'h1af == _T_378[9:0] ? 4'hd : _GEN_19063; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19065 = 10'h1b0 == _T_378[9:0] ? 4'hd : _GEN_19064; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19066 = 10'h1b1 == _T_378[9:0] ? 4'hd : _GEN_19065; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19067 = 10'h1b2 == _T_378[9:0] ? 4'hd : _GEN_19066; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19068 = 10'h1b3 == _T_378[9:0] ? 4'hd : _GEN_19067; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19069 = 10'h1b4 == _T_378[9:0] ? 4'hd : _GEN_19068; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19070 = 10'h1b5 == _T_378[9:0] ? 4'hd : _GEN_19069; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19071 = 10'h1b6 == _T_378[9:0] ? 4'hf : _GEN_19070; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19072 = 10'h1b7 == _T_378[9:0] ? 4'hd : _GEN_19071; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19073 = 10'h1b8 == _T_378[9:0] ? 4'hf : _GEN_19072; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19074 = 10'h1b9 == _T_378[9:0] ? 4'hd : _GEN_19073; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19075 = 10'h1ba == _T_378[9:0] ? 4'hd : _GEN_19074; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19076 = 10'h1bb == _T_378[9:0] ? 4'hd : _GEN_19075; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19077 = 10'h1bc == _T_378[9:0] ? 4'h2 : _GEN_19076; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19078 = 10'h1bd == _T_378[9:0] ? 4'h3 : _GEN_19077; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19079 = 10'h1be == _T_378[9:0] ? 4'hd : _GEN_19078; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19080 = 10'h1bf == _T_378[9:0] ? 4'h0 : _GEN_19079; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19081 = 10'h1c0 == _T_378[9:0] ? 4'hd : _GEN_19080; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19082 = 10'h1c1 == _T_378[9:0] ? 4'hd : _GEN_19081; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19083 = 10'h1c2 == _T_378[9:0] ? 4'hd : _GEN_19082; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19084 = 10'h1c3 == _T_378[9:0] ? 4'h2 : _GEN_19083; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19085 = 10'h1c4 == _T_378[9:0] ? 4'h2 : _GEN_19084; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19086 = 10'h1c5 == _T_378[9:0] ? 4'hd : _GEN_19085; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19087 = 10'h1c6 == _T_378[9:0] ? 4'hd : _GEN_19086; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19088 = 10'h1c7 == _T_378[9:0] ? 4'hd : _GEN_19087; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19089 = 10'h1c8 == _T_378[9:0] ? 4'hd : _GEN_19088; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19090 = 10'h1c9 == _T_378[9:0] ? 4'hb : _GEN_19089; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19091 = 10'h1ca == _T_378[9:0] ? 4'hb : _GEN_19090; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19092 = 10'h1cb == _T_378[9:0] ? 4'hb : _GEN_19091; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19093 = 10'h1cc == _T_378[9:0] ? 4'hb : _GEN_19092; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19094 = 10'h1cd == _T_378[9:0] ? 4'hb : _GEN_19093; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19095 = 10'h1ce == _T_378[9:0] ? 4'hb : _GEN_19094; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19096 = 10'h1cf == _T_378[9:0] ? 4'hb : _GEN_19095; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19097 = 10'h1d0 == _T_378[9:0] ? 4'hb : _GEN_19096; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19098 = 10'h1d1 == _T_378[9:0] ? 4'hb : _GEN_19097; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19099 = 10'h1d2 == _T_378[9:0] ? 4'hb : _GEN_19098; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19100 = 10'h1d3 == _T_378[9:0] ? 4'hb : _GEN_19099; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19101 = 10'h1d4 == _T_378[9:0] ? 4'hb : _GEN_19100; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19102 = 10'h1d5 == _T_378[9:0] ? 4'hb : _GEN_19101; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19103 = 10'h1d6 == _T_378[9:0] ? 4'hd : _GEN_19102; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19104 = 10'h1d7 == _T_378[9:0] ? 4'hd : _GEN_19103; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19105 = 10'h1d8 == _T_378[9:0] ? 4'hd : _GEN_19104; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19106 = 10'h1d9 == _T_378[9:0] ? 4'hd : _GEN_19105; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19107 = 10'h1da == _T_378[9:0] ? 4'hd : _GEN_19106; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19108 = 10'h1db == _T_378[9:0] ? 4'hd : _GEN_19107; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19109 = 10'h1dc == _T_378[9:0] ? 4'hd : _GEN_19108; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19110 = 10'h1dd == _T_378[9:0] ? 4'h3 : _GEN_19109; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19111 = 10'h1de == _T_378[9:0] ? 4'hd : _GEN_19110; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19112 = 10'h1df == _T_378[9:0] ? 4'h0 : _GEN_19111; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19113 = 10'h1e0 == _T_378[9:0] ? 4'h9 : _GEN_19112; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19114 = 10'h1e1 == _T_378[9:0] ? 4'hd : _GEN_19113; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19115 = 10'h1e2 == _T_378[9:0] ? 4'h2 : _GEN_19114; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19116 = 10'h1e3 == _T_378[9:0] ? 4'h2 : _GEN_19115; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19117 = 10'h1e4 == _T_378[9:0] ? 4'hd : _GEN_19116; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19118 = 10'h1e5 == _T_378[9:0] ? 4'hd : _GEN_19117; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19119 = 10'h1e6 == _T_378[9:0] ? 4'hd : _GEN_19118; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19120 = 10'h1e7 == _T_378[9:0] ? 4'hd : _GEN_19119; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19121 = 10'h1e8 == _T_378[9:0] ? 4'hb : _GEN_19120; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19122 = 10'h1e9 == _T_378[9:0] ? 4'hd : _GEN_19121; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19123 = 10'h1ea == _T_378[9:0] ? 4'hd : _GEN_19122; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19124 = 10'h1eb == _T_378[9:0] ? 4'hb : _GEN_19123; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19125 = 10'h1ec == _T_378[9:0] ? 4'hd : _GEN_19124; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19126 = 10'h1ed == _T_378[9:0] ? 4'hb : _GEN_19125; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19127 = 10'h1ee == _T_378[9:0] ? 4'hd : _GEN_19126; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19128 = 10'h1ef == _T_378[9:0] ? 4'hb : _GEN_19127; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19129 = 10'h1f0 == _T_378[9:0] ? 4'hd : _GEN_19128; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19130 = 10'h1f1 == _T_378[9:0] ? 4'hb : _GEN_19129; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19131 = 10'h1f2 == _T_378[9:0] ? 4'hb : _GEN_19130; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19132 = 10'h1f3 == _T_378[9:0] ? 4'hd : _GEN_19131; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19133 = 10'h1f4 == _T_378[9:0] ? 4'hb : _GEN_19132; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19134 = 10'h1f5 == _T_378[9:0] ? 4'hb : _GEN_19133; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19135 = 10'h1f6 == _T_378[9:0] ? 4'hd : _GEN_19134; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19136 = 10'h1f7 == _T_378[9:0] ? 4'hd : _GEN_19135; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19137 = 10'h1f8 == _T_378[9:0] ? 4'hd : _GEN_19136; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19138 = 10'h1f9 == _T_378[9:0] ? 4'hd : _GEN_19137; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19139 = 10'h1fa == _T_378[9:0] ? 4'h9 : _GEN_19138; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19140 = 10'h1fb == _T_378[9:0] ? 4'hd : _GEN_19139; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19141 = 10'h1fc == _T_378[9:0] ? 4'hd : _GEN_19140; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19142 = 10'h1fd == _T_378[9:0] ? 4'h2 : _GEN_19141; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19143 = 10'h1fe == _T_378[9:0] ? 4'hd : _GEN_19142; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19144 = 10'h1ff == _T_378[9:0] ? 4'h0 : _GEN_19143; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19145 = 10'h200 == _T_378[9:0] ? 4'hd : _GEN_19144; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19146 = 10'h201 == _T_378[9:0] ? 4'hd : _GEN_19145; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19147 = 10'h202 == _T_378[9:0] ? 4'h3 : _GEN_19146; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19148 = 10'h203 == _T_378[9:0] ? 4'hd : _GEN_19147; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19149 = 10'h204 == _T_378[9:0] ? 4'hd : _GEN_19148; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19150 = 10'h205 == _T_378[9:0] ? 4'hd : _GEN_19149; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19151 = 10'h206 == _T_378[9:0] ? 4'hb : _GEN_19150; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19152 = 10'h207 == _T_378[9:0] ? 4'hb : _GEN_19151; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19153 = 10'h208 == _T_378[9:0] ? 4'hd : _GEN_19152; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19154 = 10'h209 == _T_378[9:0] ? 4'hd : _GEN_19153; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19155 = 10'h20a == _T_378[9:0] ? 4'hd : _GEN_19154; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19156 = 10'h20b == _T_378[9:0] ? 4'hb : _GEN_19155; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19157 = 10'h20c == _T_378[9:0] ? 4'hd : _GEN_19156; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19158 = 10'h20d == _T_378[9:0] ? 4'hb : _GEN_19157; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19159 = 10'h20e == _T_378[9:0] ? 4'hd : _GEN_19158; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19160 = 10'h20f == _T_378[9:0] ? 4'hb : _GEN_19159; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19161 = 10'h210 == _T_378[9:0] ? 4'hd : _GEN_19160; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19162 = 10'h211 == _T_378[9:0] ? 4'hd : _GEN_19161; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19163 = 10'h212 == _T_378[9:0] ? 4'hb : _GEN_19162; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19164 = 10'h213 == _T_378[9:0] ? 4'hb : _GEN_19163; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19165 = 10'h214 == _T_378[9:0] ? 4'hb : _GEN_19164; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19166 = 10'h215 == _T_378[9:0] ? 4'hd : _GEN_19165; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19167 = 10'h216 == _T_378[9:0] ? 4'hd : _GEN_19166; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19168 = 10'h217 == _T_378[9:0] ? 4'hd : _GEN_19167; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19169 = 10'h218 == _T_378[9:0] ? 4'hd : _GEN_19168; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19170 = 10'h219 == _T_378[9:0] ? 4'hd : _GEN_19169; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19171 = 10'h21a == _T_378[9:0] ? 4'hd : _GEN_19170; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19172 = 10'h21b == _T_378[9:0] ? 4'hd : _GEN_19171; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19173 = 10'h21c == _T_378[9:0] ? 4'h3 : _GEN_19172; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19174 = 10'h21d == _T_378[9:0] ? 4'h2 : _GEN_19173; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19175 = 10'h21e == _T_378[9:0] ? 4'hd : _GEN_19174; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19176 = 10'h21f == _T_378[9:0] ? 4'h0 : _GEN_19175; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19177 = 10'h220 == _T_378[9:0] ? 4'h0 : _GEN_19176; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19178 = 10'h221 == _T_378[9:0] ? 4'h0 : _GEN_19177; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19179 = 10'h222 == _T_378[9:0] ? 4'h0 : _GEN_19178; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19180 = 10'h223 == _T_378[9:0] ? 4'h0 : _GEN_19179; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19181 = 10'h224 == _T_378[9:0] ? 4'h0 : _GEN_19180; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19182 = 10'h225 == _T_378[9:0] ? 4'h0 : _GEN_19181; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19183 = 10'h226 == _T_378[9:0] ? 4'h0 : _GEN_19182; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19184 = 10'h227 == _T_378[9:0] ? 4'h0 : _GEN_19183; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19185 = 10'h228 == _T_378[9:0] ? 4'h0 : _GEN_19184; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19186 = 10'h229 == _T_378[9:0] ? 4'h0 : _GEN_19185; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19187 = 10'h22a == _T_378[9:0] ? 4'h0 : _GEN_19186; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19188 = 10'h22b == _T_378[9:0] ? 4'h0 : _GEN_19187; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19189 = 10'h22c == _T_378[9:0] ? 4'h0 : _GEN_19188; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19190 = 10'h22d == _T_378[9:0] ? 4'h0 : _GEN_19189; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19191 = 10'h22e == _T_378[9:0] ? 4'h0 : _GEN_19190; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19192 = 10'h22f == _T_378[9:0] ? 4'h0 : _GEN_19191; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19193 = 10'h230 == _T_378[9:0] ? 4'h0 : _GEN_19192; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19194 = 10'h231 == _T_378[9:0] ? 4'h0 : _GEN_19193; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19195 = 10'h232 == _T_378[9:0] ? 4'h0 : _GEN_19194; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19196 = 10'h233 == _T_378[9:0] ? 4'h0 : _GEN_19195; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19197 = 10'h234 == _T_378[9:0] ? 4'h0 : _GEN_19196; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19198 = 10'h235 == _T_378[9:0] ? 4'h0 : _GEN_19197; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19199 = 10'h236 == _T_378[9:0] ? 4'h0 : _GEN_19198; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19200 = 10'h237 == _T_378[9:0] ? 4'h0 : _GEN_19199; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19201 = 10'h238 == _T_378[9:0] ? 4'h0 : _GEN_19200; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19202 = 10'h239 == _T_378[9:0] ? 4'h0 : _GEN_19201; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19203 = 10'h23a == _T_378[9:0] ? 4'h0 : _GEN_19202; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19204 = 10'h23b == _T_378[9:0] ? 4'h0 : _GEN_19203; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19205 = 10'h23c == _T_378[9:0] ? 4'h0 : _GEN_19204; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19206 = 10'h23d == _T_378[9:0] ? 4'h0 : _GEN_19205; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19207 = 10'h23e == _T_378[9:0] ? 4'h0 : _GEN_19206; // @[Filter.scala 191:142]
  wire [3:0] _GEN_19208 = 10'h23f == _T_378[9:0] ? 4'h0 : _GEN_19207; // @[Filter.scala 191:142]
  wire [7:0] _T_392 = _GEN_19208 * 4'ha; // @[Filter.scala 191:142]
  wire [10:0] _GEN_28363 = {{3'd0}, _T_392}; // @[Filter.scala 191:109]
  wire [10:0] _T_394 = _T_387 + _GEN_28363; // @[Filter.scala 191:109]
  wire [10:0] _T_395 = _T_394 / 11'h64; // @[Filter.scala 191:150]
  wire  _T_397 = _T_368 >= 6'h20; // @[Filter.scala 194:31]
  wire  _T_401 = _T_375 >= 32'h12; // @[Filter.scala 194:63]
  wire  _T_402 = _T_397 | _T_401; // @[Filter.scala 194:58]
  wire [10:0] _GEN_19785 = io_SPI_distort ? _T_395 : {{7'd0}, _GEN_18056}; // @[Filter.scala 196:35]
  wire [10:0] _GEN_19786 = _T_402 ? 11'h0 : _GEN_19785; // @[Filter.scala 194:80]
  wire [10:0] _GEN_20363 = io_SPI_distort ? _T_395 : {{7'd0}, _GEN_18632}; // @[Filter.scala 196:35]
  wire [10:0] _GEN_20364 = _T_402 ? 11'h0 : _GEN_20363; // @[Filter.scala 194:80]
  wire [10:0] _GEN_20941 = io_SPI_distort ? _T_395 : {{7'd0}, _GEN_19208}; // @[Filter.scala 196:35]
  wire [10:0] _GEN_20942 = _T_402 ? 11'h0 : _GEN_20941; // @[Filter.scala 194:80]
  wire [31:0] _T_430 = pixelIndex + 32'h6; // @[Filter.scala 189:31]
  wire [31:0] _GEN_6 = _T_430 % 32'h20; // @[Filter.scala 189:38]
  wire [5:0] _T_431 = _GEN_6[5:0]; // @[Filter.scala 189:38]
  wire [5:0] _T_433 = _T_431 + _GEN_28295; // @[Filter.scala 189:53]
  wire [5:0] _T_435 = _T_433 - 6'h1; // @[Filter.scala 189:69]
  wire [31:0] _T_438 = _T_430 / 32'h20; // @[Filter.scala 190:38]
  wire [31:0] _T_440 = _T_438 + _GEN_28296; // @[Filter.scala 190:53]
  wire [31:0] _T_442 = _T_440 - 32'h1; // @[Filter.scala 190:69]
  wire [37:0] _T_443 = _T_442 * 32'h20; // @[Filter.scala 191:42]
  wire [37:0] _GEN_28369 = {{32'd0}, _T_435}; // @[Filter.scala 191:57]
  wire [37:0] _T_445 = _T_443 + _GEN_28369; // @[Filter.scala 191:57]
  wire [3:0] _GEN_20946 = 10'h3 == _T_445[9:0] ? 4'h3 : 4'ha; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20947 = 10'h4 == _T_445[9:0] ? 4'ha : _GEN_20946; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20948 = 10'h5 == _T_445[9:0] ? 4'ha : _GEN_20947; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20949 = 10'h6 == _T_445[9:0] ? 4'ha : _GEN_20948; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20950 = 10'h7 == _T_445[9:0] ? 4'ha : _GEN_20949; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20951 = 10'h8 == _T_445[9:0] ? 4'ha : _GEN_20950; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20952 = 10'h9 == _T_445[9:0] ? 4'ha : _GEN_20951; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20953 = 10'ha == _T_445[9:0] ? 4'ha : _GEN_20952; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20954 = 10'hb == _T_445[9:0] ? 4'ha : _GEN_20953; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20955 = 10'hc == _T_445[9:0] ? 4'ha : _GEN_20954; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20956 = 10'hd == _T_445[9:0] ? 4'ha : _GEN_20955; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20957 = 10'he == _T_445[9:0] ? 4'ha : _GEN_20956; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20958 = 10'hf == _T_445[9:0] ? 4'ha : _GEN_20957; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20959 = 10'h10 == _T_445[9:0] ? 4'ha : _GEN_20958; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20960 = 10'h11 == _T_445[9:0] ? 4'ha : _GEN_20959; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20961 = 10'h12 == _T_445[9:0] ? 4'ha : _GEN_20960; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20962 = 10'h13 == _T_445[9:0] ? 4'ha : _GEN_20961; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20963 = 10'h14 == _T_445[9:0] ? 4'ha : _GEN_20962; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20964 = 10'h15 == _T_445[9:0] ? 4'ha : _GEN_20963; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20965 = 10'h16 == _T_445[9:0] ? 4'ha : _GEN_20964; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20966 = 10'h17 == _T_445[9:0] ? 4'ha : _GEN_20965; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20967 = 10'h18 == _T_445[9:0] ? 4'ha : _GEN_20966; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20968 = 10'h19 == _T_445[9:0] ? 4'ha : _GEN_20967; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20969 = 10'h1a == _T_445[9:0] ? 4'ha : _GEN_20968; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20970 = 10'h1b == _T_445[9:0] ? 4'ha : _GEN_20969; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20971 = 10'h1c == _T_445[9:0] ? 4'ha : _GEN_20970; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20972 = 10'h1d == _T_445[9:0] ? 4'ha : _GEN_20971; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20973 = 10'h1e == _T_445[9:0] ? 4'ha : _GEN_20972; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20974 = 10'h1f == _T_445[9:0] ? 4'h0 : _GEN_20973; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20975 = 10'h20 == _T_445[9:0] ? 4'ha : _GEN_20974; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20976 = 10'h21 == _T_445[9:0] ? 4'ha : _GEN_20975; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20977 = 10'h22 == _T_445[9:0] ? 4'ha : _GEN_20976; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20978 = 10'h23 == _T_445[9:0] ? 4'h3 : _GEN_20977; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20979 = 10'h24 == _T_445[9:0] ? 4'ha : _GEN_20978; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20980 = 10'h25 == _T_445[9:0] ? 4'ha : _GEN_20979; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20981 = 10'h26 == _T_445[9:0] ? 4'ha : _GEN_20980; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20982 = 10'h27 == _T_445[9:0] ? 4'h1 : _GEN_20981; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20983 = 10'h28 == _T_445[9:0] ? 4'h1 : _GEN_20982; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20984 = 10'h29 == _T_445[9:0] ? 4'ha : _GEN_20983; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20985 = 10'h2a == _T_445[9:0] ? 4'ha : _GEN_20984; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20986 = 10'h2b == _T_445[9:0] ? 4'ha : _GEN_20985; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20987 = 10'h2c == _T_445[9:0] ? 4'ha : _GEN_20986; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20988 = 10'h2d == _T_445[9:0] ? 4'ha : _GEN_20987; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20989 = 10'h2e == _T_445[9:0] ? 4'ha : _GEN_20988; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20990 = 10'h2f == _T_445[9:0] ? 4'ha : _GEN_20989; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20991 = 10'h30 == _T_445[9:0] ? 4'ha : _GEN_20990; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20992 = 10'h31 == _T_445[9:0] ? 4'ha : _GEN_20991; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20993 = 10'h32 == _T_445[9:0] ? 4'ha : _GEN_20992; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20994 = 10'h33 == _T_445[9:0] ? 4'ha : _GEN_20993; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20995 = 10'h34 == _T_445[9:0] ? 4'ha : _GEN_20994; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20996 = 10'h35 == _T_445[9:0] ? 4'ha : _GEN_20995; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20997 = 10'h36 == _T_445[9:0] ? 4'ha : _GEN_20996; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20998 = 10'h37 == _T_445[9:0] ? 4'h1 : _GEN_20997; // @[Filter.scala 191:62]
  wire [3:0] _GEN_20999 = 10'h38 == _T_445[9:0] ? 4'h1 : _GEN_20998; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21000 = 10'h39 == _T_445[9:0] ? 4'ha : _GEN_20999; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21001 = 10'h3a == _T_445[9:0] ? 4'ha : _GEN_21000; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21002 = 10'h3b == _T_445[9:0] ? 4'ha : _GEN_21001; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21003 = 10'h3c == _T_445[9:0] ? 4'ha : _GEN_21002; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21004 = 10'h3d == _T_445[9:0] ? 4'h3 : _GEN_21003; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21005 = 10'h3e == _T_445[9:0] ? 4'ha : _GEN_21004; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21006 = 10'h3f == _T_445[9:0] ? 4'h0 : _GEN_21005; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21007 = 10'h40 == _T_445[9:0] ? 4'ha : _GEN_21006; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21008 = 10'h41 == _T_445[9:0] ? 4'ha : _GEN_21007; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21009 = 10'h42 == _T_445[9:0] ? 4'ha : _GEN_21008; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21010 = 10'h43 == _T_445[9:0] ? 4'h2 : _GEN_21009; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21011 = 10'h44 == _T_445[9:0] ? 4'h3 : _GEN_21010; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21012 = 10'h45 == _T_445[9:0] ? 4'h0 : _GEN_21011; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21013 = 10'h46 == _T_445[9:0] ? 4'h0 : _GEN_21012; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21014 = 10'h47 == _T_445[9:0] ? 4'h0 : _GEN_21013; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21015 = 10'h48 == _T_445[9:0] ? 4'h0 : _GEN_21014; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21016 = 10'h49 == _T_445[9:0] ? 4'ha : _GEN_21015; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21017 = 10'h4a == _T_445[9:0] ? 4'ha : _GEN_21016; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21018 = 10'h4b == _T_445[9:0] ? 4'ha : _GEN_21017; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21019 = 10'h4c == _T_445[9:0] ? 4'ha : _GEN_21018; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21020 = 10'h4d == _T_445[9:0] ? 4'ha : _GEN_21019; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21021 = 10'h4e == _T_445[9:0] ? 4'ha : _GEN_21020; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21022 = 10'h4f == _T_445[9:0] ? 4'ha : _GEN_21021; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21023 = 10'h50 == _T_445[9:0] ? 4'ha : _GEN_21022; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21024 = 10'h51 == _T_445[9:0] ? 4'ha : _GEN_21023; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21025 = 10'h52 == _T_445[9:0] ? 4'ha : _GEN_21024; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21026 = 10'h53 == _T_445[9:0] ? 4'ha : _GEN_21025; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21027 = 10'h54 == _T_445[9:0] ? 4'h1 : _GEN_21026; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21028 = 10'h55 == _T_445[9:0] ? 4'h1 : _GEN_21027; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21029 = 10'h56 == _T_445[9:0] ? 4'h1 : _GEN_21028; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21030 = 10'h57 == _T_445[9:0] ? 4'h0 : _GEN_21029; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21031 = 10'h58 == _T_445[9:0] ? 4'ha : _GEN_21030; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21032 = 10'h59 == _T_445[9:0] ? 4'h0 : _GEN_21031; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21033 = 10'h5a == _T_445[9:0] ? 4'ha : _GEN_21032; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21034 = 10'h5b == _T_445[9:0] ? 4'ha : _GEN_21033; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21035 = 10'h5c == _T_445[9:0] ? 4'ha : _GEN_21034; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21036 = 10'h5d == _T_445[9:0] ? 4'h3 : _GEN_21035; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21037 = 10'h5e == _T_445[9:0] ? 4'ha : _GEN_21036; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21038 = 10'h5f == _T_445[9:0] ? 4'h0 : _GEN_21037; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21039 = 10'h60 == _T_445[9:0] ? 4'ha : _GEN_21038; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21040 = 10'h61 == _T_445[9:0] ? 4'ha : _GEN_21039; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21041 = 10'h62 == _T_445[9:0] ? 4'ha : _GEN_21040; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21042 = 10'h63 == _T_445[9:0] ? 4'ha : _GEN_21041; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21043 = 10'h64 == _T_445[9:0] ? 4'h3 : _GEN_21042; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21044 = 10'h65 == _T_445[9:0] ? 4'h0 : _GEN_21043; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21045 = 10'h66 == _T_445[9:0] ? 4'ha : _GEN_21044; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21046 = 10'h67 == _T_445[9:0] ? 4'ha : _GEN_21045; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21047 = 10'h68 == _T_445[9:0] ? 4'ha : _GEN_21046; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21048 = 10'h69 == _T_445[9:0] ? 4'h0 : _GEN_21047; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21049 = 10'h6a == _T_445[9:0] ? 4'h1 : _GEN_21048; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21050 = 10'h6b == _T_445[9:0] ? 4'h1 : _GEN_21049; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21051 = 10'h6c == _T_445[9:0] ? 4'ha : _GEN_21050; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21052 = 10'h6d == _T_445[9:0] ? 4'ha : _GEN_21051; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21053 = 10'h6e == _T_445[9:0] ? 4'ha : _GEN_21052; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21054 = 10'h6f == _T_445[9:0] ? 4'ha : _GEN_21053; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21055 = 10'h70 == _T_445[9:0] ? 4'ha : _GEN_21054; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21056 = 10'h71 == _T_445[9:0] ? 4'ha : _GEN_21055; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21057 = 10'h72 == _T_445[9:0] ? 4'ha : _GEN_21056; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21058 = 10'h73 == _T_445[9:0] ? 4'h1 : _GEN_21057; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21059 = 10'h74 == _T_445[9:0] ? 4'h0 : _GEN_21058; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21060 = 10'h75 == _T_445[9:0] ? 4'h0 : _GEN_21059; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21061 = 10'h76 == _T_445[9:0] ? 4'h0 : _GEN_21060; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21062 = 10'h77 == _T_445[9:0] ? 4'ha : _GEN_21061; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21063 = 10'h78 == _T_445[9:0] ? 4'ha : _GEN_21062; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21064 = 10'h79 == _T_445[9:0] ? 4'ha : _GEN_21063; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21065 = 10'h7a == _T_445[9:0] ? 4'h0 : _GEN_21064; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21066 = 10'h7b == _T_445[9:0] ? 4'ha : _GEN_21065; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21067 = 10'h7c == _T_445[9:0] ? 4'ha : _GEN_21066; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21068 = 10'h7d == _T_445[9:0] ? 4'h2 : _GEN_21067; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21069 = 10'h7e == _T_445[9:0] ? 4'h3 : _GEN_21068; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21070 = 10'h7f == _T_445[9:0] ? 4'h0 : _GEN_21069; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21071 = 10'h80 == _T_445[9:0] ? 4'ha : _GEN_21070; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21072 = 10'h81 == _T_445[9:0] ? 4'ha : _GEN_21071; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21073 = 10'h82 == _T_445[9:0] ? 4'h1 : _GEN_21072; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21074 = 10'h83 == _T_445[9:0] ? 4'h0 : _GEN_21073; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21075 = 10'h84 == _T_445[9:0] ? 4'h2 : _GEN_21074; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21076 = 10'h85 == _T_445[9:0] ? 4'h1 : _GEN_21075; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21077 = 10'h86 == _T_445[9:0] ? 4'h1 : _GEN_21076; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21078 = 10'h87 == _T_445[9:0] ? 4'ha : _GEN_21077; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21079 = 10'h88 == _T_445[9:0] ? 4'ha : _GEN_21078; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21080 = 10'h89 == _T_445[9:0] ? 4'h0 : _GEN_21079; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21081 = 10'h8a == _T_445[9:0] ? 4'h0 : _GEN_21080; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21082 = 10'h8b == _T_445[9:0] ? 4'h1 : _GEN_21081; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21083 = 10'h8c == _T_445[9:0] ? 4'h1 : _GEN_21082; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21084 = 10'h8d == _T_445[9:0] ? 4'h1 : _GEN_21083; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21085 = 10'h8e == _T_445[9:0] ? 4'h1 : _GEN_21084; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21086 = 10'h8f == _T_445[9:0] ? 4'h1 : _GEN_21085; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21087 = 10'h90 == _T_445[9:0] ? 4'h1 : _GEN_21086; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21088 = 10'h91 == _T_445[9:0] ? 4'h1 : _GEN_21087; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21089 = 10'h92 == _T_445[9:0] ? 4'h1 : _GEN_21088; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21090 = 10'h93 == _T_445[9:0] ? 4'h0 : _GEN_21089; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21091 = 10'h94 == _T_445[9:0] ? 4'h0 : _GEN_21090; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21092 = 10'h95 == _T_445[9:0] ? 4'ha : _GEN_21091; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21093 = 10'h96 == _T_445[9:0] ? 4'ha : _GEN_21092; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21094 = 10'h97 == _T_445[9:0] ? 4'ha : _GEN_21093; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21095 = 10'h98 == _T_445[9:0] ? 4'h1 : _GEN_21094; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21096 = 10'h99 == _T_445[9:0] ? 4'h0 : _GEN_21095; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21097 = 10'h9a == _T_445[9:0] ? 4'h1 : _GEN_21096; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21098 = 10'h9b == _T_445[9:0] ? 4'h1 : _GEN_21097; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21099 = 10'h9c == _T_445[9:0] ? 4'ha : _GEN_21098; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21100 = 10'h9d == _T_445[9:0] ? 4'ha : _GEN_21099; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21101 = 10'h9e == _T_445[9:0] ? 4'h3 : _GEN_21100; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21102 = 10'h9f == _T_445[9:0] ? 4'h0 : _GEN_21101; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21103 = 10'ha0 == _T_445[9:0] ? 4'ha : _GEN_21102; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21104 = 10'ha1 == _T_445[9:0] ? 4'h1 : _GEN_21103; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21105 = 10'ha2 == _T_445[9:0] ? 4'h0 : _GEN_21104; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21106 = 10'ha3 == _T_445[9:0] ? 4'h3 : _GEN_21105; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21107 = 10'ha4 == _T_445[9:0] ? 4'ha : _GEN_21106; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21108 = 10'ha5 == _T_445[9:0] ? 4'ha : _GEN_21107; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21109 = 10'ha6 == _T_445[9:0] ? 4'ha : _GEN_21108; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21110 = 10'ha7 == _T_445[9:0] ? 4'h0 : _GEN_21109; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21111 = 10'ha8 == _T_445[9:0] ? 4'ha : _GEN_21110; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21112 = 10'ha9 == _T_445[9:0] ? 4'h1 : _GEN_21111; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21113 = 10'haa == _T_445[9:0] ? 4'h0 : _GEN_21112; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21114 = 10'hab == _T_445[9:0] ? 4'h0 : _GEN_21113; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21115 = 10'hac == _T_445[9:0] ? 4'h0 : _GEN_21114; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21116 = 10'had == _T_445[9:0] ? 4'h0 : _GEN_21115; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21117 = 10'hae == _T_445[9:0] ? 4'h0 : _GEN_21116; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21118 = 10'haf == _T_445[9:0] ? 4'h0 : _GEN_21117; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21119 = 10'hb0 == _T_445[9:0] ? 4'h0 : _GEN_21118; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21120 = 10'hb1 == _T_445[9:0] ? 4'h0 : _GEN_21119; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21121 = 10'hb2 == _T_445[9:0] ? 4'h0 : _GEN_21120; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21122 = 10'hb3 == _T_445[9:0] ? 4'h0 : _GEN_21121; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21123 = 10'hb4 == _T_445[9:0] ? 4'h1 : _GEN_21122; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21124 = 10'hb5 == _T_445[9:0] ? 4'h1 : _GEN_21123; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21125 = 10'hb6 == _T_445[9:0] ? 4'ha : _GEN_21124; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21126 = 10'hb7 == _T_445[9:0] ? 4'h0 : _GEN_21125; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21127 = 10'hb8 == _T_445[9:0] ? 4'ha : _GEN_21126; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21128 = 10'hb9 == _T_445[9:0] ? 4'ha : _GEN_21127; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21129 = 10'hba == _T_445[9:0] ? 4'ha : _GEN_21128; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21130 = 10'hbb == _T_445[9:0] ? 4'h0 : _GEN_21129; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21131 = 10'hbc == _T_445[9:0] ? 4'ha : _GEN_21130; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21132 = 10'hbd == _T_445[9:0] ? 4'ha : _GEN_21131; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21133 = 10'hbe == _T_445[9:0] ? 4'h3 : _GEN_21132; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21134 = 10'hbf == _T_445[9:0] ? 4'h0 : _GEN_21133; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21135 = 10'hc0 == _T_445[9:0] ? 4'ha : _GEN_21134; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21136 = 10'hc1 == _T_445[9:0] ? 4'ha : _GEN_21135; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21137 = 10'hc2 == _T_445[9:0] ? 4'h3 : _GEN_21136; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21138 = 10'hc3 == _T_445[9:0] ? 4'h2 : _GEN_21137; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21139 = 10'hc4 == _T_445[9:0] ? 4'h0 : _GEN_21138; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21140 = 10'hc5 == _T_445[9:0] ? 4'h0 : _GEN_21139; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21141 = 10'hc6 == _T_445[9:0] ? 4'h0 : _GEN_21140; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21142 = 10'hc7 == _T_445[9:0] ? 4'ha : _GEN_21141; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21143 = 10'hc8 == _T_445[9:0] ? 4'h1 : _GEN_21142; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21144 = 10'hc9 == _T_445[9:0] ? 4'h0 : _GEN_21143; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21145 = 10'hca == _T_445[9:0] ? 4'h0 : _GEN_21144; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21146 = 10'hcb == _T_445[9:0] ? 4'h0 : _GEN_21145; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21147 = 10'hcc == _T_445[9:0] ? 4'h0 : _GEN_21146; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21148 = 10'hcd == _T_445[9:0] ? 4'h0 : _GEN_21147; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21149 = 10'hce == _T_445[9:0] ? 4'h0 : _GEN_21148; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21150 = 10'hcf == _T_445[9:0] ? 4'h0 : _GEN_21149; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21151 = 10'hd0 == _T_445[9:0] ? 4'h0 : _GEN_21150; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21152 = 10'hd1 == _T_445[9:0] ? 4'h0 : _GEN_21151; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21153 = 10'hd2 == _T_445[9:0] ? 4'h0 : _GEN_21152; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21154 = 10'hd3 == _T_445[9:0] ? 4'h0 : _GEN_21153; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21155 = 10'hd4 == _T_445[9:0] ? 4'h0 : _GEN_21154; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21156 = 10'hd5 == _T_445[9:0] ? 4'h0 : _GEN_21155; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21157 = 10'hd6 == _T_445[9:0] ? 4'h1 : _GEN_21156; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21158 = 10'hd7 == _T_445[9:0] ? 4'ha : _GEN_21157; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21159 = 10'hd8 == _T_445[9:0] ? 4'h0 : _GEN_21158; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21160 = 10'hd9 == _T_445[9:0] ? 4'ha : _GEN_21159; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21161 = 10'hda == _T_445[9:0] ? 4'ha : _GEN_21160; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21162 = 10'hdb == _T_445[9:0] ? 4'ha : _GEN_21161; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21163 = 10'hdc == _T_445[9:0] ? 4'ha : _GEN_21162; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21164 = 10'hdd == _T_445[9:0] ? 4'h3 : _GEN_21163; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21165 = 10'hde == _T_445[9:0] ? 4'h2 : _GEN_21164; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21166 = 10'hdf == _T_445[9:0] ? 4'h0 : _GEN_21165; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21167 = 10'he0 == _T_445[9:0] ? 4'ha : _GEN_21166; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21168 = 10'he1 == _T_445[9:0] ? 4'ha : _GEN_21167; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21169 = 10'he2 == _T_445[9:0] ? 4'h3 : _GEN_21168; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21170 = 10'he3 == _T_445[9:0] ? 4'ha : _GEN_21169; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21171 = 10'he4 == _T_445[9:0] ? 4'ha : _GEN_21170; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21172 = 10'he5 == _T_445[9:0] ? 4'ha : _GEN_21171; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21173 = 10'he6 == _T_445[9:0] ? 4'ha : _GEN_21172; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21174 = 10'he7 == _T_445[9:0] ? 4'h1 : _GEN_21173; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21175 = 10'he8 == _T_445[9:0] ? 4'h1 : _GEN_21174; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21176 = 10'he9 == _T_445[9:0] ? 4'h1 : _GEN_21175; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21177 = 10'hea == _T_445[9:0] ? 4'h0 : _GEN_21176; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21178 = 10'heb == _T_445[9:0] ? 4'h0 : _GEN_21177; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21179 = 10'hec == _T_445[9:0] ? 4'h0 : _GEN_21178; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21180 = 10'hed == _T_445[9:0] ? 4'h0 : _GEN_21179; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21181 = 10'hee == _T_445[9:0] ? 4'h0 : _GEN_21180; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21182 = 10'hef == _T_445[9:0] ? 4'h0 : _GEN_21181; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21183 = 10'hf0 == _T_445[9:0] ? 4'h0 : _GEN_21182; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21184 = 10'hf1 == _T_445[9:0] ? 4'h0 : _GEN_21183; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21185 = 10'hf2 == _T_445[9:0] ? 4'h0 : _GEN_21184; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21186 = 10'hf3 == _T_445[9:0] ? 4'h0 : _GEN_21185; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21187 = 10'hf4 == _T_445[9:0] ? 4'h0 : _GEN_21186; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21188 = 10'hf5 == _T_445[9:0] ? 4'h1 : _GEN_21187; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21189 = 10'hf6 == _T_445[9:0] ? 4'h0 : _GEN_21188; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21190 = 10'hf7 == _T_445[9:0] ? 4'h0 : _GEN_21189; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21191 = 10'hf8 == _T_445[9:0] ? 4'h1 : _GEN_21190; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21192 = 10'hf9 == _T_445[9:0] ? 4'h0 : _GEN_21191; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21193 = 10'hfa == _T_445[9:0] ? 4'ha : _GEN_21192; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21194 = 10'hfb == _T_445[9:0] ? 4'ha : _GEN_21193; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21195 = 10'hfc == _T_445[9:0] ? 4'ha : _GEN_21194; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21196 = 10'hfd == _T_445[9:0] ? 4'h3 : _GEN_21195; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21197 = 10'hfe == _T_445[9:0] ? 4'ha : _GEN_21196; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21198 = 10'hff == _T_445[9:0] ? 4'h0 : _GEN_21197; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21199 = 10'h100 == _T_445[9:0] ? 4'ha : _GEN_21198; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21200 = 10'h101 == _T_445[9:0] ? 4'h0 : _GEN_21199; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21201 = 10'h102 == _T_445[9:0] ? 4'h3 : _GEN_21200; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21202 = 10'h103 == _T_445[9:0] ? 4'ha : _GEN_21201; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21203 = 10'h104 == _T_445[9:0] ? 4'ha : _GEN_21202; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21204 = 10'h105 == _T_445[9:0] ? 4'ha : _GEN_21203; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21205 = 10'h106 == _T_445[9:0] ? 4'ha : _GEN_21204; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21206 = 10'h107 == _T_445[9:0] ? 4'ha : _GEN_21205; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21207 = 10'h108 == _T_445[9:0] ? 4'h1 : _GEN_21206; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21208 = 10'h109 == _T_445[9:0] ? 4'h0 : _GEN_21207; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21209 = 10'h10a == _T_445[9:0] ? 4'h0 : _GEN_21208; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21210 = 10'h10b == _T_445[9:0] ? 4'h0 : _GEN_21209; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21211 = 10'h10c == _T_445[9:0] ? 4'h0 : _GEN_21210; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21212 = 10'h10d == _T_445[9:0] ? 4'h0 : _GEN_21211; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21213 = 10'h10e == _T_445[9:0] ? 4'h0 : _GEN_21212; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21214 = 10'h10f == _T_445[9:0] ? 4'h0 : _GEN_21213; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21215 = 10'h110 == _T_445[9:0] ? 4'h0 : _GEN_21214; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21216 = 10'h111 == _T_445[9:0] ? 4'h0 : _GEN_21215; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21217 = 10'h112 == _T_445[9:0] ? 4'h0 : _GEN_21216; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21218 = 10'h113 == _T_445[9:0] ? 4'h0 : _GEN_21217; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21219 = 10'h114 == _T_445[9:0] ? 4'h0 : _GEN_21218; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21220 = 10'h115 == _T_445[9:0] ? 4'h0 : _GEN_21219; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21221 = 10'h116 == _T_445[9:0] ? 4'h1 : _GEN_21220; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21222 = 10'h117 == _T_445[9:0] ? 4'ha : _GEN_21221; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21223 = 10'h118 == _T_445[9:0] ? 4'ha : _GEN_21222; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21224 = 10'h119 == _T_445[9:0] ? 4'ha : _GEN_21223; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21225 = 10'h11a == _T_445[9:0] ? 4'h0 : _GEN_21224; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21226 = 10'h11b == _T_445[9:0] ? 4'ha : _GEN_21225; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21227 = 10'h11c == _T_445[9:0] ? 4'ha : _GEN_21226; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21228 = 10'h11d == _T_445[9:0] ? 4'h2 : _GEN_21227; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21229 = 10'h11e == _T_445[9:0] ? 4'h3 : _GEN_21228; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21230 = 10'h11f == _T_445[9:0] ? 4'h0 : _GEN_21229; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21231 = 10'h120 == _T_445[9:0] ? 4'ha : _GEN_21230; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21232 = 10'h121 == _T_445[9:0] ? 4'ha : _GEN_21231; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21233 = 10'h122 == _T_445[9:0] ? 4'h3 : _GEN_21232; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21234 = 10'h123 == _T_445[9:0] ? 4'ha : _GEN_21233; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21235 = 10'h124 == _T_445[9:0] ? 4'ha : _GEN_21234; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21236 = 10'h125 == _T_445[9:0] ? 4'ha : _GEN_21235; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21237 = 10'h126 == _T_445[9:0] ? 4'ha : _GEN_21236; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21238 = 10'h127 == _T_445[9:0] ? 4'h1 : _GEN_21237; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21239 = 10'h128 == _T_445[9:0] ? 4'h0 : _GEN_21238; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21240 = 10'h129 == _T_445[9:0] ? 4'ha : _GEN_21239; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21241 = 10'h12a == _T_445[9:0] ? 4'ha : _GEN_21240; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21242 = 10'h12b == _T_445[9:0] ? 4'h0 : _GEN_21241; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21243 = 10'h12c == _T_445[9:0] ? 4'h0 : _GEN_21242; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21244 = 10'h12d == _T_445[9:0] ? 4'h0 : _GEN_21243; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21245 = 10'h12e == _T_445[9:0] ? 4'h0 : _GEN_21244; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21246 = 10'h12f == _T_445[9:0] ? 4'h0 : _GEN_21245; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21247 = 10'h130 == _T_445[9:0] ? 4'h0 : _GEN_21246; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21248 = 10'h131 == _T_445[9:0] ? 4'h0 : _GEN_21247; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21249 = 10'h132 == _T_445[9:0] ? 4'h0 : _GEN_21248; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21250 = 10'h133 == _T_445[9:0] ? 4'h0 : _GEN_21249; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21251 = 10'h134 == _T_445[9:0] ? 4'ha : _GEN_21250; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21252 = 10'h135 == _T_445[9:0] ? 4'ha : _GEN_21251; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21253 = 10'h136 == _T_445[9:0] ? 4'h0 : _GEN_21252; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21254 = 10'h137 == _T_445[9:0] ? 4'h1 : _GEN_21253; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21255 = 10'h138 == _T_445[9:0] ? 4'ha : _GEN_21254; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21256 = 10'h139 == _T_445[9:0] ? 4'ha : _GEN_21255; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21257 = 10'h13a == _T_445[9:0] ? 4'ha : _GEN_21256; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21258 = 10'h13b == _T_445[9:0] ? 4'ha : _GEN_21257; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21259 = 10'h13c == _T_445[9:0] ? 4'ha : _GEN_21258; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21260 = 10'h13d == _T_445[9:0] ? 4'ha : _GEN_21259; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21261 = 10'h13e == _T_445[9:0] ? 4'h3 : _GEN_21260; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21262 = 10'h13f == _T_445[9:0] ? 4'h0 : _GEN_21261; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21263 = 10'h140 == _T_445[9:0] ? 4'ha : _GEN_21262; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21264 = 10'h141 == _T_445[9:0] ? 4'ha : _GEN_21263; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21265 = 10'h142 == _T_445[9:0] ? 4'h2 : _GEN_21264; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21266 = 10'h143 == _T_445[9:0] ? 4'h3 : _GEN_21265; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21267 = 10'h144 == _T_445[9:0] ? 4'ha : _GEN_21266; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21268 = 10'h145 == _T_445[9:0] ? 4'ha : _GEN_21267; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21269 = 10'h146 == _T_445[9:0] ? 4'h1 : _GEN_21268; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21270 = 10'h147 == _T_445[9:0] ? 4'h0 : _GEN_21269; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21271 = 10'h148 == _T_445[9:0] ? 4'ha : _GEN_21270; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21272 = 10'h149 == _T_445[9:0] ? 4'ha : _GEN_21271; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21273 = 10'h14a == _T_445[9:0] ? 4'ha : _GEN_21272; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21274 = 10'h14b == _T_445[9:0] ? 4'ha : _GEN_21273; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21275 = 10'h14c == _T_445[9:0] ? 4'ha : _GEN_21274; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21276 = 10'h14d == _T_445[9:0] ? 4'ha : _GEN_21275; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21277 = 10'h14e == _T_445[9:0] ? 4'ha : _GEN_21276; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21278 = 10'h14f == _T_445[9:0] ? 4'ha : _GEN_21277; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21279 = 10'h150 == _T_445[9:0] ? 4'ha : _GEN_21278; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21280 = 10'h151 == _T_445[9:0] ? 4'ha : _GEN_21279; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21281 = 10'h152 == _T_445[9:0] ? 4'ha : _GEN_21280; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21282 = 10'h153 == _T_445[9:0] ? 4'ha : _GEN_21281; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21283 = 10'h154 == _T_445[9:0] ? 4'ha : _GEN_21282; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21284 = 10'h155 == _T_445[9:0] ? 4'ha : _GEN_21283; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21285 = 10'h156 == _T_445[9:0] ? 4'ha : _GEN_21284; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21286 = 10'h157 == _T_445[9:0] ? 4'h0 : _GEN_21285; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21287 = 10'h158 == _T_445[9:0] ? 4'ha : _GEN_21286; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21288 = 10'h159 == _T_445[9:0] ? 4'ha : _GEN_21287; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21289 = 10'h15a == _T_445[9:0] ? 4'ha : _GEN_21288; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21290 = 10'h15b == _T_445[9:0] ? 4'ha : _GEN_21289; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21291 = 10'h15c == _T_445[9:0] ? 4'ha : _GEN_21290; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21292 = 10'h15d == _T_445[9:0] ? 4'h3 : _GEN_21291; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21293 = 10'h15e == _T_445[9:0] ? 4'h2 : _GEN_21292; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21294 = 10'h15f == _T_445[9:0] ? 4'h0 : _GEN_21293; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21295 = 10'h160 == _T_445[9:0] ? 4'ha : _GEN_21294; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21296 = 10'h161 == _T_445[9:0] ? 4'ha : _GEN_21295; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21297 = 10'h162 == _T_445[9:0] ? 4'ha : _GEN_21296; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21298 = 10'h163 == _T_445[9:0] ? 4'h2 : _GEN_21297; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21299 = 10'h164 == _T_445[9:0] ? 4'h3 : _GEN_21298; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21300 = 10'h165 == _T_445[9:0] ? 4'h1 : _GEN_21299; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21301 = 10'h166 == _T_445[9:0] ? 4'h0 : _GEN_21300; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21302 = 10'h167 == _T_445[9:0] ? 4'h0 : _GEN_21301; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21303 = 10'h168 == _T_445[9:0] ? 4'h5 : _GEN_21302; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21304 = 10'h169 == _T_445[9:0] ? 4'h3 : _GEN_21303; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21305 = 10'h16a == _T_445[9:0] ? 4'h5 : _GEN_21304; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21306 = 10'h16b == _T_445[9:0] ? 4'h5 : _GEN_21305; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21307 = 10'h16c == _T_445[9:0] ? 4'ha : _GEN_21306; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21308 = 10'h16d == _T_445[9:0] ? 4'ha : _GEN_21307; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21309 = 10'h16e == _T_445[9:0] ? 4'ha : _GEN_21308; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21310 = 10'h16f == _T_445[9:0] ? 4'ha : _GEN_21309; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21311 = 10'h170 == _T_445[9:0] ? 4'ha : _GEN_21310; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21312 = 10'h171 == _T_445[9:0] ? 4'ha : _GEN_21311; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21313 = 10'h172 == _T_445[9:0] ? 4'ha : _GEN_21312; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21314 = 10'h173 == _T_445[9:0] ? 4'ha : _GEN_21313; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21315 = 10'h174 == _T_445[9:0] ? 4'ha : _GEN_21314; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21316 = 10'h175 == _T_445[9:0] ? 4'ha : _GEN_21315; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21317 = 10'h176 == _T_445[9:0] ? 4'h0 : _GEN_21316; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21318 = 10'h177 == _T_445[9:0] ? 4'h0 : _GEN_21317; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21319 = 10'h178 == _T_445[9:0] ? 4'h1 : _GEN_21318; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21320 = 10'h179 == _T_445[9:0] ? 4'ha : _GEN_21319; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21321 = 10'h17a == _T_445[9:0] ? 4'ha : _GEN_21320; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21322 = 10'h17b == _T_445[9:0] ? 4'ha : _GEN_21321; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21323 = 10'h17c == _T_445[9:0] ? 4'h3 : _GEN_21322; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21324 = 10'h17d == _T_445[9:0] ? 4'h2 : _GEN_21323; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21325 = 10'h17e == _T_445[9:0] ? 4'ha : _GEN_21324; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21326 = 10'h17f == _T_445[9:0] ? 4'h0 : _GEN_21325; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21327 = 10'h180 == _T_445[9:0] ? 4'h5 : _GEN_21326; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21328 = 10'h181 == _T_445[9:0] ? 4'h5 : _GEN_21327; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21329 = 10'h182 == _T_445[9:0] ? 4'h5 : _GEN_21328; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21330 = 10'h183 == _T_445[9:0] ? 4'h5 : _GEN_21329; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21331 = 10'h184 == _T_445[9:0] ? 4'h3 : _GEN_21330; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21332 = 10'h185 == _T_445[9:0] ? 4'h1 : _GEN_21331; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21333 = 10'h186 == _T_445[9:0] ? 4'hb : _GEN_21332; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21334 = 10'h187 == _T_445[9:0] ? 4'h0 : _GEN_21333; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21335 = 10'h188 == _T_445[9:0] ? 4'h5 : _GEN_21334; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21336 = 10'h189 == _T_445[9:0] ? 4'h5 : _GEN_21335; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21337 = 10'h18a == _T_445[9:0] ? 4'h5 : _GEN_21336; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21338 = 10'h18b == _T_445[9:0] ? 4'h5 : _GEN_21337; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21339 = 10'h18c == _T_445[9:0] ? 4'h5 : _GEN_21338; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21340 = 10'h18d == _T_445[9:0] ? 4'h5 : _GEN_21339; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21341 = 10'h18e == _T_445[9:0] ? 4'h5 : _GEN_21340; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21342 = 10'h18f == _T_445[9:0] ? 4'h5 : _GEN_21341; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21343 = 10'h190 == _T_445[9:0] ? 4'h5 : _GEN_21342; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21344 = 10'h191 == _T_445[9:0] ? 4'h5 : _GEN_21343; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21345 = 10'h192 == _T_445[9:0] ? 4'h3 : _GEN_21344; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21346 = 10'h193 == _T_445[9:0] ? 4'h5 : _GEN_21345; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21347 = 10'h194 == _T_445[9:0] ? 4'h5 : _GEN_21346; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21348 = 10'h195 == _T_445[9:0] ? 4'h5 : _GEN_21347; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21349 = 10'h196 == _T_445[9:0] ? 4'h0 : _GEN_21348; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21350 = 10'h197 == _T_445[9:0] ? 4'ha : _GEN_21349; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21351 = 10'h198 == _T_445[9:0] ? 4'h1 : _GEN_21350; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21352 = 10'h199 == _T_445[9:0] ? 4'ha : _GEN_21351; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21353 = 10'h19a == _T_445[9:0] ? 4'ha : _GEN_21352; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21354 = 10'h19b == _T_445[9:0] ? 4'ha : _GEN_21353; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21355 = 10'h19c == _T_445[9:0] ? 4'h3 : _GEN_21354; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21356 = 10'h19d == _T_445[9:0] ? 4'ha : _GEN_21355; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21357 = 10'h19e == _T_445[9:0] ? 4'ha : _GEN_21356; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21358 = 10'h19f == _T_445[9:0] ? 4'h0 : _GEN_21357; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21359 = 10'h1a0 == _T_445[9:0] ? 4'h5 : _GEN_21358; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21360 = 10'h1a1 == _T_445[9:0] ? 4'h5 : _GEN_21359; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21361 = 10'h1a2 == _T_445[9:0] ? 4'h3 : _GEN_21360; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21362 = 10'h1a3 == _T_445[9:0] ? 4'h5 : _GEN_21361; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21363 = 10'h1a4 == _T_445[9:0] ? 4'h3 : _GEN_21362; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21364 = 10'h1a5 == _T_445[9:0] ? 4'h0 : _GEN_21363; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21365 = 10'h1a6 == _T_445[9:0] ? 4'h5 : _GEN_21364; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21366 = 10'h1a7 == _T_445[9:0] ? 4'h0 : _GEN_21365; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21367 = 10'h1a8 == _T_445[9:0] ? 4'hb : _GEN_21366; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21368 = 10'h1a9 == _T_445[9:0] ? 4'h5 : _GEN_21367; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21369 = 10'h1aa == _T_445[9:0] ? 4'h5 : _GEN_21368; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21370 = 10'h1ab == _T_445[9:0] ? 4'h3 : _GEN_21369; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21371 = 10'h1ac == _T_445[9:0] ? 4'h5 : _GEN_21370; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21372 = 10'h1ad == _T_445[9:0] ? 4'h5 : _GEN_21371; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21373 = 10'h1ae == _T_445[9:0] ? 4'h5 : _GEN_21372; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21374 = 10'h1af == _T_445[9:0] ? 4'h5 : _GEN_21373; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21375 = 10'h1b0 == _T_445[9:0] ? 4'h5 : _GEN_21374; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21376 = 10'h1b1 == _T_445[9:0] ? 4'h5 : _GEN_21375; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21377 = 10'h1b2 == _T_445[9:0] ? 4'h5 : _GEN_21376; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21378 = 10'h1b3 == _T_445[9:0] ? 4'h5 : _GEN_21377; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21379 = 10'h1b4 == _T_445[9:0] ? 4'h5 : _GEN_21378; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21380 = 10'h1b5 == _T_445[9:0] ? 4'h5 : _GEN_21379; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21381 = 10'h1b6 == _T_445[9:0] ? 4'h0 : _GEN_21380; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21382 = 10'h1b7 == _T_445[9:0] ? 4'h5 : _GEN_21381; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21383 = 10'h1b8 == _T_445[9:0] ? 4'h0 : _GEN_21382; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21384 = 10'h1b9 == _T_445[9:0] ? 4'h5 : _GEN_21383; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21385 = 10'h1ba == _T_445[9:0] ? 4'h5 : _GEN_21384; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21386 = 10'h1bb == _T_445[9:0] ? 4'h5 : _GEN_21385; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21387 = 10'h1bc == _T_445[9:0] ? 4'h2 : _GEN_21386; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21388 = 10'h1bd == _T_445[9:0] ? 4'h3 : _GEN_21387; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21389 = 10'h1be == _T_445[9:0] ? 4'h5 : _GEN_21388; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21390 = 10'h1bf == _T_445[9:0] ? 4'h0 : _GEN_21389; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21391 = 10'h1c0 == _T_445[9:0] ? 4'h5 : _GEN_21390; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21392 = 10'h1c1 == _T_445[9:0] ? 4'h5 : _GEN_21391; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21393 = 10'h1c2 == _T_445[9:0] ? 4'h5 : _GEN_21392; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21394 = 10'h1c3 == _T_445[9:0] ? 4'h2 : _GEN_21393; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21395 = 10'h1c4 == _T_445[9:0] ? 4'h2 : _GEN_21394; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21396 = 10'h1c5 == _T_445[9:0] ? 4'h5 : _GEN_21395; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21397 = 10'h1c6 == _T_445[9:0] ? 4'h5 : _GEN_21396; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21398 = 10'h1c7 == _T_445[9:0] ? 4'h5 : _GEN_21397; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21399 = 10'h1c8 == _T_445[9:0] ? 4'h5 : _GEN_21398; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21400 = 10'h1c9 == _T_445[9:0] ? 4'hb : _GEN_21399; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21401 = 10'h1ca == _T_445[9:0] ? 4'hb : _GEN_21400; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21402 = 10'h1cb == _T_445[9:0] ? 4'hb : _GEN_21401; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21403 = 10'h1cc == _T_445[9:0] ? 4'hb : _GEN_21402; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21404 = 10'h1cd == _T_445[9:0] ? 4'hb : _GEN_21403; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21405 = 10'h1ce == _T_445[9:0] ? 4'hb : _GEN_21404; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21406 = 10'h1cf == _T_445[9:0] ? 4'hb : _GEN_21405; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21407 = 10'h1d0 == _T_445[9:0] ? 4'hb : _GEN_21406; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21408 = 10'h1d1 == _T_445[9:0] ? 4'hb : _GEN_21407; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21409 = 10'h1d2 == _T_445[9:0] ? 4'hb : _GEN_21408; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21410 = 10'h1d3 == _T_445[9:0] ? 4'hb : _GEN_21409; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21411 = 10'h1d4 == _T_445[9:0] ? 4'hb : _GEN_21410; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21412 = 10'h1d5 == _T_445[9:0] ? 4'hb : _GEN_21411; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21413 = 10'h1d6 == _T_445[9:0] ? 4'h5 : _GEN_21412; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21414 = 10'h1d7 == _T_445[9:0] ? 4'h5 : _GEN_21413; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21415 = 10'h1d8 == _T_445[9:0] ? 4'h5 : _GEN_21414; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21416 = 10'h1d9 == _T_445[9:0] ? 4'h5 : _GEN_21415; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21417 = 10'h1da == _T_445[9:0] ? 4'h5 : _GEN_21416; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21418 = 10'h1db == _T_445[9:0] ? 4'h5 : _GEN_21417; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21419 = 10'h1dc == _T_445[9:0] ? 4'h5 : _GEN_21418; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21420 = 10'h1dd == _T_445[9:0] ? 4'h3 : _GEN_21419; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21421 = 10'h1de == _T_445[9:0] ? 4'h5 : _GEN_21420; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21422 = 10'h1df == _T_445[9:0] ? 4'h0 : _GEN_21421; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21423 = 10'h1e0 == _T_445[9:0] ? 4'h3 : _GEN_21422; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21424 = 10'h1e1 == _T_445[9:0] ? 4'h5 : _GEN_21423; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21425 = 10'h1e2 == _T_445[9:0] ? 4'h2 : _GEN_21424; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21426 = 10'h1e3 == _T_445[9:0] ? 4'h2 : _GEN_21425; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21427 = 10'h1e4 == _T_445[9:0] ? 4'h5 : _GEN_21426; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21428 = 10'h1e5 == _T_445[9:0] ? 4'h5 : _GEN_21427; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21429 = 10'h1e6 == _T_445[9:0] ? 4'h5 : _GEN_21428; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21430 = 10'h1e7 == _T_445[9:0] ? 4'h5 : _GEN_21429; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21431 = 10'h1e8 == _T_445[9:0] ? 4'hb : _GEN_21430; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21432 = 10'h1e9 == _T_445[9:0] ? 4'h5 : _GEN_21431; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21433 = 10'h1ea == _T_445[9:0] ? 4'h5 : _GEN_21432; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21434 = 10'h1eb == _T_445[9:0] ? 4'hb : _GEN_21433; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21435 = 10'h1ec == _T_445[9:0] ? 4'h5 : _GEN_21434; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21436 = 10'h1ed == _T_445[9:0] ? 4'hb : _GEN_21435; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21437 = 10'h1ee == _T_445[9:0] ? 4'h5 : _GEN_21436; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21438 = 10'h1ef == _T_445[9:0] ? 4'hb : _GEN_21437; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21439 = 10'h1f0 == _T_445[9:0] ? 4'h5 : _GEN_21438; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21440 = 10'h1f1 == _T_445[9:0] ? 4'hb : _GEN_21439; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21441 = 10'h1f2 == _T_445[9:0] ? 4'hb : _GEN_21440; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21442 = 10'h1f3 == _T_445[9:0] ? 4'h5 : _GEN_21441; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21443 = 10'h1f4 == _T_445[9:0] ? 4'hb : _GEN_21442; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21444 = 10'h1f5 == _T_445[9:0] ? 4'hb : _GEN_21443; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21445 = 10'h1f6 == _T_445[9:0] ? 4'h5 : _GEN_21444; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21446 = 10'h1f7 == _T_445[9:0] ? 4'h5 : _GEN_21445; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21447 = 10'h1f8 == _T_445[9:0] ? 4'h5 : _GEN_21446; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21448 = 10'h1f9 == _T_445[9:0] ? 4'h5 : _GEN_21447; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21449 = 10'h1fa == _T_445[9:0] ? 4'h3 : _GEN_21448; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21450 = 10'h1fb == _T_445[9:0] ? 4'h5 : _GEN_21449; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21451 = 10'h1fc == _T_445[9:0] ? 4'h5 : _GEN_21450; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21452 = 10'h1fd == _T_445[9:0] ? 4'h2 : _GEN_21451; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21453 = 10'h1fe == _T_445[9:0] ? 4'h5 : _GEN_21452; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21454 = 10'h1ff == _T_445[9:0] ? 4'h0 : _GEN_21453; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21455 = 10'h200 == _T_445[9:0] ? 4'h5 : _GEN_21454; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21456 = 10'h201 == _T_445[9:0] ? 4'h5 : _GEN_21455; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21457 = 10'h202 == _T_445[9:0] ? 4'h3 : _GEN_21456; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21458 = 10'h203 == _T_445[9:0] ? 4'h5 : _GEN_21457; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21459 = 10'h204 == _T_445[9:0] ? 4'h5 : _GEN_21458; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21460 = 10'h205 == _T_445[9:0] ? 4'h5 : _GEN_21459; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21461 = 10'h206 == _T_445[9:0] ? 4'hb : _GEN_21460; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21462 = 10'h207 == _T_445[9:0] ? 4'hb : _GEN_21461; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21463 = 10'h208 == _T_445[9:0] ? 4'h5 : _GEN_21462; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21464 = 10'h209 == _T_445[9:0] ? 4'h5 : _GEN_21463; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21465 = 10'h20a == _T_445[9:0] ? 4'h5 : _GEN_21464; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21466 = 10'h20b == _T_445[9:0] ? 4'hb : _GEN_21465; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21467 = 10'h20c == _T_445[9:0] ? 4'h5 : _GEN_21466; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21468 = 10'h20d == _T_445[9:0] ? 4'hb : _GEN_21467; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21469 = 10'h20e == _T_445[9:0] ? 4'h5 : _GEN_21468; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21470 = 10'h20f == _T_445[9:0] ? 4'hb : _GEN_21469; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21471 = 10'h210 == _T_445[9:0] ? 4'h5 : _GEN_21470; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21472 = 10'h211 == _T_445[9:0] ? 4'h5 : _GEN_21471; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21473 = 10'h212 == _T_445[9:0] ? 4'hb : _GEN_21472; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21474 = 10'h213 == _T_445[9:0] ? 4'hb : _GEN_21473; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21475 = 10'h214 == _T_445[9:0] ? 4'hb : _GEN_21474; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21476 = 10'h215 == _T_445[9:0] ? 4'h5 : _GEN_21475; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21477 = 10'h216 == _T_445[9:0] ? 4'h5 : _GEN_21476; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21478 = 10'h217 == _T_445[9:0] ? 4'h5 : _GEN_21477; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21479 = 10'h218 == _T_445[9:0] ? 4'h5 : _GEN_21478; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21480 = 10'h219 == _T_445[9:0] ? 4'h5 : _GEN_21479; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21481 = 10'h21a == _T_445[9:0] ? 4'h5 : _GEN_21480; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21482 = 10'h21b == _T_445[9:0] ? 4'h5 : _GEN_21481; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21483 = 10'h21c == _T_445[9:0] ? 4'h3 : _GEN_21482; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21484 = 10'h21d == _T_445[9:0] ? 4'h2 : _GEN_21483; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21485 = 10'h21e == _T_445[9:0] ? 4'h5 : _GEN_21484; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21486 = 10'h21f == _T_445[9:0] ? 4'h0 : _GEN_21485; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21487 = 10'h220 == _T_445[9:0] ? 4'h0 : _GEN_21486; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21488 = 10'h221 == _T_445[9:0] ? 4'h0 : _GEN_21487; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21489 = 10'h222 == _T_445[9:0] ? 4'h0 : _GEN_21488; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21490 = 10'h223 == _T_445[9:0] ? 4'h0 : _GEN_21489; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21491 = 10'h224 == _T_445[9:0] ? 4'h0 : _GEN_21490; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21492 = 10'h225 == _T_445[9:0] ? 4'h0 : _GEN_21491; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21493 = 10'h226 == _T_445[9:0] ? 4'h0 : _GEN_21492; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21494 = 10'h227 == _T_445[9:0] ? 4'h0 : _GEN_21493; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21495 = 10'h228 == _T_445[9:0] ? 4'h0 : _GEN_21494; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21496 = 10'h229 == _T_445[9:0] ? 4'h0 : _GEN_21495; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21497 = 10'h22a == _T_445[9:0] ? 4'h0 : _GEN_21496; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21498 = 10'h22b == _T_445[9:0] ? 4'h0 : _GEN_21497; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21499 = 10'h22c == _T_445[9:0] ? 4'h0 : _GEN_21498; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21500 = 10'h22d == _T_445[9:0] ? 4'h0 : _GEN_21499; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21501 = 10'h22e == _T_445[9:0] ? 4'h0 : _GEN_21500; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21502 = 10'h22f == _T_445[9:0] ? 4'h0 : _GEN_21501; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21503 = 10'h230 == _T_445[9:0] ? 4'h0 : _GEN_21502; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21504 = 10'h231 == _T_445[9:0] ? 4'h0 : _GEN_21503; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21505 = 10'h232 == _T_445[9:0] ? 4'h0 : _GEN_21504; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21506 = 10'h233 == _T_445[9:0] ? 4'h0 : _GEN_21505; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21507 = 10'h234 == _T_445[9:0] ? 4'h0 : _GEN_21506; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21508 = 10'h235 == _T_445[9:0] ? 4'h0 : _GEN_21507; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21509 = 10'h236 == _T_445[9:0] ? 4'h0 : _GEN_21508; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21510 = 10'h237 == _T_445[9:0] ? 4'h0 : _GEN_21509; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21511 = 10'h238 == _T_445[9:0] ? 4'h0 : _GEN_21510; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21512 = 10'h239 == _T_445[9:0] ? 4'h0 : _GEN_21511; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21513 = 10'h23a == _T_445[9:0] ? 4'h0 : _GEN_21512; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21514 = 10'h23b == _T_445[9:0] ? 4'h0 : _GEN_21513; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21515 = 10'h23c == _T_445[9:0] ? 4'h0 : _GEN_21514; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21516 = 10'h23d == _T_445[9:0] ? 4'h0 : _GEN_21515; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21517 = 10'h23e == _T_445[9:0] ? 4'h0 : _GEN_21516; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21518 = 10'h23f == _T_445[9:0] ? 4'h0 : _GEN_21517; // @[Filter.scala 191:62]
  wire [4:0] _GEN_28370 = {{1'd0}, _GEN_21518}; // @[Filter.scala 191:62]
  wire [8:0] _T_447 = _GEN_28370 * 5'h14; // @[Filter.scala 191:62]
  wire [3:0] _GEN_21522 = 10'h3 == _T_445[9:0] ? 4'ha : 4'h3; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21523 = 10'h4 == _T_445[9:0] ? 4'h3 : _GEN_21522; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21524 = 10'h5 == _T_445[9:0] ? 4'h3 : _GEN_21523; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21525 = 10'h6 == _T_445[9:0] ? 4'h3 : _GEN_21524; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21526 = 10'h7 == _T_445[9:0] ? 4'h3 : _GEN_21525; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21527 = 10'h8 == _T_445[9:0] ? 4'h3 : _GEN_21526; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21528 = 10'h9 == _T_445[9:0] ? 4'h3 : _GEN_21527; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21529 = 10'ha == _T_445[9:0] ? 4'h3 : _GEN_21528; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21530 = 10'hb == _T_445[9:0] ? 4'h3 : _GEN_21529; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21531 = 10'hc == _T_445[9:0] ? 4'h5 : _GEN_21530; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21532 = 10'hd == _T_445[9:0] ? 4'h3 : _GEN_21531; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21533 = 10'he == _T_445[9:0] ? 4'h3 : _GEN_21532; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21534 = 10'hf == _T_445[9:0] ? 4'h3 : _GEN_21533; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21535 = 10'h10 == _T_445[9:0] ? 4'h3 : _GEN_21534; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21536 = 10'h11 == _T_445[9:0] ? 4'h3 : _GEN_21535; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21537 = 10'h12 == _T_445[9:0] ? 4'h3 : _GEN_21536; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21538 = 10'h13 == _T_445[9:0] ? 4'h3 : _GEN_21537; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21539 = 10'h14 == _T_445[9:0] ? 4'h3 : _GEN_21538; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21540 = 10'h15 == _T_445[9:0] ? 4'h3 : _GEN_21539; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21541 = 10'h16 == _T_445[9:0] ? 4'h3 : _GEN_21540; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21542 = 10'h17 == _T_445[9:0] ? 4'h3 : _GEN_21541; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21543 = 10'h18 == _T_445[9:0] ? 4'h3 : _GEN_21542; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21544 = 10'h19 == _T_445[9:0] ? 4'h3 : _GEN_21543; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21545 = 10'h1a == _T_445[9:0] ? 4'h3 : _GEN_21544; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21546 = 10'h1b == _T_445[9:0] ? 4'h3 : _GEN_21545; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21547 = 10'h1c == _T_445[9:0] ? 4'h3 : _GEN_21546; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21548 = 10'h1d == _T_445[9:0] ? 4'h3 : _GEN_21547; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21549 = 10'h1e == _T_445[9:0] ? 4'h3 : _GEN_21548; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21550 = 10'h1f == _T_445[9:0] ? 4'h0 : _GEN_21549; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21551 = 10'h20 == _T_445[9:0] ? 4'h3 : _GEN_21550; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21552 = 10'h21 == _T_445[9:0] ? 4'h5 : _GEN_21551; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21553 = 10'h22 == _T_445[9:0] ? 4'h3 : _GEN_21552; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21554 = 10'h23 == _T_445[9:0] ? 4'ha : _GEN_21553; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21555 = 10'h24 == _T_445[9:0] ? 4'h3 : _GEN_21554; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21556 = 10'h25 == _T_445[9:0] ? 4'h3 : _GEN_21555; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21557 = 10'h26 == _T_445[9:0] ? 4'h3 : _GEN_21556; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21558 = 10'h27 == _T_445[9:0] ? 4'h1 : _GEN_21557; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21559 = 10'h28 == _T_445[9:0] ? 4'h1 : _GEN_21558; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21560 = 10'h29 == _T_445[9:0] ? 4'h3 : _GEN_21559; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21561 = 10'h2a == _T_445[9:0] ? 4'h3 : _GEN_21560; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21562 = 10'h2b == _T_445[9:0] ? 4'h3 : _GEN_21561; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21563 = 10'h2c == _T_445[9:0] ? 4'h3 : _GEN_21562; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21564 = 10'h2d == _T_445[9:0] ? 4'h3 : _GEN_21563; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21565 = 10'h2e == _T_445[9:0] ? 4'h3 : _GEN_21564; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21566 = 10'h2f == _T_445[9:0] ? 4'h3 : _GEN_21565; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21567 = 10'h30 == _T_445[9:0] ? 4'h3 : _GEN_21566; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21568 = 10'h31 == _T_445[9:0] ? 4'h5 : _GEN_21567; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21569 = 10'h32 == _T_445[9:0] ? 4'h3 : _GEN_21568; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21570 = 10'h33 == _T_445[9:0] ? 4'h3 : _GEN_21569; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21571 = 10'h34 == _T_445[9:0] ? 4'h3 : _GEN_21570; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21572 = 10'h35 == _T_445[9:0] ? 4'h3 : _GEN_21571; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21573 = 10'h36 == _T_445[9:0] ? 4'h3 : _GEN_21572; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21574 = 10'h37 == _T_445[9:0] ? 4'h1 : _GEN_21573; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21575 = 10'h38 == _T_445[9:0] ? 4'h1 : _GEN_21574; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21576 = 10'h39 == _T_445[9:0] ? 4'h3 : _GEN_21575; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21577 = 10'h3a == _T_445[9:0] ? 4'h3 : _GEN_21576; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21578 = 10'h3b == _T_445[9:0] ? 4'h5 : _GEN_21577; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21579 = 10'h3c == _T_445[9:0] ? 4'h3 : _GEN_21578; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21580 = 10'h3d == _T_445[9:0] ? 4'ha : _GEN_21579; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21581 = 10'h3e == _T_445[9:0] ? 4'h3 : _GEN_21580; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21582 = 10'h3f == _T_445[9:0] ? 4'h0 : _GEN_21581; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21583 = 10'h40 == _T_445[9:0] ? 4'h3 : _GEN_21582; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21584 = 10'h41 == _T_445[9:0] ? 4'h3 : _GEN_21583; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21585 = 10'h42 == _T_445[9:0] ? 4'h3 : _GEN_21584; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21586 = 10'h43 == _T_445[9:0] ? 4'h7 : _GEN_21585; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21587 = 10'h44 == _T_445[9:0] ? 4'ha : _GEN_21586; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21588 = 10'h45 == _T_445[9:0] ? 4'h0 : _GEN_21587; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21589 = 10'h46 == _T_445[9:0] ? 4'h0 : _GEN_21588; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21590 = 10'h47 == _T_445[9:0] ? 4'h0 : _GEN_21589; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21591 = 10'h48 == _T_445[9:0] ? 4'h0 : _GEN_21590; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21592 = 10'h49 == _T_445[9:0] ? 4'h3 : _GEN_21591; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21593 = 10'h4a == _T_445[9:0] ? 4'h3 : _GEN_21592; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21594 = 10'h4b == _T_445[9:0] ? 4'h3 : _GEN_21593; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21595 = 10'h4c == _T_445[9:0] ? 4'h3 : _GEN_21594; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21596 = 10'h4d == _T_445[9:0] ? 4'h5 : _GEN_21595; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21597 = 10'h4e == _T_445[9:0] ? 4'h3 : _GEN_21596; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21598 = 10'h4f == _T_445[9:0] ? 4'h3 : _GEN_21597; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21599 = 10'h50 == _T_445[9:0] ? 4'h3 : _GEN_21598; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21600 = 10'h51 == _T_445[9:0] ? 4'h3 : _GEN_21599; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21601 = 10'h52 == _T_445[9:0] ? 4'h3 : _GEN_21600; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21602 = 10'h53 == _T_445[9:0] ? 4'h3 : _GEN_21601; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21603 = 10'h54 == _T_445[9:0] ? 4'h1 : _GEN_21602; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21604 = 10'h55 == _T_445[9:0] ? 4'h1 : _GEN_21603; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21605 = 10'h56 == _T_445[9:0] ? 4'h1 : _GEN_21604; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21606 = 10'h57 == _T_445[9:0] ? 4'h0 : _GEN_21605; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21607 = 10'h58 == _T_445[9:0] ? 4'h3 : _GEN_21606; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21608 = 10'h59 == _T_445[9:0] ? 4'h0 : _GEN_21607; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21609 = 10'h5a == _T_445[9:0] ? 4'h3 : _GEN_21608; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21610 = 10'h5b == _T_445[9:0] ? 4'h3 : _GEN_21609; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21611 = 10'h5c == _T_445[9:0] ? 4'h3 : _GEN_21610; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21612 = 10'h5d == _T_445[9:0] ? 4'ha : _GEN_21611; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21613 = 10'h5e == _T_445[9:0] ? 4'h3 : _GEN_21612; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21614 = 10'h5f == _T_445[9:0] ? 4'h0 : _GEN_21613; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21615 = 10'h60 == _T_445[9:0] ? 4'h3 : _GEN_21614; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21616 = 10'h61 == _T_445[9:0] ? 4'h3 : _GEN_21615; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21617 = 10'h62 == _T_445[9:0] ? 4'h3 : _GEN_21616; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21618 = 10'h63 == _T_445[9:0] ? 4'h3 : _GEN_21617; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21619 = 10'h64 == _T_445[9:0] ? 4'ha : _GEN_21618; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21620 = 10'h65 == _T_445[9:0] ? 4'h0 : _GEN_21619; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21621 = 10'h66 == _T_445[9:0] ? 4'h3 : _GEN_21620; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21622 = 10'h67 == _T_445[9:0] ? 4'h3 : _GEN_21621; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21623 = 10'h68 == _T_445[9:0] ? 4'h3 : _GEN_21622; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21624 = 10'h69 == _T_445[9:0] ? 4'h0 : _GEN_21623; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21625 = 10'h6a == _T_445[9:0] ? 4'h1 : _GEN_21624; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21626 = 10'h6b == _T_445[9:0] ? 4'h1 : _GEN_21625; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21627 = 10'h6c == _T_445[9:0] ? 4'h3 : _GEN_21626; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21628 = 10'h6d == _T_445[9:0] ? 4'h3 : _GEN_21627; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21629 = 10'h6e == _T_445[9:0] ? 4'h3 : _GEN_21628; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21630 = 10'h6f == _T_445[9:0] ? 4'h3 : _GEN_21629; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21631 = 10'h70 == _T_445[9:0] ? 4'h3 : _GEN_21630; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21632 = 10'h71 == _T_445[9:0] ? 4'h3 : _GEN_21631; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21633 = 10'h72 == _T_445[9:0] ? 4'h3 : _GEN_21632; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21634 = 10'h73 == _T_445[9:0] ? 4'h1 : _GEN_21633; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21635 = 10'h74 == _T_445[9:0] ? 4'h0 : _GEN_21634; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21636 = 10'h75 == _T_445[9:0] ? 4'h0 : _GEN_21635; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21637 = 10'h76 == _T_445[9:0] ? 4'h0 : _GEN_21636; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21638 = 10'h77 == _T_445[9:0] ? 4'h3 : _GEN_21637; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21639 = 10'h78 == _T_445[9:0] ? 4'h3 : _GEN_21638; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21640 = 10'h79 == _T_445[9:0] ? 4'h3 : _GEN_21639; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21641 = 10'h7a == _T_445[9:0] ? 4'h0 : _GEN_21640; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21642 = 10'h7b == _T_445[9:0] ? 4'h3 : _GEN_21641; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21643 = 10'h7c == _T_445[9:0] ? 4'h3 : _GEN_21642; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21644 = 10'h7d == _T_445[9:0] ? 4'h7 : _GEN_21643; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21645 = 10'h7e == _T_445[9:0] ? 4'ha : _GEN_21644; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21646 = 10'h7f == _T_445[9:0] ? 4'h0 : _GEN_21645; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21647 = 10'h80 == _T_445[9:0] ? 4'h3 : _GEN_21646; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21648 = 10'h81 == _T_445[9:0] ? 4'h3 : _GEN_21647; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21649 = 10'h82 == _T_445[9:0] ? 4'h1 : _GEN_21648; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21650 = 10'h83 == _T_445[9:0] ? 4'h0 : _GEN_21649; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21651 = 10'h84 == _T_445[9:0] ? 4'h7 : _GEN_21650; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21652 = 10'h85 == _T_445[9:0] ? 4'h1 : _GEN_21651; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21653 = 10'h86 == _T_445[9:0] ? 4'h1 : _GEN_21652; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21654 = 10'h87 == _T_445[9:0] ? 4'h3 : _GEN_21653; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21655 = 10'h88 == _T_445[9:0] ? 4'h3 : _GEN_21654; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21656 = 10'h89 == _T_445[9:0] ? 4'h0 : _GEN_21655; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21657 = 10'h8a == _T_445[9:0] ? 4'h0 : _GEN_21656; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21658 = 10'h8b == _T_445[9:0] ? 4'h1 : _GEN_21657; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21659 = 10'h8c == _T_445[9:0] ? 4'h1 : _GEN_21658; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21660 = 10'h8d == _T_445[9:0] ? 4'h1 : _GEN_21659; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21661 = 10'h8e == _T_445[9:0] ? 4'h1 : _GEN_21660; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21662 = 10'h8f == _T_445[9:0] ? 4'h1 : _GEN_21661; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21663 = 10'h90 == _T_445[9:0] ? 4'h1 : _GEN_21662; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21664 = 10'h91 == _T_445[9:0] ? 4'h1 : _GEN_21663; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21665 = 10'h92 == _T_445[9:0] ? 4'h1 : _GEN_21664; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21666 = 10'h93 == _T_445[9:0] ? 4'h0 : _GEN_21665; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21667 = 10'h94 == _T_445[9:0] ? 4'h0 : _GEN_21666; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21668 = 10'h95 == _T_445[9:0] ? 4'h3 : _GEN_21667; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21669 = 10'h96 == _T_445[9:0] ? 4'h3 : _GEN_21668; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21670 = 10'h97 == _T_445[9:0] ? 4'h3 : _GEN_21669; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21671 = 10'h98 == _T_445[9:0] ? 4'h1 : _GEN_21670; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21672 = 10'h99 == _T_445[9:0] ? 4'h0 : _GEN_21671; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21673 = 10'h9a == _T_445[9:0] ? 4'h1 : _GEN_21672; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21674 = 10'h9b == _T_445[9:0] ? 4'h1 : _GEN_21673; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21675 = 10'h9c == _T_445[9:0] ? 4'h3 : _GEN_21674; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21676 = 10'h9d == _T_445[9:0] ? 4'h3 : _GEN_21675; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21677 = 10'h9e == _T_445[9:0] ? 4'ha : _GEN_21676; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21678 = 10'h9f == _T_445[9:0] ? 4'h0 : _GEN_21677; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21679 = 10'ha0 == _T_445[9:0] ? 4'h3 : _GEN_21678; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21680 = 10'ha1 == _T_445[9:0] ? 4'h1 : _GEN_21679; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21681 = 10'ha2 == _T_445[9:0] ? 4'h0 : _GEN_21680; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21682 = 10'ha3 == _T_445[9:0] ? 4'ha : _GEN_21681; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21683 = 10'ha4 == _T_445[9:0] ? 4'h3 : _GEN_21682; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21684 = 10'ha5 == _T_445[9:0] ? 4'h3 : _GEN_21683; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21685 = 10'ha6 == _T_445[9:0] ? 4'h3 : _GEN_21684; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21686 = 10'ha7 == _T_445[9:0] ? 4'h0 : _GEN_21685; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21687 = 10'ha8 == _T_445[9:0] ? 4'h3 : _GEN_21686; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21688 = 10'ha9 == _T_445[9:0] ? 4'h1 : _GEN_21687; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21689 = 10'haa == _T_445[9:0] ? 4'h0 : _GEN_21688; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21690 = 10'hab == _T_445[9:0] ? 4'h0 : _GEN_21689; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21691 = 10'hac == _T_445[9:0] ? 4'h0 : _GEN_21690; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21692 = 10'had == _T_445[9:0] ? 4'h0 : _GEN_21691; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21693 = 10'hae == _T_445[9:0] ? 4'h0 : _GEN_21692; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21694 = 10'haf == _T_445[9:0] ? 4'h0 : _GEN_21693; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21695 = 10'hb0 == _T_445[9:0] ? 4'h0 : _GEN_21694; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21696 = 10'hb1 == _T_445[9:0] ? 4'h0 : _GEN_21695; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21697 = 10'hb2 == _T_445[9:0] ? 4'h0 : _GEN_21696; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21698 = 10'hb3 == _T_445[9:0] ? 4'h0 : _GEN_21697; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21699 = 10'hb4 == _T_445[9:0] ? 4'h1 : _GEN_21698; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21700 = 10'hb5 == _T_445[9:0] ? 4'h1 : _GEN_21699; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21701 = 10'hb6 == _T_445[9:0] ? 4'h3 : _GEN_21700; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21702 = 10'hb7 == _T_445[9:0] ? 4'h0 : _GEN_21701; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21703 = 10'hb8 == _T_445[9:0] ? 4'h3 : _GEN_21702; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21704 = 10'hb9 == _T_445[9:0] ? 4'h3 : _GEN_21703; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21705 = 10'hba == _T_445[9:0] ? 4'h3 : _GEN_21704; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21706 = 10'hbb == _T_445[9:0] ? 4'h0 : _GEN_21705; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21707 = 10'hbc == _T_445[9:0] ? 4'h3 : _GEN_21706; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21708 = 10'hbd == _T_445[9:0] ? 4'h3 : _GEN_21707; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21709 = 10'hbe == _T_445[9:0] ? 4'ha : _GEN_21708; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21710 = 10'hbf == _T_445[9:0] ? 4'h0 : _GEN_21709; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21711 = 10'hc0 == _T_445[9:0] ? 4'h3 : _GEN_21710; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21712 = 10'hc1 == _T_445[9:0] ? 4'h3 : _GEN_21711; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21713 = 10'hc2 == _T_445[9:0] ? 4'ha : _GEN_21712; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21714 = 10'hc3 == _T_445[9:0] ? 4'h7 : _GEN_21713; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21715 = 10'hc4 == _T_445[9:0] ? 4'h0 : _GEN_21714; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21716 = 10'hc5 == _T_445[9:0] ? 4'h0 : _GEN_21715; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21717 = 10'hc6 == _T_445[9:0] ? 4'h0 : _GEN_21716; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21718 = 10'hc7 == _T_445[9:0] ? 4'h3 : _GEN_21717; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21719 = 10'hc8 == _T_445[9:0] ? 4'h1 : _GEN_21718; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21720 = 10'hc9 == _T_445[9:0] ? 4'h0 : _GEN_21719; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21721 = 10'hca == _T_445[9:0] ? 4'h0 : _GEN_21720; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21722 = 10'hcb == _T_445[9:0] ? 4'h0 : _GEN_21721; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21723 = 10'hcc == _T_445[9:0] ? 4'h0 : _GEN_21722; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21724 = 10'hcd == _T_445[9:0] ? 4'h0 : _GEN_21723; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21725 = 10'hce == _T_445[9:0] ? 4'h0 : _GEN_21724; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21726 = 10'hcf == _T_445[9:0] ? 4'h0 : _GEN_21725; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21727 = 10'hd0 == _T_445[9:0] ? 4'h0 : _GEN_21726; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21728 = 10'hd1 == _T_445[9:0] ? 4'h0 : _GEN_21727; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21729 = 10'hd2 == _T_445[9:0] ? 4'h0 : _GEN_21728; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21730 = 10'hd3 == _T_445[9:0] ? 4'h0 : _GEN_21729; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21731 = 10'hd4 == _T_445[9:0] ? 4'h0 : _GEN_21730; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21732 = 10'hd5 == _T_445[9:0] ? 4'h0 : _GEN_21731; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21733 = 10'hd6 == _T_445[9:0] ? 4'h1 : _GEN_21732; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21734 = 10'hd7 == _T_445[9:0] ? 4'h3 : _GEN_21733; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21735 = 10'hd8 == _T_445[9:0] ? 4'h0 : _GEN_21734; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21736 = 10'hd9 == _T_445[9:0] ? 4'h3 : _GEN_21735; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21737 = 10'hda == _T_445[9:0] ? 4'h3 : _GEN_21736; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21738 = 10'hdb == _T_445[9:0] ? 4'h3 : _GEN_21737; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21739 = 10'hdc == _T_445[9:0] ? 4'h3 : _GEN_21738; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21740 = 10'hdd == _T_445[9:0] ? 4'ha : _GEN_21739; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21741 = 10'hde == _T_445[9:0] ? 4'h7 : _GEN_21740; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21742 = 10'hdf == _T_445[9:0] ? 4'h0 : _GEN_21741; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21743 = 10'he0 == _T_445[9:0] ? 4'h3 : _GEN_21742; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21744 = 10'he1 == _T_445[9:0] ? 4'h3 : _GEN_21743; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21745 = 10'he2 == _T_445[9:0] ? 4'ha : _GEN_21744; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21746 = 10'he3 == _T_445[9:0] ? 4'h3 : _GEN_21745; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21747 = 10'he4 == _T_445[9:0] ? 4'h3 : _GEN_21746; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21748 = 10'he5 == _T_445[9:0] ? 4'h3 : _GEN_21747; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21749 = 10'he6 == _T_445[9:0] ? 4'h3 : _GEN_21748; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21750 = 10'he7 == _T_445[9:0] ? 4'h1 : _GEN_21749; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21751 = 10'he8 == _T_445[9:0] ? 4'h1 : _GEN_21750; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21752 = 10'he9 == _T_445[9:0] ? 4'h1 : _GEN_21751; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21753 = 10'hea == _T_445[9:0] ? 4'h0 : _GEN_21752; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21754 = 10'heb == _T_445[9:0] ? 4'h0 : _GEN_21753; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21755 = 10'hec == _T_445[9:0] ? 4'h0 : _GEN_21754; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21756 = 10'hed == _T_445[9:0] ? 4'h0 : _GEN_21755; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21757 = 10'hee == _T_445[9:0] ? 4'h0 : _GEN_21756; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21758 = 10'hef == _T_445[9:0] ? 4'h0 : _GEN_21757; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21759 = 10'hf0 == _T_445[9:0] ? 4'h0 : _GEN_21758; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21760 = 10'hf1 == _T_445[9:0] ? 4'h0 : _GEN_21759; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21761 = 10'hf2 == _T_445[9:0] ? 4'h0 : _GEN_21760; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21762 = 10'hf3 == _T_445[9:0] ? 4'h0 : _GEN_21761; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21763 = 10'hf4 == _T_445[9:0] ? 4'h0 : _GEN_21762; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21764 = 10'hf5 == _T_445[9:0] ? 4'h1 : _GEN_21763; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21765 = 10'hf6 == _T_445[9:0] ? 4'h0 : _GEN_21764; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21766 = 10'hf7 == _T_445[9:0] ? 4'h0 : _GEN_21765; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21767 = 10'hf8 == _T_445[9:0] ? 4'h1 : _GEN_21766; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21768 = 10'hf9 == _T_445[9:0] ? 4'h0 : _GEN_21767; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21769 = 10'hfa == _T_445[9:0] ? 4'h3 : _GEN_21768; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21770 = 10'hfb == _T_445[9:0] ? 4'h3 : _GEN_21769; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21771 = 10'hfc == _T_445[9:0] ? 4'h3 : _GEN_21770; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21772 = 10'hfd == _T_445[9:0] ? 4'ha : _GEN_21771; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21773 = 10'hfe == _T_445[9:0] ? 4'h3 : _GEN_21772; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21774 = 10'hff == _T_445[9:0] ? 4'h0 : _GEN_21773; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21775 = 10'h100 == _T_445[9:0] ? 4'h3 : _GEN_21774; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21776 = 10'h101 == _T_445[9:0] ? 4'h0 : _GEN_21775; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21777 = 10'h102 == _T_445[9:0] ? 4'ha : _GEN_21776; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21778 = 10'h103 == _T_445[9:0] ? 4'h3 : _GEN_21777; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21779 = 10'h104 == _T_445[9:0] ? 4'h3 : _GEN_21778; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21780 = 10'h105 == _T_445[9:0] ? 4'h3 : _GEN_21779; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21781 = 10'h106 == _T_445[9:0] ? 4'h3 : _GEN_21780; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21782 = 10'h107 == _T_445[9:0] ? 4'h3 : _GEN_21781; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21783 = 10'h108 == _T_445[9:0] ? 4'h1 : _GEN_21782; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21784 = 10'h109 == _T_445[9:0] ? 4'h0 : _GEN_21783; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21785 = 10'h10a == _T_445[9:0] ? 4'h0 : _GEN_21784; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21786 = 10'h10b == _T_445[9:0] ? 4'h0 : _GEN_21785; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21787 = 10'h10c == _T_445[9:0] ? 4'h0 : _GEN_21786; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21788 = 10'h10d == _T_445[9:0] ? 4'h0 : _GEN_21787; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21789 = 10'h10e == _T_445[9:0] ? 4'h0 : _GEN_21788; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21790 = 10'h10f == _T_445[9:0] ? 4'h0 : _GEN_21789; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21791 = 10'h110 == _T_445[9:0] ? 4'h0 : _GEN_21790; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21792 = 10'h111 == _T_445[9:0] ? 4'h0 : _GEN_21791; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21793 = 10'h112 == _T_445[9:0] ? 4'h0 : _GEN_21792; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21794 = 10'h113 == _T_445[9:0] ? 4'h0 : _GEN_21793; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21795 = 10'h114 == _T_445[9:0] ? 4'h0 : _GEN_21794; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21796 = 10'h115 == _T_445[9:0] ? 4'h0 : _GEN_21795; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21797 = 10'h116 == _T_445[9:0] ? 4'h1 : _GEN_21796; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21798 = 10'h117 == _T_445[9:0] ? 4'h3 : _GEN_21797; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21799 = 10'h118 == _T_445[9:0] ? 4'h3 : _GEN_21798; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21800 = 10'h119 == _T_445[9:0] ? 4'h3 : _GEN_21799; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21801 = 10'h11a == _T_445[9:0] ? 4'h0 : _GEN_21800; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21802 = 10'h11b == _T_445[9:0] ? 4'h3 : _GEN_21801; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21803 = 10'h11c == _T_445[9:0] ? 4'h3 : _GEN_21802; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21804 = 10'h11d == _T_445[9:0] ? 4'h7 : _GEN_21803; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21805 = 10'h11e == _T_445[9:0] ? 4'ha : _GEN_21804; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21806 = 10'h11f == _T_445[9:0] ? 4'h0 : _GEN_21805; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21807 = 10'h120 == _T_445[9:0] ? 4'h3 : _GEN_21806; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21808 = 10'h121 == _T_445[9:0] ? 4'h3 : _GEN_21807; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21809 = 10'h122 == _T_445[9:0] ? 4'ha : _GEN_21808; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21810 = 10'h123 == _T_445[9:0] ? 4'h3 : _GEN_21809; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21811 = 10'h124 == _T_445[9:0] ? 4'h3 : _GEN_21810; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21812 = 10'h125 == _T_445[9:0] ? 4'h3 : _GEN_21811; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21813 = 10'h126 == _T_445[9:0] ? 4'h3 : _GEN_21812; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21814 = 10'h127 == _T_445[9:0] ? 4'h1 : _GEN_21813; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21815 = 10'h128 == _T_445[9:0] ? 4'h0 : _GEN_21814; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21816 = 10'h129 == _T_445[9:0] ? 4'h3 : _GEN_21815; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21817 = 10'h12a == _T_445[9:0] ? 4'h3 : _GEN_21816; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21818 = 10'h12b == _T_445[9:0] ? 4'h0 : _GEN_21817; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21819 = 10'h12c == _T_445[9:0] ? 4'h0 : _GEN_21818; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21820 = 10'h12d == _T_445[9:0] ? 4'h0 : _GEN_21819; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21821 = 10'h12e == _T_445[9:0] ? 4'h0 : _GEN_21820; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21822 = 10'h12f == _T_445[9:0] ? 4'h0 : _GEN_21821; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21823 = 10'h130 == _T_445[9:0] ? 4'h0 : _GEN_21822; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21824 = 10'h131 == _T_445[9:0] ? 4'h0 : _GEN_21823; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21825 = 10'h132 == _T_445[9:0] ? 4'h0 : _GEN_21824; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21826 = 10'h133 == _T_445[9:0] ? 4'h0 : _GEN_21825; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21827 = 10'h134 == _T_445[9:0] ? 4'h3 : _GEN_21826; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21828 = 10'h135 == _T_445[9:0] ? 4'h3 : _GEN_21827; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21829 = 10'h136 == _T_445[9:0] ? 4'h0 : _GEN_21828; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21830 = 10'h137 == _T_445[9:0] ? 4'h1 : _GEN_21829; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21831 = 10'h138 == _T_445[9:0] ? 4'h3 : _GEN_21830; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21832 = 10'h139 == _T_445[9:0] ? 4'h3 : _GEN_21831; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21833 = 10'h13a == _T_445[9:0] ? 4'h3 : _GEN_21832; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21834 = 10'h13b == _T_445[9:0] ? 4'h3 : _GEN_21833; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21835 = 10'h13c == _T_445[9:0] ? 4'h3 : _GEN_21834; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21836 = 10'h13d == _T_445[9:0] ? 4'h3 : _GEN_21835; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21837 = 10'h13e == _T_445[9:0] ? 4'ha : _GEN_21836; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21838 = 10'h13f == _T_445[9:0] ? 4'h0 : _GEN_21837; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21839 = 10'h140 == _T_445[9:0] ? 4'h5 : _GEN_21838; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21840 = 10'h141 == _T_445[9:0] ? 4'h3 : _GEN_21839; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21841 = 10'h142 == _T_445[9:0] ? 4'h7 : _GEN_21840; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21842 = 10'h143 == _T_445[9:0] ? 4'ha : _GEN_21841; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21843 = 10'h144 == _T_445[9:0] ? 4'h3 : _GEN_21842; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21844 = 10'h145 == _T_445[9:0] ? 4'h3 : _GEN_21843; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21845 = 10'h146 == _T_445[9:0] ? 4'h1 : _GEN_21844; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21846 = 10'h147 == _T_445[9:0] ? 4'h0 : _GEN_21845; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21847 = 10'h148 == _T_445[9:0] ? 4'h3 : _GEN_21846; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21848 = 10'h149 == _T_445[9:0] ? 4'h3 : _GEN_21847; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21849 = 10'h14a == _T_445[9:0] ? 4'h3 : _GEN_21848; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21850 = 10'h14b == _T_445[9:0] ? 4'h3 : _GEN_21849; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21851 = 10'h14c == _T_445[9:0] ? 4'h3 : _GEN_21850; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21852 = 10'h14d == _T_445[9:0] ? 4'h3 : _GEN_21851; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21853 = 10'h14e == _T_445[9:0] ? 4'h3 : _GEN_21852; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21854 = 10'h14f == _T_445[9:0] ? 4'h3 : _GEN_21853; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21855 = 10'h150 == _T_445[9:0] ? 4'h3 : _GEN_21854; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21856 = 10'h151 == _T_445[9:0] ? 4'h3 : _GEN_21855; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21857 = 10'h152 == _T_445[9:0] ? 4'h3 : _GEN_21856; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21858 = 10'h153 == _T_445[9:0] ? 4'h3 : _GEN_21857; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21859 = 10'h154 == _T_445[9:0] ? 4'h3 : _GEN_21858; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21860 = 10'h155 == _T_445[9:0] ? 4'h3 : _GEN_21859; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21861 = 10'h156 == _T_445[9:0] ? 4'h3 : _GEN_21860; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21862 = 10'h157 == _T_445[9:0] ? 4'h0 : _GEN_21861; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21863 = 10'h158 == _T_445[9:0] ? 4'h3 : _GEN_21862; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21864 = 10'h159 == _T_445[9:0] ? 4'h3 : _GEN_21863; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21865 = 10'h15a == _T_445[9:0] ? 4'h3 : _GEN_21864; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21866 = 10'h15b == _T_445[9:0] ? 4'h3 : _GEN_21865; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21867 = 10'h15c == _T_445[9:0] ? 4'h3 : _GEN_21866; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21868 = 10'h15d == _T_445[9:0] ? 4'ha : _GEN_21867; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21869 = 10'h15e == _T_445[9:0] ? 4'h7 : _GEN_21868; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21870 = 10'h15f == _T_445[9:0] ? 4'h0 : _GEN_21869; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21871 = 10'h160 == _T_445[9:0] ? 4'h3 : _GEN_21870; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21872 = 10'h161 == _T_445[9:0] ? 4'h3 : _GEN_21871; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21873 = 10'h162 == _T_445[9:0] ? 4'h3 : _GEN_21872; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21874 = 10'h163 == _T_445[9:0] ? 4'h7 : _GEN_21873; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21875 = 10'h164 == _T_445[9:0] ? 4'ha : _GEN_21874; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21876 = 10'h165 == _T_445[9:0] ? 4'h1 : _GEN_21875; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21877 = 10'h166 == _T_445[9:0] ? 4'h0 : _GEN_21876; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21878 = 10'h167 == _T_445[9:0] ? 4'h0 : _GEN_21877; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21879 = 10'h168 == _T_445[9:0] ? 4'hc : _GEN_21878; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21880 = 10'h169 == _T_445[9:0] ? 4'h9 : _GEN_21879; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21881 = 10'h16a == _T_445[9:0] ? 4'hc : _GEN_21880; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21882 = 10'h16b == _T_445[9:0] ? 4'hc : _GEN_21881; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21883 = 10'h16c == _T_445[9:0] ? 4'h3 : _GEN_21882; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21884 = 10'h16d == _T_445[9:0] ? 4'h3 : _GEN_21883; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21885 = 10'h16e == _T_445[9:0] ? 4'h3 : _GEN_21884; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21886 = 10'h16f == _T_445[9:0] ? 4'h3 : _GEN_21885; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21887 = 10'h170 == _T_445[9:0] ? 4'h5 : _GEN_21886; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21888 = 10'h171 == _T_445[9:0] ? 4'h3 : _GEN_21887; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21889 = 10'h172 == _T_445[9:0] ? 4'h3 : _GEN_21888; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21890 = 10'h173 == _T_445[9:0] ? 4'h3 : _GEN_21889; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21891 = 10'h174 == _T_445[9:0] ? 4'h3 : _GEN_21890; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21892 = 10'h175 == _T_445[9:0] ? 4'h3 : _GEN_21891; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21893 = 10'h176 == _T_445[9:0] ? 4'h0 : _GEN_21892; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21894 = 10'h177 == _T_445[9:0] ? 4'h0 : _GEN_21893; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21895 = 10'h178 == _T_445[9:0] ? 4'h1 : _GEN_21894; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21896 = 10'h179 == _T_445[9:0] ? 4'h3 : _GEN_21895; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21897 = 10'h17a == _T_445[9:0] ? 4'h5 : _GEN_21896; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21898 = 10'h17b == _T_445[9:0] ? 4'h3 : _GEN_21897; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21899 = 10'h17c == _T_445[9:0] ? 4'ha : _GEN_21898; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21900 = 10'h17d == _T_445[9:0] ? 4'h7 : _GEN_21899; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21901 = 10'h17e == _T_445[9:0] ? 4'h3 : _GEN_21900; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21902 = 10'h17f == _T_445[9:0] ? 4'h0 : _GEN_21901; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21903 = 10'h180 == _T_445[9:0] ? 4'hc : _GEN_21902; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21904 = 10'h181 == _T_445[9:0] ? 4'hc : _GEN_21903; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21905 = 10'h182 == _T_445[9:0] ? 4'hc : _GEN_21904; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21906 = 10'h183 == _T_445[9:0] ? 4'hc : _GEN_21905; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21907 = 10'h184 == _T_445[9:0] ? 4'ha : _GEN_21906; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21908 = 10'h185 == _T_445[9:0] ? 4'h1 : _GEN_21907; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21909 = 10'h186 == _T_445[9:0] ? 4'hc : _GEN_21908; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21910 = 10'h187 == _T_445[9:0] ? 4'h0 : _GEN_21909; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21911 = 10'h188 == _T_445[9:0] ? 4'hc : _GEN_21910; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21912 = 10'h189 == _T_445[9:0] ? 4'hc : _GEN_21911; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21913 = 10'h18a == _T_445[9:0] ? 4'hc : _GEN_21912; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21914 = 10'h18b == _T_445[9:0] ? 4'hc : _GEN_21913; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21915 = 10'h18c == _T_445[9:0] ? 4'hc : _GEN_21914; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21916 = 10'h18d == _T_445[9:0] ? 4'hc : _GEN_21915; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21917 = 10'h18e == _T_445[9:0] ? 4'hc : _GEN_21916; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21918 = 10'h18f == _T_445[9:0] ? 4'hc : _GEN_21917; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21919 = 10'h190 == _T_445[9:0] ? 4'hc : _GEN_21918; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21920 = 10'h191 == _T_445[9:0] ? 4'hc : _GEN_21919; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21921 = 10'h192 == _T_445[9:0] ? 4'h9 : _GEN_21920; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21922 = 10'h193 == _T_445[9:0] ? 4'hc : _GEN_21921; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21923 = 10'h194 == _T_445[9:0] ? 4'hc : _GEN_21922; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21924 = 10'h195 == _T_445[9:0] ? 4'hc : _GEN_21923; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21925 = 10'h196 == _T_445[9:0] ? 4'h0 : _GEN_21924; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21926 = 10'h197 == _T_445[9:0] ? 4'h3 : _GEN_21925; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21927 = 10'h198 == _T_445[9:0] ? 4'h1 : _GEN_21926; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21928 = 10'h199 == _T_445[9:0] ? 4'h3 : _GEN_21927; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21929 = 10'h19a == _T_445[9:0] ? 4'h3 : _GEN_21928; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21930 = 10'h19b == _T_445[9:0] ? 4'h3 : _GEN_21929; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21931 = 10'h19c == _T_445[9:0] ? 4'ha : _GEN_21930; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21932 = 10'h19d == _T_445[9:0] ? 4'h3 : _GEN_21931; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21933 = 10'h19e == _T_445[9:0] ? 4'h3 : _GEN_21932; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21934 = 10'h19f == _T_445[9:0] ? 4'h0 : _GEN_21933; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21935 = 10'h1a0 == _T_445[9:0] ? 4'hc : _GEN_21934; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21936 = 10'h1a1 == _T_445[9:0] ? 4'hc : _GEN_21935; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21937 = 10'h1a2 == _T_445[9:0] ? 4'h9 : _GEN_21936; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21938 = 10'h1a3 == _T_445[9:0] ? 4'hc : _GEN_21937; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21939 = 10'h1a4 == _T_445[9:0] ? 4'ha : _GEN_21938; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21940 = 10'h1a5 == _T_445[9:0] ? 4'h0 : _GEN_21939; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21941 = 10'h1a6 == _T_445[9:0] ? 4'hc : _GEN_21940; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21942 = 10'h1a7 == _T_445[9:0] ? 4'h0 : _GEN_21941; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21943 = 10'h1a8 == _T_445[9:0] ? 4'hc : _GEN_21942; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21944 = 10'h1a9 == _T_445[9:0] ? 4'hc : _GEN_21943; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21945 = 10'h1aa == _T_445[9:0] ? 4'hc : _GEN_21944; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21946 = 10'h1ab == _T_445[9:0] ? 4'h9 : _GEN_21945; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21947 = 10'h1ac == _T_445[9:0] ? 4'hc : _GEN_21946; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21948 = 10'h1ad == _T_445[9:0] ? 4'hc : _GEN_21947; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21949 = 10'h1ae == _T_445[9:0] ? 4'hc : _GEN_21948; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21950 = 10'h1af == _T_445[9:0] ? 4'hc : _GEN_21949; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21951 = 10'h1b0 == _T_445[9:0] ? 4'hc : _GEN_21950; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21952 = 10'h1b1 == _T_445[9:0] ? 4'hc : _GEN_21951; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21953 = 10'h1b2 == _T_445[9:0] ? 4'hc : _GEN_21952; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21954 = 10'h1b3 == _T_445[9:0] ? 4'hc : _GEN_21953; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21955 = 10'h1b4 == _T_445[9:0] ? 4'hc : _GEN_21954; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21956 = 10'h1b5 == _T_445[9:0] ? 4'hc : _GEN_21955; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21957 = 10'h1b6 == _T_445[9:0] ? 4'h0 : _GEN_21956; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21958 = 10'h1b7 == _T_445[9:0] ? 4'hc : _GEN_21957; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21959 = 10'h1b8 == _T_445[9:0] ? 4'h0 : _GEN_21958; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21960 = 10'h1b9 == _T_445[9:0] ? 4'hc : _GEN_21959; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21961 = 10'h1ba == _T_445[9:0] ? 4'hc : _GEN_21960; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21962 = 10'h1bb == _T_445[9:0] ? 4'hc : _GEN_21961; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21963 = 10'h1bc == _T_445[9:0] ? 4'h7 : _GEN_21962; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21964 = 10'h1bd == _T_445[9:0] ? 4'ha : _GEN_21963; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21965 = 10'h1be == _T_445[9:0] ? 4'hc : _GEN_21964; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21966 = 10'h1bf == _T_445[9:0] ? 4'h0 : _GEN_21965; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21967 = 10'h1c0 == _T_445[9:0] ? 4'hc : _GEN_21966; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21968 = 10'h1c1 == _T_445[9:0] ? 4'hc : _GEN_21967; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21969 = 10'h1c2 == _T_445[9:0] ? 4'hc : _GEN_21968; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21970 = 10'h1c3 == _T_445[9:0] ? 4'h7 : _GEN_21969; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21971 = 10'h1c4 == _T_445[9:0] ? 4'h7 : _GEN_21970; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21972 = 10'h1c5 == _T_445[9:0] ? 4'hc : _GEN_21971; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21973 = 10'h1c6 == _T_445[9:0] ? 4'hc : _GEN_21972; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21974 = 10'h1c7 == _T_445[9:0] ? 4'hc : _GEN_21973; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21975 = 10'h1c8 == _T_445[9:0] ? 4'hc : _GEN_21974; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21976 = 10'h1c9 == _T_445[9:0] ? 4'hc : _GEN_21975; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21977 = 10'h1ca == _T_445[9:0] ? 4'hc : _GEN_21976; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21978 = 10'h1cb == _T_445[9:0] ? 4'hc : _GEN_21977; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21979 = 10'h1cc == _T_445[9:0] ? 4'hc : _GEN_21978; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21980 = 10'h1cd == _T_445[9:0] ? 4'hc : _GEN_21979; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21981 = 10'h1ce == _T_445[9:0] ? 4'hc : _GEN_21980; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21982 = 10'h1cf == _T_445[9:0] ? 4'hc : _GEN_21981; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21983 = 10'h1d0 == _T_445[9:0] ? 4'hc : _GEN_21982; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21984 = 10'h1d1 == _T_445[9:0] ? 4'hc : _GEN_21983; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21985 = 10'h1d2 == _T_445[9:0] ? 4'hc : _GEN_21984; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21986 = 10'h1d3 == _T_445[9:0] ? 4'hc : _GEN_21985; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21987 = 10'h1d4 == _T_445[9:0] ? 4'hc : _GEN_21986; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21988 = 10'h1d5 == _T_445[9:0] ? 4'hc : _GEN_21987; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21989 = 10'h1d6 == _T_445[9:0] ? 4'hc : _GEN_21988; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21990 = 10'h1d7 == _T_445[9:0] ? 4'hc : _GEN_21989; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21991 = 10'h1d8 == _T_445[9:0] ? 4'hc : _GEN_21990; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21992 = 10'h1d9 == _T_445[9:0] ? 4'hc : _GEN_21991; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21993 = 10'h1da == _T_445[9:0] ? 4'hc : _GEN_21992; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21994 = 10'h1db == _T_445[9:0] ? 4'hc : _GEN_21993; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21995 = 10'h1dc == _T_445[9:0] ? 4'hc : _GEN_21994; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21996 = 10'h1dd == _T_445[9:0] ? 4'ha : _GEN_21995; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21997 = 10'h1de == _T_445[9:0] ? 4'hc : _GEN_21996; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21998 = 10'h1df == _T_445[9:0] ? 4'h0 : _GEN_21997; // @[Filter.scala 191:102]
  wire [3:0] _GEN_21999 = 10'h1e0 == _T_445[9:0] ? 4'h9 : _GEN_21998; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22000 = 10'h1e1 == _T_445[9:0] ? 4'hc : _GEN_21999; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22001 = 10'h1e2 == _T_445[9:0] ? 4'h7 : _GEN_22000; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22002 = 10'h1e3 == _T_445[9:0] ? 4'h7 : _GEN_22001; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22003 = 10'h1e4 == _T_445[9:0] ? 4'hc : _GEN_22002; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22004 = 10'h1e5 == _T_445[9:0] ? 4'hc : _GEN_22003; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22005 = 10'h1e6 == _T_445[9:0] ? 4'hc : _GEN_22004; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22006 = 10'h1e7 == _T_445[9:0] ? 4'hc : _GEN_22005; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22007 = 10'h1e8 == _T_445[9:0] ? 4'hc : _GEN_22006; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22008 = 10'h1e9 == _T_445[9:0] ? 4'hc : _GEN_22007; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22009 = 10'h1ea == _T_445[9:0] ? 4'hc : _GEN_22008; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22010 = 10'h1eb == _T_445[9:0] ? 4'hc : _GEN_22009; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22011 = 10'h1ec == _T_445[9:0] ? 4'hc : _GEN_22010; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22012 = 10'h1ed == _T_445[9:0] ? 4'hc : _GEN_22011; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22013 = 10'h1ee == _T_445[9:0] ? 4'hc : _GEN_22012; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22014 = 10'h1ef == _T_445[9:0] ? 4'hc : _GEN_22013; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22015 = 10'h1f0 == _T_445[9:0] ? 4'hc : _GEN_22014; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22016 = 10'h1f1 == _T_445[9:0] ? 4'hc : _GEN_22015; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22017 = 10'h1f2 == _T_445[9:0] ? 4'hc : _GEN_22016; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22018 = 10'h1f3 == _T_445[9:0] ? 4'hc : _GEN_22017; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22019 = 10'h1f4 == _T_445[9:0] ? 4'hc : _GEN_22018; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22020 = 10'h1f5 == _T_445[9:0] ? 4'hc : _GEN_22019; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22021 = 10'h1f6 == _T_445[9:0] ? 4'hc : _GEN_22020; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22022 = 10'h1f7 == _T_445[9:0] ? 4'hc : _GEN_22021; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22023 = 10'h1f8 == _T_445[9:0] ? 4'hc : _GEN_22022; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22024 = 10'h1f9 == _T_445[9:0] ? 4'hc : _GEN_22023; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22025 = 10'h1fa == _T_445[9:0] ? 4'h9 : _GEN_22024; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22026 = 10'h1fb == _T_445[9:0] ? 4'hc : _GEN_22025; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22027 = 10'h1fc == _T_445[9:0] ? 4'hc : _GEN_22026; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22028 = 10'h1fd == _T_445[9:0] ? 4'h7 : _GEN_22027; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22029 = 10'h1fe == _T_445[9:0] ? 4'hc : _GEN_22028; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22030 = 10'h1ff == _T_445[9:0] ? 4'h0 : _GEN_22029; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22031 = 10'h200 == _T_445[9:0] ? 4'hc : _GEN_22030; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22032 = 10'h201 == _T_445[9:0] ? 4'hc : _GEN_22031; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22033 = 10'h202 == _T_445[9:0] ? 4'ha : _GEN_22032; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22034 = 10'h203 == _T_445[9:0] ? 4'hc : _GEN_22033; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22035 = 10'h204 == _T_445[9:0] ? 4'hc : _GEN_22034; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22036 = 10'h205 == _T_445[9:0] ? 4'hc : _GEN_22035; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22037 = 10'h206 == _T_445[9:0] ? 4'hc : _GEN_22036; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22038 = 10'h207 == _T_445[9:0] ? 4'hc : _GEN_22037; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22039 = 10'h208 == _T_445[9:0] ? 4'hc : _GEN_22038; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22040 = 10'h209 == _T_445[9:0] ? 4'hc : _GEN_22039; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22041 = 10'h20a == _T_445[9:0] ? 4'hc : _GEN_22040; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22042 = 10'h20b == _T_445[9:0] ? 4'hc : _GEN_22041; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22043 = 10'h20c == _T_445[9:0] ? 4'hc : _GEN_22042; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22044 = 10'h20d == _T_445[9:0] ? 4'hc : _GEN_22043; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22045 = 10'h20e == _T_445[9:0] ? 4'hc : _GEN_22044; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22046 = 10'h20f == _T_445[9:0] ? 4'hc : _GEN_22045; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22047 = 10'h210 == _T_445[9:0] ? 4'hc : _GEN_22046; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22048 = 10'h211 == _T_445[9:0] ? 4'hc : _GEN_22047; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22049 = 10'h212 == _T_445[9:0] ? 4'hc : _GEN_22048; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22050 = 10'h213 == _T_445[9:0] ? 4'hc : _GEN_22049; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22051 = 10'h214 == _T_445[9:0] ? 4'hc : _GEN_22050; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22052 = 10'h215 == _T_445[9:0] ? 4'hc : _GEN_22051; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22053 = 10'h216 == _T_445[9:0] ? 4'hc : _GEN_22052; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22054 = 10'h217 == _T_445[9:0] ? 4'hc : _GEN_22053; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22055 = 10'h218 == _T_445[9:0] ? 4'hc : _GEN_22054; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22056 = 10'h219 == _T_445[9:0] ? 4'hc : _GEN_22055; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22057 = 10'h21a == _T_445[9:0] ? 4'hc : _GEN_22056; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22058 = 10'h21b == _T_445[9:0] ? 4'hc : _GEN_22057; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22059 = 10'h21c == _T_445[9:0] ? 4'ha : _GEN_22058; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22060 = 10'h21d == _T_445[9:0] ? 4'h7 : _GEN_22059; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22061 = 10'h21e == _T_445[9:0] ? 4'hc : _GEN_22060; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22062 = 10'h21f == _T_445[9:0] ? 4'h0 : _GEN_22061; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22063 = 10'h220 == _T_445[9:0] ? 4'h0 : _GEN_22062; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22064 = 10'h221 == _T_445[9:0] ? 4'h0 : _GEN_22063; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22065 = 10'h222 == _T_445[9:0] ? 4'h0 : _GEN_22064; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22066 = 10'h223 == _T_445[9:0] ? 4'h0 : _GEN_22065; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22067 = 10'h224 == _T_445[9:0] ? 4'h0 : _GEN_22066; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22068 = 10'h225 == _T_445[9:0] ? 4'h0 : _GEN_22067; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22069 = 10'h226 == _T_445[9:0] ? 4'h0 : _GEN_22068; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22070 = 10'h227 == _T_445[9:0] ? 4'h0 : _GEN_22069; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22071 = 10'h228 == _T_445[9:0] ? 4'h0 : _GEN_22070; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22072 = 10'h229 == _T_445[9:0] ? 4'h0 : _GEN_22071; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22073 = 10'h22a == _T_445[9:0] ? 4'h0 : _GEN_22072; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22074 = 10'h22b == _T_445[9:0] ? 4'h0 : _GEN_22073; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22075 = 10'h22c == _T_445[9:0] ? 4'h0 : _GEN_22074; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22076 = 10'h22d == _T_445[9:0] ? 4'h0 : _GEN_22075; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22077 = 10'h22e == _T_445[9:0] ? 4'h0 : _GEN_22076; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22078 = 10'h22f == _T_445[9:0] ? 4'h0 : _GEN_22077; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22079 = 10'h230 == _T_445[9:0] ? 4'h0 : _GEN_22078; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22080 = 10'h231 == _T_445[9:0] ? 4'h0 : _GEN_22079; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22081 = 10'h232 == _T_445[9:0] ? 4'h0 : _GEN_22080; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22082 = 10'h233 == _T_445[9:0] ? 4'h0 : _GEN_22081; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22083 = 10'h234 == _T_445[9:0] ? 4'h0 : _GEN_22082; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22084 = 10'h235 == _T_445[9:0] ? 4'h0 : _GEN_22083; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22085 = 10'h236 == _T_445[9:0] ? 4'h0 : _GEN_22084; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22086 = 10'h237 == _T_445[9:0] ? 4'h0 : _GEN_22085; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22087 = 10'h238 == _T_445[9:0] ? 4'h0 : _GEN_22086; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22088 = 10'h239 == _T_445[9:0] ? 4'h0 : _GEN_22087; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22089 = 10'h23a == _T_445[9:0] ? 4'h0 : _GEN_22088; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22090 = 10'h23b == _T_445[9:0] ? 4'h0 : _GEN_22089; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22091 = 10'h23c == _T_445[9:0] ? 4'h0 : _GEN_22090; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22092 = 10'h23d == _T_445[9:0] ? 4'h0 : _GEN_22091; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22093 = 10'h23e == _T_445[9:0] ? 4'h0 : _GEN_22092; // @[Filter.scala 191:102]
  wire [3:0] _GEN_22094 = 10'h23f == _T_445[9:0] ? 4'h0 : _GEN_22093; // @[Filter.scala 191:102]
  wire [6:0] _GEN_28372 = {{3'd0}, _GEN_22094}; // @[Filter.scala 191:102]
  wire [10:0] _T_452 = _GEN_28372 * 7'h46; // @[Filter.scala 191:102]
  wire [10:0] _GEN_28373 = {{2'd0}, _T_447}; // @[Filter.scala 191:69]
  wire [10:0] _T_454 = _GEN_28373 + _T_452; // @[Filter.scala 191:69]
  wire [3:0] _GEN_22126 = 10'h1f == _T_445[9:0] ? 4'h0 : 4'h3; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22127 = 10'h20 == _T_445[9:0] ? 4'h3 : _GEN_22126; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22128 = 10'h21 == _T_445[9:0] ? 4'h3 : _GEN_22127; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22129 = 10'h22 == _T_445[9:0] ? 4'h3 : _GEN_22128; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22130 = 10'h23 == _T_445[9:0] ? 4'h3 : _GEN_22129; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22131 = 10'h24 == _T_445[9:0] ? 4'h3 : _GEN_22130; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22132 = 10'h25 == _T_445[9:0] ? 4'h3 : _GEN_22131; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22133 = 10'h26 == _T_445[9:0] ? 4'h3 : _GEN_22132; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22134 = 10'h27 == _T_445[9:0] ? 4'h9 : _GEN_22133; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22135 = 10'h28 == _T_445[9:0] ? 4'h9 : _GEN_22134; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22136 = 10'h29 == _T_445[9:0] ? 4'h3 : _GEN_22135; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22137 = 10'h2a == _T_445[9:0] ? 4'h3 : _GEN_22136; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22138 = 10'h2b == _T_445[9:0] ? 4'h3 : _GEN_22137; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22139 = 10'h2c == _T_445[9:0] ? 4'h3 : _GEN_22138; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22140 = 10'h2d == _T_445[9:0] ? 4'h3 : _GEN_22139; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22141 = 10'h2e == _T_445[9:0] ? 4'h3 : _GEN_22140; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22142 = 10'h2f == _T_445[9:0] ? 4'h3 : _GEN_22141; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22143 = 10'h30 == _T_445[9:0] ? 4'h3 : _GEN_22142; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22144 = 10'h31 == _T_445[9:0] ? 4'h3 : _GEN_22143; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22145 = 10'h32 == _T_445[9:0] ? 4'h3 : _GEN_22144; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22146 = 10'h33 == _T_445[9:0] ? 4'h3 : _GEN_22145; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22147 = 10'h34 == _T_445[9:0] ? 4'h3 : _GEN_22146; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22148 = 10'h35 == _T_445[9:0] ? 4'h3 : _GEN_22147; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22149 = 10'h36 == _T_445[9:0] ? 4'h3 : _GEN_22148; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22150 = 10'h37 == _T_445[9:0] ? 4'h9 : _GEN_22149; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22151 = 10'h38 == _T_445[9:0] ? 4'h9 : _GEN_22150; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22152 = 10'h39 == _T_445[9:0] ? 4'h3 : _GEN_22151; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22153 = 10'h3a == _T_445[9:0] ? 4'h3 : _GEN_22152; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22154 = 10'h3b == _T_445[9:0] ? 4'h3 : _GEN_22153; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22155 = 10'h3c == _T_445[9:0] ? 4'h3 : _GEN_22154; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22156 = 10'h3d == _T_445[9:0] ? 4'h3 : _GEN_22155; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22157 = 10'h3e == _T_445[9:0] ? 4'h3 : _GEN_22156; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22158 = 10'h3f == _T_445[9:0] ? 4'h0 : _GEN_22157; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22159 = 10'h40 == _T_445[9:0] ? 4'h3 : _GEN_22158; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22160 = 10'h41 == _T_445[9:0] ? 4'h3 : _GEN_22159; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22161 = 10'h42 == _T_445[9:0] ? 4'h3 : _GEN_22160; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22162 = 10'h43 == _T_445[9:0] ? 4'h2 : _GEN_22161; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22163 = 10'h44 == _T_445[9:0] ? 4'h3 : _GEN_22162; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22164 = 10'h45 == _T_445[9:0] ? 4'hf : _GEN_22163; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22165 = 10'h46 == _T_445[9:0] ? 4'hf : _GEN_22164; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22166 = 10'h47 == _T_445[9:0] ? 4'hf : _GEN_22165; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22167 = 10'h48 == _T_445[9:0] ? 4'hf : _GEN_22166; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22168 = 10'h49 == _T_445[9:0] ? 4'h3 : _GEN_22167; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22169 = 10'h4a == _T_445[9:0] ? 4'h3 : _GEN_22168; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22170 = 10'h4b == _T_445[9:0] ? 4'h3 : _GEN_22169; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22171 = 10'h4c == _T_445[9:0] ? 4'h3 : _GEN_22170; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22172 = 10'h4d == _T_445[9:0] ? 4'h3 : _GEN_22171; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22173 = 10'h4e == _T_445[9:0] ? 4'h3 : _GEN_22172; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22174 = 10'h4f == _T_445[9:0] ? 4'h3 : _GEN_22173; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22175 = 10'h50 == _T_445[9:0] ? 4'h3 : _GEN_22174; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22176 = 10'h51 == _T_445[9:0] ? 4'h3 : _GEN_22175; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22177 = 10'h52 == _T_445[9:0] ? 4'h3 : _GEN_22176; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22178 = 10'h53 == _T_445[9:0] ? 4'h3 : _GEN_22177; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22179 = 10'h54 == _T_445[9:0] ? 4'h9 : _GEN_22178; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22180 = 10'h55 == _T_445[9:0] ? 4'h9 : _GEN_22179; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22181 = 10'h56 == _T_445[9:0] ? 4'h9 : _GEN_22180; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22182 = 10'h57 == _T_445[9:0] ? 4'hf : _GEN_22181; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22183 = 10'h58 == _T_445[9:0] ? 4'h3 : _GEN_22182; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22184 = 10'h59 == _T_445[9:0] ? 4'hf : _GEN_22183; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22185 = 10'h5a == _T_445[9:0] ? 4'h3 : _GEN_22184; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22186 = 10'h5b == _T_445[9:0] ? 4'h3 : _GEN_22185; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22187 = 10'h5c == _T_445[9:0] ? 4'h3 : _GEN_22186; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22188 = 10'h5d == _T_445[9:0] ? 4'h3 : _GEN_22187; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22189 = 10'h5e == _T_445[9:0] ? 4'h3 : _GEN_22188; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22190 = 10'h5f == _T_445[9:0] ? 4'h0 : _GEN_22189; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22191 = 10'h60 == _T_445[9:0] ? 4'h3 : _GEN_22190; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22192 = 10'h61 == _T_445[9:0] ? 4'h3 : _GEN_22191; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22193 = 10'h62 == _T_445[9:0] ? 4'h3 : _GEN_22192; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22194 = 10'h63 == _T_445[9:0] ? 4'h3 : _GEN_22193; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22195 = 10'h64 == _T_445[9:0] ? 4'h3 : _GEN_22194; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22196 = 10'h65 == _T_445[9:0] ? 4'hf : _GEN_22195; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22197 = 10'h66 == _T_445[9:0] ? 4'h3 : _GEN_22196; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22198 = 10'h67 == _T_445[9:0] ? 4'h3 : _GEN_22197; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22199 = 10'h68 == _T_445[9:0] ? 4'h3 : _GEN_22198; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22200 = 10'h69 == _T_445[9:0] ? 4'hf : _GEN_22199; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22201 = 10'h6a == _T_445[9:0] ? 4'h9 : _GEN_22200; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22202 = 10'h6b == _T_445[9:0] ? 4'h9 : _GEN_22201; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22203 = 10'h6c == _T_445[9:0] ? 4'h3 : _GEN_22202; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22204 = 10'h6d == _T_445[9:0] ? 4'h3 : _GEN_22203; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22205 = 10'h6e == _T_445[9:0] ? 4'h3 : _GEN_22204; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22206 = 10'h6f == _T_445[9:0] ? 4'h3 : _GEN_22205; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22207 = 10'h70 == _T_445[9:0] ? 4'h3 : _GEN_22206; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22208 = 10'h71 == _T_445[9:0] ? 4'h3 : _GEN_22207; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22209 = 10'h72 == _T_445[9:0] ? 4'h3 : _GEN_22208; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22210 = 10'h73 == _T_445[9:0] ? 4'h9 : _GEN_22209; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22211 = 10'h74 == _T_445[9:0] ? 4'hf : _GEN_22210; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22212 = 10'h75 == _T_445[9:0] ? 4'hf : _GEN_22211; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22213 = 10'h76 == _T_445[9:0] ? 4'hf : _GEN_22212; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22214 = 10'h77 == _T_445[9:0] ? 4'h3 : _GEN_22213; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22215 = 10'h78 == _T_445[9:0] ? 4'h3 : _GEN_22214; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22216 = 10'h79 == _T_445[9:0] ? 4'h3 : _GEN_22215; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22217 = 10'h7a == _T_445[9:0] ? 4'hf : _GEN_22216; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22218 = 10'h7b == _T_445[9:0] ? 4'h3 : _GEN_22217; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22219 = 10'h7c == _T_445[9:0] ? 4'h3 : _GEN_22218; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22220 = 10'h7d == _T_445[9:0] ? 4'h2 : _GEN_22219; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22221 = 10'h7e == _T_445[9:0] ? 4'h3 : _GEN_22220; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22222 = 10'h7f == _T_445[9:0] ? 4'h0 : _GEN_22221; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22223 = 10'h80 == _T_445[9:0] ? 4'h3 : _GEN_22222; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22224 = 10'h81 == _T_445[9:0] ? 4'h3 : _GEN_22223; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22225 = 10'h82 == _T_445[9:0] ? 4'h9 : _GEN_22224; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22226 = 10'h83 == _T_445[9:0] ? 4'hf : _GEN_22225; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22227 = 10'h84 == _T_445[9:0] ? 4'h2 : _GEN_22226; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22228 = 10'h85 == _T_445[9:0] ? 4'h9 : _GEN_22227; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22229 = 10'h86 == _T_445[9:0] ? 4'h9 : _GEN_22228; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22230 = 10'h87 == _T_445[9:0] ? 4'h3 : _GEN_22229; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22231 = 10'h88 == _T_445[9:0] ? 4'h3 : _GEN_22230; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22232 = 10'h89 == _T_445[9:0] ? 4'hf : _GEN_22231; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22233 = 10'h8a == _T_445[9:0] ? 4'hf : _GEN_22232; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22234 = 10'h8b == _T_445[9:0] ? 4'h9 : _GEN_22233; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22235 = 10'h8c == _T_445[9:0] ? 4'h9 : _GEN_22234; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22236 = 10'h8d == _T_445[9:0] ? 4'h9 : _GEN_22235; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22237 = 10'h8e == _T_445[9:0] ? 4'h9 : _GEN_22236; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22238 = 10'h8f == _T_445[9:0] ? 4'h9 : _GEN_22237; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22239 = 10'h90 == _T_445[9:0] ? 4'h9 : _GEN_22238; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22240 = 10'h91 == _T_445[9:0] ? 4'h9 : _GEN_22239; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22241 = 10'h92 == _T_445[9:0] ? 4'h9 : _GEN_22240; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22242 = 10'h93 == _T_445[9:0] ? 4'hf : _GEN_22241; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22243 = 10'h94 == _T_445[9:0] ? 4'hf : _GEN_22242; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22244 = 10'h95 == _T_445[9:0] ? 4'h3 : _GEN_22243; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22245 = 10'h96 == _T_445[9:0] ? 4'h3 : _GEN_22244; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22246 = 10'h97 == _T_445[9:0] ? 4'h3 : _GEN_22245; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22247 = 10'h98 == _T_445[9:0] ? 4'h9 : _GEN_22246; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22248 = 10'h99 == _T_445[9:0] ? 4'hf : _GEN_22247; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22249 = 10'h9a == _T_445[9:0] ? 4'h9 : _GEN_22248; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22250 = 10'h9b == _T_445[9:0] ? 4'h9 : _GEN_22249; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22251 = 10'h9c == _T_445[9:0] ? 4'h3 : _GEN_22250; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22252 = 10'h9d == _T_445[9:0] ? 4'h3 : _GEN_22251; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22253 = 10'h9e == _T_445[9:0] ? 4'h3 : _GEN_22252; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22254 = 10'h9f == _T_445[9:0] ? 4'h0 : _GEN_22253; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22255 = 10'ha0 == _T_445[9:0] ? 4'h3 : _GEN_22254; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22256 = 10'ha1 == _T_445[9:0] ? 4'h9 : _GEN_22255; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22257 = 10'ha2 == _T_445[9:0] ? 4'hf : _GEN_22256; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22258 = 10'ha3 == _T_445[9:0] ? 4'h3 : _GEN_22257; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22259 = 10'ha4 == _T_445[9:0] ? 4'h3 : _GEN_22258; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22260 = 10'ha5 == _T_445[9:0] ? 4'h3 : _GEN_22259; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22261 = 10'ha6 == _T_445[9:0] ? 4'h3 : _GEN_22260; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22262 = 10'ha7 == _T_445[9:0] ? 4'hf : _GEN_22261; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22263 = 10'ha8 == _T_445[9:0] ? 4'h3 : _GEN_22262; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22264 = 10'ha9 == _T_445[9:0] ? 4'h9 : _GEN_22263; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22265 = 10'haa == _T_445[9:0] ? 4'hf : _GEN_22264; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22266 = 10'hab == _T_445[9:0] ? 4'hf : _GEN_22265; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22267 = 10'hac == _T_445[9:0] ? 4'hf : _GEN_22266; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22268 = 10'had == _T_445[9:0] ? 4'hf : _GEN_22267; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22269 = 10'hae == _T_445[9:0] ? 4'hf : _GEN_22268; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22270 = 10'haf == _T_445[9:0] ? 4'hf : _GEN_22269; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22271 = 10'hb0 == _T_445[9:0] ? 4'hf : _GEN_22270; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22272 = 10'hb1 == _T_445[9:0] ? 4'hf : _GEN_22271; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22273 = 10'hb2 == _T_445[9:0] ? 4'hf : _GEN_22272; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22274 = 10'hb3 == _T_445[9:0] ? 4'hf : _GEN_22273; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22275 = 10'hb4 == _T_445[9:0] ? 4'h9 : _GEN_22274; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22276 = 10'hb5 == _T_445[9:0] ? 4'h9 : _GEN_22275; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22277 = 10'hb6 == _T_445[9:0] ? 4'h3 : _GEN_22276; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22278 = 10'hb7 == _T_445[9:0] ? 4'hf : _GEN_22277; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22279 = 10'hb8 == _T_445[9:0] ? 4'h3 : _GEN_22278; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22280 = 10'hb9 == _T_445[9:0] ? 4'h3 : _GEN_22279; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22281 = 10'hba == _T_445[9:0] ? 4'h3 : _GEN_22280; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22282 = 10'hbb == _T_445[9:0] ? 4'hf : _GEN_22281; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22283 = 10'hbc == _T_445[9:0] ? 4'h3 : _GEN_22282; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22284 = 10'hbd == _T_445[9:0] ? 4'h3 : _GEN_22283; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22285 = 10'hbe == _T_445[9:0] ? 4'h3 : _GEN_22284; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22286 = 10'hbf == _T_445[9:0] ? 4'h0 : _GEN_22285; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22287 = 10'hc0 == _T_445[9:0] ? 4'h3 : _GEN_22286; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22288 = 10'hc1 == _T_445[9:0] ? 4'h3 : _GEN_22287; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22289 = 10'hc2 == _T_445[9:0] ? 4'h3 : _GEN_22288; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22290 = 10'hc3 == _T_445[9:0] ? 4'h2 : _GEN_22289; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22291 = 10'hc4 == _T_445[9:0] ? 4'hf : _GEN_22290; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22292 = 10'hc5 == _T_445[9:0] ? 4'hf : _GEN_22291; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22293 = 10'hc6 == _T_445[9:0] ? 4'hf : _GEN_22292; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22294 = 10'hc7 == _T_445[9:0] ? 4'h3 : _GEN_22293; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22295 = 10'hc8 == _T_445[9:0] ? 4'h9 : _GEN_22294; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22296 = 10'hc9 == _T_445[9:0] ? 4'hf : _GEN_22295; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22297 = 10'hca == _T_445[9:0] ? 4'hf : _GEN_22296; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22298 = 10'hcb == _T_445[9:0] ? 4'hf : _GEN_22297; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22299 = 10'hcc == _T_445[9:0] ? 4'hf : _GEN_22298; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22300 = 10'hcd == _T_445[9:0] ? 4'hf : _GEN_22299; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22301 = 10'hce == _T_445[9:0] ? 4'hf : _GEN_22300; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22302 = 10'hcf == _T_445[9:0] ? 4'hf : _GEN_22301; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22303 = 10'hd0 == _T_445[9:0] ? 4'hf : _GEN_22302; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22304 = 10'hd1 == _T_445[9:0] ? 4'hf : _GEN_22303; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22305 = 10'hd2 == _T_445[9:0] ? 4'hf : _GEN_22304; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22306 = 10'hd3 == _T_445[9:0] ? 4'hf : _GEN_22305; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22307 = 10'hd4 == _T_445[9:0] ? 4'hf : _GEN_22306; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22308 = 10'hd5 == _T_445[9:0] ? 4'hf : _GEN_22307; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22309 = 10'hd6 == _T_445[9:0] ? 4'h9 : _GEN_22308; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22310 = 10'hd7 == _T_445[9:0] ? 4'h3 : _GEN_22309; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22311 = 10'hd8 == _T_445[9:0] ? 4'hf : _GEN_22310; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22312 = 10'hd9 == _T_445[9:0] ? 4'h3 : _GEN_22311; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22313 = 10'hda == _T_445[9:0] ? 4'h3 : _GEN_22312; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22314 = 10'hdb == _T_445[9:0] ? 4'h3 : _GEN_22313; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22315 = 10'hdc == _T_445[9:0] ? 4'h3 : _GEN_22314; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22316 = 10'hdd == _T_445[9:0] ? 4'h3 : _GEN_22315; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22317 = 10'hde == _T_445[9:0] ? 4'h2 : _GEN_22316; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22318 = 10'hdf == _T_445[9:0] ? 4'h0 : _GEN_22317; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22319 = 10'he0 == _T_445[9:0] ? 4'h3 : _GEN_22318; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22320 = 10'he1 == _T_445[9:0] ? 4'h3 : _GEN_22319; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22321 = 10'he2 == _T_445[9:0] ? 4'h3 : _GEN_22320; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22322 = 10'he3 == _T_445[9:0] ? 4'h3 : _GEN_22321; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22323 = 10'he4 == _T_445[9:0] ? 4'h3 : _GEN_22322; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22324 = 10'he5 == _T_445[9:0] ? 4'h3 : _GEN_22323; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22325 = 10'he6 == _T_445[9:0] ? 4'h3 : _GEN_22324; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22326 = 10'he7 == _T_445[9:0] ? 4'h9 : _GEN_22325; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22327 = 10'he8 == _T_445[9:0] ? 4'h9 : _GEN_22326; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22328 = 10'he9 == _T_445[9:0] ? 4'h9 : _GEN_22327; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22329 = 10'hea == _T_445[9:0] ? 4'hf : _GEN_22328; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22330 = 10'heb == _T_445[9:0] ? 4'hf : _GEN_22329; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22331 = 10'hec == _T_445[9:0] ? 4'hf : _GEN_22330; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22332 = 10'hed == _T_445[9:0] ? 4'hf : _GEN_22331; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22333 = 10'hee == _T_445[9:0] ? 4'hf : _GEN_22332; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22334 = 10'hef == _T_445[9:0] ? 4'hf : _GEN_22333; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22335 = 10'hf0 == _T_445[9:0] ? 4'hf : _GEN_22334; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22336 = 10'hf1 == _T_445[9:0] ? 4'hf : _GEN_22335; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22337 = 10'hf2 == _T_445[9:0] ? 4'hf : _GEN_22336; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22338 = 10'hf3 == _T_445[9:0] ? 4'hf : _GEN_22337; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22339 = 10'hf4 == _T_445[9:0] ? 4'hf : _GEN_22338; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22340 = 10'hf5 == _T_445[9:0] ? 4'h9 : _GEN_22339; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22341 = 10'hf6 == _T_445[9:0] ? 4'hf : _GEN_22340; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22342 = 10'hf7 == _T_445[9:0] ? 4'hf : _GEN_22341; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22343 = 10'hf8 == _T_445[9:0] ? 4'h9 : _GEN_22342; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22344 = 10'hf9 == _T_445[9:0] ? 4'hf : _GEN_22343; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22345 = 10'hfa == _T_445[9:0] ? 4'h3 : _GEN_22344; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22346 = 10'hfb == _T_445[9:0] ? 4'h3 : _GEN_22345; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22347 = 10'hfc == _T_445[9:0] ? 4'h3 : _GEN_22346; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22348 = 10'hfd == _T_445[9:0] ? 4'h3 : _GEN_22347; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22349 = 10'hfe == _T_445[9:0] ? 4'h3 : _GEN_22348; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22350 = 10'hff == _T_445[9:0] ? 4'h0 : _GEN_22349; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22351 = 10'h100 == _T_445[9:0] ? 4'h3 : _GEN_22350; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22352 = 10'h101 == _T_445[9:0] ? 4'hf : _GEN_22351; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22353 = 10'h102 == _T_445[9:0] ? 4'h3 : _GEN_22352; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22354 = 10'h103 == _T_445[9:0] ? 4'h3 : _GEN_22353; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22355 = 10'h104 == _T_445[9:0] ? 4'h3 : _GEN_22354; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22356 = 10'h105 == _T_445[9:0] ? 4'h3 : _GEN_22355; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22357 = 10'h106 == _T_445[9:0] ? 4'h3 : _GEN_22356; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22358 = 10'h107 == _T_445[9:0] ? 4'h3 : _GEN_22357; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22359 = 10'h108 == _T_445[9:0] ? 4'h9 : _GEN_22358; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22360 = 10'h109 == _T_445[9:0] ? 4'hf : _GEN_22359; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22361 = 10'h10a == _T_445[9:0] ? 4'hf : _GEN_22360; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22362 = 10'h10b == _T_445[9:0] ? 4'hf : _GEN_22361; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22363 = 10'h10c == _T_445[9:0] ? 4'hf : _GEN_22362; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22364 = 10'h10d == _T_445[9:0] ? 4'h0 : _GEN_22363; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22365 = 10'h10e == _T_445[9:0] ? 4'hf : _GEN_22364; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22366 = 10'h10f == _T_445[9:0] ? 4'hf : _GEN_22365; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22367 = 10'h110 == _T_445[9:0] ? 4'hf : _GEN_22366; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22368 = 10'h111 == _T_445[9:0] ? 4'h0 : _GEN_22367; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22369 = 10'h112 == _T_445[9:0] ? 4'hf : _GEN_22368; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22370 = 10'h113 == _T_445[9:0] ? 4'hf : _GEN_22369; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22371 = 10'h114 == _T_445[9:0] ? 4'hf : _GEN_22370; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22372 = 10'h115 == _T_445[9:0] ? 4'hf : _GEN_22371; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22373 = 10'h116 == _T_445[9:0] ? 4'h9 : _GEN_22372; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22374 = 10'h117 == _T_445[9:0] ? 4'h3 : _GEN_22373; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22375 = 10'h118 == _T_445[9:0] ? 4'h3 : _GEN_22374; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22376 = 10'h119 == _T_445[9:0] ? 4'h3 : _GEN_22375; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22377 = 10'h11a == _T_445[9:0] ? 4'hf : _GEN_22376; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22378 = 10'h11b == _T_445[9:0] ? 4'h3 : _GEN_22377; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22379 = 10'h11c == _T_445[9:0] ? 4'h3 : _GEN_22378; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22380 = 10'h11d == _T_445[9:0] ? 4'h2 : _GEN_22379; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22381 = 10'h11e == _T_445[9:0] ? 4'h3 : _GEN_22380; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22382 = 10'h11f == _T_445[9:0] ? 4'h0 : _GEN_22381; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22383 = 10'h120 == _T_445[9:0] ? 4'h3 : _GEN_22382; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22384 = 10'h121 == _T_445[9:0] ? 4'h3 : _GEN_22383; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22385 = 10'h122 == _T_445[9:0] ? 4'h3 : _GEN_22384; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22386 = 10'h123 == _T_445[9:0] ? 4'h3 : _GEN_22385; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22387 = 10'h124 == _T_445[9:0] ? 4'h3 : _GEN_22386; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22388 = 10'h125 == _T_445[9:0] ? 4'h3 : _GEN_22387; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22389 = 10'h126 == _T_445[9:0] ? 4'h3 : _GEN_22388; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22390 = 10'h127 == _T_445[9:0] ? 4'h9 : _GEN_22389; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22391 = 10'h128 == _T_445[9:0] ? 4'hf : _GEN_22390; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22392 = 10'h129 == _T_445[9:0] ? 4'h3 : _GEN_22391; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22393 = 10'h12a == _T_445[9:0] ? 4'h3 : _GEN_22392; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22394 = 10'h12b == _T_445[9:0] ? 4'hf : _GEN_22393; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22395 = 10'h12c == _T_445[9:0] ? 4'hf : _GEN_22394; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22396 = 10'h12d == _T_445[9:0] ? 4'hf : _GEN_22395; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22397 = 10'h12e == _T_445[9:0] ? 4'hf : _GEN_22396; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22398 = 10'h12f == _T_445[9:0] ? 4'hf : _GEN_22397; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22399 = 10'h130 == _T_445[9:0] ? 4'hf : _GEN_22398; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22400 = 10'h131 == _T_445[9:0] ? 4'hf : _GEN_22399; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22401 = 10'h132 == _T_445[9:0] ? 4'hf : _GEN_22400; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22402 = 10'h133 == _T_445[9:0] ? 4'hf : _GEN_22401; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22403 = 10'h134 == _T_445[9:0] ? 4'h3 : _GEN_22402; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22404 = 10'h135 == _T_445[9:0] ? 4'h3 : _GEN_22403; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22405 = 10'h136 == _T_445[9:0] ? 4'hf : _GEN_22404; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22406 = 10'h137 == _T_445[9:0] ? 4'h9 : _GEN_22405; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22407 = 10'h138 == _T_445[9:0] ? 4'h3 : _GEN_22406; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22408 = 10'h139 == _T_445[9:0] ? 4'h3 : _GEN_22407; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22409 = 10'h13a == _T_445[9:0] ? 4'h3 : _GEN_22408; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22410 = 10'h13b == _T_445[9:0] ? 4'h3 : _GEN_22409; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22411 = 10'h13c == _T_445[9:0] ? 4'h3 : _GEN_22410; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22412 = 10'h13d == _T_445[9:0] ? 4'h3 : _GEN_22411; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22413 = 10'h13e == _T_445[9:0] ? 4'h3 : _GEN_22412; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22414 = 10'h13f == _T_445[9:0] ? 4'h0 : _GEN_22413; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22415 = 10'h140 == _T_445[9:0] ? 4'h3 : _GEN_22414; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22416 = 10'h141 == _T_445[9:0] ? 4'h3 : _GEN_22415; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22417 = 10'h142 == _T_445[9:0] ? 4'h2 : _GEN_22416; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22418 = 10'h143 == _T_445[9:0] ? 4'h3 : _GEN_22417; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22419 = 10'h144 == _T_445[9:0] ? 4'h3 : _GEN_22418; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22420 = 10'h145 == _T_445[9:0] ? 4'h3 : _GEN_22419; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22421 = 10'h146 == _T_445[9:0] ? 4'h9 : _GEN_22420; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22422 = 10'h147 == _T_445[9:0] ? 4'hf : _GEN_22421; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22423 = 10'h148 == _T_445[9:0] ? 4'h3 : _GEN_22422; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22424 = 10'h149 == _T_445[9:0] ? 4'h3 : _GEN_22423; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22425 = 10'h14a == _T_445[9:0] ? 4'h3 : _GEN_22424; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22426 = 10'h14b == _T_445[9:0] ? 4'h3 : _GEN_22425; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22427 = 10'h14c == _T_445[9:0] ? 4'h3 : _GEN_22426; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22428 = 10'h14d == _T_445[9:0] ? 4'h3 : _GEN_22427; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22429 = 10'h14e == _T_445[9:0] ? 4'h3 : _GEN_22428; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22430 = 10'h14f == _T_445[9:0] ? 4'h3 : _GEN_22429; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22431 = 10'h150 == _T_445[9:0] ? 4'h3 : _GEN_22430; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22432 = 10'h151 == _T_445[9:0] ? 4'h3 : _GEN_22431; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22433 = 10'h152 == _T_445[9:0] ? 4'h3 : _GEN_22432; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22434 = 10'h153 == _T_445[9:0] ? 4'h3 : _GEN_22433; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22435 = 10'h154 == _T_445[9:0] ? 4'h3 : _GEN_22434; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22436 = 10'h155 == _T_445[9:0] ? 4'h3 : _GEN_22435; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22437 = 10'h156 == _T_445[9:0] ? 4'h3 : _GEN_22436; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22438 = 10'h157 == _T_445[9:0] ? 4'hf : _GEN_22437; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22439 = 10'h158 == _T_445[9:0] ? 4'h3 : _GEN_22438; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22440 = 10'h159 == _T_445[9:0] ? 4'h3 : _GEN_22439; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22441 = 10'h15a == _T_445[9:0] ? 4'h3 : _GEN_22440; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22442 = 10'h15b == _T_445[9:0] ? 4'h3 : _GEN_22441; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22443 = 10'h15c == _T_445[9:0] ? 4'h3 : _GEN_22442; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22444 = 10'h15d == _T_445[9:0] ? 4'h3 : _GEN_22443; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22445 = 10'h15e == _T_445[9:0] ? 4'h2 : _GEN_22444; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22446 = 10'h15f == _T_445[9:0] ? 4'h0 : _GEN_22445; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22447 = 10'h160 == _T_445[9:0] ? 4'h3 : _GEN_22446; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22448 = 10'h161 == _T_445[9:0] ? 4'h3 : _GEN_22447; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22449 = 10'h162 == _T_445[9:0] ? 4'h3 : _GEN_22448; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22450 = 10'h163 == _T_445[9:0] ? 4'h2 : _GEN_22449; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22451 = 10'h164 == _T_445[9:0] ? 4'h3 : _GEN_22450; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22452 = 10'h165 == _T_445[9:0] ? 4'h9 : _GEN_22451; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22453 = 10'h166 == _T_445[9:0] ? 4'hf : _GEN_22452; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22454 = 10'h167 == _T_445[9:0] ? 4'hf : _GEN_22453; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22455 = 10'h168 == _T_445[9:0] ? 4'hd : _GEN_22454; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22456 = 10'h169 == _T_445[9:0] ? 4'h9 : _GEN_22455; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22457 = 10'h16a == _T_445[9:0] ? 4'hd : _GEN_22456; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22458 = 10'h16b == _T_445[9:0] ? 4'hd : _GEN_22457; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22459 = 10'h16c == _T_445[9:0] ? 4'h3 : _GEN_22458; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22460 = 10'h16d == _T_445[9:0] ? 4'h3 : _GEN_22459; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22461 = 10'h16e == _T_445[9:0] ? 4'h3 : _GEN_22460; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22462 = 10'h16f == _T_445[9:0] ? 4'h3 : _GEN_22461; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22463 = 10'h170 == _T_445[9:0] ? 4'h3 : _GEN_22462; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22464 = 10'h171 == _T_445[9:0] ? 4'h3 : _GEN_22463; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22465 = 10'h172 == _T_445[9:0] ? 4'h3 : _GEN_22464; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22466 = 10'h173 == _T_445[9:0] ? 4'h3 : _GEN_22465; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22467 = 10'h174 == _T_445[9:0] ? 4'h3 : _GEN_22466; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22468 = 10'h175 == _T_445[9:0] ? 4'h3 : _GEN_22467; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22469 = 10'h176 == _T_445[9:0] ? 4'hf : _GEN_22468; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22470 = 10'h177 == _T_445[9:0] ? 4'hf : _GEN_22469; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22471 = 10'h178 == _T_445[9:0] ? 4'h9 : _GEN_22470; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22472 = 10'h179 == _T_445[9:0] ? 4'h3 : _GEN_22471; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22473 = 10'h17a == _T_445[9:0] ? 4'h3 : _GEN_22472; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22474 = 10'h17b == _T_445[9:0] ? 4'h3 : _GEN_22473; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22475 = 10'h17c == _T_445[9:0] ? 4'h3 : _GEN_22474; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22476 = 10'h17d == _T_445[9:0] ? 4'h2 : _GEN_22475; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22477 = 10'h17e == _T_445[9:0] ? 4'h3 : _GEN_22476; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22478 = 10'h17f == _T_445[9:0] ? 4'h0 : _GEN_22477; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22479 = 10'h180 == _T_445[9:0] ? 4'hd : _GEN_22478; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22480 = 10'h181 == _T_445[9:0] ? 4'hd : _GEN_22479; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22481 = 10'h182 == _T_445[9:0] ? 4'hd : _GEN_22480; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22482 = 10'h183 == _T_445[9:0] ? 4'hd : _GEN_22481; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22483 = 10'h184 == _T_445[9:0] ? 4'h3 : _GEN_22482; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22484 = 10'h185 == _T_445[9:0] ? 4'h9 : _GEN_22483; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22485 = 10'h186 == _T_445[9:0] ? 4'hb : _GEN_22484; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22486 = 10'h187 == _T_445[9:0] ? 4'hf : _GEN_22485; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22487 = 10'h188 == _T_445[9:0] ? 4'hd : _GEN_22486; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22488 = 10'h189 == _T_445[9:0] ? 4'hd : _GEN_22487; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22489 = 10'h18a == _T_445[9:0] ? 4'hd : _GEN_22488; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22490 = 10'h18b == _T_445[9:0] ? 4'hd : _GEN_22489; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22491 = 10'h18c == _T_445[9:0] ? 4'hd : _GEN_22490; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22492 = 10'h18d == _T_445[9:0] ? 4'hd : _GEN_22491; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22493 = 10'h18e == _T_445[9:0] ? 4'hd : _GEN_22492; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22494 = 10'h18f == _T_445[9:0] ? 4'hd : _GEN_22493; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22495 = 10'h190 == _T_445[9:0] ? 4'hd : _GEN_22494; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22496 = 10'h191 == _T_445[9:0] ? 4'hd : _GEN_22495; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22497 = 10'h192 == _T_445[9:0] ? 4'h9 : _GEN_22496; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22498 = 10'h193 == _T_445[9:0] ? 4'hd : _GEN_22497; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22499 = 10'h194 == _T_445[9:0] ? 4'hd : _GEN_22498; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22500 = 10'h195 == _T_445[9:0] ? 4'hd : _GEN_22499; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22501 = 10'h196 == _T_445[9:0] ? 4'hf : _GEN_22500; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22502 = 10'h197 == _T_445[9:0] ? 4'h3 : _GEN_22501; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22503 = 10'h198 == _T_445[9:0] ? 4'h9 : _GEN_22502; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22504 = 10'h199 == _T_445[9:0] ? 4'h3 : _GEN_22503; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22505 = 10'h19a == _T_445[9:0] ? 4'h3 : _GEN_22504; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22506 = 10'h19b == _T_445[9:0] ? 4'h3 : _GEN_22505; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22507 = 10'h19c == _T_445[9:0] ? 4'h3 : _GEN_22506; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22508 = 10'h19d == _T_445[9:0] ? 4'h3 : _GEN_22507; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22509 = 10'h19e == _T_445[9:0] ? 4'h3 : _GEN_22508; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22510 = 10'h19f == _T_445[9:0] ? 4'h0 : _GEN_22509; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22511 = 10'h1a0 == _T_445[9:0] ? 4'hd : _GEN_22510; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22512 = 10'h1a1 == _T_445[9:0] ? 4'hd : _GEN_22511; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22513 = 10'h1a2 == _T_445[9:0] ? 4'h9 : _GEN_22512; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22514 = 10'h1a3 == _T_445[9:0] ? 4'hd : _GEN_22513; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22515 = 10'h1a4 == _T_445[9:0] ? 4'h3 : _GEN_22514; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22516 = 10'h1a5 == _T_445[9:0] ? 4'hf : _GEN_22515; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22517 = 10'h1a6 == _T_445[9:0] ? 4'hd : _GEN_22516; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22518 = 10'h1a7 == _T_445[9:0] ? 4'hf : _GEN_22517; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22519 = 10'h1a8 == _T_445[9:0] ? 4'hb : _GEN_22518; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22520 = 10'h1a9 == _T_445[9:0] ? 4'hd : _GEN_22519; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22521 = 10'h1aa == _T_445[9:0] ? 4'hd : _GEN_22520; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22522 = 10'h1ab == _T_445[9:0] ? 4'h9 : _GEN_22521; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22523 = 10'h1ac == _T_445[9:0] ? 4'hd : _GEN_22522; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22524 = 10'h1ad == _T_445[9:0] ? 4'hd : _GEN_22523; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22525 = 10'h1ae == _T_445[9:0] ? 4'hd : _GEN_22524; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22526 = 10'h1af == _T_445[9:0] ? 4'hd : _GEN_22525; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22527 = 10'h1b0 == _T_445[9:0] ? 4'hd : _GEN_22526; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22528 = 10'h1b1 == _T_445[9:0] ? 4'hd : _GEN_22527; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22529 = 10'h1b2 == _T_445[9:0] ? 4'hd : _GEN_22528; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22530 = 10'h1b3 == _T_445[9:0] ? 4'hd : _GEN_22529; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22531 = 10'h1b4 == _T_445[9:0] ? 4'hd : _GEN_22530; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22532 = 10'h1b5 == _T_445[9:0] ? 4'hd : _GEN_22531; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22533 = 10'h1b6 == _T_445[9:0] ? 4'hf : _GEN_22532; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22534 = 10'h1b7 == _T_445[9:0] ? 4'hd : _GEN_22533; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22535 = 10'h1b8 == _T_445[9:0] ? 4'hf : _GEN_22534; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22536 = 10'h1b9 == _T_445[9:0] ? 4'hd : _GEN_22535; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22537 = 10'h1ba == _T_445[9:0] ? 4'hd : _GEN_22536; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22538 = 10'h1bb == _T_445[9:0] ? 4'hd : _GEN_22537; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22539 = 10'h1bc == _T_445[9:0] ? 4'h2 : _GEN_22538; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22540 = 10'h1bd == _T_445[9:0] ? 4'h3 : _GEN_22539; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22541 = 10'h1be == _T_445[9:0] ? 4'hd : _GEN_22540; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22542 = 10'h1bf == _T_445[9:0] ? 4'h0 : _GEN_22541; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22543 = 10'h1c0 == _T_445[9:0] ? 4'hd : _GEN_22542; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22544 = 10'h1c1 == _T_445[9:0] ? 4'hd : _GEN_22543; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22545 = 10'h1c2 == _T_445[9:0] ? 4'hd : _GEN_22544; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22546 = 10'h1c3 == _T_445[9:0] ? 4'h2 : _GEN_22545; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22547 = 10'h1c4 == _T_445[9:0] ? 4'h2 : _GEN_22546; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22548 = 10'h1c5 == _T_445[9:0] ? 4'hd : _GEN_22547; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22549 = 10'h1c6 == _T_445[9:0] ? 4'hd : _GEN_22548; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22550 = 10'h1c7 == _T_445[9:0] ? 4'hd : _GEN_22549; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22551 = 10'h1c8 == _T_445[9:0] ? 4'hd : _GEN_22550; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22552 = 10'h1c9 == _T_445[9:0] ? 4'hb : _GEN_22551; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22553 = 10'h1ca == _T_445[9:0] ? 4'hb : _GEN_22552; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22554 = 10'h1cb == _T_445[9:0] ? 4'hb : _GEN_22553; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22555 = 10'h1cc == _T_445[9:0] ? 4'hb : _GEN_22554; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22556 = 10'h1cd == _T_445[9:0] ? 4'hb : _GEN_22555; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22557 = 10'h1ce == _T_445[9:0] ? 4'hb : _GEN_22556; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22558 = 10'h1cf == _T_445[9:0] ? 4'hb : _GEN_22557; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22559 = 10'h1d0 == _T_445[9:0] ? 4'hb : _GEN_22558; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22560 = 10'h1d1 == _T_445[9:0] ? 4'hb : _GEN_22559; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22561 = 10'h1d2 == _T_445[9:0] ? 4'hb : _GEN_22560; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22562 = 10'h1d3 == _T_445[9:0] ? 4'hb : _GEN_22561; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22563 = 10'h1d4 == _T_445[9:0] ? 4'hb : _GEN_22562; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22564 = 10'h1d5 == _T_445[9:0] ? 4'hb : _GEN_22563; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22565 = 10'h1d6 == _T_445[9:0] ? 4'hd : _GEN_22564; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22566 = 10'h1d7 == _T_445[9:0] ? 4'hd : _GEN_22565; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22567 = 10'h1d8 == _T_445[9:0] ? 4'hd : _GEN_22566; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22568 = 10'h1d9 == _T_445[9:0] ? 4'hd : _GEN_22567; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22569 = 10'h1da == _T_445[9:0] ? 4'hd : _GEN_22568; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22570 = 10'h1db == _T_445[9:0] ? 4'hd : _GEN_22569; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22571 = 10'h1dc == _T_445[9:0] ? 4'hd : _GEN_22570; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22572 = 10'h1dd == _T_445[9:0] ? 4'h3 : _GEN_22571; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22573 = 10'h1de == _T_445[9:0] ? 4'hd : _GEN_22572; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22574 = 10'h1df == _T_445[9:0] ? 4'h0 : _GEN_22573; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22575 = 10'h1e0 == _T_445[9:0] ? 4'h9 : _GEN_22574; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22576 = 10'h1e1 == _T_445[9:0] ? 4'hd : _GEN_22575; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22577 = 10'h1e2 == _T_445[9:0] ? 4'h2 : _GEN_22576; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22578 = 10'h1e3 == _T_445[9:0] ? 4'h2 : _GEN_22577; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22579 = 10'h1e4 == _T_445[9:0] ? 4'hd : _GEN_22578; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22580 = 10'h1e5 == _T_445[9:0] ? 4'hd : _GEN_22579; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22581 = 10'h1e6 == _T_445[9:0] ? 4'hd : _GEN_22580; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22582 = 10'h1e7 == _T_445[9:0] ? 4'hd : _GEN_22581; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22583 = 10'h1e8 == _T_445[9:0] ? 4'hb : _GEN_22582; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22584 = 10'h1e9 == _T_445[9:0] ? 4'hd : _GEN_22583; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22585 = 10'h1ea == _T_445[9:0] ? 4'hd : _GEN_22584; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22586 = 10'h1eb == _T_445[9:0] ? 4'hb : _GEN_22585; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22587 = 10'h1ec == _T_445[9:0] ? 4'hd : _GEN_22586; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22588 = 10'h1ed == _T_445[9:0] ? 4'hb : _GEN_22587; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22589 = 10'h1ee == _T_445[9:0] ? 4'hd : _GEN_22588; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22590 = 10'h1ef == _T_445[9:0] ? 4'hb : _GEN_22589; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22591 = 10'h1f0 == _T_445[9:0] ? 4'hd : _GEN_22590; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22592 = 10'h1f1 == _T_445[9:0] ? 4'hb : _GEN_22591; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22593 = 10'h1f2 == _T_445[9:0] ? 4'hb : _GEN_22592; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22594 = 10'h1f3 == _T_445[9:0] ? 4'hd : _GEN_22593; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22595 = 10'h1f4 == _T_445[9:0] ? 4'hb : _GEN_22594; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22596 = 10'h1f5 == _T_445[9:0] ? 4'hb : _GEN_22595; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22597 = 10'h1f6 == _T_445[9:0] ? 4'hd : _GEN_22596; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22598 = 10'h1f7 == _T_445[9:0] ? 4'hd : _GEN_22597; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22599 = 10'h1f8 == _T_445[9:0] ? 4'hd : _GEN_22598; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22600 = 10'h1f9 == _T_445[9:0] ? 4'hd : _GEN_22599; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22601 = 10'h1fa == _T_445[9:0] ? 4'h9 : _GEN_22600; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22602 = 10'h1fb == _T_445[9:0] ? 4'hd : _GEN_22601; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22603 = 10'h1fc == _T_445[9:0] ? 4'hd : _GEN_22602; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22604 = 10'h1fd == _T_445[9:0] ? 4'h2 : _GEN_22603; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22605 = 10'h1fe == _T_445[9:0] ? 4'hd : _GEN_22604; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22606 = 10'h1ff == _T_445[9:0] ? 4'h0 : _GEN_22605; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22607 = 10'h200 == _T_445[9:0] ? 4'hd : _GEN_22606; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22608 = 10'h201 == _T_445[9:0] ? 4'hd : _GEN_22607; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22609 = 10'h202 == _T_445[9:0] ? 4'h3 : _GEN_22608; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22610 = 10'h203 == _T_445[9:0] ? 4'hd : _GEN_22609; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22611 = 10'h204 == _T_445[9:0] ? 4'hd : _GEN_22610; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22612 = 10'h205 == _T_445[9:0] ? 4'hd : _GEN_22611; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22613 = 10'h206 == _T_445[9:0] ? 4'hb : _GEN_22612; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22614 = 10'h207 == _T_445[9:0] ? 4'hb : _GEN_22613; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22615 = 10'h208 == _T_445[9:0] ? 4'hd : _GEN_22614; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22616 = 10'h209 == _T_445[9:0] ? 4'hd : _GEN_22615; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22617 = 10'h20a == _T_445[9:0] ? 4'hd : _GEN_22616; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22618 = 10'h20b == _T_445[9:0] ? 4'hb : _GEN_22617; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22619 = 10'h20c == _T_445[9:0] ? 4'hd : _GEN_22618; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22620 = 10'h20d == _T_445[9:0] ? 4'hb : _GEN_22619; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22621 = 10'h20e == _T_445[9:0] ? 4'hd : _GEN_22620; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22622 = 10'h20f == _T_445[9:0] ? 4'hb : _GEN_22621; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22623 = 10'h210 == _T_445[9:0] ? 4'hd : _GEN_22622; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22624 = 10'h211 == _T_445[9:0] ? 4'hd : _GEN_22623; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22625 = 10'h212 == _T_445[9:0] ? 4'hb : _GEN_22624; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22626 = 10'h213 == _T_445[9:0] ? 4'hb : _GEN_22625; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22627 = 10'h214 == _T_445[9:0] ? 4'hb : _GEN_22626; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22628 = 10'h215 == _T_445[9:0] ? 4'hd : _GEN_22627; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22629 = 10'h216 == _T_445[9:0] ? 4'hd : _GEN_22628; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22630 = 10'h217 == _T_445[9:0] ? 4'hd : _GEN_22629; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22631 = 10'h218 == _T_445[9:0] ? 4'hd : _GEN_22630; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22632 = 10'h219 == _T_445[9:0] ? 4'hd : _GEN_22631; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22633 = 10'h21a == _T_445[9:0] ? 4'hd : _GEN_22632; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22634 = 10'h21b == _T_445[9:0] ? 4'hd : _GEN_22633; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22635 = 10'h21c == _T_445[9:0] ? 4'h3 : _GEN_22634; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22636 = 10'h21d == _T_445[9:0] ? 4'h2 : _GEN_22635; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22637 = 10'h21e == _T_445[9:0] ? 4'hd : _GEN_22636; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22638 = 10'h21f == _T_445[9:0] ? 4'h0 : _GEN_22637; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22639 = 10'h220 == _T_445[9:0] ? 4'h0 : _GEN_22638; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22640 = 10'h221 == _T_445[9:0] ? 4'h0 : _GEN_22639; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22641 = 10'h222 == _T_445[9:0] ? 4'h0 : _GEN_22640; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22642 = 10'h223 == _T_445[9:0] ? 4'h0 : _GEN_22641; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22643 = 10'h224 == _T_445[9:0] ? 4'h0 : _GEN_22642; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22644 = 10'h225 == _T_445[9:0] ? 4'h0 : _GEN_22643; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22645 = 10'h226 == _T_445[9:0] ? 4'h0 : _GEN_22644; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22646 = 10'h227 == _T_445[9:0] ? 4'h0 : _GEN_22645; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22647 = 10'h228 == _T_445[9:0] ? 4'h0 : _GEN_22646; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22648 = 10'h229 == _T_445[9:0] ? 4'h0 : _GEN_22647; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22649 = 10'h22a == _T_445[9:0] ? 4'h0 : _GEN_22648; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22650 = 10'h22b == _T_445[9:0] ? 4'h0 : _GEN_22649; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22651 = 10'h22c == _T_445[9:0] ? 4'h0 : _GEN_22650; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22652 = 10'h22d == _T_445[9:0] ? 4'h0 : _GEN_22651; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22653 = 10'h22e == _T_445[9:0] ? 4'h0 : _GEN_22652; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22654 = 10'h22f == _T_445[9:0] ? 4'h0 : _GEN_22653; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22655 = 10'h230 == _T_445[9:0] ? 4'h0 : _GEN_22654; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22656 = 10'h231 == _T_445[9:0] ? 4'h0 : _GEN_22655; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22657 = 10'h232 == _T_445[9:0] ? 4'h0 : _GEN_22656; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22658 = 10'h233 == _T_445[9:0] ? 4'h0 : _GEN_22657; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22659 = 10'h234 == _T_445[9:0] ? 4'h0 : _GEN_22658; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22660 = 10'h235 == _T_445[9:0] ? 4'h0 : _GEN_22659; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22661 = 10'h236 == _T_445[9:0] ? 4'h0 : _GEN_22660; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22662 = 10'h237 == _T_445[9:0] ? 4'h0 : _GEN_22661; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22663 = 10'h238 == _T_445[9:0] ? 4'h0 : _GEN_22662; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22664 = 10'h239 == _T_445[9:0] ? 4'h0 : _GEN_22663; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22665 = 10'h23a == _T_445[9:0] ? 4'h0 : _GEN_22664; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22666 = 10'h23b == _T_445[9:0] ? 4'h0 : _GEN_22665; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22667 = 10'h23c == _T_445[9:0] ? 4'h0 : _GEN_22666; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22668 = 10'h23d == _T_445[9:0] ? 4'h0 : _GEN_22667; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22669 = 10'h23e == _T_445[9:0] ? 4'h0 : _GEN_22668; // @[Filter.scala 191:142]
  wire [3:0] _GEN_22670 = 10'h23f == _T_445[9:0] ? 4'h0 : _GEN_22669; // @[Filter.scala 191:142]
  wire [7:0] _T_459 = _GEN_22670 * 4'ha; // @[Filter.scala 191:142]
  wire [10:0] _GEN_28375 = {{3'd0}, _T_459}; // @[Filter.scala 191:109]
  wire [10:0] _T_461 = _T_454 + _GEN_28375; // @[Filter.scala 191:109]
  wire [10:0] _T_462 = _T_461 / 11'h64; // @[Filter.scala 191:150]
  wire  _T_464 = _T_435 >= 6'h20; // @[Filter.scala 194:31]
  wire  _T_468 = _T_442 >= 32'h12; // @[Filter.scala 194:63]
  wire  _T_469 = _T_464 | _T_468; // @[Filter.scala 194:58]
  wire [10:0] _GEN_23247 = io_SPI_distort ? _T_462 : {{7'd0}, _GEN_21518}; // @[Filter.scala 196:35]
  wire [10:0] _GEN_23248 = _T_469 ? 11'h0 : _GEN_23247; // @[Filter.scala 194:80]
  wire [10:0] _GEN_23825 = io_SPI_distort ? _T_462 : {{7'd0}, _GEN_22094}; // @[Filter.scala 196:35]
  wire [10:0] _GEN_23826 = _T_469 ? 11'h0 : _GEN_23825; // @[Filter.scala 194:80]
  wire [10:0] _GEN_24403 = io_SPI_distort ? _T_462 : {{7'd0}, _GEN_22670}; // @[Filter.scala 196:35]
  wire [10:0] _GEN_24404 = _T_469 ? 11'h0 : _GEN_24403; // @[Filter.scala 194:80]
  wire [31:0] _T_497 = pixelIndex + 32'h7; // @[Filter.scala 189:31]
  wire [31:0] _GEN_56 = _T_497 % 32'h20; // @[Filter.scala 189:38]
  wire [5:0] _T_498 = _GEN_56[5:0]; // @[Filter.scala 189:38]
  wire [5:0] _T_500 = _T_498 + _GEN_28295; // @[Filter.scala 189:53]
  wire [5:0] _T_502 = _T_500 - 6'h1; // @[Filter.scala 189:69]
  wire [31:0] _T_505 = _T_497 / 32'h20; // @[Filter.scala 190:38]
  wire [31:0] _T_507 = _T_505 + _GEN_28296; // @[Filter.scala 190:53]
  wire [31:0] _T_509 = _T_507 - 32'h1; // @[Filter.scala 190:69]
  wire [37:0] _T_510 = _T_509 * 32'h20; // @[Filter.scala 191:42]
  wire [37:0] _GEN_28381 = {{32'd0}, _T_502}; // @[Filter.scala 191:57]
  wire [37:0] _T_512 = _T_510 + _GEN_28381; // @[Filter.scala 191:57]
  wire [3:0] _GEN_24408 = 10'h3 == _T_512[9:0] ? 4'h3 : 4'ha; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24409 = 10'h4 == _T_512[9:0] ? 4'ha : _GEN_24408; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24410 = 10'h5 == _T_512[9:0] ? 4'ha : _GEN_24409; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24411 = 10'h6 == _T_512[9:0] ? 4'ha : _GEN_24410; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24412 = 10'h7 == _T_512[9:0] ? 4'ha : _GEN_24411; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24413 = 10'h8 == _T_512[9:0] ? 4'ha : _GEN_24412; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24414 = 10'h9 == _T_512[9:0] ? 4'ha : _GEN_24413; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24415 = 10'ha == _T_512[9:0] ? 4'ha : _GEN_24414; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24416 = 10'hb == _T_512[9:0] ? 4'ha : _GEN_24415; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24417 = 10'hc == _T_512[9:0] ? 4'ha : _GEN_24416; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24418 = 10'hd == _T_512[9:0] ? 4'ha : _GEN_24417; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24419 = 10'he == _T_512[9:0] ? 4'ha : _GEN_24418; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24420 = 10'hf == _T_512[9:0] ? 4'ha : _GEN_24419; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24421 = 10'h10 == _T_512[9:0] ? 4'ha : _GEN_24420; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24422 = 10'h11 == _T_512[9:0] ? 4'ha : _GEN_24421; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24423 = 10'h12 == _T_512[9:0] ? 4'ha : _GEN_24422; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24424 = 10'h13 == _T_512[9:0] ? 4'ha : _GEN_24423; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24425 = 10'h14 == _T_512[9:0] ? 4'ha : _GEN_24424; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24426 = 10'h15 == _T_512[9:0] ? 4'ha : _GEN_24425; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24427 = 10'h16 == _T_512[9:0] ? 4'ha : _GEN_24426; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24428 = 10'h17 == _T_512[9:0] ? 4'ha : _GEN_24427; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24429 = 10'h18 == _T_512[9:0] ? 4'ha : _GEN_24428; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24430 = 10'h19 == _T_512[9:0] ? 4'ha : _GEN_24429; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24431 = 10'h1a == _T_512[9:0] ? 4'ha : _GEN_24430; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24432 = 10'h1b == _T_512[9:0] ? 4'ha : _GEN_24431; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24433 = 10'h1c == _T_512[9:0] ? 4'ha : _GEN_24432; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24434 = 10'h1d == _T_512[9:0] ? 4'ha : _GEN_24433; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24435 = 10'h1e == _T_512[9:0] ? 4'ha : _GEN_24434; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24436 = 10'h1f == _T_512[9:0] ? 4'h0 : _GEN_24435; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24437 = 10'h20 == _T_512[9:0] ? 4'ha : _GEN_24436; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24438 = 10'h21 == _T_512[9:0] ? 4'ha : _GEN_24437; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24439 = 10'h22 == _T_512[9:0] ? 4'ha : _GEN_24438; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24440 = 10'h23 == _T_512[9:0] ? 4'h3 : _GEN_24439; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24441 = 10'h24 == _T_512[9:0] ? 4'ha : _GEN_24440; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24442 = 10'h25 == _T_512[9:0] ? 4'ha : _GEN_24441; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24443 = 10'h26 == _T_512[9:0] ? 4'ha : _GEN_24442; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24444 = 10'h27 == _T_512[9:0] ? 4'h1 : _GEN_24443; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24445 = 10'h28 == _T_512[9:0] ? 4'h1 : _GEN_24444; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24446 = 10'h29 == _T_512[9:0] ? 4'ha : _GEN_24445; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24447 = 10'h2a == _T_512[9:0] ? 4'ha : _GEN_24446; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24448 = 10'h2b == _T_512[9:0] ? 4'ha : _GEN_24447; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24449 = 10'h2c == _T_512[9:0] ? 4'ha : _GEN_24448; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24450 = 10'h2d == _T_512[9:0] ? 4'ha : _GEN_24449; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24451 = 10'h2e == _T_512[9:0] ? 4'ha : _GEN_24450; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24452 = 10'h2f == _T_512[9:0] ? 4'ha : _GEN_24451; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24453 = 10'h30 == _T_512[9:0] ? 4'ha : _GEN_24452; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24454 = 10'h31 == _T_512[9:0] ? 4'ha : _GEN_24453; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24455 = 10'h32 == _T_512[9:0] ? 4'ha : _GEN_24454; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24456 = 10'h33 == _T_512[9:0] ? 4'ha : _GEN_24455; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24457 = 10'h34 == _T_512[9:0] ? 4'ha : _GEN_24456; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24458 = 10'h35 == _T_512[9:0] ? 4'ha : _GEN_24457; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24459 = 10'h36 == _T_512[9:0] ? 4'ha : _GEN_24458; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24460 = 10'h37 == _T_512[9:0] ? 4'h1 : _GEN_24459; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24461 = 10'h38 == _T_512[9:0] ? 4'h1 : _GEN_24460; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24462 = 10'h39 == _T_512[9:0] ? 4'ha : _GEN_24461; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24463 = 10'h3a == _T_512[9:0] ? 4'ha : _GEN_24462; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24464 = 10'h3b == _T_512[9:0] ? 4'ha : _GEN_24463; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24465 = 10'h3c == _T_512[9:0] ? 4'ha : _GEN_24464; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24466 = 10'h3d == _T_512[9:0] ? 4'h3 : _GEN_24465; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24467 = 10'h3e == _T_512[9:0] ? 4'ha : _GEN_24466; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24468 = 10'h3f == _T_512[9:0] ? 4'h0 : _GEN_24467; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24469 = 10'h40 == _T_512[9:0] ? 4'ha : _GEN_24468; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24470 = 10'h41 == _T_512[9:0] ? 4'ha : _GEN_24469; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24471 = 10'h42 == _T_512[9:0] ? 4'ha : _GEN_24470; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24472 = 10'h43 == _T_512[9:0] ? 4'h2 : _GEN_24471; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24473 = 10'h44 == _T_512[9:0] ? 4'h3 : _GEN_24472; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24474 = 10'h45 == _T_512[9:0] ? 4'h0 : _GEN_24473; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24475 = 10'h46 == _T_512[9:0] ? 4'h0 : _GEN_24474; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24476 = 10'h47 == _T_512[9:0] ? 4'h0 : _GEN_24475; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24477 = 10'h48 == _T_512[9:0] ? 4'h0 : _GEN_24476; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24478 = 10'h49 == _T_512[9:0] ? 4'ha : _GEN_24477; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24479 = 10'h4a == _T_512[9:0] ? 4'ha : _GEN_24478; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24480 = 10'h4b == _T_512[9:0] ? 4'ha : _GEN_24479; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24481 = 10'h4c == _T_512[9:0] ? 4'ha : _GEN_24480; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24482 = 10'h4d == _T_512[9:0] ? 4'ha : _GEN_24481; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24483 = 10'h4e == _T_512[9:0] ? 4'ha : _GEN_24482; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24484 = 10'h4f == _T_512[9:0] ? 4'ha : _GEN_24483; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24485 = 10'h50 == _T_512[9:0] ? 4'ha : _GEN_24484; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24486 = 10'h51 == _T_512[9:0] ? 4'ha : _GEN_24485; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24487 = 10'h52 == _T_512[9:0] ? 4'ha : _GEN_24486; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24488 = 10'h53 == _T_512[9:0] ? 4'ha : _GEN_24487; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24489 = 10'h54 == _T_512[9:0] ? 4'h1 : _GEN_24488; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24490 = 10'h55 == _T_512[9:0] ? 4'h1 : _GEN_24489; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24491 = 10'h56 == _T_512[9:0] ? 4'h1 : _GEN_24490; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24492 = 10'h57 == _T_512[9:0] ? 4'h0 : _GEN_24491; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24493 = 10'h58 == _T_512[9:0] ? 4'ha : _GEN_24492; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24494 = 10'h59 == _T_512[9:0] ? 4'h0 : _GEN_24493; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24495 = 10'h5a == _T_512[9:0] ? 4'ha : _GEN_24494; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24496 = 10'h5b == _T_512[9:0] ? 4'ha : _GEN_24495; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24497 = 10'h5c == _T_512[9:0] ? 4'ha : _GEN_24496; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24498 = 10'h5d == _T_512[9:0] ? 4'h3 : _GEN_24497; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24499 = 10'h5e == _T_512[9:0] ? 4'ha : _GEN_24498; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24500 = 10'h5f == _T_512[9:0] ? 4'h0 : _GEN_24499; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24501 = 10'h60 == _T_512[9:0] ? 4'ha : _GEN_24500; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24502 = 10'h61 == _T_512[9:0] ? 4'ha : _GEN_24501; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24503 = 10'h62 == _T_512[9:0] ? 4'ha : _GEN_24502; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24504 = 10'h63 == _T_512[9:0] ? 4'ha : _GEN_24503; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24505 = 10'h64 == _T_512[9:0] ? 4'h3 : _GEN_24504; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24506 = 10'h65 == _T_512[9:0] ? 4'h0 : _GEN_24505; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24507 = 10'h66 == _T_512[9:0] ? 4'ha : _GEN_24506; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24508 = 10'h67 == _T_512[9:0] ? 4'ha : _GEN_24507; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24509 = 10'h68 == _T_512[9:0] ? 4'ha : _GEN_24508; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24510 = 10'h69 == _T_512[9:0] ? 4'h0 : _GEN_24509; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24511 = 10'h6a == _T_512[9:0] ? 4'h1 : _GEN_24510; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24512 = 10'h6b == _T_512[9:0] ? 4'h1 : _GEN_24511; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24513 = 10'h6c == _T_512[9:0] ? 4'ha : _GEN_24512; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24514 = 10'h6d == _T_512[9:0] ? 4'ha : _GEN_24513; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24515 = 10'h6e == _T_512[9:0] ? 4'ha : _GEN_24514; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24516 = 10'h6f == _T_512[9:0] ? 4'ha : _GEN_24515; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24517 = 10'h70 == _T_512[9:0] ? 4'ha : _GEN_24516; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24518 = 10'h71 == _T_512[9:0] ? 4'ha : _GEN_24517; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24519 = 10'h72 == _T_512[9:0] ? 4'ha : _GEN_24518; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24520 = 10'h73 == _T_512[9:0] ? 4'h1 : _GEN_24519; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24521 = 10'h74 == _T_512[9:0] ? 4'h0 : _GEN_24520; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24522 = 10'h75 == _T_512[9:0] ? 4'h0 : _GEN_24521; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24523 = 10'h76 == _T_512[9:0] ? 4'h0 : _GEN_24522; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24524 = 10'h77 == _T_512[9:0] ? 4'ha : _GEN_24523; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24525 = 10'h78 == _T_512[9:0] ? 4'ha : _GEN_24524; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24526 = 10'h79 == _T_512[9:0] ? 4'ha : _GEN_24525; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24527 = 10'h7a == _T_512[9:0] ? 4'h0 : _GEN_24526; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24528 = 10'h7b == _T_512[9:0] ? 4'ha : _GEN_24527; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24529 = 10'h7c == _T_512[9:0] ? 4'ha : _GEN_24528; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24530 = 10'h7d == _T_512[9:0] ? 4'h2 : _GEN_24529; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24531 = 10'h7e == _T_512[9:0] ? 4'h3 : _GEN_24530; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24532 = 10'h7f == _T_512[9:0] ? 4'h0 : _GEN_24531; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24533 = 10'h80 == _T_512[9:0] ? 4'ha : _GEN_24532; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24534 = 10'h81 == _T_512[9:0] ? 4'ha : _GEN_24533; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24535 = 10'h82 == _T_512[9:0] ? 4'h1 : _GEN_24534; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24536 = 10'h83 == _T_512[9:0] ? 4'h0 : _GEN_24535; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24537 = 10'h84 == _T_512[9:0] ? 4'h2 : _GEN_24536; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24538 = 10'h85 == _T_512[9:0] ? 4'h1 : _GEN_24537; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24539 = 10'h86 == _T_512[9:0] ? 4'h1 : _GEN_24538; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24540 = 10'h87 == _T_512[9:0] ? 4'ha : _GEN_24539; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24541 = 10'h88 == _T_512[9:0] ? 4'ha : _GEN_24540; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24542 = 10'h89 == _T_512[9:0] ? 4'h0 : _GEN_24541; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24543 = 10'h8a == _T_512[9:0] ? 4'h0 : _GEN_24542; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24544 = 10'h8b == _T_512[9:0] ? 4'h1 : _GEN_24543; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24545 = 10'h8c == _T_512[9:0] ? 4'h1 : _GEN_24544; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24546 = 10'h8d == _T_512[9:0] ? 4'h1 : _GEN_24545; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24547 = 10'h8e == _T_512[9:0] ? 4'h1 : _GEN_24546; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24548 = 10'h8f == _T_512[9:0] ? 4'h1 : _GEN_24547; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24549 = 10'h90 == _T_512[9:0] ? 4'h1 : _GEN_24548; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24550 = 10'h91 == _T_512[9:0] ? 4'h1 : _GEN_24549; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24551 = 10'h92 == _T_512[9:0] ? 4'h1 : _GEN_24550; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24552 = 10'h93 == _T_512[9:0] ? 4'h0 : _GEN_24551; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24553 = 10'h94 == _T_512[9:0] ? 4'h0 : _GEN_24552; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24554 = 10'h95 == _T_512[9:0] ? 4'ha : _GEN_24553; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24555 = 10'h96 == _T_512[9:0] ? 4'ha : _GEN_24554; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24556 = 10'h97 == _T_512[9:0] ? 4'ha : _GEN_24555; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24557 = 10'h98 == _T_512[9:0] ? 4'h1 : _GEN_24556; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24558 = 10'h99 == _T_512[9:0] ? 4'h0 : _GEN_24557; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24559 = 10'h9a == _T_512[9:0] ? 4'h1 : _GEN_24558; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24560 = 10'h9b == _T_512[9:0] ? 4'h1 : _GEN_24559; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24561 = 10'h9c == _T_512[9:0] ? 4'ha : _GEN_24560; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24562 = 10'h9d == _T_512[9:0] ? 4'ha : _GEN_24561; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24563 = 10'h9e == _T_512[9:0] ? 4'h3 : _GEN_24562; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24564 = 10'h9f == _T_512[9:0] ? 4'h0 : _GEN_24563; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24565 = 10'ha0 == _T_512[9:0] ? 4'ha : _GEN_24564; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24566 = 10'ha1 == _T_512[9:0] ? 4'h1 : _GEN_24565; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24567 = 10'ha2 == _T_512[9:0] ? 4'h0 : _GEN_24566; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24568 = 10'ha3 == _T_512[9:0] ? 4'h3 : _GEN_24567; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24569 = 10'ha4 == _T_512[9:0] ? 4'ha : _GEN_24568; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24570 = 10'ha5 == _T_512[9:0] ? 4'ha : _GEN_24569; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24571 = 10'ha6 == _T_512[9:0] ? 4'ha : _GEN_24570; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24572 = 10'ha7 == _T_512[9:0] ? 4'h0 : _GEN_24571; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24573 = 10'ha8 == _T_512[9:0] ? 4'ha : _GEN_24572; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24574 = 10'ha9 == _T_512[9:0] ? 4'h1 : _GEN_24573; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24575 = 10'haa == _T_512[9:0] ? 4'h0 : _GEN_24574; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24576 = 10'hab == _T_512[9:0] ? 4'h0 : _GEN_24575; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24577 = 10'hac == _T_512[9:0] ? 4'h0 : _GEN_24576; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24578 = 10'had == _T_512[9:0] ? 4'h0 : _GEN_24577; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24579 = 10'hae == _T_512[9:0] ? 4'h0 : _GEN_24578; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24580 = 10'haf == _T_512[9:0] ? 4'h0 : _GEN_24579; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24581 = 10'hb0 == _T_512[9:0] ? 4'h0 : _GEN_24580; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24582 = 10'hb1 == _T_512[9:0] ? 4'h0 : _GEN_24581; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24583 = 10'hb2 == _T_512[9:0] ? 4'h0 : _GEN_24582; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24584 = 10'hb3 == _T_512[9:0] ? 4'h0 : _GEN_24583; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24585 = 10'hb4 == _T_512[9:0] ? 4'h1 : _GEN_24584; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24586 = 10'hb5 == _T_512[9:0] ? 4'h1 : _GEN_24585; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24587 = 10'hb6 == _T_512[9:0] ? 4'ha : _GEN_24586; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24588 = 10'hb7 == _T_512[9:0] ? 4'h0 : _GEN_24587; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24589 = 10'hb8 == _T_512[9:0] ? 4'ha : _GEN_24588; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24590 = 10'hb9 == _T_512[9:0] ? 4'ha : _GEN_24589; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24591 = 10'hba == _T_512[9:0] ? 4'ha : _GEN_24590; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24592 = 10'hbb == _T_512[9:0] ? 4'h0 : _GEN_24591; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24593 = 10'hbc == _T_512[9:0] ? 4'ha : _GEN_24592; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24594 = 10'hbd == _T_512[9:0] ? 4'ha : _GEN_24593; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24595 = 10'hbe == _T_512[9:0] ? 4'h3 : _GEN_24594; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24596 = 10'hbf == _T_512[9:0] ? 4'h0 : _GEN_24595; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24597 = 10'hc0 == _T_512[9:0] ? 4'ha : _GEN_24596; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24598 = 10'hc1 == _T_512[9:0] ? 4'ha : _GEN_24597; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24599 = 10'hc2 == _T_512[9:0] ? 4'h3 : _GEN_24598; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24600 = 10'hc3 == _T_512[9:0] ? 4'h2 : _GEN_24599; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24601 = 10'hc4 == _T_512[9:0] ? 4'h0 : _GEN_24600; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24602 = 10'hc5 == _T_512[9:0] ? 4'h0 : _GEN_24601; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24603 = 10'hc6 == _T_512[9:0] ? 4'h0 : _GEN_24602; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24604 = 10'hc7 == _T_512[9:0] ? 4'ha : _GEN_24603; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24605 = 10'hc8 == _T_512[9:0] ? 4'h1 : _GEN_24604; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24606 = 10'hc9 == _T_512[9:0] ? 4'h0 : _GEN_24605; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24607 = 10'hca == _T_512[9:0] ? 4'h0 : _GEN_24606; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24608 = 10'hcb == _T_512[9:0] ? 4'h0 : _GEN_24607; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24609 = 10'hcc == _T_512[9:0] ? 4'h0 : _GEN_24608; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24610 = 10'hcd == _T_512[9:0] ? 4'h0 : _GEN_24609; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24611 = 10'hce == _T_512[9:0] ? 4'h0 : _GEN_24610; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24612 = 10'hcf == _T_512[9:0] ? 4'h0 : _GEN_24611; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24613 = 10'hd0 == _T_512[9:0] ? 4'h0 : _GEN_24612; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24614 = 10'hd1 == _T_512[9:0] ? 4'h0 : _GEN_24613; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24615 = 10'hd2 == _T_512[9:0] ? 4'h0 : _GEN_24614; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24616 = 10'hd3 == _T_512[9:0] ? 4'h0 : _GEN_24615; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24617 = 10'hd4 == _T_512[9:0] ? 4'h0 : _GEN_24616; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24618 = 10'hd5 == _T_512[9:0] ? 4'h0 : _GEN_24617; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24619 = 10'hd6 == _T_512[9:0] ? 4'h1 : _GEN_24618; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24620 = 10'hd7 == _T_512[9:0] ? 4'ha : _GEN_24619; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24621 = 10'hd8 == _T_512[9:0] ? 4'h0 : _GEN_24620; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24622 = 10'hd9 == _T_512[9:0] ? 4'ha : _GEN_24621; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24623 = 10'hda == _T_512[9:0] ? 4'ha : _GEN_24622; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24624 = 10'hdb == _T_512[9:0] ? 4'ha : _GEN_24623; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24625 = 10'hdc == _T_512[9:0] ? 4'ha : _GEN_24624; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24626 = 10'hdd == _T_512[9:0] ? 4'h3 : _GEN_24625; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24627 = 10'hde == _T_512[9:0] ? 4'h2 : _GEN_24626; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24628 = 10'hdf == _T_512[9:0] ? 4'h0 : _GEN_24627; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24629 = 10'he0 == _T_512[9:0] ? 4'ha : _GEN_24628; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24630 = 10'he1 == _T_512[9:0] ? 4'ha : _GEN_24629; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24631 = 10'he2 == _T_512[9:0] ? 4'h3 : _GEN_24630; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24632 = 10'he3 == _T_512[9:0] ? 4'ha : _GEN_24631; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24633 = 10'he4 == _T_512[9:0] ? 4'ha : _GEN_24632; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24634 = 10'he5 == _T_512[9:0] ? 4'ha : _GEN_24633; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24635 = 10'he6 == _T_512[9:0] ? 4'ha : _GEN_24634; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24636 = 10'he7 == _T_512[9:0] ? 4'h1 : _GEN_24635; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24637 = 10'he8 == _T_512[9:0] ? 4'h1 : _GEN_24636; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24638 = 10'he9 == _T_512[9:0] ? 4'h1 : _GEN_24637; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24639 = 10'hea == _T_512[9:0] ? 4'h0 : _GEN_24638; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24640 = 10'heb == _T_512[9:0] ? 4'h0 : _GEN_24639; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24641 = 10'hec == _T_512[9:0] ? 4'h0 : _GEN_24640; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24642 = 10'hed == _T_512[9:0] ? 4'h0 : _GEN_24641; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24643 = 10'hee == _T_512[9:0] ? 4'h0 : _GEN_24642; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24644 = 10'hef == _T_512[9:0] ? 4'h0 : _GEN_24643; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24645 = 10'hf0 == _T_512[9:0] ? 4'h0 : _GEN_24644; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24646 = 10'hf1 == _T_512[9:0] ? 4'h0 : _GEN_24645; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24647 = 10'hf2 == _T_512[9:0] ? 4'h0 : _GEN_24646; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24648 = 10'hf3 == _T_512[9:0] ? 4'h0 : _GEN_24647; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24649 = 10'hf4 == _T_512[9:0] ? 4'h0 : _GEN_24648; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24650 = 10'hf5 == _T_512[9:0] ? 4'h1 : _GEN_24649; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24651 = 10'hf6 == _T_512[9:0] ? 4'h0 : _GEN_24650; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24652 = 10'hf7 == _T_512[9:0] ? 4'h0 : _GEN_24651; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24653 = 10'hf8 == _T_512[9:0] ? 4'h1 : _GEN_24652; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24654 = 10'hf9 == _T_512[9:0] ? 4'h0 : _GEN_24653; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24655 = 10'hfa == _T_512[9:0] ? 4'ha : _GEN_24654; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24656 = 10'hfb == _T_512[9:0] ? 4'ha : _GEN_24655; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24657 = 10'hfc == _T_512[9:0] ? 4'ha : _GEN_24656; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24658 = 10'hfd == _T_512[9:0] ? 4'h3 : _GEN_24657; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24659 = 10'hfe == _T_512[9:0] ? 4'ha : _GEN_24658; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24660 = 10'hff == _T_512[9:0] ? 4'h0 : _GEN_24659; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24661 = 10'h100 == _T_512[9:0] ? 4'ha : _GEN_24660; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24662 = 10'h101 == _T_512[9:0] ? 4'h0 : _GEN_24661; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24663 = 10'h102 == _T_512[9:0] ? 4'h3 : _GEN_24662; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24664 = 10'h103 == _T_512[9:0] ? 4'ha : _GEN_24663; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24665 = 10'h104 == _T_512[9:0] ? 4'ha : _GEN_24664; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24666 = 10'h105 == _T_512[9:0] ? 4'ha : _GEN_24665; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24667 = 10'h106 == _T_512[9:0] ? 4'ha : _GEN_24666; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24668 = 10'h107 == _T_512[9:0] ? 4'ha : _GEN_24667; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24669 = 10'h108 == _T_512[9:0] ? 4'h1 : _GEN_24668; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24670 = 10'h109 == _T_512[9:0] ? 4'h0 : _GEN_24669; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24671 = 10'h10a == _T_512[9:0] ? 4'h0 : _GEN_24670; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24672 = 10'h10b == _T_512[9:0] ? 4'h0 : _GEN_24671; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24673 = 10'h10c == _T_512[9:0] ? 4'h0 : _GEN_24672; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24674 = 10'h10d == _T_512[9:0] ? 4'h0 : _GEN_24673; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24675 = 10'h10e == _T_512[9:0] ? 4'h0 : _GEN_24674; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24676 = 10'h10f == _T_512[9:0] ? 4'h0 : _GEN_24675; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24677 = 10'h110 == _T_512[9:0] ? 4'h0 : _GEN_24676; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24678 = 10'h111 == _T_512[9:0] ? 4'h0 : _GEN_24677; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24679 = 10'h112 == _T_512[9:0] ? 4'h0 : _GEN_24678; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24680 = 10'h113 == _T_512[9:0] ? 4'h0 : _GEN_24679; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24681 = 10'h114 == _T_512[9:0] ? 4'h0 : _GEN_24680; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24682 = 10'h115 == _T_512[9:0] ? 4'h0 : _GEN_24681; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24683 = 10'h116 == _T_512[9:0] ? 4'h1 : _GEN_24682; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24684 = 10'h117 == _T_512[9:0] ? 4'ha : _GEN_24683; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24685 = 10'h118 == _T_512[9:0] ? 4'ha : _GEN_24684; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24686 = 10'h119 == _T_512[9:0] ? 4'ha : _GEN_24685; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24687 = 10'h11a == _T_512[9:0] ? 4'h0 : _GEN_24686; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24688 = 10'h11b == _T_512[9:0] ? 4'ha : _GEN_24687; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24689 = 10'h11c == _T_512[9:0] ? 4'ha : _GEN_24688; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24690 = 10'h11d == _T_512[9:0] ? 4'h2 : _GEN_24689; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24691 = 10'h11e == _T_512[9:0] ? 4'h3 : _GEN_24690; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24692 = 10'h11f == _T_512[9:0] ? 4'h0 : _GEN_24691; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24693 = 10'h120 == _T_512[9:0] ? 4'ha : _GEN_24692; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24694 = 10'h121 == _T_512[9:0] ? 4'ha : _GEN_24693; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24695 = 10'h122 == _T_512[9:0] ? 4'h3 : _GEN_24694; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24696 = 10'h123 == _T_512[9:0] ? 4'ha : _GEN_24695; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24697 = 10'h124 == _T_512[9:0] ? 4'ha : _GEN_24696; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24698 = 10'h125 == _T_512[9:0] ? 4'ha : _GEN_24697; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24699 = 10'h126 == _T_512[9:0] ? 4'ha : _GEN_24698; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24700 = 10'h127 == _T_512[9:0] ? 4'h1 : _GEN_24699; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24701 = 10'h128 == _T_512[9:0] ? 4'h0 : _GEN_24700; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24702 = 10'h129 == _T_512[9:0] ? 4'ha : _GEN_24701; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24703 = 10'h12a == _T_512[9:0] ? 4'ha : _GEN_24702; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24704 = 10'h12b == _T_512[9:0] ? 4'h0 : _GEN_24703; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24705 = 10'h12c == _T_512[9:0] ? 4'h0 : _GEN_24704; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24706 = 10'h12d == _T_512[9:0] ? 4'h0 : _GEN_24705; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24707 = 10'h12e == _T_512[9:0] ? 4'h0 : _GEN_24706; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24708 = 10'h12f == _T_512[9:0] ? 4'h0 : _GEN_24707; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24709 = 10'h130 == _T_512[9:0] ? 4'h0 : _GEN_24708; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24710 = 10'h131 == _T_512[9:0] ? 4'h0 : _GEN_24709; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24711 = 10'h132 == _T_512[9:0] ? 4'h0 : _GEN_24710; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24712 = 10'h133 == _T_512[9:0] ? 4'h0 : _GEN_24711; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24713 = 10'h134 == _T_512[9:0] ? 4'ha : _GEN_24712; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24714 = 10'h135 == _T_512[9:0] ? 4'ha : _GEN_24713; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24715 = 10'h136 == _T_512[9:0] ? 4'h0 : _GEN_24714; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24716 = 10'h137 == _T_512[9:0] ? 4'h1 : _GEN_24715; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24717 = 10'h138 == _T_512[9:0] ? 4'ha : _GEN_24716; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24718 = 10'h139 == _T_512[9:0] ? 4'ha : _GEN_24717; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24719 = 10'h13a == _T_512[9:0] ? 4'ha : _GEN_24718; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24720 = 10'h13b == _T_512[9:0] ? 4'ha : _GEN_24719; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24721 = 10'h13c == _T_512[9:0] ? 4'ha : _GEN_24720; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24722 = 10'h13d == _T_512[9:0] ? 4'ha : _GEN_24721; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24723 = 10'h13e == _T_512[9:0] ? 4'h3 : _GEN_24722; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24724 = 10'h13f == _T_512[9:0] ? 4'h0 : _GEN_24723; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24725 = 10'h140 == _T_512[9:0] ? 4'ha : _GEN_24724; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24726 = 10'h141 == _T_512[9:0] ? 4'ha : _GEN_24725; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24727 = 10'h142 == _T_512[9:0] ? 4'h2 : _GEN_24726; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24728 = 10'h143 == _T_512[9:0] ? 4'h3 : _GEN_24727; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24729 = 10'h144 == _T_512[9:0] ? 4'ha : _GEN_24728; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24730 = 10'h145 == _T_512[9:0] ? 4'ha : _GEN_24729; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24731 = 10'h146 == _T_512[9:0] ? 4'h1 : _GEN_24730; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24732 = 10'h147 == _T_512[9:0] ? 4'h0 : _GEN_24731; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24733 = 10'h148 == _T_512[9:0] ? 4'ha : _GEN_24732; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24734 = 10'h149 == _T_512[9:0] ? 4'ha : _GEN_24733; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24735 = 10'h14a == _T_512[9:0] ? 4'ha : _GEN_24734; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24736 = 10'h14b == _T_512[9:0] ? 4'ha : _GEN_24735; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24737 = 10'h14c == _T_512[9:0] ? 4'ha : _GEN_24736; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24738 = 10'h14d == _T_512[9:0] ? 4'ha : _GEN_24737; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24739 = 10'h14e == _T_512[9:0] ? 4'ha : _GEN_24738; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24740 = 10'h14f == _T_512[9:0] ? 4'ha : _GEN_24739; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24741 = 10'h150 == _T_512[9:0] ? 4'ha : _GEN_24740; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24742 = 10'h151 == _T_512[9:0] ? 4'ha : _GEN_24741; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24743 = 10'h152 == _T_512[9:0] ? 4'ha : _GEN_24742; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24744 = 10'h153 == _T_512[9:0] ? 4'ha : _GEN_24743; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24745 = 10'h154 == _T_512[9:0] ? 4'ha : _GEN_24744; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24746 = 10'h155 == _T_512[9:0] ? 4'ha : _GEN_24745; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24747 = 10'h156 == _T_512[9:0] ? 4'ha : _GEN_24746; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24748 = 10'h157 == _T_512[9:0] ? 4'h0 : _GEN_24747; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24749 = 10'h158 == _T_512[9:0] ? 4'ha : _GEN_24748; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24750 = 10'h159 == _T_512[9:0] ? 4'ha : _GEN_24749; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24751 = 10'h15a == _T_512[9:0] ? 4'ha : _GEN_24750; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24752 = 10'h15b == _T_512[9:0] ? 4'ha : _GEN_24751; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24753 = 10'h15c == _T_512[9:0] ? 4'ha : _GEN_24752; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24754 = 10'h15d == _T_512[9:0] ? 4'h3 : _GEN_24753; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24755 = 10'h15e == _T_512[9:0] ? 4'h2 : _GEN_24754; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24756 = 10'h15f == _T_512[9:0] ? 4'h0 : _GEN_24755; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24757 = 10'h160 == _T_512[9:0] ? 4'ha : _GEN_24756; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24758 = 10'h161 == _T_512[9:0] ? 4'ha : _GEN_24757; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24759 = 10'h162 == _T_512[9:0] ? 4'ha : _GEN_24758; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24760 = 10'h163 == _T_512[9:0] ? 4'h2 : _GEN_24759; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24761 = 10'h164 == _T_512[9:0] ? 4'h3 : _GEN_24760; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24762 = 10'h165 == _T_512[9:0] ? 4'h1 : _GEN_24761; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24763 = 10'h166 == _T_512[9:0] ? 4'h0 : _GEN_24762; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24764 = 10'h167 == _T_512[9:0] ? 4'h0 : _GEN_24763; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24765 = 10'h168 == _T_512[9:0] ? 4'h5 : _GEN_24764; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24766 = 10'h169 == _T_512[9:0] ? 4'h3 : _GEN_24765; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24767 = 10'h16a == _T_512[9:0] ? 4'h5 : _GEN_24766; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24768 = 10'h16b == _T_512[9:0] ? 4'h5 : _GEN_24767; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24769 = 10'h16c == _T_512[9:0] ? 4'ha : _GEN_24768; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24770 = 10'h16d == _T_512[9:0] ? 4'ha : _GEN_24769; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24771 = 10'h16e == _T_512[9:0] ? 4'ha : _GEN_24770; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24772 = 10'h16f == _T_512[9:0] ? 4'ha : _GEN_24771; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24773 = 10'h170 == _T_512[9:0] ? 4'ha : _GEN_24772; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24774 = 10'h171 == _T_512[9:0] ? 4'ha : _GEN_24773; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24775 = 10'h172 == _T_512[9:0] ? 4'ha : _GEN_24774; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24776 = 10'h173 == _T_512[9:0] ? 4'ha : _GEN_24775; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24777 = 10'h174 == _T_512[9:0] ? 4'ha : _GEN_24776; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24778 = 10'h175 == _T_512[9:0] ? 4'ha : _GEN_24777; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24779 = 10'h176 == _T_512[9:0] ? 4'h0 : _GEN_24778; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24780 = 10'h177 == _T_512[9:0] ? 4'h0 : _GEN_24779; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24781 = 10'h178 == _T_512[9:0] ? 4'h1 : _GEN_24780; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24782 = 10'h179 == _T_512[9:0] ? 4'ha : _GEN_24781; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24783 = 10'h17a == _T_512[9:0] ? 4'ha : _GEN_24782; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24784 = 10'h17b == _T_512[9:0] ? 4'ha : _GEN_24783; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24785 = 10'h17c == _T_512[9:0] ? 4'h3 : _GEN_24784; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24786 = 10'h17d == _T_512[9:0] ? 4'h2 : _GEN_24785; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24787 = 10'h17e == _T_512[9:0] ? 4'ha : _GEN_24786; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24788 = 10'h17f == _T_512[9:0] ? 4'h0 : _GEN_24787; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24789 = 10'h180 == _T_512[9:0] ? 4'h5 : _GEN_24788; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24790 = 10'h181 == _T_512[9:0] ? 4'h5 : _GEN_24789; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24791 = 10'h182 == _T_512[9:0] ? 4'h5 : _GEN_24790; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24792 = 10'h183 == _T_512[9:0] ? 4'h5 : _GEN_24791; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24793 = 10'h184 == _T_512[9:0] ? 4'h3 : _GEN_24792; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24794 = 10'h185 == _T_512[9:0] ? 4'h1 : _GEN_24793; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24795 = 10'h186 == _T_512[9:0] ? 4'hb : _GEN_24794; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24796 = 10'h187 == _T_512[9:0] ? 4'h0 : _GEN_24795; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24797 = 10'h188 == _T_512[9:0] ? 4'h5 : _GEN_24796; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24798 = 10'h189 == _T_512[9:0] ? 4'h5 : _GEN_24797; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24799 = 10'h18a == _T_512[9:0] ? 4'h5 : _GEN_24798; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24800 = 10'h18b == _T_512[9:0] ? 4'h5 : _GEN_24799; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24801 = 10'h18c == _T_512[9:0] ? 4'h5 : _GEN_24800; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24802 = 10'h18d == _T_512[9:0] ? 4'h5 : _GEN_24801; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24803 = 10'h18e == _T_512[9:0] ? 4'h5 : _GEN_24802; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24804 = 10'h18f == _T_512[9:0] ? 4'h5 : _GEN_24803; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24805 = 10'h190 == _T_512[9:0] ? 4'h5 : _GEN_24804; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24806 = 10'h191 == _T_512[9:0] ? 4'h5 : _GEN_24805; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24807 = 10'h192 == _T_512[9:0] ? 4'h3 : _GEN_24806; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24808 = 10'h193 == _T_512[9:0] ? 4'h5 : _GEN_24807; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24809 = 10'h194 == _T_512[9:0] ? 4'h5 : _GEN_24808; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24810 = 10'h195 == _T_512[9:0] ? 4'h5 : _GEN_24809; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24811 = 10'h196 == _T_512[9:0] ? 4'h0 : _GEN_24810; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24812 = 10'h197 == _T_512[9:0] ? 4'ha : _GEN_24811; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24813 = 10'h198 == _T_512[9:0] ? 4'h1 : _GEN_24812; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24814 = 10'h199 == _T_512[9:0] ? 4'ha : _GEN_24813; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24815 = 10'h19a == _T_512[9:0] ? 4'ha : _GEN_24814; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24816 = 10'h19b == _T_512[9:0] ? 4'ha : _GEN_24815; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24817 = 10'h19c == _T_512[9:0] ? 4'h3 : _GEN_24816; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24818 = 10'h19d == _T_512[9:0] ? 4'ha : _GEN_24817; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24819 = 10'h19e == _T_512[9:0] ? 4'ha : _GEN_24818; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24820 = 10'h19f == _T_512[9:0] ? 4'h0 : _GEN_24819; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24821 = 10'h1a0 == _T_512[9:0] ? 4'h5 : _GEN_24820; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24822 = 10'h1a1 == _T_512[9:0] ? 4'h5 : _GEN_24821; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24823 = 10'h1a2 == _T_512[9:0] ? 4'h3 : _GEN_24822; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24824 = 10'h1a3 == _T_512[9:0] ? 4'h5 : _GEN_24823; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24825 = 10'h1a4 == _T_512[9:0] ? 4'h3 : _GEN_24824; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24826 = 10'h1a5 == _T_512[9:0] ? 4'h0 : _GEN_24825; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24827 = 10'h1a6 == _T_512[9:0] ? 4'h5 : _GEN_24826; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24828 = 10'h1a7 == _T_512[9:0] ? 4'h0 : _GEN_24827; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24829 = 10'h1a8 == _T_512[9:0] ? 4'hb : _GEN_24828; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24830 = 10'h1a9 == _T_512[9:0] ? 4'h5 : _GEN_24829; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24831 = 10'h1aa == _T_512[9:0] ? 4'h5 : _GEN_24830; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24832 = 10'h1ab == _T_512[9:0] ? 4'h3 : _GEN_24831; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24833 = 10'h1ac == _T_512[9:0] ? 4'h5 : _GEN_24832; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24834 = 10'h1ad == _T_512[9:0] ? 4'h5 : _GEN_24833; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24835 = 10'h1ae == _T_512[9:0] ? 4'h5 : _GEN_24834; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24836 = 10'h1af == _T_512[9:0] ? 4'h5 : _GEN_24835; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24837 = 10'h1b0 == _T_512[9:0] ? 4'h5 : _GEN_24836; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24838 = 10'h1b1 == _T_512[9:0] ? 4'h5 : _GEN_24837; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24839 = 10'h1b2 == _T_512[9:0] ? 4'h5 : _GEN_24838; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24840 = 10'h1b3 == _T_512[9:0] ? 4'h5 : _GEN_24839; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24841 = 10'h1b4 == _T_512[9:0] ? 4'h5 : _GEN_24840; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24842 = 10'h1b5 == _T_512[9:0] ? 4'h5 : _GEN_24841; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24843 = 10'h1b6 == _T_512[9:0] ? 4'h0 : _GEN_24842; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24844 = 10'h1b7 == _T_512[9:0] ? 4'h5 : _GEN_24843; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24845 = 10'h1b8 == _T_512[9:0] ? 4'h0 : _GEN_24844; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24846 = 10'h1b9 == _T_512[9:0] ? 4'h5 : _GEN_24845; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24847 = 10'h1ba == _T_512[9:0] ? 4'h5 : _GEN_24846; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24848 = 10'h1bb == _T_512[9:0] ? 4'h5 : _GEN_24847; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24849 = 10'h1bc == _T_512[9:0] ? 4'h2 : _GEN_24848; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24850 = 10'h1bd == _T_512[9:0] ? 4'h3 : _GEN_24849; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24851 = 10'h1be == _T_512[9:0] ? 4'h5 : _GEN_24850; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24852 = 10'h1bf == _T_512[9:0] ? 4'h0 : _GEN_24851; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24853 = 10'h1c0 == _T_512[9:0] ? 4'h5 : _GEN_24852; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24854 = 10'h1c1 == _T_512[9:0] ? 4'h5 : _GEN_24853; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24855 = 10'h1c2 == _T_512[9:0] ? 4'h5 : _GEN_24854; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24856 = 10'h1c3 == _T_512[9:0] ? 4'h2 : _GEN_24855; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24857 = 10'h1c4 == _T_512[9:0] ? 4'h2 : _GEN_24856; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24858 = 10'h1c5 == _T_512[9:0] ? 4'h5 : _GEN_24857; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24859 = 10'h1c6 == _T_512[9:0] ? 4'h5 : _GEN_24858; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24860 = 10'h1c7 == _T_512[9:0] ? 4'h5 : _GEN_24859; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24861 = 10'h1c8 == _T_512[9:0] ? 4'h5 : _GEN_24860; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24862 = 10'h1c9 == _T_512[9:0] ? 4'hb : _GEN_24861; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24863 = 10'h1ca == _T_512[9:0] ? 4'hb : _GEN_24862; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24864 = 10'h1cb == _T_512[9:0] ? 4'hb : _GEN_24863; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24865 = 10'h1cc == _T_512[9:0] ? 4'hb : _GEN_24864; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24866 = 10'h1cd == _T_512[9:0] ? 4'hb : _GEN_24865; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24867 = 10'h1ce == _T_512[9:0] ? 4'hb : _GEN_24866; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24868 = 10'h1cf == _T_512[9:0] ? 4'hb : _GEN_24867; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24869 = 10'h1d0 == _T_512[9:0] ? 4'hb : _GEN_24868; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24870 = 10'h1d1 == _T_512[9:0] ? 4'hb : _GEN_24869; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24871 = 10'h1d2 == _T_512[9:0] ? 4'hb : _GEN_24870; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24872 = 10'h1d3 == _T_512[9:0] ? 4'hb : _GEN_24871; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24873 = 10'h1d4 == _T_512[9:0] ? 4'hb : _GEN_24872; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24874 = 10'h1d5 == _T_512[9:0] ? 4'hb : _GEN_24873; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24875 = 10'h1d6 == _T_512[9:0] ? 4'h5 : _GEN_24874; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24876 = 10'h1d7 == _T_512[9:0] ? 4'h5 : _GEN_24875; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24877 = 10'h1d8 == _T_512[9:0] ? 4'h5 : _GEN_24876; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24878 = 10'h1d9 == _T_512[9:0] ? 4'h5 : _GEN_24877; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24879 = 10'h1da == _T_512[9:0] ? 4'h5 : _GEN_24878; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24880 = 10'h1db == _T_512[9:0] ? 4'h5 : _GEN_24879; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24881 = 10'h1dc == _T_512[9:0] ? 4'h5 : _GEN_24880; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24882 = 10'h1dd == _T_512[9:0] ? 4'h3 : _GEN_24881; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24883 = 10'h1de == _T_512[9:0] ? 4'h5 : _GEN_24882; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24884 = 10'h1df == _T_512[9:0] ? 4'h0 : _GEN_24883; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24885 = 10'h1e0 == _T_512[9:0] ? 4'h3 : _GEN_24884; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24886 = 10'h1e1 == _T_512[9:0] ? 4'h5 : _GEN_24885; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24887 = 10'h1e2 == _T_512[9:0] ? 4'h2 : _GEN_24886; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24888 = 10'h1e3 == _T_512[9:0] ? 4'h2 : _GEN_24887; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24889 = 10'h1e4 == _T_512[9:0] ? 4'h5 : _GEN_24888; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24890 = 10'h1e5 == _T_512[9:0] ? 4'h5 : _GEN_24889; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24891 = 10'h1e6 == _T_512[9:0] ? 4'h5 : _GEN_24890; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24892 = 10'h1e7 == _T_512[9:0] ? 4'h5 : _GEN_24891; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24893 = 10'h1e8 == _T_512[9:0] ? 4'hb : _GEN_24892; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24894 = 10'h1e9 == _T_512[9:0] ? 4'h5 : _GEN_24893; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24895 = 10'h1ea == _T_512[9:0] ? 4'h5 : _GEN_24894; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24896 = 10'h1eb == _T_512[9:0] ? 4'hb : _GEN_24895; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24897 = 10'h1ec == _T_512[9:0] ? 4'h5 : _GEN_24896; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24898 = 10'h1ed == _T_512[9:0] ? 4'hb : _GEN_24897; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24899 = 10'h1ee == _T_512[9:0] ? 4'h5 : _GEN_24898; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24900 = 10'h1ef == _T_512[9:0] ? 4'hb : _GEN_24899; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24901 = 10'h1f0 == _T_512[9:0] ? 4'h5 : _GEN_24900; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24902 = 10'h1f1 == _T_512[9:0] ? 4'hb : _GEN_24901; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24903 = 10'h1f2 == _T_512[9:0] ? 4'hb : _GEN_24902; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24904 = 10'h1f3 == _T_512[9:0] ? 4'h5 : _GEN_24903; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24905 = 10'h1f4 == _T_512[9:0] ? 4'hb : _GEN_24904; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24906 = 10'h1f5 == _T_512[9:0] ? 4'hb : _GEN_24905; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24907 = 10'h1f6 == _T_512[9:0] ? 4'h5 : _GEN_24906; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24908 = 10'h1f7 == _T_512[9:0] ? 4'h5 : _GEN_24907; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24909 = 10'h1f8 == _T_512[9:0] ? 4'h5 : _GEN_24908; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24910 = 10'h1f9 == _T_512[9:0] ? 4'h5 : _GEN_24909; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24911 = 10'h1fa == _T_512[9:0] ? 4'h3 : _GEN_24910; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24912 = 10'h1fb == _T_512[9:0] ? 4'h5 : _GEN_24911; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24913 = 10'h1fc == _T_512[9:0] ? 4'h5 : _GEN_24912; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24914 = 10'h1fd == _T_512[9:0] ? 4'h2 : _GEN_24913; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24915 = 10'h1fe == _T_512[9:0] ? 4'h5 : _GEN_24914; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24916 = 10'h1ff == _T_512[9:0] ? 4'h0 : _GEN_24915; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24917 = 10'h200 == _T_512[9:0] ? 4'h5 : _GEN_24916; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24918 = 10'h201 == _T_512[9:0] ? 4'h5 : _GEN_24917; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24919 = 10'h202 == _T_512[9:0] ? 4'h3 : _GEN_24918; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24920 = 10'h203 == _T_512[9:0] ? 4'h5 : _GEN_24919; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24921 = 10'h204 == _T_512[9:0] ? 4'h5 : _GEN_24920; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24922 = 10'h205 == _T_512[9:0] ? 4'h5 : _GEN_24921; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24923 = 10'h206 == _T_512[9:0] ? 4'hb : _GEN_24922; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24924 = 10'h207 == _T_512[9:0] ? 4'hb : _GEN_24923; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24925 = 10'h208 == _T_512[9:0] ? 4'h5 : _GEN_24924; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24926 = 10'h209 == _T_512[9:0] ? 4'h5 : _GEN_24925; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24927 = 10'h20a == _T_512[9:0] ? 4'h5 : _GEN_24926; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24928 = 10'h20b == _T_512[9:0] ? 4'hb : _GEN_24927; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24929 = 10'h20c == _T_512[9:0] ? 4'h5 : _GEN_24928; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24930 = 10'h20d == _T_512[9:0] ? 4'hb : _GEN_24929; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24931 = 10'h20e == _T_512[9:0] ? 4'h5 : _GEN_24930; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24932 = 10'h20f == _T_512[9:0] ? 4'hb : _GEN_24931; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24933 = 10'h210 == _T_512[9:0] ? 4'h5 : _GEN_24932; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24934 = 10'h211 == _T_512[9:0] ? 4'h5 : _GEN_24933; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24935 = 10'h212 == _T_512[9:0] ? 4'hb : _GEN_24934; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24936 = 10'h213 == _T_512[9:0] ? 4'hb : _GEN_24935; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24937 = 10'h214 == _T_512[9:0] ? 4'hb : _GEN_24936; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24938 = 10'h215 == _T_512[9:0] ? 4'h5 : _GEN_24937; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24939 = 10'h216 == _T_512[9:0] ? 4'h5 : _GEN_24938; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24940 = 10'h217 == _T_512[9:0] ? 4'h5 : _GEN_24939; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24941 = 10'h218 == _T_512[9:0] ? 4'h5 : _GEN_24940; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24942 = 10'h219 == _T_512[9:0] ? 4'h5 : _GEN_24941; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24943 = 10'h21a == _T_512[9:0] ? 4'h5 : _GEN_24942; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24944 = 10'h21b == _T_512[9:0] ? 4'h5 : _GEN_24943; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24945 = 10'h21c == _T_512[9:0] ? 4'h3 : _GEN_24944; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24946 = 10'h21d == _T_512[9:0] ? 4'h2 : _GEN_24945; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24947 = 10'h21e == _T_512[9:0] ? 4'h5 : _GEN_24946; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24948 = 10'h21f == _T_512[9:0] ? 4'h0 : _GEN_24947; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24949 = 10'h220 == _T_512[9:0] ? 4'h0 : _GEN_24948; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24950 = 10'h221 == _T_512[9:0] ? 4'h0 : _GEN_24949; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24951 = 10'h222 == _T_512[9:0] ? 4'h0 : _GEN_24950; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24952 = 10'h223 == _T_512[9:0] ? 4'h0 : _GEN_24951; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24953 = 10'h224 == _T_512[9:0] ? 4'h0 : _GEN_24952; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24954 = 10'h225 == _T_512[9:0] ? 4'h0 : _GEN_24953; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24955 = 10'h226 == _T_512[9:0] ? 4'h0 : _GEN_24954; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24956 = 10'h227 == _T_512[9:0] ? 4'h0 : _GEN_24955; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24957 = 10'h228 == _T_512[9:0] ? 4'h0 : _GEN_24956; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24958 = 10'h229 == _T_512[9:0] ? 4'h0 : _GEN_24957; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24959 = 10'h22a == _T_512[9:0] ? 4'h0 : _GEN_24958; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24960 = 10'h22b == _T_512[9:0] ? 4'h0 : _GEN_24959; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24961 = 10'h22c == _T_512[9:0] ? 4'h0 : _GEN_24960; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24962 = 10'h22d == _T_512[9:0] ? 4'h0 : _GEN_24961; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24963 = 10'h22e == _T_512[9:0] ? 4'h0 : _GEN_24962; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24964 = 10'h22f == _T_512[9:0] ? 4'h0 : _GEN_24963; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24965 = 10'h230 == _T_512[9:0] ? 4'h0 : _GEN_24964; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24966 = 10'h231 == _T_512[9:0] ? 4'h0 : _GEN_24965; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24967 = 10'h232 == _T_512[9:0] ? 4'h0 : _GEN_24966; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24968 = 10'h233 == _T_512[9:0] ? 4'h0 : _GEN_24967; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24969 = 10'h234 == _T_512[9:0] ? 4'h0 : _GEN_24968; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24970 = 10'h235 == _T_512[9:0] ? 4'h0 : _GEN_24969; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24971 = 10'h236 == _T_512[9:0] ? 4'h0 : _GEN_24970; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24972 = 10'h237 == _T_512[9:0] ? 4'h0 : _GEN_24971; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24973 = 10'h238 == _T_512[9:0] ? 4'h0 : _GEN_24972; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24974 = 10'h239 == _T_512[9:0] ? 4'h0 : _GEN_24973; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24975 = 10'h23a == _T_512[9:0] ? 4'h0 : _GEN_24974; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24976 = 10'h23b == _T_512[9:0] ? 4'h0 : _GEN_24975; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24977 = 10'h23c == _T_512[9:0] ? 4'h0 : _GEN_24976; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24978 = 10'h23d == _T_512[9:0] ? 4'h0 : _GEN_24977; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24979 = 10'h23e == _T_512[9:0] ? 4'h0 : _GEN_24978; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24980 = 10'h23f == _T_512[9:0] ? 4'h0 : _GEN_24979; // @[Filter.scala 191:62]
  wire [4:0] _GEN_28382 = {{1'd0}, _GEN_24980}; // @[Filter.scala 191:62]
  wire [8:0] _T_514 = _GEN_28382 * 5'h14; // @[Filter.scala 191:62]
  wire [3:0] _GEN_24984 = 10'h3 == _T_512[9:0] ? 4'ha : 4'h3; // @[Filter.scala 191:102]
  wire [3:0] _GEN_24985 = 10'h4 == _T_512[9:0] ? 4'h3 : _GEN_24984; // @[Filter.scala 191:102]
  wire [3:0] _GEN_24986 = 10'h5 == _T_512[9:0] ? 4'h3 : _GEN_24985; // @[Filter.scala 191:102]
  wire [3:0] _GEN_24987 = 10'h6 == _T_512[9:0] ? 4'h3 : _GEN_24986; // @[Filter.scala 191:102]
  wire [3:0] _GEN_24988 = 10'h7 == _T_512[9:0] ? 4'h3 : _GEN_24987; // @[Filter.scala 191:102]
  wire [3:0] _GEN_24989 = 10'h8 == _T_512[9:0] ? 4'h3 : _GEN_24988; // @[Filter.scala 191:102]
  wire [3:0] _GEN_24990 = 10'h9 == _T_512[9:0] ? 4'h3 : _GEN_24989; // @[Filter.scala 191:102]
  wire [3:0] _GEN_24991 = 10'ha == _T_512[9:0] ? 4'h3 : _GEN_24990; // @[Filter.scala 191:102]
  wire [3:0] _GEN_24992 = 10'hb == _T_512[9:0] ? 4'h3 : _GEN_24991; // @[Filter.scala 191:102]
  wire [3:0] _GEN_24993 = 10'hc == _T_512[9:0] ? 4'h5 : _GEN_24992; // @[Filter.scala 191:102]
  wire [3:0] _GEN_24994 = 10'hd == _T_512[9:0] ? 4'h3 : _GEN_24993; // @[Filter.scala 191:102]
  wire [3:0] _GEN_24995 = 10'he == _T_512[9:0] ? 4'h3 : _GEN_24994; // @[Filter.scala 191:102]
  wire [3:0] _GEN_24996 = 10'hf == _T_512[9:0] ? 4'h3 : _GEN_24995; // @[Filter.scala 191:102]
  wire [3:0] _GEN_24997 = 10'h10 == _T_512[9:0] ? 4'h3 : _GEN_24996; // @[Filter.scala 191:102]
  wire [3:0] _GEN_24998 = 10'h11 == _T_512[9:0] ? 4'h3 : _GEN_24997; // @[Filter.scala 191:102]
  wire [3:0] _GEN_24999 = 10'h12 == _T_512[9:0] ? 4'h3 : _GEN_24998; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25000 = 10'h13 == _T_512[9:0] ? 4'h3 : _GEN_24999; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25001 = 10'h14 == _T_512[9:0] ? 4'h3 : _GEN_25000; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25002 = 10'h15 == _T_512[9:0] ? 4'h3 : _GEN_25001; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25003 = 10'h16 == _T_512[9:0] ? 4'h3 : _GEN_25002; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25004 = 10'h17 == _T_512[9:0] ? 4'h3 : _GEN_25003; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25005 = 10'h18 == _T_512[9:0] ? 4'h3 : _GEN_25004; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25006 = 10'h19 == _T_512[9:0] ? 4'h3 : _GEN_25005; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25007 = 10'h1a == _T_512[9:0] ? 4'h3 : _GEN_25006; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25008 = 10'h1b == _T_512[9:0] ? 4'h3 : _GEN_25007; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25009 = 10'h1c == _T_512[9:0] ? 4'h3 : _GEN_25008; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25010 = 10'h1d == _T_512[9:0] ? 4'h3 : _GEN_25009; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25011 = 10'h1e == _T_512[9:0] ? 4'h3 : _GEN_25010; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25012 = 10'h1f == _T_512[9:0] ? 4'h0 : _GEN_25011; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25013 = 10'h20 == _T_512[9:0] ? 4'h3 : _GEN_25012; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25014 = 10'h21 == _T_512[9:0] ? 4'h5 : _GEN_25013; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25015 = 10'h22 == _T_512[9:0] ? 4'h3 : _GEN_25014; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25016 = 10'h23 == _T_512[9:0] ? 4'ha : _GEN_25015; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25017 = 10'h24 == _T_512[9:0] ? 4'h3 : _GEN_25016; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25018 = 10'h25 == _T_512[9:0] ? 4'h3 : _GEN_25017; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25019 = 10'h26 == _T_512[9:0] ? 4'h3 : _GEN_25018; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25020 = 10'h27 == _T_512[9:0] ? 4'h1 : _GEN_25019; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25021 = 10'h28 == _T_512[9:0] ? 4'h1 : _GEN_25020; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25022 = 10'h29 == _T_512[9:0] ? 4'h3 : _GEN_25021; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25023 = 10'h2a == _T_512[9:0] ? 4'h3 : _GEN_25022; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25024 = 10'h2b == _T_512[9:0] ? 4'h3 : _GEN_25023; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25025 = 10'h2c == _T_512[9:0] ? 4'h3 : _GEN_25024; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25026 = 10'h2d == _T_512[9:0] ? 4'h3 : _GEN_25025; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25027 = 10'h2e == _T_512[9:0] ? 4'h3 : _GEN_25026; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25028 = 10'h2f == _T_512[9:0] ? 4'h3 : _GEN_25027; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25029 = 10'h30 == _T_512[9:0] ? 4'h3 : _GEN_25028; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25030 = 10'h31 == _T_512[9:0] ? 4'h5 : _GEN_25029; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25031 = 10'h32 == _T_512[9:0] ? 4'h3 : _GEN_25030; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25032 = 10'h33 == _T_512[9:0] ? 4'h3 : _GEN_25031; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25033 = 10'h34 == _T_512[9:0] ? 4'h3 : _GEN_25032; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25034 = 10'h35 == _T_512[9:0] ? 4'h3 : _GEN_25033; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25035 = 10'h36 == _T_512[9:0] ? 4'h3 : _GEN_25034; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25036 = 10'h37 == _T_512[9:0] ? 4'h1 : _GEN_25035; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25037 = 10'h38 == _T_512[9:0] ? 4'h1 : _GEN_25036; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25038 = 10'h39 == _T_512[9:0] ? 4'h3 : _GEN_25037; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25039 = 10'h3a == _T_512[9:0] ? 4'h3 : _GEN_25038; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25040 = 10'h3b == _T_512[9:0] ? 4'h5 : _GEN_25039; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25041 = 10'h3c == _T_512[9:0] ? 4'h3 : _GEN_25040; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25042 = 10'h3d == _T_512[9:0] ? 4'ha : _GEN_25041; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25043 = 10'h3e == _T_512[9:0] ? 4'h3 : _GEN_25042; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25044 = 10'h3f == _T_512[9:0] ? 4'h0 : _GEN_25043; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25045 = 10'h40 == _T_512[9:0] ? 4'h3 : _GEN_25044; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25046 = 10'h41 == _T_512[9:0] ? 4'h3 : _GEN_25045; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25047 = 10'h42 == _T_512[9:0] ? 4'h3 : _GEN_25046; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25048 = 10'h43 == _T_512[9:0] ? 4'h7 : _GEN_25047; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25049 = 10'h44 == _T_512[9:0] ? 4'ha : _GEN_25048; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25050 = 10'h45 == _T_512[9:0] ? 4'h0 : _GEN_25049; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25051 = 10'h46 == _T_512[9:0] ? 4'h0 : _GEN_25050; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25052 = 10'h47 == _T_512[9:0] ? 4'h0 : _GEN_25051; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25053 = 10'h48 == _T_512[9:0] ? 4'h0 : _GEN_25052; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25054 = 10'h49 == _T_512[9:0] ? 4'h3 : _GEN_25053; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25055 = 10'h4a == _T_512[9:0] ? 4'h3 : _GEN_25054; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25056 = 10'h4b == _T_512[9:0] ? 4'h3 : _GEN_25055; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25057 = 10'h4c == _T_512[9:0] ? 4'h3 : _GEN_25056; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25058 = 10'h4d == _T_512[9:0] ? 4'h5 : _GEN_25057; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25059 = 10'h4e == _T_512[9:0] ? 4'h3 : _GEN_25058; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25060 = 10'h4f == _T_512[9:0] ? 4'h3 : _GEN_25059; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25061 = 10'h50 == _T_512[9:0] ? 4'h3 : _GEN_25060; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25062 = 10'h51 == _T_512[9:0] ? 4'h3 : _GEN_25061; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25063 = 10'h52 == _T_512[9:0] ? 4'h3 : _GEN_25062; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25064 = 10'h53 == _T_512[9:0] ? 4'h3 : _GEN_25063; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25065 = 10'h54 == _T_512[9:0] ? 4'h1 : _GEN_25064; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25066 = 10'h55 == _T_512[9:0] ? 4'h1 : _GEN_25065; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25067 = 10'h56 == _T_512[9:0] ? 4'h1 : _GEN_25066; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25068 = 10'h57 == _T_512[9:0] ? 4'h0 : _GEN_25067; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25069 = 10'h58 == _T_512[9:0] ? 4'h3 : _GEN_25068; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25070 = 10'h59 == _T_512[9:0] ? 4'h0 : _GEN_25069; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25071 = 10'h5a == _T_512[9:0] ? 4'h3 : _GEN_25070; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25072 = 10'h5b == _T_512[9:0] ? 4'h3 : _GEN_25071; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25073 = 10'h5c == _T_512[9:0] ? 4'h3 : _GEN_25072; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25074 = 10'h5d == _T_512[9:0] ? 4'ha : _GEN_25073; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25075 = 10'h5e == _T_512[9:0] ? 4'h3 : _GEN_25074; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25076 = 10'h5f == _T_512[9:0] ? 4'h0 : _GEN_25075; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25077 = 10'h60 == _T_512[9:0] ? 4'h3 : _GEN_25076; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25078 = 10'h61 == _T_512[9:0] ? 4'h3 : _GEN_25077; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25079 = 10'h62 == _T_512[9:0] ? 4'h3 : _GEN_25078; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25080 = 10'h63 == _T_512[9:0] ? 4'h3 : _GEN_25079; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25081 = 10'h64 == _T_512[9:0] ? 4'ha : _GEN_25080; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25082 = 10'h65 == _T_512[9:0] ? 4'h0 : _GEN_25081; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25083 = 10'h66 == _T_512[9:0] ? 4'h3 : _GEN_25082; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25084 = 10'h67 == _T_512[9:0] ? 4'h3 : _GEN_25083; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25085 = 10'h68 == _T_512[9:0] ? 4'h3 : _GEN_25084; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25086 = 10'h69 == _T_512[9:0] ? 4'h0 : _GEN_25085; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25087 = 10'h6a == _T_512[9:0] ? 4'h1 : _GEN_25086; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25088 = 10'h6b == _T_512[9:0] ? 4'h1 : _GEN_25087; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25089 = 10'h6c == _T_512[9:0] ? 4'h3 : _GEN_25088; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25090 = 10'h6d == _T_512[9:0] ? 4'h3 : _GEN_25089; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25091 = 10'h6e == _T_512[9:0] ? 4'h3 : _GEN_25090; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25092 = 10'h6f == _T_512[9:0] ? 4'h3 : _GEN_25091; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25093 = 10'h70 == _T_512[9:0] ? 4'h3 : _GEN_25092; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25094 = 10'h71 == _T_512[9:0] ? 4'h3 : _GEN_25093; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25095 = 10'h72 == _T_512[9:0] ? 4'h3 : _GEN_25094; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25096 = 10'h73 == _T_512[9:0] ? 4'h1 : _GEN_25095; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25097 = 10'h74 == _T_512[9:0] ? 4'h0 : _GEN_25096; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25098 = 10'h75 == _T_512[9:0] ? 4'h0 : _GEN_25097; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25099 = 10'h76 == _T_512[9:0] ? 4'h0 : _GEN_25098; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25100 = 10'h77 == _T_512[9:0] ? 4'h3 : _GEN_25099; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25101 = 10'h78 == _T_512[9:0] ? 4'h3 : _GEN_25100; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25102 = 10'h79 == _T_512[9:0] ? 4'h3 : _GEN_25101; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25103 = 10'h7a == _T_512[9:0] ? 4'h0 : _GEN_25102; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25104 = 10'h7b == _T_512[9:0] ? 4'h3 : _GEN_25103; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25105 = 10'h7c == _T_512[9:0] ? 4'h3 : _GEN_25104; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25106 = 10'h7d == _T_512[9:0] ? 4'h7 : _GEN_25105; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25107 = 10'h7e == _T_512[9:0] ? 4'ha : _GEN_25106; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25108 = 10'h7f == _T_512[9:0] ? 4'h0 : _GEN_25107; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25109 = 10'h80 == _T_512[9:0] ? 4'h3 : _GEN_25108; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25110 = 10'h81 == _T_512[9:0] ? 4'h3 : _GEN_25109; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25111 = 10'h82 == _T_512[9:0] ? 4'h1 : _GEN_25110; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25112 = 10'h83 == _T_512[9:0] ? 4'h0 : _GEN_25111; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25113 = 10'h84 == _T_512[9:0] ? 4'h7 : _GEN_25112; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25114 = 10'h85 == _T_512[9:0] ? 4'h1 : _GEN_25113; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25115 = 10'h86 == _T_512[9:0] ? 4'h1 : _GEN_25114; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25116 = 10'h87 == _T_512[9:0] ? 4'h3 : _GEN_25115; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25117 = 10'h88 == _T_512[9:0] ? 4'h3 : _GEN_25116; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25118 = 10'h89 == _T_512[9:0] ? 4'h0 : _GEN_25117; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25119 = 10'h8a == _T_512[9:0] ? 4'h0 : _GEN_25118; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25120 = 10'h8b == _T_512[9:0] ? 4'h1 : _GEN_25119; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25121 = 10'h8c == _T_512[9:0] ? 4'h1 : _GEN_25120; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25122 = 10'h8d == _T_512[9:0] ? 4'h1 : _GEN_25121; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25123 = 10'h8e == _T_512[9:0] ? 4'h1 : _GEN_25122; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25124 = 10'h8f == _T_512[9:0] ? 4'h1 : _GEN_25123; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25125 = 10'h90 == _T_512[9:0] ? 4'h1 : _GEN_25124; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25126 = 10'h91 == _T_512[9:0] ? 4'h1 : _GEN_25125; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25127 = 10'h92 == _T_512[9:0] ? 4'h1 : _GEN_25126; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25128 = 10'h93 == _T_512[9:0] ? 4'h0 : _GEN_25127; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25129 = 10'h94 == _T_512[9:0] ? 4'h0 : _GEN_25128; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25130 = 10'h95 == _T_512[9:0] ? 4'h3 : _GEN_25129; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25131 = 10'h96 == _T_512[9:0] ? 4'h3 : _GEN_25130; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25132 = 10'h97 == _T_512[9:0] ? 4'h3 : _GEN_25131; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25133 = 10'h98 == _T_512[9:0] ? 4'h1 : _GEN_25132; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25134 = 10'h99 == _T_512[9:0] ? 4'h0 : _GEN_25133; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25135 = 10'h9a == _T_512[9:0] ? 4'h1 : _GEN_25134; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25136 = 10'h9b == _T_512[9:0] ? 4'h1 : _GEN_25135; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25137 = 10'h9c == _T_512[9:0] ? 4'h3 : _GEN_25136; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25138 = 10'h9d == _T_512[9:0] ? 4'h3 : _GEN_25137; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25139 = 10'h9e == _T_512[9:0] ? 4'ha : _GEN_25138; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25140 = 10'h9f == _T_512[9:0] ? 4'h0 : _GEN_25139; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25141 = 10'ha0 == _T_512[9:0] ? 4'h3 : _GEN_25140; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25142 = 10'ha1 == _T_512[9:0] ? 4'h1 : _GEN_25141; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25143 = 10'ha2 == _T_512[9:0] ? 4'h0 : _GEN_25142; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25144 = 10'ha3 == _T_512[9:0] ? 4'ha : _GEN_25143; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25145 = 10'ha4 == _T_512[9:0] ? 4'h3 : _GEN_25144; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25146 = 10'ha5 == _T_512[9:0] ? 4'h3 : _GEN_25145; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25147 = 10'ha6 == _T_512[9:0] ? 4'h3 : _GEN_25146; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25148 = 10'ha7 == _T_512[9:0] ? 4'h0 : _GEN_25147; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25149 = 10'ha8 == _T_512[9:0] ? 4'h3 : _GEN_25148; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25150 = 10'ha9 == _T_512[9:0] ? 4'h1 : _GEN_25149; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25151 = 10'haa == _T_512[9:0] ? 4'h0 : _GEN_25150; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25152 = 10'hab == _T_512[9:0] ? 4'h0 : _GEN_25151; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25153 = 10'hac == _T_512[9:0] ? 4'h0 : _GEN_25152; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25154 = 10'had == _T_512[9:0] ? 4'h0 : _GEN_25153; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25155 = 10'hae == _T_512[9:0] ? 4'h0 : _GEN_25154; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25156 = 10'haf == _T_512[9:0] ? 4'h0 : _GEN_25155; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25157 = 10'hb0 == _T_512[9:0] ? 4'h0 : _GEN_25156; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25158 = 10'hb1 == _T_512[9:0] ? 4'h0 : _GEN_25157; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25159 = 10'hb2 == _T_512[9:0] ? 4'h0 : _GEN_25158; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25160 = 10'hb3 == _T_512[9:0] ? 4'h0 : _GEN_25159; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25161 = 10'hb4 == _T_512[9:0] ? 4'h1 : _GEN_25160; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25162 = 10'hb5 == _T_512[9:0] ? 4'h1 : _GEN_25161; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25163 = 10'hb6 == _T_512[9:0] ? 4'h3 : _GEN_25162; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25164 = 10'hb7 == _T_512[9:0] ? 4'h0 : _GEN_25163; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25165 = 10'hb8 == _T_512[9:0] ? 4'h3 : _GEN_25164; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25166 = 10'hb9 == _T_512[9:0] ? 4'h3 : _GEN_25165; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25167 = 10'hba == _T_512[9:0] ? 4'h3 : _GEN_25166; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25168 = 10'hbb == _T_512[9:0] ? 4'h0 : _GEN_25167; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25169 = 10'hbc == _T_512[9:0] ? 4'h3 : _GEN_25168; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25170 = 10'hbd == _T_512[9:0] ? 4'h3 : _GEN_25169; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25171 = 10'hbe == _T_512[9:0] ? 4'ha : _GEN_25170; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25172 = 10'hbf == _T_512[9:0] ? 4'h0 : _GEN_25171; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25173 = 10'hc0 == _T_512[9:0] ? 4'h3 : _GEN_25172; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25174 = 10'hc1 == _T_512[9:0] ? 4'h3 : _GEN_25173; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25175 = 10'hc2 == _T_512[9:0] ? 4'ha : _GEN_25174; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25176 = 10'hc3 == _T_512[9:0] ? 4'h7 : _GEN_25175; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25177 = 10'hc4 == _T_512[9:0] ? 4'h0 : _GEN_25176; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25178 = 10'hc5 == _T_512[9:0] ? 4'h0 : _GEN_25177; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25179 = 10'hc6 == _T_512[9:0] ? 4'h0 : _GEN_25178; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25180 = 10'hc7 == _T_512[9:0] ? 4'h3 : _GEN_25179; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25181 = 10'hc8 == _T_512[9:0] ? 4'h1 : _GEN_25180; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25182 = 10'hc9 == _T_512[9:0] ? 4'h0 : _GEN_25181; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25183 = 10'hca == _T_512[9:0] ? 4'h0 : _GEN_25182; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25184 = 10'hcb == _T_512[9:0] ? 4'h0 : _GEN_25183; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25185 = 10'hcc == _T_512[9:0] ? 4'h0 : _GEN_25184; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25186 = 10'hcd == _T_512[9:0] ? 4'h0 : _GEN_25185; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25187 = 10'hce == _T_512[9:0] ? 4'h0 : _GEN_25186; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25188 = 10'hcf == _T_512[9:0] ? 4'h0 : _GEN_25187; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25189 = 10'hd0 == _T_512[9:0] ? 4'h0 : _GEN_25188; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25190 = 10'hd1 == _T_512[9:0] ? 4'h0 : _GEN_25189; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25191 = 10'hd2 == _T_512[9:0] ? 4'h0 : _GEN_25190; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25192 = 10'hd3 == _T_512[9:0] ? 4'h0 : _GEN_25191; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25193 = 10'hd4 == _T_512[9:0] ? 4'h0 : _GEN_25192; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25194 = 10'hd5 == _T_512[9:0] ? 4'h0 : _GEN_25193; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25195 = 10'hd6 == _T_512[9:0] ? 4'h1 : _GEN_25194; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25196 = 10'hd7 == _T_512[9:0] ? 4'h3 : _GEN_25195; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25197 = 10'hd8 == _T_512[9:0] ? 4'h0 : _GEN_25196; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25198 = 10'hd9 == _T_512[9:0] ? 4'h3 : _GEN_25197; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25199 = 10'hda == _T_512[9:0] ? 4'h3 : _GEN_25198; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25200 = 10'hdb == _T_512[9:0] ? 4'h3 : _GEN_25199; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25201 = 10'hdc == _T_512[9:0] ? 4'h3 : _GEN_25200; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25202 = 10'hdd == _T_512[9:0] ? 4'ha : _GEN_25201; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25203 = 10'hde == _T_512[9:0] ? 4'h7 : _GEN_25202; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25204 = 10'hdf == _T_512[9:0] ? 4'h0 : _GEN_25203; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25205 = 10'he0 == _T_512[9:0] ? 4'h3 : _GEN_25204; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25206 = 10'he1 == _T_512[9:0] ? 4'h3 : _GEN_25205; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25207 = 10'he2 == _T_512[9:0] ? 4'ha : _GEN_25206; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25208 = 10'he3 == _T_512[9:0] ? 4'h3 : _GEN_25207; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25209 = 10'he4 == _T_512[9:0] ? 4'h3 : _GEN_25208; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25210 = 10'he5 == _T_512[9:0] ? 4'h3 : _GEN_25209; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25211 = 10'he6 == _T_512[9:0] ? 4'h3 : _GEN_25210; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25212 = 10'he7 == _T_512[9:0] ? 4'h1 : _GEN_25211; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25213 = 10'he8 == _T_512[9:0] ? 4'h1 : _GEN_25212; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25214 = 10'he9 == _T_512[9:0] ? 4'h1 : _GEN_25213; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25215 = 10'hea == _T_512[9:0] ? 4'h0 : _GEN_25214; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25216 = 10'heb == _T_512[9:0] ? 4'h0 : _GEN_25215; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25217 = 10'hec == _T_512[9:0] ? 4'h0 : _GEN_25216; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25218 = 10'hed == _T_512[9:0] ? 4'h0 : _GEN_25217; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25219 = 10'hee == _T_512[9:0] ? 4'h0 : _GEN_25218; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25220 = 10'hef == _T_512[9:0] ? 4'h0 : _GEN_25219; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25221 = 10'hf0 == _T_512[9:0] ? 4'h0 : _GEN_25220; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25222 = 10'hf1 == _T_512[9:0] ? 4'h0 : _GEN_25221; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25223 = 10'hf2 == _T_512[9:0] ? 4'h0 : _GEN_25222; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25224 = 10'hf3 == _T_512[9:0] ? 4'h0 : _GEN_25223; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25225 = 10'hf4 == _T_512[9:0] ? 4'h0 : _GEN_25224; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25226 = 10'hf5 == _T_512[9:0] ? 4'h1 : _GEN_25225; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25227 = 10'hf6 == _T_512[9:0] ? 4'h0 : _GEN_25226; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25228 = 10'hf7 == _T_512[9:0] ? 4'h0 : _GEN_25227; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25229 = 10'hf8 == _T_512[9:0] ? 4'h1 : _GEN_25228; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25230 = 10'hf9 == _T_512[9:0] ? 4'h0 : _GEN_25229; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25231 = 10'hfa == _T_512[9:0] ? 4'h3 : _GEN_25230; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25232 = 10'hfb == _T_512[9:0] ? 4'h3 : _GEN_25231; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25233 = 10'hfc == _T_512[9:0] ? 4'h3 : _GEN_25232; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25234 = 10'hfd == _T_512[9:0] ? 4'ha : _GEN_25233; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25235 = 10'hfe == _T_512[9:0] ? 4'h3 : _GEN_25234; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25236 = 10'hff == _T_512[9:0] ? 4'h0 : _GEN_25235; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25237 = 10'h100 == _T_512[9:0] ? 4'h3 : _GEN_25236; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25238 = 10'h101 == _T_512[9:0] ? 4'h0 : _GEN_25237; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25239 = 10'h102 == _T_512[9:0] ? 4'ha : _GEN_25238; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25240 = 10'h103 == _T_512[9:0] ? 4'h3 : _GEN_25239; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25241 = 10'h104 == _T_512[9:0] ? 4'h3 : _GEN_25240; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25242 = 10'h105 == _T_512[9:0] ? 4'h3 : _GEN_25241; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25243 = 10'h106 == _T_512[9:0] ? 4'h3 : _GEN_25242; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25244 = 10'h107 == _T_512[9:0] ? 4'h3 : _GEN_25243; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25245 = 10'h108 == _T_512[9:0] ? 4'h1 : _GEN_25244; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25246 = 10'h109 == _T_512[9:0] ? 4'h0 : _GEN_25245; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25247 = 10'h10a == _T_512[9:0] ? 4'h0 : _GEN_25246; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25248 = 10'h10b == _T_512[9:0] ? 4'h0 : _GEN_25247; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25249 = 10'h10c == _T_512[9:0] ? 4'h0 : _GEN_25248; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25250 = 10'h10d == _T_512[9:0] ? 4'h0 : _GEN_25249; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25251 = 10'h10e == _T_512[9:0] ? 4'h0 : _GEN_25250; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25252 = 10'h10f == _T_512[9:0] ? 4'h0 : _GEN_25251; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25253 = 10'h110 == _T_512[9:0] ? 4'h0 : _GEN_25252; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25254 = 10'h111 == _T_512[9:0] ? 4'h0 : _GEN_25253; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25255 = 10'h112 == _T_512[9:0] ? 4'h0 : _GEN_25254; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25256 = 10'h113 == _T_512[9:0] ? 4'h0 : _GEN_25255; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25257 = 10'h114 == _T_512[9:0] ? 4'h0 : _GEN_25256; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25258 = 10'h115 == _T_512[9:0] ? 4'h0 : _GEN_25257; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25259 = 10'h116 == _T_512[9:0] ? 4'h1 : _GEN_25258; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25260 = 10'h117 == _T_512[9:0] ? 4'h3 : _GEN_25259; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25261 = 10'h118 == _T_512[9:0] ? 4'h3 : _GEN_25260; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25262 = 10'h119 == _T_512[9:0] ? 4'h3 : _GEN_25261; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25263 = 10'h11a == _T_512[9:0] ? 4'h0 : _GEN_25262; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25264 = 10'h11b == _T_512[9:0] ? 4'h3 : _GEN_25263; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25265 = 10'h11c == _T_512[9:0] ? 4'h3 : _GEN_25264; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25266 = 10'h11d == _T_512[9:0] ? 4'h7 : _GEN_25265; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25267 = 10'h11e == _T_512[9:0] ? 4'ha : _GEN_25266; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25268 = 10'h11f == _T_512[9:0] ? 4'h0 : _GEN_25267; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25269 = 10'h120 == _T_512[9:0] ? 4'h3 : _GEN_25268; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25270 = 10'h121 == _T_512[9:0] ? 4'h3 : _GEN_25269; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25271 = 10'h122 == _T_512[9:0] ? 4'ha : _GEN_25270; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25272 = 10'h123 == _T_512[9:0] ? 4'h3 : _GEN_25271; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25273 = 10'h124 == _T_512[9:0] ? 4'h3 : _GEN_25272; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25274 = 10'h125 == _T_512[9:0] ? 4'h3 : _GEN_25273; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25275 = 10'h126 == _T_512[9:0] ? 4'h3 : _GEN_25274; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25276 = 10'h127 == _T_512[9:0] ? 4'h1 : _GEN_25275; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25277 = 10'h128 == _T_512[9:0] ? 4'h0 : _GEN_25276; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25278 = 10'h129 == _T_512[9:0] ? 4'h3 : _GEN_25277; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25279 = 10'h12a == _T_512[9:0] ? 4'h3 : _GEN_25278; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25280 = 10'h12b == _T_512[9:0] ? 4'h0 : _GEN_25279; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25281 = 10'h12c == _T_512[9:0] ? 4'h0 : _GEN_25280; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25282 = 10'h12d == _T_512[9:0] ? 4'h0 : _GEN_25281; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25283 = 10'h12e == _T_512[9:0] ? 4'h0 : _GEN_25282; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25284 = 10'h12f == _T_512[9:0] ? 4'h0 : _GEN_25283; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25285 = 10'h130 == _T_512[9:0] ? 4'h0 : _GEN_25284; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25286 = 10'h131 == _T_512[9:0] ? 4'h0 : _GEN_25285; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25287 = 10'h132 == _T_512[9:0] ? 4'h0 : _GEN_25286; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25288 = 10'h133 == _T_512[9:0] ? 4'h0 : _GEN_25287; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25289 = 10'h134 == _T_512[9:0] ? 4'h3 : _GEN_25288; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25290 = 10'h135 == _T_512[9:0] ? 4'h3 : _GEN_25289; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25291 = 10'h136 == _T_512[9:0] ? 4'h0 : _GEN_25290; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25292 = 10'h137 == _T_512[9:0] ? 4'h1 : _GEN_25291; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25293 = 10'h138 == _T_512[9:0] ? 4'h3 : _GEN_25292; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25294 = 10'h139 == _T_512[9:0] ? 4'h3 : _GEN_25293; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25295 = 10'h13a == _T_512[9:0] ? 4'h3 : _GEN_25294; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25296 = 10'h13b == _T_512[9:0] ? 4'h3 : _GEN_25295; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25297 = 10'h13c == _T_512[9:0] ? 4'h3 : _GEN_25296; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25298 = 10'h13d == _T_512[9:0] ? 4'h3 : _GEN_25297; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25299 = 10'h13e == _T_512[9:0] ? 4'ha : _GEN_25298; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25300 = 10'h13f == _T_512[9:0] ? 4'h0 : _GEN_25299; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25301 = 10'h140 == _T_512[9:0] ? 4'h5 : _GEN_25300; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25302 = 10'h141 == _T_512[9:0] ? 4'h3 : _GEN_25301; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25303 = 10'h142 == _T_512[9:0] ? 4'h7 : _GEN_25302; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25304 = 10'h143 == _T_512[9:0] ? 4'ha : _GEN_25303; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25305 = 10'h144 == _T_512[9:0] ? 4'h3 : _GEN_25304; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25306 = 10'h145 == _T_512[9:0] ? 4'h3 : _GEN_25305; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25307 = 10'h146 == _T_512[9:0] ? 4'h1 : _GEN_25306; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25308 = 10'h147 == _T_512[9:0] ? 4'h0 : _GEN_25307; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25309 = 10'h148 == _T_512[9:0] ? 4'h3 : _GEN_25308; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25310 = 10'h149 == _T_512[9:0] ? 4'h3 : _GEN_25309; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25311 = 10'h14a == _T_512[9:0] ? 4'h3 : _GEN_25310; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25312 = 10'h14b == _T_512[9:0] ? 4'h3 : _GEN_25311; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25313 = 10'h14c == _T_512[9:0] ? 4'h3 : _GEN_25312; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25314 = 10'h14d == _T_512[9:0] ? 4'h3 : _GEN_25313; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25315 = 10'h14e == _T_512[9:0] ? 4'h3 : _GEN_25314; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25316 = 10'h14f == _T_512[9:0] ? 4'h3 : _GEN_25315; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25317 = 10'h150 == _T_512[9:0] ? 4'h3 : _GEN_25316; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25318 = 10'h151 == _T_512[9:0] ? 4'h3 : _GEN_25317; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25319 = 10'h152 == _T_512[9:0] ? 4'h3 : _GEN_25318; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25320 = 10'h153 == _T_512[9:0] ? 4'h3 : _GEN_25319; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25321 = 10'h154 == _T_512[9:0] ? 4'h3 : _GEN_25320; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25322 = 10'h155 == _T_512[9:0] ? 4'h3 : _GEN_25321; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25323 = 10'h156 == _T_512[9:0] ? 4'h3 : _GEN_25322; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25324 = 10'h157 == _T_512[9:0] ? 4'h0 : _GEN_25323; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25325 = 10'h158 == _T_512[9:0] ? 4'h3 : _GEN_25324; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25326 = 10'h159 == _T_512[9:0] ? 4'h3 : _GEN_25325; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25327 = 10'h15a == _T_512[9:0] ? 4'h3 : _GEN_25326; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25328 = 10'h15b == _T_512[9:0] ? 4'h3 : _GEN_25327; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25329 = 10'h15c == _T_512[9:0] ? 4'h3 : _GEN_25328; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25330 = 10'h15d == _T_512[9:0] ? 4'ha : _GEN_25329; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25331 = 10'h15e == _T_512[9:0] ? 4'h7 : _GEN_25330; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25332 = 10'h15f == _T_512[9:0] ? 4'h0 : _GEN_25331; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25333 = 10'h160 == _T_512[9:0] ? 4'h3 : _GEN_25332; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25334 = 10'h161 == _T_512[9:0] ? 4'h3 : _GEN_25333; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25335 = 10'h162 == _T_512[9:0] ? 4'h3 : _GEN_25334; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25336 = 10'h163 == _T_512[9:0] ? 4'h7 : _GEN_25335; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25337 = 10'h164 == _T_512[9:0] ? 4'ha : _GEN_25336; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25338 = 10'h165 == _T_512[9:0] ? 4'h1 : _GEN_25337; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25339 = 10'h166 == _T_512[9:0] ? 4'h0 : _GEN_25338; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25340 = 10'h167 == _T_512[9:0] ? 4'h0 : _GEN_25339; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25341 = 10'h168 == _T_512[9:0] ? 4'hc : _GEN_25340; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25342 = 10'h169 == _T_512[9:0] ? 4'h9 : _GEN_25341; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25343 = 10'h16a == _T_512[9:0] ? 4'hc : _GEN_25342; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25344 = 10'h16b == _T_512[9:0] ? 4'hc : _GEN_25343; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25345 = 10'h16c == _T_512[9:0] ? 4'h3 : _GEN_25344; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25346 = 10'h16d == _T_512[9:0] ? 4'h3 : _GEN_25345; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25347 = 10'h16e == _T_512[9:0] ? 4'h3 : _GEN_25346; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25348 = 10'h16f == _T_512[9:0] ? 4'h3 : _GEN_25347; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25349 = 10'h170 == _T_512[9:0] ? 4'h5 : _GEN_25348; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25350 = 10'h171 == _T_512[9:0] ? 4'h3 : _GEN_25349; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25351 = 10'h172 == _T_512[9:0] ? 4'h3 : _GEN_25350; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25352 = 10'h173 == _T_512[9:0] ? 4'h3 : _GEN_25351; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25353 = 10'h174 == _T_512[9:0] ? 4'h3 : _GEN_25352; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25354 = 10'h175 == _T_512[9:0] ? 4'h3 : _GEN_25353; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25355 = 10'h176 == _T_512[9:0] ? 4'h0 : _GEN_25354; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25356 = 10'h177 == _T_512[9:0] ? 4'h0 : _GEN_25355; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25357 = 10'h178 == _T_512[9:0] ? 4'h1 : _GEN_25356; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25358 = 10'h179 == _T_512[9:0] ? 4'h3 : _GEN_25357; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25359 = 10'h17a == _T_512[9:0] ? 4'h5 : _GEN_25358; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25360 = 10'h17b == _T_512[9:0] ? 4'h3 : _GEN_25359; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25361 = 10'h17c == _T_512[9:0] ? 4'ha : _GEN_25360; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25362 = 10'h17d == _T_512[9:0] ? 4'h7 : _GEN_25361; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25363 = 10'h17e == _T_512[9:0] ? 4'h3 : _GEN_25362; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25364 = 10'h17f == _T_512[9:0] ? 4'h0 : _GEN_25363; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25365 = 10'h180 == _T_512[9:0] ? 4'hc : _GEN_25364; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25366 = 10'h181 == _T_512[9:0] ? 4'hc : _GEN_25365; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25367 = 10'h182 == _T_512[9:0] ? 4'hc : _GEN_25366; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25368 = 10'h183 == _T_512[9:0] ? 4'hc : _GEN_25367; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25369 = 10'h184 == _T_512[9:0] ? 4'ha : _GEN_25368; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25370 = 10'h185 == _T_512[9:0] ? 4'h1 : _GEN_25369; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25371 = 10'h186 == _T_512[9:0] ? 4'hc : _GEN_25370; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25372 = 10'h187 == _T_512[9:0] ? 4'h0 : _GEN_25371; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25373 = 10'h188 == _T_512[9:0] ? 4'hc : _GEN_25372; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25374 = 10'h189 == _T_512[9:0] ? 4'hc : _GEN_25373; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25375 = 10'h18a == _T_512[9:0] ? 4'hc : _GEN_25374; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25376 = 10'h18b == _T_512[9:0] ? 4'hc : _GEN_25375; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25377 = 10'h18c == _T_512[9:0] ? 4'hc : _GEN_25376; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25378 = 10'h18d == _T_512[9:0] ? 4'hc : _GEN_25377; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25379 = 10'h18e == _T_512[9:0] ? 4'hc : _GEN_25378; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25380 = 10'h18f == _T_512[9:0] ? 4'hc : _GEN_25379; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25381 = 10'h190 == _T_512[9:0] ? 4'hc : _GEN_25380; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25382 = 10'h191 == _T_512[9:0] ? 4'hc : _GEN_25381; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25383 = 10'h192 == _T_512[9:0] ? 4'h9 : _GEN_25382; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25384 = 10'h193 == _T_512[9:0] ? 4'hc : _GEN_25383; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25385 = 10'h194 == _T_512[9:0] ? 4'hc : _GEN_25384; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25386 = 10'h195 == _T_512[9:0] ? 4'hc : _GEN_25385; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25387 = 10'h196 == _T_512[9:0] ? 4'h0 : _GEN_25386; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25388 = 10'h197 == _T_512[9:0] ? 4'h3 : _GEN_25387; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25389 = 10'h198 == _T_512[9:0] ? 4'h1 : _GEN_25388; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25390 = 10'h199 == _T_512[9:0] ? 4'h3 : _GEN_25389; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25391 = 10'h19a == _T_512[9:0] ? 4'h3 : _GEN_25390; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25392 = 10'h19b == _T_512[9:0] ? 4'h3 : _GEN_25391; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25393 = 10'h19c == _T_512[9:0] ? 4'ha : _GEN_25392; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25394 = 10'h19d == _T_512[9:0] ? 4'h3 : _GEN_25393; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25395 = 10'h19e == _T_512[9:0] ? 4'h3 : _GEN_25394; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25396 = 10'h19f == _T_512[9:0] ? 4'h0 : _GEN_25395; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25397 = 10'h1a0 == _T_512[9:0] ? 4'hc : _GEN_25396; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25398 = 10'h1a1 == _T_512[9:0] ? 4'hc : _GEN_25397; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25399 = 10'h1a2 == _T_512[9:0] ? 4'h9 : _GEN_25398; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25400 = 10'h1a3 == _T_512[9:0] ? 4'hc : _GEN_25399; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25401 = 10'h1a4 == _T_512[9:0] ? 4'ha : _GEN_25400; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25402 = 10'h1a5 == _T_512[9:0] ? 4'h0 : _GEN_25401; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25403 = 10'h1a6 == _T_512[9:0] ? 4'hc : _GEN_25402; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25404 = 10'h1a7 == _T_512[9:0] ? 4'h0 : _GEN_25403; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25405 = 10'h1a8 == _T_512[9:0] ? 4'hc : _GEN_25404; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25406 = 10'h1a9 == _T_512[9:0] ? 4'hc : _GEN_25405; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25407 = 10'h1aa == _T_512[9:0] ? 4'hc : _GEN_25406; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25408 = 10'h1ab == _T_512[9:0] ? 4'h9 : _GEN_25407; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25409 = 10'h1ac == _T_512[9:0] ? 4'hc : _GEN_25408; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25410 = 10'h1ad == _T_512[9:0] ? 4'hc : _GEN_25409; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25411 = 10'h1ae == _T_512[9:0] ? 4'hc : _GEN_25410; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25412 = 10'h1af == _T_512[9:0] ? 4'hc : _GEN_25411; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25413 = 10'h1b0 == _T_512[9:0] ? 4'hc : _GEN_25412; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25414 = 10'h1b1 == _T_512[9:0] ? 4'hc : _GEN_25413; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25415 = 10'h1b2 == _T_512[9:0] ? 4'hc : _GEN_25414; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25416 = 10'h1b3 == _T_512[9:0] ? 4'hc : _GEN_25415; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25417 = 10'h1b4 == _T_512[9:0] ? 4'hc : _GEN_25416; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25418 = 10'h1b5 == _T_512[9:0] ? 4'hc : _GEN_25417; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25419 = 10'h1b6 == _T_512[9:0] ? 4'h0 : _GEN_25418; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25420 = 10'h1b7 == _T_512[9:0] ? 4'hc : _GEN_25419; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25421 = 10'h1b8 == _T_512[9:0] ? 4'h0 : _GEN_25420; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25422 = 10'h1b9 == _T_512[9:0] ? 4'hc : _GEN_25421; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25423 = 10'h1ba == _T_512[9:0] ? 4'hc : _GEN_25422; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25424 = 10'h1bb == _T_512[9:0] ? 4'hc : _GEN_25423; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25425 = 10'h1bc == _T_512[9:0] ? 4'h7 : _GEN_25424; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25426 = 10'h1bd == _T_512[9:0] ? 4'ha : _GEN_25425; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25427 = 10'h1be == _T_512[9:0] ? 4'hc : _GEN_25426; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25428 = 10'h1bf == _T_512[9:0] ? 4'h0 : _GEN_25427; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25429 = 10'h1c0 == _T_512[9:0] ? 4'hc : _GEN_25428; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25430 = 10'h1c1 == _T_512[9:0] ? 4'hc : _GEN_25429; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25431 = 10'h1c2 == _T_512[9:0] ? 4'hc : _GEN_25430; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25432 = 10'h1c3 == _T_512[9:0] ? 4'h7 : _GEN_25431; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25433 = 10'h1c4 == _T_512[9:0] ? 4'h7 : _GEN_25432; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25434 = 10'h1c5 == _T_512[9:0] ? 4'hc : _GEN_25433; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25435 = 10'h1c6 == _T_512[9:0] ? 4'hc : _GEN_25434; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25436 = 10'h1c7 == _T_512[9:0] ? 4'hc : _GEN_25435; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25437 = 10'h1c8 == _T_512[9:0] ? 4'hc : _GEN_25436; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25438 = 10'h1c9 == _T_512[9:0] ? 4'hc : _GEN_25437; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25439 = 10'h1ca == _T_512[9:0] ? 4'hc : _GEN_25438; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25440 = 10'h1cb == _T_512[9:0] ? 4'hc : _GEN_25439; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25441 = 10'h1cc == _T_512[9:0] ? 4'hc : _GEN_25440; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25442 = 10'h1cd == _T_512[9:0] ? 4'hc : _GEN_25441; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25443 = 10'h1ce == _T_512[9:0] ? 4'hc : _GEN_25442; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25444 = 10'h1cf == _T_512[9:0] ? 4'hc : _GEN_25443; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25445 = 10'h1d0 == _T_512[9:0] ? 4'hc : _GEN_25444; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25446 = 10'h1d1 == _T_512[9:0] ? 4'hc : _GEN_25445; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25447 = 10'h1d2 == _T_512[9:0] ? 4'hc : _GEN_25446; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25448 = 10'h1d3 == _T_512[9:0] ? 4'hc : _GEN_25447; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25449 = 10'h1d4 == _T_512[9:0] ? 4'hc : _GEN_25448; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25450 = 10'h1d5 == _T_512[9:0] ? 4'hc : _GEN_25449; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25451 = 10'h1d6 == _T_512[9:0] ? 4'hc : _GEN_25450; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25452 = 10'h1d7 == _T_512[9:0] ? 4'hc : _GEN_25451; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25453 = 10'h1d8 == _T_512[9:0] ? 4'hc : _GEN_25452; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25454 = 10'h1d9 == _T_512[9:0] ? 4'hc : _GEN_25453; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25455 = 10'h1da == _T_512[9:0] ? 4'hc : _GEN_25454; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25456 = 10'h1db == _T_512[9:0] ? 4'hc : _GEN_25455; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25457 = 10'h1dc == _T_512[9:0] ? 4'hc : _GEN_25456; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25458 = 10'h1dd == _T_512[9:0] ? 4'ha : _GEN_25457; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25459 = 10'h1de == _T_512[9:0] ? 4'hc : _GEN_25458; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25460 = 10'h1df == _T_512[9:0] ? 4'h0 : _GEN_25459; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25461 = 10'h1e0 == _T_512[9:0] ? 4'h9 : _GEN_25460; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25462 = 10'h1e1 == _T_512[9:0] ? 4'hc : _GEN_25461; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25463 = 10'h1e2 == _T_512[9:0] ? 4'h7 : _GEN_25462; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25464 = 10'h1e3 == _T_512[9:0] ? 4'h7 : _GEN_25463; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25465 = 10'h1e4 == _T_512[9:0] ? 4'hc : _GEN_25464; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25466 = 10'h1e5 == _T_512[9:0] ? 4'hc : _GEN_25465; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25467 = 10'h1e6 == _T_512[9:0] ? 4'hc : _GEN_25466; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25468 = 10'h1e7 == _T_512[9:0] ? 4'hc : _GEN_25467; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25469 = 10'h1e8 == _T_512[9:0] ? 4'hc : _GEN_25468; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25470 = 10'h1e9 == _T_512[9:0] ? 4'hc : _GEN_25469; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25471 = 10'h1ea == _T_512[9:0] ? 4'hc : _GEN_25470; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25472 = 10'h1eb == _T_512[9:0] ? 4'hc : _GEN_25471; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25473 = 10'h1ec == _T_512[9:0] ? 4'hc : _GEN_25472; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25474 = 10'h1ed == _T_512[9:0] ? 4'hc : _GEN_25473; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25475 = 10'h1ee == _T_512[9:0] ? 4'hc : _GEN_25474; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25476 = 10'h1ef == _T_512[9:0] ? 4'hc : _GEN_25475; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25477 = 10'h1f0 == _T_512[9:0] ? 4'hc : _GEN_25476; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25478 = 10'h1f1 == _T_512[9:0] ? 4'hc : _GEN_25477; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25479 = 10'h1f2 == _T_512[9:0] ? 4'hc : _GEN_25478; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25480 = 10'h1f3 == _T_512[9:0] ? 4'hc : _GEN_25479; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25481 = 10'h1f4 == _T_512[9:0] ? 4'hc : _GEN_25480; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25482 = 10'h1f5 == _T_512[9:0] ? 4'hc : _GEN_25481; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25483 = 10'h1f6 == _T_512[9:0] ? 4'hc : _GEN_25482; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25484 = 10'h1f7 == _T_512[9:0] ? 4'hc : _GEN_25483; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25485 = 10'h1f8 == _T_512[9:0] ? 4'hc : _GEN_25484; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25486 = 10'h1f9 == _T_512[9:0] ? 4'hc : _GEN_25485; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25487 = 10'h1fa == _T_512[9:0] ? 4'h9 : _GEN_25486; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25488 = 10'h1fb == _T_512[9:0] ? 4'hc : _GEN_25487; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25489 = 10'h1fc == _T_512[9:0] ? 4'hc : _GEN_25488; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25490 = 10'h1fd == _T_512[9:0] ? 4'h7 : _GEN_25489; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25491 = 10'h1fe == _T_512[9:0] ? 4'hc : _GEN_25490; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25492 = 10'h1ff == _T_512[9:0] ? 4'h0 : _GEN_25491; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25493 = 10'h200 == _T_512[9:0] ? 4'hc : _GEN_25492; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25494 = 10'h201 == _T_512[9:0] ? 4'hc : _GEN_25493; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25495 = 10'h202 == _T_512[9:0] ? 4'ha : _GEN_25494; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25496 = 10'h203 == _T_512[9:0] ? 4'hc : _GEN_25495; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25497 = 10'h204 == _T_512[9:0] ? 4'hc : _GEN_25496; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25498 = 10'h205 == _T_512[9:0] ? 4'hc : _GEN_25497; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25499 = 10'h206 == _T_512[9:0] ? 4'hc : _GEN_25498; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25500 = 10'h207 == _T_512[9:0] ? 4'hc : _GEN_25499; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25501 = 10'h208 == _T_512[9:0] ? 4'hc : _GEN_25500; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25502 = 10'h209 == _T_512[9:0] ? 4'hc : _GEN_25501; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25503 = 10'h20a == _T_512[9:0] ? 4'hc : _GEN_25502; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25504 = 10'h20b == _T_512[9:0] ? 4'hc : _GEN_25503; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25505 = 10'h20c == _T_512[9:0] ? 4'hc : _GEN_25504; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25506 = 10'h20d == _T_512[9:0] ? 4'hc : _GEN_25505; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25507 = 10'h20e == _T_512[9:0] ? 4'hc : _GEN_25506; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25508 = 10'h20f == _T_512[9:0] ? 4'hc : _GEN_25507; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25509 = 10'h210 == _T_512[9:0] ? 4'hc : _GEN_25508; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25510 = 10'h211 == _T_512[9:0] ? 4'hc : _GEN_25509; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25511 = 10'h212 == _T_512[9:0] ? 4'hc : _GEN_25510; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25512 = 10'h213 == _T_512[9:0] ? 4'hc : _GEN_25511; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25513 = 10'h214 == _T_512[9:0] ? 4'hc : _GEN_25512; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25514 = 10'h215 == _T_512[9:0] ? 4'hc : _GEN_25513; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25515 = 10'h216 == _T_512[9:0] ? 4'hc : _GEN_25514; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25516 = 10'h217 == _T_512[9:0] ? 4'hc : _GEN_25515; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25517 = 10'h218 == _T_512[9:0] ? 4'hc : _GEN_25516; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25518 = 10'h219 == _T_512[9:0] ? 4'hc : _GEN_25517; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25519 = 10'h21a == _T_512[9:0] ? 4'hc : _GEN_25518; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25520 = 10'h21b == _T_512[9:0] ? 4'hc : _GEN_25519; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25521 = 10'h21c == _T_512[9:0] ? 4'ha : _GEN_25520; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25522 = 10'h21d == _T_512[9:0] ? 4'h7 : _GEN_25521; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25523 = 10'h21e == _T_512[9:0] ? 4'hc : _GEN_25522; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25524 = 10'h21f == _T_512[9:0] ? 4'h0 : _GEN_25523; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25525 = 10'h220 == _T_512[9:0] ? 4'h0 : _GEN_25524; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25526 = 10'h221 == _T_512[9:0] ? 4'h0 : _GEN_25525; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25527 = 10'h222 == _T_512[9:0] ? 4'h0 : _GEN_25526; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25528 = 10'h223 == _T_512[9:0] ? 4'h0 : _GEN_25527; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25529 = 10'h224 == _T_512[9:0] ? 4'h0 : _GEN_25528; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25530 = 10'h225 == _T_512[9:0] ? 4'h0 : _GEN_25529; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25531 = 10'h226 == _T_512[9:0] ? 4'h0 : _GEN_25530; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25532 = 10'h227 == _T_512[9:0] ? 4'h0 : _GEN_25531; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25533 = 10'h228 == _T_512[9:0] ? 4'h0 : _GEN_25532; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25534 = 10'h229 == _T_512[9:0] ? 4'h0 : _GEN_25533; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25535 = 10'h22a == _T_512[9:0] ? 4'h0 : _GEN_25534; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25536 = 10'h22b == _T_512[9:0] ? 4'h0 : _GEN_25535; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25537 = 10'h22c == _T_512[9:0] ? 4'h0 : _GEN_25536; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25538 = 10'h22d == _T_512[9:0] ? 4'h0 : _GEN_25537; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25539 = 10'h22e == _T_512[9:0] ? 4'h0 : _GEN_25538; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25540 = 10'h22f == _T_512[9:0] ? 4'h0 : _GEN_25539; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25541 = 10'h230 == _T_512[9:0] ? 4'h0 : _GEN_25540; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25542 = 10'h231 == _T_512[9:0] ? 4'h0 : _GEN_25541; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25543 = 10'h232 == _T_512[9:0] ? 4'h0 : _GEN_25542; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25544 = 10'h233 == _T_512[9:0] ? 4'h0 : _GEN_25543; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25545 = 10'h234 == _T_512[9:0] ? 4'h0 : _GEN_25544; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25546 = 10'h235 == _T_512[9:0] ? 4'h0 : _GEN_25545; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25547 = 10'h236 == _T_512[9:0] ? 4'h0 : _GEN_25546; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25548 = 10'h237 == _T_512[9:0] ? 4'h0 : _GEN_25547; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25549 = 10'h238 == _T_512[9:0] ? 4'h0 : _GEN_25548; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25550 = 10'h239 == _T_512[9:0] ? 4'h0 : _GEN_25549; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25551 = 10'h23a == _T_512[9:0] ? 4'h0 : _GEN_25550; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25552 = 10'h23b == _T_512[9:0] ? 4'h0 : _GEN_25551; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25553 = 10'h23c == _T_512[9:0] ? 4'h0 : _GEN_25552; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25554 = 10'h23d == _T_512[9:0] ? 4'h0 : _GEN_25553; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25555 = 10'h23e == _T_512[9:0] ? 4'h0 : _GEN_25554; // @[Filter.scala 191:102]
  wire [3:0] _GEN_25556 = 10'h23f == _T_512[9:0] ? 4'h0 : _GEN_25555; // @[Filter.scala 191:102]
  wire [6:0] _GEN_28384 = {{3'd0}, _GEN_25556}; // @[Filter.scala 191:102]
  wire [10:0] _T_519 = _GEN_28384 * 7'h46; // @[Filter.scala 191:102]
  wire [10:0] _GEN_28385 = {{2'd0}, _T_514}; // @[Filter.scala 191:69]
  wire [10:0] _T_521 = _GEN_28385 + _T_519; // @[Filter.scala 191:69]
  wire [3:0] _GEN_25588 = 10'h1f == _T_512[9:0] ? 4'h0 : 4'h3; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25589 = 10'h20 == _T_512[9:0] ? 4'h3 : _GEN_25588; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25590 = 10'h21 == _T_512[9:0] ? 4'h3 : _GEN_25589; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25591 = 10'h22 == _T_512[9:0] ? 4'h3 : _GEN_25590; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25592 = 10'h23 == _T_512[9:0] ? 4'h3 : _GEN_25591; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25593 = 10'h24 == _T_512[9:0] ? 4'h3 : _GEN_25592; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25594 = 10'h25 == _T_512[9:0] ? 4'h3 : _GEN_25593; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25595 = 10'h26 == _T_512[9:0] ? 4'h3 : _GEN_25594; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25596 = 10'h27 == _T_512[9:0] ? 4'h9 : _GEN_25595; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25597 = 10'h28 == _T_512[9:0] ? 4'h9 : _GEN_25596; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25598 = 10'h29 == _T_512[9:0] ? 4'h3 : _GEN_25597; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25599 = 10'h2a == _T_512[9:0] ? 4'h3 : _GEN_25598; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25600 = 10'h2b == _T_512[9:0] ? 4'h3 : _GEN_25599; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25601 = 10'h2c == _T_512[9:0] ? 4'h3 : _GEN_25600; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25602 = 10'h2d == _T_512[9:0] ? 4'h3 : _GEN_25601; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25603 = 10'h2e == _T_512[9:0] ? 4'h3 : _GEN_25602; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25604 = 10'h2f == _T_512[9:0] ? 4'h3 : _GEN_25603; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25605 = 10'h30 == _T_512[9:0] ? 4'h3 : _GEN_25604; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25606 = 10'h31 == _T_512[9:0] ? 4'h3 : _GEN_25605; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25607 = 10'h32 == _T_512[9:0] ? 4'h3 : _GEN_25606; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25608 = 10'h33 == _T_512[9:0] ? 4'h3 : _GEN_25607; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25609 = 10'h34 == _T_512[9:0] ? 4'h3 : _GEN_25608; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25610 = 10'h35 == _T_512[9:0] ? 4'h3 : _GEN_25609; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25611 = 10'h36 == _T_512[9:0] ? 4'h3 : _GEN_25610; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25612 = 10'h37 == _T_512[9:0] ? 4'h9 : _GEN_25611; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25613 = 10'h38 == _T_512[9:0] ? 4'h9 : _GEN_25612; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25614 = 10'h39 == _T_512[9:0] ? 4'h3 : _GEN_25613; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25615 = 10'h3a == _T_512[9:0] ? 4'h3 : _GEN_25614; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25616 = 10'h3b == _T_512[9:0] ? 4'h3 : _GEN_25615; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25617 = 10'h3c == _T_512[9:0] ? 4'h3 : _GEN_25616; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25618 = 10'h3d == _T_512[9:0] ? 4'h3 : _GEN_25617; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25619 = 10'h3e == _T_512[9:0] ? 4'h3 : _GEN_25618; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25620 = 10'h3f == _T_512[9:0] ? 4'h0 : _GEN_25619; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25621 = 10'h40 == _T_512[9:0] ? 4'h3 : _GEN_25620; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25622 = 10'h41 == _T_512[9:0] ? 4'h3 : _GEN_25621; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25623 = 10'h42 == _T_512[9:0] ? 4'h3 : _GEN_25622; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25624 = 10'h43 == _T_512[9:0] ? 4'h2 : _GEN_25623; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25625 = 10'h44 == _T_512[9:0] ? 4'h3 : _GEN_25624; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25626 = 10'h45 == _T_512[9:0] ? 4'hf : _GEN_25625; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25627 = 10'h46 == _T_512[9:0] ? 4'hf : _GEN_25626; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25628 = 10'h47 == _T_512[9:0] ? 4'hf : _GEN_25627; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25629 = 10'h48 == _T_512[9:0] ? 4'hf : _GEN_25628; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25630 = 10'h49 == _T_512[9:0] ? 4'h3 : _GEN_25629; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25631 = 10'h4a == _T_512[9:0] ? 4'h3 : _GEN_25630; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25632 = 10'h4b == _T_512[9:0] ? 4'h3 : _GEN_25631; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25633 = 10'h4c == _T_512[9:0] ? 4'h3 : _GEN_25632; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25634 = 10'h4d == _T_512[9:0] ? 4'h3 : _GEN_25633; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25635 = 10'h4e == _T_512[9:0] ? 4'h3 : _GEN_25634; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25636 = 10'h4f == _T_512[9:0] ? 4'h3 : _GEN_25635; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25637 = 10'h50 == _T_512[9:0] ? 4'h3 : _GEN_25636; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25638 = 10'h51 == _T_512[9:0] ? 4'h3 : _GEN_25637; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25639 = 10'h52 == _T_512[9:0] ? 4'h3 : _GEN_25638; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25640 = 10'h53 == _T_512[9:0] ? 4'h3 : _GEN_25639; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25641 = 10'h54 == _T_512[9:0] ? 4'h9 : _GEN_25640; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25642 = 10'h55 == _T_512[9:0] ? 4'h9 : _GEN_25641; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25643 = 10'h56 == _T_512[9:0] ? 4'h9 : _GEN_25642; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25644 = 10'h57 == _T_512[9:0] ? 4'hf : _GEN_25643; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25645 = 10'h58 == _T_512[9:0] ? 4'h3 : _GEN_25644; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25646 = 10'h59 == _T_512[9:0] ? 4'hf : _GEN_25645; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25647 = 10'h5a == _T_512[9:0] ? 4'h3 : _GEN_25646; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25648 = 10'h5b == _T_512[9:0] ? 4'h3 : _GEN_25647; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25649 = 10'h5c == _T_512[9:0] ? 4'h3 : _GEN_25648; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25650 = 10'h5d == _T_512[9:0] ? 4'h3 : _GEN_25649; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25651 = 10'h5e == _T_512[9:0] ? 4'h3 : _GEN_25650; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25652 = 10'h5f == _T_512[9:0] ? 4'h0 : _GEN_25651; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25653 = 10'h60 == _T_512[9:0] ? 4'h3 : _GEN_25652; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25654 = 10'h61 == _T_512[9:0] ? 4'h3 : _GEN_25653; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25655 = 10'h62 == _T_512[9:0] ? 4'h3 : _GEN_25654; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25656 = 10'h63 == _T_512[9:0] ? 4'h3 : _GEN_25655; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25657 = 10'h64 == _T_512[9:0] ? 4'h3 : _GEN_25656; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25658 = 10'h65 == _T_512[9:0] ? 4'hf : _GEN_25657; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25659 = 10'h66 == _T_512[9:0] ? 4'h3 : _GEN_25658; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25660 = 10'h67 == _T_512[9:0] ? 4'h3 : _GEN_25659; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25661 = 10'h68 == _T_512[9:0] ? 4'h3 : _GEN_25660; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25662 = 10'h69 == _T_512[9:0] ? 4'hf : _GEN_25661; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25663 = 10'h6a == _T_512[9:0] ? 4'h9 : _GEN_25662; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25664 = 10'h6b == _T_512[9:0] ? 4'h9 : _GEN_25663; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25665 = 10'h6c == _T_512[9:0] ? 4'h3 : _GEN_25664; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25666 = 10'h6d == _T_512[9:0] ? 4'h3 : _GEN_25665; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25667 = 10'h6e == _T_512[9:0] ? 4'h3 : _GEN_25666; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25668 = 10'h6f == _T_512[9:0] ? 4'h3 : _GEN_25667; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25669 = 10'h70 == _T_512[9:0] ? 4'h3 : _GEN_25668; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25670 = 10'h71 == _T_512[9:0] ? 4'h3 : _GEN_25669; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25671 = 10'h72 == _T_512[9:0] ? 4'h3 : _GEN_25670; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25672 = 10'h73 == _T_512[9:0] ? 4'h9 : _GEN_25671; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25673 = 10'h74 == _T_512[9:0] ? 4'hf : _GEN_25672; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25674 = 10'h75 == _T_512[9:0] ? 4'hf : _GEN_25673; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25675 = 10'h76 == _T_512[9:0] ? 4'hf : _GEN_25674; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25676 = 10'h77 == _T_512[9:0] ? 4'h3 : _GEN_25675; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25677 = 10'h78 == _T_512[9:0] ? 4'h3 : _GEN_25676; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25678 = 10'h79 == _T_512[9:0] ? 4'h3 : _GEN_25677; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25679 = 10'h7a == _T_512[9:0] ? 4'hf : _GEN_25678; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25680 = 10'h7b == _T_512[9:0] ? 4'h3 : _GEN_25679; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25681 = 10'h7c == _T_512[9:0] ? 4'h3 : _GEN_25680; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25682 = 10'h7d == _T_512[9:0] ? 4'h2 : _GEN_25681; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25683 = 10'h7e == _T_512[9:0] ? 4'h3 : _GEN_25682; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25684 = 10'h7f == _T_512[9:0] ? 4'h0 : _GEN_25683; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25685 = 10'h80 == _T_512[9:0] ? 4'h3 : _GEN_25684; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25686 = 10'h81 == _T_512[9:0] ? 4'h3 : _GEN_25685; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25687 = 10'h82 == _T_512[9:0] ? 4'h9 : _GEN_25686; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25688 = 10'h83 == _T_512[9:0] ? 4'hf : _GEN_25687; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25689 = 10'h84 == _T_512[9:0] ? 4'h2 : _GEN_25688; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25690 = 10'h85 == _T_512[9:0] ? 4'h9 : _GEN_25689; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25691 = 10'h86 == _T_512[9:0] ? 4'h9 : _GEN_25690; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25692 = 10'h87 == _T_512[9:0] ? 4'h3 : _GEN_25691; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25693 = 10'h88 == _T_512[9:0] ? 4'h3 : _GEN_25692; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25694 = 10'h89 == _T_512[9:0] ? 4'hf : _GEN_25693; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25695 = 10'h8a == _T_512[9:0] ? 4'hf : _GEN_25694; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25696 = 10'h8b == _T_512[9:0] ? 4'h9 : _GEN_25695; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25697 = 10'h8c == _T_512[9:0] ? 4'h9 : _GEN_25696; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25698 = 10'h8d == _T_512[9:0] ? 4'h9 : _GEN_25697; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25699 = 10'h8e == _T_512[9:0] ? 4'h9 : _GEN_25698; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25700 = 10'h8f == _T_512[9:0] ? 4'h9 : _GEN_25699; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25701 = 10'h90 == _T_512[9:0] ? 4'h9 : _GEN_25700; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25702 = 10'h91 == _T_512[9:0] ? 4'h9 : _GEN_25701; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25703 = 10'h92 == _T_512[9:0] ? 4'h9 : _GEN_25702; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25704 = 10'h93 == _T_512[9:0] ? 4'hf : _GEN_25703; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25705 = 10'h94 == _T_512[9:0] ? 4'hf : _GEN_25704; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25706 = 10'h95 == _T_512[9:0] ? 4'h3 : _GEN_25705; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25707 = 10'h96 == _T_512[9:0] ? 4'h3 : _GEN_25706; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25708 = 10'h97 == _T_512[9:0] ? 4'h3 : _GEN_25707; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25709 = 10'h98 == _T_512[9:0] ? 4'h9 : _GEN_25708; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25710 = 10'h99 == _T_512[9:0] ? 4'hf : _GEN_25709; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25711 = 10'h9a == _T_512[9:0] ? 4'h9 : _GEN_25710; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25712 = 10'h9b == _T_512[9:0] ? 4'h9 : _GEN_25711; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25713 = 10'h9c == _T_512[9:0] ? 4'h3 : _GEN_25712; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25714 = 10'h9d == _T_512[9:0] ? 4'h3 : _GEN_25713; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25715 = 10'h9e == _T_512[9:0] ? 4'h3 : _GEN_25714; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25716 = 10'h9f == _T_512[9:0] ? 4'h0 : _GEN_25715; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25717 = 10'ha0 == _T_512[9:0] ? 4'h3 : _GEN_25716; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25718 = 10'ha1 == _T_512[9:0] ? 4'h9 : _GEN_25717; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25719 = 10'ha2 == _T_512[9:0] ? 4'hf : _GEN_25718; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25720 = 10'ha3 == _T_512[9:0] ? 4'h3 : _GEN_25719; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25721 = 10'ha4 == _T_512[9:0] ? 4'h3 : _GEN_25720; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25722 = 10'ha5 == _T_512[9:0] ? 4'h3 : _GEN_25721; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25723 = 10'ha6 == _T_512[9:0] ? 4'h3 : _GEN_25722; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25724 = 10'ha7 == _T_512[9:0] ? 4'hf : _GEN_25723; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25725 = 10'ha8 == _T_512[9:0] ? 4'h3 : _GEN_25724; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25726 = 10'ha9 == _T_512[9:0] ? 4'h9 : _GEN_25725; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25727 = 10'haa == _T_512[9:0] ? 4'hf : _GEN_25726; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25728 = 10'hab == _T_512[9:0] ? 4'hf : _GEN_25727; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25729 = 10'hac == _T_512[9:0] ? 4'hf : _GEN_25728; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25730 = 10'had == _T_512[9:0] ? 4'hf : _GEN_25729; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25731 = 10'hae == _T_512[9:0] ? 4'hf : _GEN_25730; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25732 = 10'haf == _T_512[9:0] ? 4'hf : _GEN_25731; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25733 = 10'hb0 == _T_512[9:0] ? 4'hf : _GEN_25732; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25734 = 10'hb1 == _T_512[9:0] ? 4'hf : _GEN_25733; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25735 = 10'hb2 == _T_512[9:0] ? 4'hf : _GEN_25734; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25736 = 10'hb3 == _T_512[9:0] ? 4'hf : _GEN_25735; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25737 = 10'hb4 == _T_512[9:0] ? 4'h9 : _GEN_25736; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25738 = 10'hb5 == _T_512[9:0] ? 4'h9 : _GEN_25737; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25739 = 10'hb6 == _T_512[9:0] ? 4'h3 : _GEN_25738; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25740 = 10'hb7 == _T_512[9:0] ? 4'hf : _GEN_25739; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25741 = 10'hb8 == _T_512[9:0] ? 4'h3 : _GEN_25740; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25742 = 10'hb9 == _T_512[9:0] ? 4'h3 : _GEN_25741; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25743 = 10'hba == _T_512[9:0] ? 4'h3 : _GEN_25742; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25744 = 10'hbb == _T_512[9:0] ? 4'hf : _GEN_25743; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25745 = 10'hbc == _T_512[9:0] ? 4'h3 : _GEN_25744; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25746 = 10'hbd == _T_512[9:0] ? 4'h3 : _GEN_25745; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25747 = 10'hbe == _T_512[9:0] ? 4'h3 : _GEN_25746; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25748 = 10'hbf == _T_512[9:0] ? 4'h0 : _GEN_25747; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25749 = 10'hc0 == _T_512[9:0] ? 4'h3 : _GEN_25748; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25750 = 10'hc1 == _T_512[9:0] ? 4'h3 : _GEN_25749; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25751 = 10'hc2 == _T_512[9:0] ? 4'h3 : _GEN_25750; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25752 = 10'hc3 == _T_512[9:0] ? 4'h2 : _GEN_25751; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25753 = 10'hc4 == _T_512[9:0] ? 4'hf : _GEN_25752; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25754 = 10'hc5 == _T_512[9:0] ? 4'hf : _GEN_25753; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25755 = 10'hc6 == _T_512[9:0] ? 4'hf : _GEN_25754; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25756 = 10'hc7 == _T_512[9:0] ? 4'h3 : _GEN_25755; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25757 = 10'hc8 == _T_512[9:0] ? 4'h9 : _GEN_25756; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25758 = 10'hc9 == _T_512[9:0] ? 4'hf : _GEN_25757; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25759 = 10'hca == _T_512[9:0] ? 4'hf : _GEN_25758; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25760 = 10'hcb == _T_512[9:0] ? 4'hf : _GEN_25759; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25761 = 10'hcc == _T_512[9:0] ? 4'hf : _GEN_25760; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25762 = 10'hcd == _T_512[9:0] ? 4'hf : _GEN_25761; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25763 = 10'hce == _T_512[9:0] ? 4'hf : _GEN_25762; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25764 = 10'hcf == _T_512[9:0] ? 4'hf : _GEN_25763; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25765 = 10'hd0 == _T_512[9:0] ? 4'hf : _GEN_25764; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25766 = 10'hd1 == _T_512[9:0] ? 4'hf : _GEN_25765; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25767 = 10'hd2 == _T_512[9:0] ? 4'hf : _GEN_25766; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25768 = 10'hd3 == _T_512[9:0] ? 4'hf : _GEN_25767; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25769 = 10'hd4 == _T_512[9:0] ? 4'hf : _GEN_25768; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25770 = 10'hd5 == _T_512[9:0] ? 4'hf : _GEN_25769; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25771 = 10'hd6 == _T_512[9:0] ? 4'h9 : _GEN_25770; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25772 = 10'hd7 == _T_512[9:0] ? 4'h3 : _GEN_25771; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25773 = 10'hd8 == _T_512[9:0] ? 4'hf : _GEN_25772; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25774 = 10'hd9 == _T_512[9:0] ? 4'h3 : _GEN_25773; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25775 = 10'hda == _T_512[9:0] ? 4'h3 : _GEN_25774; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25776 = 10'hdb == _T_512[9:0] ? 4'h3 : _GEN_25775; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25777 = 10'hdc == _T_512[9:0] ? 4'h3 : _GEN_25776; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25778 = 10'hdd == _T_512[9:0] ? 4'h3 : _GEN_25777; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25779 = 10'hde == _T_512[9:0] ? 4'h2 : _GEN_25778; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25780 = 10'hdf == _T_512[9:0] ? 4'h0 : _GEN_25779; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25781 = 10'he0 == _T_512[9:0] ? 4'h3 : _GEN_25780; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25782 = 10'he1 == _T_512[9:0] ? 4'h3 : _GEN_25781; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25783 = 10'he2 == _T_512[9:0] ? 4'h3 : _GEN_25782; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25784 = 10'he3 == _T_512[9:0] ? 4'h3 : _GEN_25783; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25785 = 10'he4 == _T_512[9:0] ? 4'h3 : _GEN_25784; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25786 = 10'he5 == _T_512[9:0] ? 4'h3 : _GEN_25785; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25787 = 10'he6 == _T_512[9:0] ? 4'h3 : _GEN_25786; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25788 = 10'he7 == _T_512[9:0] ? 4'h9 : _GEN_25787; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25789 = 10'he8 == _T_512[9:0] ? 4'h9 : _GEN_25788; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25790 = 10'he9 == _T_512[9:0] ? 4'h9 : _GEN_25789; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25791 = 10'hea == _T_512[9:0] ? 4'hf : _GEN_25790; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25792 = 10'heb == _T_512[9:0] ? 4'hf : _GEN_25791; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25793 = 10'hec == _T_512[9:0] ? 4'hf : _GEN_25792; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25794 = 10'hed == _T_512[9:0] ? 4'hf : _GEN_25793; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25795 = 10'hee == _T_512[9:0] ? 4'hf : _GEN_25794; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25796 = 10'hef == _T_512[9:0] ? 4'hf : _GEN_25795; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25797 = 10'hf0 == _T_512[9:0] ? 4'hf : _GEN_25796; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25798 = 10'hf1 == _T_512[9:0] ? 4'hf : _GEN_25797; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25799 = 10'hf2 == _T_512[9:0] ? 4'hf : _GEN_25798; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25800 = 10'hf3 == _T_512[9:0] ? 4'hf : _GEN_25799; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25801 = 10'hf4 == _T_512[9:0] ? 4'hf : _GEN_25800; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25802 = 10'hf5 == _T_512[9:0] ? 4'h9 : _GEN_25801; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25803 = 10'hf6 == _T_512[9:0] ? 4'hf : _GEN_25802; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25804 = 10'hf7 == _T_512[9:0] ? 4'hf : _GEN_25803; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25805 = 10'hf8 == _T_512[9:0] ? 4'h9 : _GEN_25804; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25806 = 10'hf9 == _T_512[9:0] ? 4'hf : _GEN_25805; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25807 = 10'hfa == _T_512[9:0] ? 4'h3 : _GEN_25806; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25808 = 10'hfb == _T_512[9:0] ? 4'h3 : _GEN_25807; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25809 = 10'hfc == _T_512[9:0] ? 4'h3 : _GEN_25808; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25810 = 10'hfd == _T_512[9:0] ? 4'h3 : _GEN_25809; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25811 = 10'hfe == _T_512[9:0] ? 4'h3 : _GEN_25810; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25812 = 10'hff == _T_512[9:0] ? 4'h0 : _GEN_25811; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25813 = 10'h100 == _T_512[9:0] ? 4'h3 : _GEN_25812; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25814 = 10'h101 == _T_512[9:0] ? 4'hf : _GEN_25813; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25815 = 10'h102 == _T_512[9:0] ? 4'h3 : _GEN_25814; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25816 = 10'h103 == _T_512[9:0] ? 4'h3 : _GEN_25815; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25817 = 10'h104 == _T_512[9:0] ? 4'h3 : _GEN_25816; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25818 = 10'h105 == _T_512[9:0] ? 4'h3 : _GEN_25817; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25819 = 10'h106 == _T_512[9:0] ? 4'h3 : _GEN_25818; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25820 = 10'h107 == _T_512[9:0] ? 4'h3 : _GEN_25819; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25821 = 10'h108 == _T_512[9:0] ? 4'h9 : _GEN_25820; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25822 = 10'h109 == _T_512[9:0] ? 4'hf : _GEN_25821; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25823 = 10'h10a == _T_512[9:0] ? 4'hf : _GEN_25822; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25824 = 10'h10b == _T_512[9:0] ? 4'hf : _GEN_25823; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25825 = 10'h10c == _T_512[9:0] ? 4'hf : _GEN_25824; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25826 = 10'h10d == _T_512[9:0] ? 4'h0 : _GEN_25825; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25827 = 10'h10e == _T_512[9:0] ? 4'hf : _GEN_25826; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25828 = 10'h10f == _T_512[9:0] ? 4'hf : _GEN_25827; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25829 = 10'h110 == _T_512[9:0] ? 4'hf : _GEN_25828; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25830 = 10'h111 == _T_512[9:0] ? 4'h0 : _GEN_25829; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25831 = 10'h112 == _T_512[9:0] ? 4'hf : _GEN_25830; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25832 = 10'h113 == _T_512[9:0] ? 4'hf : _GEN_25831; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25833 = 10'h114 == _T_512[9:0] ? 4'hf : _GEN_25832; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25834 = 10'h115 == _T_512[9:0] ? 4'hf : _GEN_25833; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25835 = 10'h116 == _T_512[9:0] ? 4'h9 : _GEN_25834; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25836 = 10'h117 == _T_512[9:0] ? 4'h3 : _GEN_25835; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25837 = 10'h118 == _T_512[9:0] ? 4'h3 : _GEN_25836; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25838 = 10'h119 == _T_512[9:0] ? 4'h3 : _GEN_25837; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25839 = 10'h11a == _T_512[9:0] ? 4'hf : _GEN_25838; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25840 = 10'h11b == _T_512[9:0] ? 4'h3 : _GEN_25839; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25841 = 10'h11c == _T_512[9:0] ? 4'h3 : _GEN_25840; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25842 = 10'h11d == _T_512[9:0] ? 4'h2 : _GEN_25841; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25843 = 10'h11e == _T_512[9:0] ? 4'h3 : _GEN_25842; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25844 = 10'h11f == _T_512[9:0] ? 4'h0 : _GEN_25843; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25845 = 10'h120 == _T_512[9:0] ? 4'h3 : _GEN_25844; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25846 = 10'h121 == _T_512[9:0] ? 4'h3 : _GEN_25845; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25847 = 10'h122 == _T_512[9:0] ? 4'h3 : _GEN_25846; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25848 = 10'h123 == _T_512[9:0] ? 4'h3 : _GEN_25847; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25849 = 10'h124 == _T_512[9:0] ? 4'h3 : _GEN_25848; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25850 = 10'h125 == _T_512[9:0] ? 4'h3 : _GEN_25849; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25851 = 10'h126 == _T_512[9:0] ? 4'h3 : _GEN_25850; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25852 = 10'h127 == _T_512[9:0] ? 4'h9 : _GEN_25851; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25853 = 10'h128 == _T_512[9:0] ? 4'hf : _GEN_25852; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25854 = 10'h129 == _T_512[9:0] ? 4'h3 : _GEN_25853; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25855 = 10'h12a == _T_512[9:0] ? 4'h3 : _GEN_25854; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25856 = 10'h12b == _T_512[9:0] ? 4'hf : _GEN_25855; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25857 = 10'h12c == _T_512[9:0] ? 4'hf : _GEN_25856; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25858 = 10'h12d == _T_512[9:0] ? 4'hf : _GEN_25857; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25859 = 10'h12e == _T_512[9:0] ? 4'hf : _GEN_25858; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25860 = 10'h12f == _T_512[9:0] ? 4'hf : _GEN_25859; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25861 = 10'h130 == _T_512[9:0] ? 4'hf : _GEN_25860; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25862 = 10'h131 == _T_512[9:0] ? 4'hf : _GEN_25861; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25863 = 10'h132 == _T_512[9:0] ? 4'hf : _GEN_25862; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25864 = 10'h133 == _T_512[9:0] ? 4'hf : _GEN_25863; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25865 = 10'h134 == _T_512[9:0] ? 4'h3 : _GEN_25864; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25866 = 10'h135 == _T_512[9:0] ? 4'h3 : _GEN_25865; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25867 = 10'h136 == _T_512[9:0] ? 4'hf : _GEN_25866; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25868 = 10'h137 == _T_512[9:0] ? 4'h9 : _GEN_25867; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25869 = 10'h138 == _T_512[9:0] ? 4'h3 : _GEN_25868; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25870 = 10'h139 == _T_512[9:0] ? 4'h3 : _GEN_25869; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25871 = 10'h13a == _T_512[9:0] ? 4'h3 : _GEN_25870; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25872 = 10'h13b == _T_512[9:0] ? 4'h3 : _GEN_25871; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25873 = 10'h13c == _T_512[9:0] ? 4'h3 : _GEN_25872; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25874 = 10'h13d == _T_512[9:0] ? 4'h3 : _GEN_25873; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25875 = 10'h13e == _T_512[9:0] ? 4'h3 : _GEN_25874; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25876 = 10'h13f == _T_512[9:0] ? 4'h0 : _GEN_25875; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25877 = 10'h140 == _T_512[9:0] ? 4'h3 : _GEN_25876; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25878 = 10'h141 == _T_512[9:0] ? 4'h3 : _GEN_25877; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25879 = 10'h142 == _T_512[9:0] ? 4'h2 : _GEN_25878; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25880 = 10'h143 == _T_512[9:0] ? 4'h3 : _GEN_25879; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25881 = 10'h144 == _T_512[9:0] ? 4'h3 : _GEN_25880; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25882 = 10'h145 == _T_512[9:0] ? 4'h3 : _GEN_25881; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25883 = 10'h146 == _T_512[9:0] ? 4'h9 : _GEN_25882; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25884 = 10'h147 == _T_512[9:0] ? 4'hf : _GEN_25883; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25885 = 10'h148 == _T_512[9:0] ? 4'h3 : _GEN_25884; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25886 = 10'h149 == _T_512[9:0] ? 4'h3 : _GEN_25885; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25887 = 10'h14a == _T_512[9:0] ? 4'h3 : _GEN_25886; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25888 = 10'h14b == _T_512[9:0] ? 4'h3 : _GEN_25887; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25889 = 10'h14c == _T_512[9:0] ? 4'h3 : _GEN_25888; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25890 = 10'h14d == _T_512[9:0] ? 4'h3 : _GEN_25889; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25891 = 10'h14e == _T_512[9:0] ? 4'h3 : _GEN_25890; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25892 = 10'h14f == _T_512[9:0] ? 4'h3 : _GEN_25891; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25893 = 10'h150 == _T_512[9:0] ? 4'h3 : _GEN_25892; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25894 = 10'h151 == _T_512[9:0] ? 4'h3 : _GEN_25893; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25895 = 10'h152 == _T_512[9:0] ? 4'h3 : _GEN_25894; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25896 = 10'h153 == _T_512[9:0] ? 4'h3 : _GEN_25895; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25897 = 10'h154 == _T_512[9:0] ? 4'h3 : _GEN_25896; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25898 = 10'h155 == _T_512[9:0] ? 4'h3 : _GEN_25897; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25899 = 10'h156 == _T_512[9:0] ? 4'h3 : _GEN_25898; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25900 = 10'h157 == _T_512[9:0] ? 4'hf : _GEN_25899; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25901 = 10'h158 == _T_512[9:0] ? 4'h3 : _GEN_25900; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25902 = 10'h159 == _T_512[9:0] ? 4'h3 : _GEN_25901; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25903 = 10'h15a == _T_512[9:0] ? 4'h3 : _GEN_25902; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25904 = 10'h15b == _T_512[9:0] ? 4'h3 : _GEN_25903; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25905 = 10'h15c == _T_512[9:0] ? 4'h3 : _GEN_25904; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25906 = 10'h15d == _T_512[9:0] ? 4'h3 : _GEN_25905; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25907 = 10'h15e == _T_512[9:0] ? 4'h2 : _GEN_25906; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25908 = 10'h15f == _T_512[9:0] ? 4'h0 : _GEN_25907; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25909 = 10'h160 == _T_512[9:0] ? 4'h3 : _GEN_25908; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25910 = 10'h161 == _T_512[9:0] ? 4'h3 : _GEN_25909; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25911 = 10'h162 == _T_512[9:0] ? 4'h3 : _GEN_25910; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25912 = 10'h163 == _T_512[9:0] ? 4'h2 : _GEN_25911; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25913 = 10'h164 == _T_512[9:0] ? 4'h3 : _GEN_25912; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25914 = 10'h165 == _T_512[9:0] ? 4'h9 : _GEN_25913; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25915 = 10'h166 == _T_512[9:0] ? 4'hf : _GEN_25914; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25916 = 10'h167 == _T_512[9:0] ? 4'hf : _GEN_25915; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25917 = 10'h168 == _T_512[9:0] ? 4'hd : _GEN_25916; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25918 = 10'h169 == _T_512[9:0] ? 4'h9 : _GEN_25917; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25919 = 10'h16a == _T_512[9:0] ? 4'hd : _GEN_25918; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25920 = 10'h16b == _T_512[9:0] ? 4'hd : _GEN_25919; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25921 = 10'h16c == _T_512[9:0] ? 4'h3 : _GEN_25920; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25922 = 10'h16d == _T_512[9:0] ? 4'h3 : _GEN_25921; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25923 = 10'h16e == _T_512[9:0] ? 4'h3 : _GEN_25922; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25924 = 10'h16f == _T_512[9:0] ? 4'h3 : _GEN_25923; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25925 = 10'h170 == _T_512[9:0] ? 4'h3 : _GEN_25924; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25926 = 10'h171 == _T_512[9:0] ? 4'h3 : _GEN_25925; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25927 = 10'h172 == _T_512[9:0] ? 4'h3 : _GEN_25926; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25928 = 10'h173 == _T_512[9:0] ? 4'h3 : _GEN_25927; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25929 = 10'h174 == _T_512[9:0] ? 4'h3 : _GEN_25928; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25930 = 10'h175 == _T_512[9:0] ? 4'h3 : _GEN_25929; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25931 = 10'h176 == _T_512[9:0] ? 4'hf : _GEN_25930; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25932 = 10'h177 == _T_512[9:0] ? 4'hf : _GEN_25931; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25933 = 10'h178 == _T_512[9:0] ? 4'h9 : _GEN_25932; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25934 = 10'h179 == _T_512[9:0] ? 4'h3 : _GEN_25933; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25935 = 10'h17a == _T_512[9:0] ? 4'h3 : _GEN_25934; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25936 = 10'h17b == _T_512[9:0] ? 4'h3 : _GEN_25935; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25937 = 10'h17c == _T_512[9:0] ? 4'h3 : _GEN_25936; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25938 = 10'h17d == _T_512[9:0] ? 4'h2 : _GEN_25937; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25939 = 10'h17e == _T_512[9:0] ? 4'h3 : _GEN_25938; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25940 = 10'h17f == _T_512[9:0] ? 4'h0 : _GEN_25939; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25941 = 10'h180 == _T_512[9:0] ? 4'hd : _GEN_25940; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25942 = 10'h181 == _T_512[9:0] ? 4'hd : _GEN_25941; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25943 = 10'h182 == _T_512[9:0] ? 4'hd : _GEN_25942; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25944 = 10'h183 == _T_512[9:0] ? 4'hd : _GEN_25943; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25945 = 10'h184 == _T_512[9:0] ? 4'h3 : _GEN_25944; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25946 = 10'h185 == _T_512[9:0] ? 4'h9 : _GEN_25945; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25947 = 10'h186 == _T_512[9:0] ? 4'hb : _GEN_25946; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25948 = 10'h187 == _T_512[9:0] ? 4'hf : _GEN_25947; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25949 = 10'h188 == _T_512[9:0] ? 4'hd : _GEN_25948; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25950 = 10'h189 == _T_512[9:0] ? 4'hd : _GEN_25949; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25951 = 10'h18a == _T_512[9:0] ? 4'hd : _GEN_25950; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25952 = 10'h18b == _T_512[9:0] ? 4'hd : _GEN_25951; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25953 = 10'h18c == _T_512[9:0] ? 4'hd : _GEN_25952; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25954 = 10'h18d == _T_512[9:0] ? 4'hd : _GEN_25953; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25955 = 10'h18e == _T_512[9:0] ? 4'hd : _GEN_25954; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25956 = 10'h18f == _T_512[9:0] ? 4'hd : _GEN_25955; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25957 = 10'h190 == _T_512[9:0] ? 4'hd : _GEN_25956; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25958 = 10'h191 == _T_512[9:0] ? 4'hd : _GEN_25957; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25959 = 10'h192 == _T_512[9:0] ? 4'h9 : _GEN_25958; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25960 = 10'h193 == _T_512[9:0] ? 4'hd : _GEN_25959; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25961 = 10'h194 == _T_512[9:0] ? 4'hd : _GEN_25960; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25962 = 10'h195 == _T_512[9:0] ? 4'hd : _GEN_25961; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25963 = 10'h196 == _T_512[9:0] ? 4'hf : _GEN_25962; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25964 = 10'h197 == _T_512[9:0] ? 4'h3 : _GEN_25963; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25965 = 10'h198 == _T_512[9:0] ? 4'h9 : _GEN_25964; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25966 = 10'h199 == _T_512[9:0] ? 4'h3 : _GEN_25965; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25967 = 10'h19a == _T_512[9:0] ? 4'h3 : _GEN_25966; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25968 = 10'h19b == _T_512[9:0] ? 4'h3 : _GEN_25967; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25969 = 10'h19c == _T_512[9:0] ? 4'h3 : _GEN_25968; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25970 = 10'h19d == _T_512[9:0] ? 4'h3 : _GEN_25969; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25971 = 10'h19e == _T_512[9:0] ? 4'h3 : _GEN_25970; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25972 = 10'h19f == _T_512[9:0] ? 4'h0 : _GEN_25971; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25973 = 10'h1a0 == _T_512[9:0] ? 4'hd : _GEN_25972; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25974 = 10'h1a1 == _T_512[9:0] ? 4'hd : _GEN_25973; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25975 = 10'h1a2 == _T_512[9:0] ? 4'h9 : _GEN_25974; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25976 = 10'h1a3 == _T_512[9:0] ? 4'hd : _GEN_25975; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25977 = 10'h1a4 == _T_512[9:0] ? 4'h3 : _GEN_25976; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25978 = 10'h1a5 == _T_512[9:0] ? 4'hf : _GEN_25977; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25979 = 10'h1a6 == _T_512[9:0] ? 4'hd : _GEN_25978; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25980 = 10'h1a7 == _T_512[9:0] ? 4'hf : _GEN_25979; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25981 = 10'h1a8 == _T_512[9:0] ? 4'hb : _GEN_25980; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25982 = 10'h1a9 == _T_512[9:0] ? 4'hd : _GEN_25981; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25983 = 10'h1aa == _T_512[9:0] ? 4'hd : _GEN_25982; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25984 = 10'h1ab == _T_512[9:0] ? 4'h9 : _GEN_25983; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25985 = 10'h1ac == _T_512[9:0] ? 4'hd : _GEN_25984; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25986 = 10'h1ad == _T_512[9:0] ? 4'hd : _GEN_25985; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25987 = 10'h1ae == _T_512[9:0] ? 4'hd : _GEN_25986; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25988 = 10'h1af == _T_512[9:0] ? 4'hd : _GEN_25987; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25989 = 10'h1b0 == _T_512[9:0] ? 4'hd : _GEN_25988; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25990 = 10'h1b1 == _T_512[9:0] ? 4'hd : _GEN_25989; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25991 = 10'h1b2 == _T_512[9:0] ? 4'hd : _GEN_25990; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25992 = 10'h1b3 == _T_512[9:0] ? 4'hd : _GEN_25991; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25993 = 10'h1b4 == _T_512[9:0] ? 4'hd : _GEN_25992; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25994 = 10'h1b5 == _T_512[9:0] ? 4'hd : _GEN_25993; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25995 = 10'h1b6 == _T_512[9:0] ? 4'hf : _GEN_25994; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25996 = 10'h1b7 == _T_512[9:0] ? 4'hd : _GEN_25995; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25997 = 10'h1b8 == _T_512[9:0] ? 4'hf : _GEN_25996; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25998 = 10'h1b9 == _T_512[9:0] ? 4'hd : _GEN_25997; // @[Filter.scala 191:142]
  wire [3:0] _GEN_25999 = 10'h1ba == _T_512[9:0] ? 4'hd : _GEN_25998; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26000 = 10'h1bb == _T_512[9:0] ? 4'hd : _GEN_25999; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26001 = 10'h1bc == _T_512[9:0] ? 4'h2 : _GEN_26000; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26002 = 10'h1bd == _T_512[9:0] ? 4'h3 : _GEN_26001; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26003 = 10'h1be == _T_512[9:0] ? 4'hd : _GEN_26002; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26004 = 10'h1bf == _T_512[9:0] ? 4'h0 : _GEN_26003; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26005 = 10'h1c0 == _T_512[9:0] ? 4'hd : _GEN_26004; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26006 = 10'h1c1 == _T_512[9:0] ? 4'hd : _GEN_26005; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26007 = 10'h1c2 == _T_512[9:0] ? 4'hd : _GEN_26006; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26008 = 10'h1c3 == _T_512[9:0] ? 4'h2 : _GEN_26007; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26009 = 10'h1c4 == _T_512[9:0] ? 4'h2 : _GEN_26008; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26010 = 10'h1c5 == _T_512[9:0] ? 4'hd : _GEN_26009; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26011 = 10'h1c6 == _T_512[9:0] ? 4'hd : _GEN_26010; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26012 = 10'h1c7 == _T_512[9:0] ? 4'hd : _GEN_26011; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26013 = 10'h1c8 == _T_512[9:0] ? 4'hd : _GEN_26012; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26014 = 10'h1c9 == _T_512[9:0] ? 4'hb : _GEN_26013; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26015 = 10'h1ca == _T_512[9:0] ? 4'hb : _GEN_26014; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26016 = 10'h1cb == _T_512[9:0] ? 4'hb : _GEN_26015; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26017 = 10'h1cc == _T_512[9:0] ? 4'hb : _GEN_26016; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26018 = 10'h1cd == _T_512[9:0] ? 4'hb : _GEN_26017; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26019 = 10'h1ce == _T_512[9:0] ? 4'hb : _GEN_26018; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26020 = 10'h1cf == _T_512[9:0] ? 4'hb : _GEN_26019; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26021 = 10'h1d0 == _T_512[9:0] ? 4'hb : _GEN_26020; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26022 = 10'h1d1 == _T_512[9:0] ? 4'hb : _GEN_26021; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26023 = 10'h1d2 == _T_512[9:0] ? 4'hb : _GEN_26022; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26024 = 10'h1d3 == _T_512[9:0] ? 4'hb : _GEN_26023; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26025 = 10'h1d4 == _T_512[9:0] ? 4'hb : _GEN_26024; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26026 = 10'h1d5 == _T_512[9:0] ? 4'hb : _GEN_26025; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26027 = 10'h1d6 == _T_512[9:0] ? 4'hd : _GEN_26026; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26028 = 10'h1d7 == _T_512[9:0] ? 4'hd : _GEN_26027; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26029 = 10'h1d8 == _T_512[9:0] ? 4'hd : _GEN_26028; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26030 = 10'h1d9 == _T_512[9:0] ? 4'hd : _GEN_26029; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26031 = 10'h1da == _T_512[9:0] ? 4'hd : _GEN_26030; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26032 = 10'h1db == _T_512[9:0] ? 4'hd : _GEN_26031; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26033 = 10'h1dc == _T_512[9:0] ? 4'hd : _GEN_26032; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26034 = 10'h1dd == _T_512[9:0] ? 4'h3 : _GEN_26033; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26035 = 10'h1de == _T_512[9:0] ? 4'hd : _GEN_26034; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26036 = 10'h1df == _T_512[9:0] ? 4'h0 : _GEN_26035; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26037 = 10'h1e0 == _T_512[9:0] ? 4'h9 : _GEN_26036; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26038 = 10'h1e1 == _T_512[9:0] ? 4'hd : _GEN_26037; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26039 = 10'h1e2 == _T_512[9:0] ? 4'h2 : _GEN_26038; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26040 = 10'h1e3 == _T_512[9:0] ? 4'h2 : _GEN_26039; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26041 = 10'h1e4 == _T_512[9:0] ? 4'hd : _GEN_26040; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26042 = 10'h1e5 == _T_512[9:0] ? 4'hd : _GEN_26041; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26043 = 10'h1e6 == _T_512[9:0] ? 4'hd : _GEN_26042; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26044 = 10'h1e7 == _T_512[9:0] ? 4'hd : _GEN_26043; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26045 = 10'h1e8 == _T_512[9:0] ? 4'hb : _GEN_26044; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26046 = 10'h1e9 == _T_512[9:0] ? 4'hd : _GEN_26045; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26047 = 10'h1ea == _T_512[9:0] ? 4'hd : _GEN_26046; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26048 = 10'h1eb == _T_512[9:0] ? 4'hb : _GEN_26047; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26049 = 10'h1ec == _T_512[9:0] ? 4'hd : _GEN_26048; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26050 = 10'h1ed == _T_512[9:0] ? 4'hb : _GEN_26049; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26051 = 10'h1ee == _T_512[9:0] ? 4'hd : _GEN_26050; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26052 = 10'h1ef == _T_512[9:0] ? 4'hb : _GEN_26051; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26053 = 10'h1f0 == _T_512[9:0] ? 4'hd : _GEN_26052; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26054 = 10'h1f1 == _T_512[9:0] ? 4'hb : _GEN_26053; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26055 = 10'h1f2 == _T_512[9:0] ? 4'hb : _GEN_26054; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26056 = 10'h1f3 == _T_512[9:0] ? 4'hd : _GEN_26055; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26057 = 10'h1f4 == _T_512[9:0] ? 4'hb : _GEN_26056; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26058 = 10'h1f5 == _T_512[9:0] ? 4'hb : _GEN_26057; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26059 = 10'h1f6 == _T_512[9:0] ? 4'hd : _GEN_26058; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26060 = 10'h1f7 == _T_512[9:0] ? 4'hd : _GEN_26059; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26061 = 10'h1f8 == _T_512[9:0] ? 4'hd : _GEN_26060; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26062 = 10'h1f9 == _T_512[9:0] ? 4'hd : _GEN_26061; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26063 = 10'h1fa == _T_512[9:0] ? 4'h9 : _GEN_26062; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26064 = 10'h1fb == _T_512[9:0] ? 4'hd : _GEN_26063; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26065 = 10'h1fc == _T_512[9:0] ? 4'hd : _GEN_26064; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26066 = 10'h1fd == _T_512[9:0] ? 4'h2 : _GEN_26065; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26067 = 10'h1fe == _T_512[9:0] ? 4'hd : _GEN_26066; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26068 = 10'h1ff == _T_512[9:0] ? 4'h0 : _GEN_26067; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26069 = 10'h200 == _T_512[9:0] ? 4'hd : _GEN_26068; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26070 = 10'h201 == _T_512[9:0] ? 4'hd : _GEN_26069; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26071 = 10'h202 == _T_512[9:0] ? 4'h3 : _GEN_26070; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26072 = 10'h203 == _T_512[9:0] ? 4'hd : _GEN_26071; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26073 = 10'h204 == _T_512[9:0] ? 4'hd : _GEN_26072; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26074 = 10'h205 == _T_512[9:0] ? 4'hd : _GEN_26073; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26075 = 10'h206 == _T_512[9:0] ? 4'hb : _GEN_26074; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26076 = 10'h207 == _T_512[9:0] ? 4'hb : _GEN_26075; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26077 = 10'h208 == _T_512[9:0] ? 4'hd : _GEN_26076; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26078 = 10'h209 == _T_512[9:0] ? 4'hd : _GEN_26077; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26079 = 10'h20a == _T_512[9:0] ? 4'hd : _GEN_26078; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26080 = 10'h20b == _T_512[9:0] ? 4'hb : _GEN_26079; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26081 = 10'h20c == _T_512[9:0] ? 4'hd : _GEN_26080; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26082 = 10'h20d == _T_512[9:0] ? 4'hb : _GEN_26081; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26083 = 10'h20e == _T_512[9:0] ? 4'hd : _GEN_26082; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26084 = 10'h20f == _T_512[9:0] ? 4'hb : _GEN_26083; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26085 = 10'h210 == _T_512[9:0] ? 4'hd : _GEN_26084; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26086 = 10'h211 == _T_512[9:0] ? 4'hd : _GEN_26085; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26087 = 10'h212 == _T_512[9:0] ? 4'hb : _GEN_26086; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26088 = 10'h213 == _T_512[9:0] ? 4'hb : _GEN_26087; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26089 = 10'h214 == _T_512[9:0] ? 4'hb : _GEN_26088; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26090 = 10'h215 == _T_512[9:0] ? 4'hd : _GEN_26089; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26091 = 10'h216 == _T_512[9:0] ? 4'hd : _GEN_26090; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26092 = 10'h217 == _T_512[9:0] ? 4'hd : _GEN_26091; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26093 = 10'h218 == _T_512[9:0] ? 4'hd : _GEN_26092; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26094 = 10'h219 == _T_512[9:0] ? 4'hd : _GEN_26093; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26095 = 10'h21a == _T_512[9:0] ? 4'hd : _GEN_26094; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26096 = 10'h21b == _T_512[9:0] ? 4'hd : _GEN_26095; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26097 = 10'h21c == _T_512[9:0] ? 4'h3 : _GEN_26096; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26098 = 10'h21d == _T_512[9:0] ? 4'h2 : _GEN_26097; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26099 = 10'h21e == _T_512[9:0] ? 4'hd : _GEN_26098; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26100 = 10'h21f == _T_512[9:0] ? 4'h0 : _GEN_26099; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26101 = 10'h220 == _T_512[9:0] ? 4'h0 : _GEN_26100; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26102 = 10'h221 == _T_512[9:0] ? 4'h0 : _GEN_26101; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26103 = 10'h222 == _T_512[9:0] ? 4'h0 : _GEN_26102; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26104 = 10'h223 == _T_512[9:0] ? 4'h0 : _GEN_26103; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26105 = 10'h224 == _T_512[9:0] ? 4'h0 : _GEN_26104; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26106 = 10'h225 == _T_512[9:0] ? 4'h0 : _GEN_26105; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26107 = 10'h226 == _T_512[9:0] ? 4'h0 : _GEN_26106; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26108 = 10'h227 == _T_512[9:0] ? 4'h0 : _GEN_26107; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26109 = 10'h228 == _T_512[9:0] ? 4'h0 : _GEN_26108; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26110 = 10'h229 == _T_512[9:0] ? 4'h0 : _GEN_26109; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26111 = 10'h22a == _T_512[9:0] ? 4'h0 : _GEN_26110; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26112 = 10'h22b == _T_512[9:0] ? 4'h0 : _GEN_26111; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26113 = 10'h22c == _T_512[9:0] ? 4'h0 : _GEN_26112; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26114 = 10'h22d == _T_512[9:0] ? 4'h0 : _GEN_26113; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26115 = 10'h22e == _T_512[9:0] ? 4'h0 : _GEN_26114; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26116 = 10'h22f == _T_512[9:0] ? 4'h0 : _GEN_26115; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26117 = 10'h230 == _T_512[9:0] ? 4'h0 : _GEN_26116; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26118 = 10'h231 == _T_512[9:0] ? 4'h0 : _GEN_26117; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26119 = 10'h232 == _T_512[9:0] ? 4'h0 : _GEN_26118; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26120 = 10'h233 == _T_512[9:0] ? 4'h0 : _GEN_26119; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26121 = 10'h234 == _T_512[9:0] ? 4'h0 : _GEN_26120; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26122 = 10'h235 == _T_512[9:0] ? 4'h0 : _GEN_26121; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26123 = 10'h236 == _T_512[9:0] ? 4'h0 : _GEN_26122; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26124 = 10'h237 == _T_512[9:0] ? 4'h0 : _GEN_26123; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26125 = 10'h238 == _T_512[9:0] ? 4'h0 : _GEN_26124; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26126 = 10'h239 == _T_512[9:0] ? 4'h0 : _GEN_26125; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26127 = 10'h23a == _T_512[9:0] ? 4'h0 : _GEN_26126; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26128 = 10'h23b == _T_512[9:0] ? 4'h0 : _GEN_26127; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26129 = 10'h23c == _T_512[9:0] ? 4'h0 : _GEN_26128; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26130 = 10'h23d == _T_512[9:0] ? 4'h0 : _GEN_26129; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26131 = 10'h23e == _T_512[9:0] ? 4'h0 : _GEN_26130; // @[Filter.scala 191:142]
  wire [3:0] _GEN_26132 = 10'h23f == _T_512[9:0] ? 4'h0 : _GEN_26131; // @[Filter.scala 191:142]
  wire [7:0] _T_526 = _GEN_26132 * 4'ha; // @[Filter.scala 191:142]
  wire [10:0] _GEN_28387 = {{3'd0}, _T_526}; // @[Filter.scala 191:109]
  wire [10:0] _T_528 = _T_521 + _GEN_28387; // @[Filter.scala 191:109]
  wire [10:0] _T_529 = _T_528 / 11'h64; // @[Filter.scala 191:150]
  wire  _T_531 = _T_502 >= 6'h20; // @[Filter.scala 194:31]
  wire  _T_535 = _T_509 >= 32'h12; // @[Filter.scala 194:63]
  wire  _T_536 = _T_531 | _T_535; // @[Filter.scala 194:58]
  wire [10:0] _GEN_26709 = io_SPI_distort ? _T_529 : {{7'd0}, _GEN_24980}; // @[Filter.scala 196:35]
  wire [10:0] _GEN_26710 = _T_536 ? 11'h0 : _GEN_26709; // @[Filter.scala 194:80]
  wire [10:0] _GEN_27287 = io_SPI_distort ? _T_529 : {{7'd0}, _GEN_25556}; // @[Filter.scala 196:35]
  wire [10:0] _GEN_27288 = _T_536 ? 11'h0 : _GEN_27287; // @[Filter.scala 194:80]
  wire [10:0] _GEN_27865 = io_SPI_distort ? _T_529 : {{7'd0}, _GEN_26132}; // @[Filter.scala 196:35]
  wire [10:0] _GEN_27866 = _T_536 ? 11'h0 : _GEN_27865; // @[Filter.scala 194:80]
  reg [8:0] pixOut_0_0; // @[Filter.scala 205:32]
  reg [8:0] pixOut_0_1; // @[Filter.scala 205:32]
  reg [8:0] pixOut_0_2; // @[Filter.scala 205:32]
  reg [8:0] pixOut_0_3; // @[Filter.scala 205:32]
  reg [8:0] pixOut_0_4; // @[Filter.scala 205:32]
  reg [8:0] pixOut_0_5; // @[Filter.scala 205:32]
  reg [8:0] pixOut_0_6; // @[Filter.scala 205:32]
  reg [8:0] pixOut_0_7; // @[Filter.scala 205:32]
  reg [8:0] pixOut_1_0; // @[Filter.scala 205:87]
  reg [8:0] pixOut_1_1; // @[Filter.scala 205:87]
  reg [8:0] pixOut_1_2; // @[Filter.scala 205:87]
  reg [8:0] pixOut_1_3; // @[Filter.scala 205:87]
  reg [8:0] pixOut_1_4; // @[Filter.scala 205:87]
  reg [8:0] pixOut_1_5; // @[Filter.scala 205:87]
  reg [8:0] pixOut_1_6; // @[Filter.scala 205:87]
  reg [8:0] pixOut_1_7; // @[Filter.scala 205:87]
  reg [8:0] pixOut_2_0; // @[Filter.scala 205:142]
  reg [8:0] pixOut_2_1; // @[Filter.scala 205:142]
  reg [8:0] pixOut_2_2; // @[Filter.scala 205:142]
  reg [8:0] pixOut_2_3; // @[Filter.scala 205:142]
  reg [8:0] pixOut_2_4; // @[Filter.scala 205:142]
  reg [8:0] pixOut_2_5; // @[Filter.scala 205:142]
  reg [8:0] pixOut_2_6; // @[Filter.scala 205:142]
  reg [8:0] pixOut_2_7; // @[Filter.scala 205:142]
  reg  validOut; // @[Filter.scala 206:29]
  wire [7:0] _GEN_27868 = 3'h1 == io_SPI_filterIndex[2:0] ? $signed(8'sh9) : $signed(8'sh1); // @[Filter.scala 210:64]
  wire [7:0] _GEN_27869 = 3'h2 == io_SPI_filterIndex[2:0] ? $signed(8'sh10) : $signed(_GEN_27868); // @[Filter.scala 210:64]
  wire [7:0] _GEN_27870 = 3'h3 == io_SPI_filterIndex[2:0] ? $signed(8'sh1) : $signed(_GEN_27869); // @[Filter.scala 210:64]
  wire [7:0] _GEN_27871 = 3'h4 == io_SPI_filterIndex[2:0] ? $signed(8'sh1) : $signed(_GEN_27870); // @[Filter.scala 210:64]
  wire [7:0] _GEN_27872 = 3'h5 == io_SPI_filterIndex[2:0] ? $signed(8'sh1) : $signed(_GEN_27871); // @[Filter.scala 210:64]
  wire [8:0] _GEN_28391 = {{1{_GEN_27872[7]}},_GEN_27872}; // @[Filter.scala 210:64]
  wire [9:0] _T_567 = $signed(KernelConvolution_io_pixelVal_out_0) / $signed(_GEN_28391); // @[Filter.scala 210:64]
  wire  _T_568 = $signed(pixOut_0_0) < 9'sh0; // @[Filter.scala 212:30]
  wire  _T_569 = _T_568 & io_SPI_invert; // @[Filter.scala 212:36]
  wire  _T_571 = $signed(pixOut_0_0) > 9'shf; // @[Filter.scala 217:36]
  wire  _T_572 = _T_571 & io_SPI_invert; // @[Filter.scala 217:43]
  wire [8:0] _T_576 = 9'hf - pixOut_0_0; // @[Filter.scala 222:43]
  wire [8:0] _GEN_27873 = io_SPI_invert ? _T_576 : pixOut_0_0; // @[Filter.scala 221:36]
  wire [8:0] _GEN_27874 = _T_571 ? 9'hf : _GEN_27873; // @[Filter.scala 219:44]
  wire [8:0] _GEN_27875 = _T_572 ? 9'h0 : _GEN_27874; // @[Filter.scala 217:59]
  wire [8:0] _GEN_27876 = _T_568 ? 9'h0 : _GEN_27875; // @[Filter.scala 214:43]
  wire [8:0] _GEN_27877 = _T_569 ? 9'hf : _GEN_27876; // @[Filter.scala 212:52]
  wire [9:0] _T_578 = $signed(KernelConvolution_io_pixelVal_out_1) / $signed(_GEN_28391); // @[Filter.scala 210:64]
  wire  _T_579 = $signed(pixOut_0_1) < 9'sh0; // @[Filter.scala 212:30]
  wire  _T_580 = _T_579 & io_SPI_invert; // @[Filter.scala 212:36]
  wire  _T_582 = $signed(pixOut_0_1) > 9'shf; // @[Filter.scala 217:36]
  wire  _T_583 = _T_582 & io_SPI_invert; // @[Filter.scala 217:43]
  wire [8:0] _T_587 = 9'hf - pixOut_0_1; // @[Filter.scala 222:43]
  wire [8:0] _GEN_27878 = io_SPI_invert ? _T_587 : pixOut_0_1; // @[Filter.scala 221:36]
  wire [8:0] _GEN_27879 = _T_582 ? 9'hf : _GEN_27878; // @[Filter.scala 219:44]
  wire [8:0] _GEN_27880 = _T_583 ? 9'h0 : _GEN_27879; // @[Filter.scala 217:59]
  wire [8:0] _GEN_27881 = _T_579 ? 9'h0 : _GEN_27880; // @[Filter.scala 214:43]
  wire [8:0] _GEN_27882 = _T_580 ? 9'hf : _GEN_27881; // @[Filter.scala 212:52]
  wire [9:0] _T_589 = $signed(KernelConvolution_io_pixelVal_out_2) / $signed(_GEN_28391); // @[Filter.scala 210:64]
  wire  _T_590 = $signed(pixOut_0_2) < 9'sh0; // @[Filter.scala 212:30]
  wire  _T_591 = _T_590 & io_SPI_invert; // @[Filter.scala 212:36]
  wire  _T_593 = $signed(pixOut_0_2) > 9'shf; // @[Filter.scala 217:36]
  wire  _T_594 = _T_593 & io_SPI_invert; // @[Filter.scala 217:43]
  wire [8:0] _T_598 = 9'hf - pixOut_0_2; // @[Filter.scala 222:43]
  wire [8:0] _GEN_27883 = io_SPI_invert ? _T_598 : pixOut_0_2; // @[Filter.scala 221:36]
  wire [8:0] _GEN_27884 = _T_593 ? 9'hf : _GEN_27883; // @[Filter.scala 219:44]
  wire [8:0] _GEN_27885 = _T_594 ? 9'h0 : _GEN_27884; // @[Filter.scala 217:59]
  wire [8:0] _GEN_27886 = _T_590 ? 9'h0 : _GEN_27885; // @[Filter.scala 214:43]
  wire [8:0] _GEN_27887 = _T_591 ? 9'hf : _GEN_27886; // @[Filter.scala 212:52]
  wire [9:0] _T_600 = $signed(KernelConvolution_io_pixelVal_out_3) / $signed(_GEN_28391); // @[Filter.scala 210:64]
  wire  _T_601 = $signed(pixOut_0_3) < 9'sh0; // @[Filter.scala 212:30]
  wire  _T_602 = _T_601 & io_SPI_invert; // @[Filter.scala 212:36]
  wire  _T_604 = $signed(pixOut_0_3) > 9'shf; // @[Filter.scala 217:36]
  wire  _T_605 = _T_604 & io_SPI_invert; // @[Filter.scala 217:43]
  wire [8:0] _T_609 = 9'hf - pixOut_0_3; // @[Filter.scala 222:43]
  wire [8:0] _GEN_27888 = io_SPI_invert ? _T_609 : pixOut_0_3; // @[Filter.scala 221:36]
  wire [8:0] _GEN_27889 = _T_604 ? 9'hf : _GEN_27888; // @[Filter.scala 219:44]
  wire [8:0] _GEN_27890 = _T_605 ? 9'h0 : _GEN_27889; // @[Filter.scala 217:59]
  wire [8:0] _GEN_27891 = _T_601 ? 9'h0 : _GEN_27890; // @[Filter.scala 214:43]
  wire [8:0] _GEN_27892 = _T_602 ? 9'hf : _GEN_27891; // @[Filter.scala 212:52]
  wire [9:0] _T_611 = $signed(KernelConvolution_io_pixelVal_out_4) / $signed(_GEN_28391); // @[Filter.scala 210:64]
  wire  _T_612 = $signed(pixOut_0_4) < 9'sh0; // @[Filter.scala 212:30]
  wire  _T_613 = _T_612 & io_SPI_invert; // @[Filter.scala 212:36]
  wire  _T_615 = $signed(pixOut_0_4) > 9'shf; // @[Filter.scala 217:36]
  wire  _T_616 = _T_615 & io_SPI_invert; // @[Filter.scala 217:43]
  wire [8:0] _T_620 = 9'hf - pixOut_0_4; // @[Filter.scala 222:43]
  wire [8:0] _GEN_27893 = io_SPI_invert ? _T_620 : pixOut_0_4; // @[Filter.scala 221:36]
  wire [8:0] _GEN_27894 = _T_615 ? 9'hf : _GEN_27893; // @[Filter.scala 219:44]
  wire [8:0] _GEN_27895 = _T_616 ? 9'h0 : _GEN_27894; // @[Filter.scala 217:59]
  wire [8:0] _GEN_27896 = _T_612 ? 9'h0 : _GEN_27895; // @[Filter.scala 214:43]
  wire [8:0] _GEN_27897 = _T_613 ? 9'hf : _GEN_27896; // @[Filter.scala 212:52]
  wire [9:0] _T_622 = $signed(KernelConvolution_io_pixelVal_out_5) / $signed(_GEN_28391); // @[Filter.scala 210:64]
  wire  _T_623 = $signed(pixOut_0_5) < 9'sh0; // @[Filter.scala 212:30]
  wire  _T_624 = _T_623 & io_SPI_invert; // @[Filter.scala 212:36]
  wire  _T_626 = $signed(pixOut_0_5) > 9'shf; // @[Filter.scala 217:36]
  wire  _T_627 = _T_626 & io_SPI_invert; // @[Filter.scala 217:43]
  wire [8:0] _T_631 = 9'hf - pixOut_0_5; // @[Filter.scala 222:43]
  wire [8:0] _GEN_27898 = io_SPI_invert ? _T_631 : pixOut_0_5; // @[Filter.scala 221:36]
  wire [8:0] _GEN_27899 = _T_626 ? 9'hf : _GEN_27898; // @[Filter.scala 219:44]
  wire [8:0] _GEN_27900 = _T_627 ? 9'h0 : _GEN_27899; // @[Filter.scala 217:59]
  wire [8:0] _GEN_27901 = _T_623 ? 9'h0 : _GEN_27900; // @[Filter.scala 214:43]
  wire [8:0] _GEN_27902 = _T_624 ? 9'hf : _GEN_27901; // @[Filter.scala 212:52]
  wire [9:0] _T_633 = $signed(KernelConvolution_io_pixelVal_out_6) / $signed(_GEN_28391); // @[Filter.scala 210:64]
  wire  _T_634 = $signed(pixOut_0_6) < 9'sh0; // @[Filter.scala 212:30]
  wire  _T_635 = _T_634 & io_SPI_invert; // @[Filter.scala 212:36]
  wire  _T_637 = $signed(pixOut_0_6) > 9'shf; // @[Filter.scala 217:36]
  wire  _T_638 = _T_637 & io_SPI_invert; // @[Filter.scala 217:43]
  wire [8:0] _T_642 = 9'hf - pixOut_0_6; // @[Filter.scala 222:43]
  wire [8:0] _GEN_27903 = io_SPI_invert ? _T_642 : pixOut_0_6; // @[Filter.scala 221:36]
  wire [8:0] _GEN_27904 = _T_637 ? 9'hf : _GEN_27903; // @[Filter.scala 219:44]
  wire [8:0] _GEN_27905 = _T_638 ? 9'h0 : _GEN_27904; // @[Filter.scala 217:59]
  wire [8:0] _GEN_27906 = _T_634 ? 9'h0 : _GEN_27905; // @[Filter.scala 214:43]
  wire [8:0] _GEN_27907 = _T_635 ? 9'hf : _GEN_27906; // @[Filter.scala 212:52]
  wire [9:0] _T_644 = $signed(KernelConvolution_io_pixelVal_out_7) / $signed(_GEN_28391); // @[Filter.scala 210:64]
  wire  _T_645 = $signed(pixOut_0_7) < 9'sh0; // @[Filter.scala 212:30]
  wire  _T_646 = _T_645 & io_SPI_invert; // @[Filter.scala 212:36]
  wire  _T_648 = $signed(pixOut_0_7) > 9'shf; // @[Filter.scala 217:36]
  wire  _T_649 = _T_648 & io_SPI_invert; // @[Filter.scala 217:43]
  wire [8:0] _T_653 = 9'hf - pixOut_0_7; // @[Filter.scala 222:43]
  wire [8:0] _GEN_27908 = io_SPI_invert ? _T_653 : pixOut_0_7; // @[Filter.scala 221:36]
  wire [8:0] _GEN_27909 = _T_648 ? 9'hf : _GEN_27908; // @[Filter.scala 219:44]
  wire [8:0] _GEN_27910 = _T_649 ? 9'h0 : _GEN_27909; // @[Filter.scala 217:59]
  wire [8:0] _GEN_27911 = _T_645 ? 9'h0 : _GEN_27910; // @[Filter.scala 214:43]
  wire [8:0] _GEN_27912 = _T_646 ? 9'hf : _GEN_27911; // @[Filter.scala 212:52]
  wire [9:0] _T_655 = $signed(KernelConvolution_1_io_pixelVal_out_0) / $signed(_GEN_28391); // @[Filter.scala 210:64]
  wire  _T_656 = $signed(pixOut_1_0) < 9'sh0; // @[Filter.scala 212:30]
  wire  _T_657 = _T_656 & io_SPI_invert; // @[Filter.scala 212:36]
  wire  _T_659 = $signed(pixOut_1_0) > 9'shf; // @[Filter.scala 217:36]
  wire  _T_660 = _T_659 & io_SPI_invert; // @[Filter.scala 217:43]
  wire [8:0] _T_664 = 9'hf - pixOut_1_0; // @[Filter.scala 222:43]
  wire [8:0] _GEN_27913 = io_SPI_invert ? _T_664 : pixOut_1_0; // @[Filter.scala 221:36]
  wire [8:0] _GEN_27914 = _T_659 ? 9'hf : _GEN_27913; // @[Filter.scala 219:44]
  wire [8:0] _GEN_27915 = _T_660 ? 9'h0 : _GEN_27914; // @[Filter.scala 217:59]
  wire [8:0] _GEN_27916 = _T_656 ? 9'h0 : _GEN_27915; // @[Filter.scala 214:43]
  wire [8:0] _GEN_27917 = _T_657 ? 9'hf : _GEN_27916; // @[Filter.scala 212:52]
  wire [9:0] _T_666 = $signed(KernelConvolution_1_io_pixelVal_out_1) / $signed(_GEN_28391); // @[Filter.scala 210:64]
  wire  _T_667 = $signed(pixOut_1_1) < 9'sh0; // @[Filter.scala 212:30]
  wire  _T_668 = _T_667 & io_SPI_invert; // @[Filter.scala 212:36]
  wire  _T_670 = $signed(pixOut_1_1) > 9'shf; // @[Filter.scala 217:36]
  wire  _T_671 = _T_670 & io_SPI_invert; // @[Filter.scala 217:43]
  wire [8:0] _T_675 = 9'hf - pixOut_1_1; // @[Filter.scala 222:43]
  wire [8:0] _GEN_27918 = io_SPI_invert ? _T_675 : pixOut_1_1; // @[Filter.scala 221:36]
  wire [8:0] _GEN_27919 = _T_670 ? 9'hf : _GEN_27918; // @[Filter.scala 219:44]
  wire [8:0] _GEN_27920 = _T_671 ? 9'h0 : _GEN_27919; // @[Filter.scala 217:59]
  wire [8:0] _GEN_27921 = _T_667 ? 9'h0 : _GEN_27920; // @[Filter.scala 214:43]
  wire [8:0] _GEN_27922 = _T_668 ? 9'hf : _GEN_27921; // @[Filter.scala 212:52]
  wire [9:0] _T_677 = $signed(KernelConvolution_1_io_pixelVal_out_2) / $signed(_GEN_28391); // @[Filter.scala 210:64]
  wire  _T_678 = $signed(pixOut_1_2) < 9'sh0; // @[Filter.scala 212:30]
  wire  _T_679 = _T_678 & io_SPI_invert; // @[Filter.scala 212:36]
  wire  _T_681 = $signed(pixOut_1_2) > 9'shf; // @[Filter.scala 217:36]
  wire  _T_682 = _T_681 & io_SPI_invert; // @[Filter.scala 217:43]
  wire [8:0] _T_686 = 9'hf - pixOut_1_2; // @[Filter.scala 222:43]
  wire [8:0] _GEN_27923 = io_SPI_invert ? _T_686 : pixOut_1_2; // @[Filter.scala 221:36]
  wire [8:0] _GEN_27924 = _T_681 ? 9'hf : _GEN_27923; // @[Filter.scala 219:44]
  wire [8:0] _GEN_27925 = _T_682 ? 9'h0 : _GEN_27924; // @[Filter.scala 217:59]
  wire [8:0] _GEN_27926 = _T_678 ? 9'h0 : _GEN_27925; // @[Filter.scala 214:43]
  wire [8:0] _GEN_27927 = _T_679 ? 9'hf : _GEN_27926; // @[Filter.scala 212:52]
  wire [9:0] _T_688 = $signed(KernelConvolution_1_io_pixelVal_out_3) / $signed(_GEN_28391); // @[Filter.scala 210:64]
  wire  _T_689 = $signed(pixOut_1_3) < 9'sh0; // @[Filter.scala 212:30]
  wire  _T_690 = _T_689 & io_SPI_invert; // @[Filter.scala 212:36]
  wire  _T_692 = $signed(pixOut_1_3) > 9'shf; // @[Filter.scala 217:36]
  wire  _T_693 = _T_692 & io_SPI_invert; // @[Filter.scala 217:43]
  wire [8:0] _T_697 = 9'hf - pixOut_1_3; // @[Filter.scala 222:43]
  wire [8:0] _GEN_27928 = io_SPI_invert ? _T_697 : pixOut_1_3; // @[Filter.scala 221:36]
  wire [8:0] _GEN_27929 = _T_692 ? 9'hf : _GEN_27928; // @[Filter.scala 219:44]
  wire [8:0] _GEN_27930 = _T_693 ? 9'h0 : _GEN_27929; // @[Filter.scala 217:59]
  wire [8:0] _GEN_27931 = _T_689 ? 9'h0 : _GEN_27930; // @[Filter.scala 214:43]
  wire [8:0] _GEN_27932 = _T_690 ? 9'hf : _GEN_27931; // @[Filter.scala 212:52]
  wire [9:0] _T_699 = $signed(KernelConvolution_1_io_pixelVal_out_4) / $signed(_GEN_28391); // @[Filter.scala 210:64]
  wire  _T_700 = $signed(pixOut_1_4) < 9'sh0; // @[Filter.scala 212:30]
  wire  _T_701 = _T_700 & io_SPI_invert; // @[Filter.scala 212:36]
  wire  _T_703 = $signed(pixOut_1_4) > 9'shf; // @[Filter.scala 217:36]
  wire  _T_704 = _T_703 & io_SPI_invert; // @[Filter.scala 217:43]
  wire [8:0] _T_708 = 9'hf - pixOut_1_4; // @[Filter.scala 222:43]
  wire [8:0] _GEN_27933 = io_SPI_invert ? _T_708 : pixOut_1_4; // @[Filter.scala 221:36]
  wire [8:0] _GEN_27934 = _T_703 ? 9'hf : _GEN_27933; // @[Filter.scala 219:44]
  wire [8:0] _GEN_27935 = _T_704 ? 9'h0 : _GEN_27934; // @[Filter.scala 217:59]
  wire [8:0] _GEN_27936 = _T_700 ? 9'h0 : _GEN_27935; // @[Filter.scala 214:43]
  wire [8:0] _GEN_27937 = _T_701 ? 9'hf : _GEN_27936; // @[Filter.scala 212:52]
  wire [9:0] _T_710 = $signed(KernelConvolution_1_io_pixelVal_out_5) / $signed(_GEN_28391); // @[Filter.scala 210:64]
  wire  _T_711 = $signed(pixOut_1_5) < 9'sh0; // @[Filter.scala 212:30]
  wire  _T_712 = _T_711 & io_SPI_invert; // @[Filter.scala 212:36]
  wire  _T_714 = $signed(pixOut_1_5) > 9'shf; // @[Filter.scala 217:36]
  wire  _T_715 = _T_714 & io_SPI_invert; // @[Filter.scala 217:43]
  wire [8:0] _T_719 = 9'hf - pixOut_1_5; // @[Filter.scala 222:43]
  wire [8:0] _GEN_27938 = io_SPI_invert ? _T_719 : pixOut_1_5; // @[Filter.scala 221:36]
  wire [8:0] _GEN_27939 = _T_714 ? 9'hf : _GEN_27938; // @[Filter.scala 219:44]
  wire [8:0] _GEN_27940 = _T_715 ? 9'h0 : _GEN_27939; // @[Filter.scala 217:59]
  wire [8:0] _GEN_27941 = _T_711 ? 9'h0 : _GEN_27940; // @[Filter.scala 214:43]
  wire [8:0] _GEN_27942 = _T_712 ? 9'hf : _GEN_27941; // @[Filter.scala 212:52]
  wire [9:0] _T_721 = $signed(KernelConvolution_1_io_pixelVal_out_6) / $signed(_GEN_28391); // @[Filter.scala 210:64]
  wire  _T_722 = $signed(pixOut_1_6) < 9'sh0; // @[Filter.scala 212:30]
  wire  _T_723 = _T_722 & io_SPI_invert; // @[Filter.scala 212:36]
  wire  _T_725 = $signed(pixOut_1_6) > 9'shf; // @[Filter.scala 217:36]
  wire  _T_726 = _T_725 & io_SPI_invert; // @[Filter.scala 217:43]
  wire [8:0] _T_730 = 9'hf - pixOut_1_6; // @[Filter.scala 222:43]
  wire [8:0] _GEN_27943 = io_SPI_invert ? _T_730 : pixOut_1_6; // @[Filter.scala 221:36]
  wire [8:0] _GEN_27944 = _T_725 ? 9'hf : _GEN_27943; // @[Filter.scala 219:44]
  wire [8:0] _GEN_27945 = _T_726 ? 9'h0 : _GEN_27944; // @[Filter.scala 217:59]
  wire [8:0] _GEN_27946 = _T_722 ? 9'h0 : _GEN_27945; // @[Filter.scala 214:43]
  wire [8:0] _GEN_27947 = _T_723 ? 9'hf : _GEN_27946; // @[Filter.scala 212:52]
  wire [9:0] _T_732 = $signed(KernelConvolution_1_io_pixelVal_out_7) / $signed(_GEN_28391); // @[Filter.scala 210:64]
  wire  _T_733 = $signed(pixOut_1_7) < 9'sh0; // @[Filter.scala 212:30]
  wire  _T_734 = _T_733 & io_SPI_invert; // @[Filter.scala 212:36]
  wire  _T_736 = $signed(pixOut_1_7) > 9'shf; // @[Filter.scala 217:36]
  wire  _T_737 = _T_736 & io_SPI_invert; // @[Filter.scala 217:43]
  wire [8:0] _T_741 = 9'hf - pixOut_1_7; // @[Filter.scala 222:43]
  wire [8:0] _GEN_27948 = io_SPI_invert ? _T_741 : pixOut_1_7; // @[Filter.scala 221:36]
  wire [8:0] _GEN_27949 = _T_736 ? 9'hf : _GEN_27948; // @[Filter.scala 219:44]
  wire [8:0] _GEN_27950 = _T_737 ? 9'h0 : _GEN_27949; // @[Filter.scala 217:59]
  wire [8:0] _GEN_27951 = _T_733 ? 9'h0 : _GEN_27950; // @[Filter.scala 214:43]
  wire [8:0] _GEN_27952 = _T_734 ? 9'hf : _GEN_27951; // @[Filter.scala 212:52]
  wire [9:0] _T_743 = $signed(KernelConvolution_2_io_pixelVal_out_0) / $signed(_GEN_28391); // @[Filter.scala 210:64]
  wire  _T_744 = $signed(pixOut_2_0) < 9'sh0; // @[Filter.scala 212:30]
  wire  _T_745 = _T_744 & io_SPI_invert; // @[Filter.scala 212:36]
  wire  _T_747 = $signed(pixOut_2_0) > 9'shf; // @[Filter.scala 217:36]
  wire  _T_748 = _T_747 & io_SPI_invert; // @[Filter.scala 217:43]
  wire [8:0] _T_752 = 9'hf - pixOut_2_0; // @[Filter.scala 222:43]
  wire [8:0] _GEN_27953 = io_SPI_invert ? _T_752 : pixOut_2_0; // @[Filter.scala 221:36]
  wire [8:0] _GEN_27954 = _T_747 ? 9'hf : _GEN_27953; // @[Filter.scala 219:44]
  wire [8:0] _GEN_27955 = _T_748 ? 9'h0 : _GEN_27954; // @[Filter.scala 217:59]
  wire [8:0] _GEN_27956 = _T_744 ? 9'h0 : _GEN_27955; // @[Filter.scala 214:43]
  wire [8:0] _GEN_27957 = _T_745 ? 9'hf : _GEN_27956; // @[Filter.scala 212:52]
  wire [9:0] _T_754 = $signed(KernelConvolution_2_io_pixelVal_out_1) / $signed(_GEN_28391); // @[Filter.scala 210:64]
  wire  _T_755 = $signed(pixOut_2_1) < 9'sh0; // @[Filter.scala 212:30]
  wire  _T_756 = _T_755 & io_SPI_invert; // @[Filter.scala 212:36]
  wire  _T_758 = $signed(pixOut_2_1) > 9'shf; // @[Filter.scala 217:36]
  wire  _T_759 = _T_758 & io_SPI_invert; // @[Filter.scala 217:43]
  wire [8:0] _T_763 = 9'hf - pixOut_2_1; // @[Filter.scala 222:43]
  wire [8:0] _GEN_27958 = io_SPI_invert ? _T_763 : pixOut_2_1; // @[Filter.scala 221:36]
  wire [8:0] _GEN_27959 = _T_758 ? 9'hf : _GEN_27958; // @[Filter.scala 219:44]
  wire [8:0] _GEN_27960 = _T_759 ? 9'h0 : _GEN_27959; // @[Filter.scala 217:59]
  wire [8:0] _GEN_27961 = _T_755 ? 9'h0 : _GEN_27960; // @[Filter.scala 214:43]
  wire [8:0] _GEN_27962 = _T_756 ? 9'hf : _GEN_27961; // @[Filter.scala 212:52]
  wire [9:0] _T_765 = $signed(KernelConvolution_2_io_pixelVal_out_2) / $signed(_GEN_28391); // @[Filter.scala 210:64]
  wire  _T_766 = $signed(pixOut_2_2) < 9'sh0; // @[Filter.scala 212:30]
  wire  _T_767 = _T_766 & io_SPI_invert; // @[Filter.scala 212:36]
  wire  _T_769 = $signed(pixOut_2_2) > 9'shf; // @[Filter.scala 217:36]
  wire  _T_770 = _T_769 & io_SPI_invert; // @[Filter.scala 217:43]
  wire [8:0] _T_774 = 9'hf - pixOut_2_2; // @[Filter.scala 222:43]
  wire [8:0] _GEN_27963 = io_SPI_invert ? _T_774 : pixOut_2_2; // @[Filter.scala 221:36]
  wire [8:0] _GEN_27964 = _T_769 ? 9'hf : _GEN_27963; // @[Filter.scala 219:44]
  wire [8:0] _GEN_27965 = _T_770 ? 9'h0 : _GEN_27964; // @[Filter.scala 217:59]
  wire [8:0] _GEN_27966 = _T_766 ? 9'h0 : _GEN_27965; // @[Filter.scala 214:43]
  wire [8:0] _GEN_27967 = _T_767 ? 9'hf : _GEN_27966; // @[Filter.scala 212:52]
  wire [9:0] _T_776 = $signed(KernelConvolution_2_io_pixelVal_out_3) / $signed(_GEN_28391); // @[Filter.scala 210:64]
  wire  _T_777 = $signed(pixOut_2_3) < 9'sh0; // @[Filter.scala 212:30]
  wire  _T_778 = _T_777 & io_SPI_invert; // @[Filter.scala 212:36]
  wire  _T_780 = $signed(pixOut_2_3) > 9'shf; // @[Filter.scala 217:36]
  wire  _T_781 = _T_780 & io_SPI_invert; // @[Filter.scala 217:43]
  wire [8:0] _T_785 = 9'hf - pixOut_2_3; // @[Filter.scala 222:43]
  wire [8:0] _GEN_27968 = io_SPI_invert ? _T_785 : pixOut_2_3; // @[Filter.scala 221:36]
  wire [8:0] _GEN_27969 = _T_780 ? 9'hf : _GEN_27968; // @[Filter.scala 219:44]
  wire [8:0] _GEN_27970 = _T_781 ? 9'h0 : _GEN_27969; // @[Filter.scala 217:59]
  wire [8:0] _GEN_27971 = _T_777 ? 9'h0 : _GEN_27970; // @[Filter.scala 214:43]
  wire [8:0] _GEN_27972 = _T_778 ? 9'hf : _GEN_27971; // @[Filter.scala 212:52]
  wire [9:0] _T_787 = $signed(KernelConvolution_2_io_pixelVal_out_4) / $signed(_GEN_28391); // @[Filter.scala 210:64]
  wire  _T_788 = $signed(pixOut_2_4) < 9'sh0; // @[Filter.scala 212:30]
  wire  _T_789 = _T_788 & io_SPI_invert; // @[Filter.scala 212:36]
  wire  _T_791 = $signed(pixOut_2_4) > 9'shf; // @[Filter.scala 217:36]
  wire  _T_792 = _T_791 & io_SPI_invert; // @[Filter.scala 217:43]
  wire [8:0] _T_796 = 9'hf - pixOut_2_4; // @[Filter.scala 222:43]
  wire [8:0] _GEN_27973 = io_SPI_invert ? _T_796 : pixOut_2_4; // @[Filter.scala 221:36]
  wire [8:0] _GEN_27974 = _T_791 ? 9'hf : _GEN_27973; // @[Filter.scala 219:44]
  wire [8:0] _GEN_27975 = _T_792 ? 9'h0 : _GEN_27974; // @[Filter.scala 217:59]
  wire [8:0] _GEN_27976 = _T_788 ? 9'h0 : _GEN_27975; // @[Filter.scala 214:43]
  wire [8:0] _GEN_27977 = _T_789 ? 9'hf : _GEN_27976; // @[Filter.scala 212:52]
  wire [9:0] _T_798 = $signed(KernelConvolution_2_io_pixelVal_out_5) / $signed(_GEN_28391); // @[Filter.scala 210:64]
  wire  _T_799 = $signed(pixOut_2_5) < 9'sh0; // @[Filter.scala 212:30]
  wire  _T_800 = _T_799 & io_SPI_invert; // @[Filter.scala 212:36]
  wire  _T_802 = $signed(pixOut_2_5) > 9'shf; // @[Filter.scala 217:36]
  wire  _T_803 = _T_802 & io_SPI_invert; // @[Filter.scala 217:43]
  wire [8:0] _T_807 = 9'hf - pixOut_2_5; // @[Filter.scala 222:43]
  wire [8:0] _GEN_27978 = io_SPI_invert ? _T_807 : pixOut_2_5; // @[Filter.scala 221:36]
  wire [8:0] _GEN_27979 = _T_802 ? 9'hf : _GEN_27978; // @[Filter.scala 219:44]
  wire [8:0] _GEN_27980 = _T_803 ? 9'h0 : _GEN_27979; // @[Filter.scala 217:59]
  wire [8:0] _GEN_27981 = _T_799 ? 9'h0 : _GEN_27980; // @[Filter.scala 214:43]
  wire [8:0] _GEN_27982 = _T_800 ? 9'hf : _GEN_27981; // @[Filter.scala 212:52]
  wire [9:0] _T_809 = $signed(KernelConvolution_2_io_pixelVal_out_6) / $signed(_GEN_28391); // @[Filter.scala 210:64]
  wire  _T_810 = $signed(pixOut_2_6) < 9'sh0; // @[Filter.scala 212:30]
  wire  _T_811 = _T_810 & io_SPI_invert; // @[Filter.scala 212:36]
  wire  _T_813 = $signed(pixOut_2_6) > 9'shf; // @[Filter.scala 217:36]
  wire  _T_814 = _T_813 & io_SPI_invert; // @[Filter.scala 217:43]
  wire [8:0] _T_818 = 9'hf - pixOut_2_6; // @[Filter.scala 222:43]
  wire [8:0] _GEN_27983 = io_SPI_invert ? _T_818 : pixOut_2_6; // @[Filter.scala 221:36]
  wire [8:0] _GEN_27984 = _T_813 ? 9'hf : _GEN_27983; // @[Filter.scala 219:44]
  wire [8:0] _GEN_27985 = _T_814 ? 9'h0 : _GEN_27984; // @[Filter.scala 217:59]
  wire [8:0] _GEN_27986 = _T_810 ? 9'h0 : _GEN_27985; // @[Filter.scala 214:43]
  wire [8:0] _GEN_27987 = _T_811 ? 9'hf : _GEN_27986; // @[Filter.scala 212:52]
  wire [9:0] _T_820 = $signed(KernelConvolution_2_io_pixelVal_out_7) / $signed(_GEN_28391); // @[Filter.scala 210:64]
  wire  _T_821 = $signed(pixOut_2_7) < 9'sh0; // @[Filter.scala 212:30]
  wire  _T_822 = _T_821 & io_SPI_invert; // @[Filter.scala 212:36]
  wire  _T_824 = $signed(pixOut_2_7) > 9'shf; // @[Filter.scala 217:36]
  wire  _T_825 = _T_824 & io_SPI_invert; // @[Filter.scala 217:43]
  wire [8:0] _T_829 = 9'hf - pixOut_2_7; // @[Filter.scala 222:43]
  wire [8:0] _GEN_27988 = io_SPI_invert ? _T_829 : pixOut_2_7; // @[Filter.scala 221:36]
  wire [8:0] _GEN_27989 = _T_824 ? 9'hf : _GEN_27988; // @[Filter.scala 219:44]
  wire [8:0] _GEN_27990 = _T_825 ? 9'h0 : _GEN_27989; // @[Filter.scala 217:59]
  wire [8:0] _GEN_27991 = _T_821 ? 9'h0 : _GEN_27990; // @[Filter.scala 214:43]
  wire [8:0] _GEN_27992 = _T_822 ? 9'hf : _GEN_27991; // @[Filter.scala 212:52]
  wire [31:0] _T_832 = pixelIndex + 32'h8; // @[Filter.scala 234:34]
  wire [10:0] _T_833 = 6'h20 * 6'h12; // @[Filter.scala 235:42]
  wire [31:0] _GEN_28415 = {{21'd0}, _T_833}; // @[Filter.scala 235:25]
  wire  _T_834 = pixelIndex == _GEN_28415; // @[Filter.scala 235:25]
  KernelConvolution KernelConvolution ( // @[Filter.scala 173:36]
    .clock(KernelConvolution_clock),
    .reset(KernelConvolution_reset),
    .io_kernelVal_in(KernelConvolution_io_kernelVal_in),
    .io_pixelVal_in_0(KernelConvolution_io_pixelVal_in_0),
    .io_pixelVal_in_1(KernelConvolution_io_pixelVal_in_1),
    .io_pixelVal_in_2(KernelConvolution_io_pixelVal_in_2),
    .io_pixelVal_in_3(KernelConvolution_io_pixelVal_in_3),
    .io_pixelVal_in_4(KernelConvolution_io_pixelVal_in_4),
    .io_pixelVal_in_5(KernelConvolution_io_pixelVal_in_5),
    .io_pixelVal_in_6(KernelConvolution_io_pixelVal_in_6),
    .io_pixelVal_in_7(KernelConvolution_io_pixelVal_in_7),
    .io_pixelVal_out_0(KernelConvolution_io_pixelVal_out_0),
    .io_pixelVal_out_1(KernelConvolution_io_pixelVal_out_1),
    .io_pixelVal_out_2(KernelConvolution_io_pixelVal_out_2),
    .io_pixelVal_out_3(KernelConvolution_io_pixelVal_out_3),
    .io_pixelVal_out_4(KernelConvolution_io_pixelVal_out_4),
    .io_pixelVal_out_5(KernelConvolution_io_pixelVal_out_5),
    .io_pixelVal_out_6(KernelConvolution_io_pixelVal_out_6),
    .io_pixelVal_out_7(KernelConvolution_io_pixelVal_out_7),
    .io_valid_out(KernelConvolution_io_valid_out)
  );
  KernelConvolution KernelConvolution_1 ( // @[Filter.scala 174:36]
    .clock(KernelConvolution_1_clock),
    .reset(KernelConvolution_1_reset),
    .io_kernelVal_in(KernelConvolution_1_io_kernelVal_in),
    .io_pixelVal_in_0(KernelConvolution_1_io_pixelVal_in_0),
    .io_pixelVal_in_1(KernelConvolution_1_io_pixelVal_in_1),
    .io_pixelVal_in_2(KernelConvolution_1_io_pixelVal_in_2),
    .io_pixelVal_in_3(KernelConvolution_1_io_pixelVal_in_3),
    .io_pixelVal_in_4(KernelConvolution_1_io_pixelVal_in_4),
    .io_pixelVal_in_5(KernelConvolution_1_io_pixelVal_in_5),
    .io_pixelVal_in_6(KernelConvolution_1_io_pixelVal_in_6),
    .io_pixelVal_in_7(KernelConvolution_1_io_pixelVal_in_7),
    .io_pixelVal_out_0(KernelConvolution_1_io_pixelVal_out_0),
    .io_pixelVal_out_1(KernelConvolution_1_io_pixelVal_out_1),
    .io_pixelVal_out_2(KernelConvolution_1_io_pixelVal_out_2),
    .io_pixelVal_out_3(KernelConvolution_1_io_pixelVal_out_3),
    .io_pixelVal_out_4(KernelConvolution_1_io_pixelVal_out_4),
    .io_pixelVal_out_5(KernelConvolution_1_io_pixelVal_out_5),
    .io_pixelVal_out_6(KernelConvolution_1_io_pixelVal_out_6),
    .io_pixelVal_out_7(KernelConvolution_1_io_pixelVal_out_7),
    .io_valid_out(KernelConvolution_1_io_valid_out)
  );
  KernelConvolution KernelConvolution_2 ( // @[Filter.scala 175:36]
    .clock(KernelConvolution_2_clock),
    .reset(KernelConvolution_2_reset),
    .io_kernelVal_in(KernelConvolution_2_io_kernelVal_in),
    .io_pixelVal_in_0(KernelConvolution_2_io_pixelVal_in_0),
    .io_pixelVal_in_1(KernelConvolution_2_io_pixelVal_in_1),
    .io_pixelVal_in_2(KernelConvolution_2_io_pixelVal_in_2),
    .io_pixelVal_in_3(KernelConvolution_2_io_pixelVal_in_3),
    .io_pixelVal_in_4(KernelConvolution_2_io_pixelVal_in_4),
    .io_pixelVal_in_5(KernelConvolution_2_io_pixelVal_in_5),
    .io_pixelVal_in_6(KernelConvolution_2_io_pixelVal_in_6),
    .io_pixelVal_in_7(KernelConvolution_2_io_pixelVal_in_7),
    .io_pixelVal_out_0(KernelConvolution_2_io_pixelVal_out_0),
    .io_pixelVal_out_1(KernelConvolution_2_io_pixelVal_out_1),
    .io_pixelVal_out_2(KernelConvolution_2_io_pixelVal_out_2),
    .io_pixelVal_out_3(KernelConvolution_2_io_pixelVal_out_3),
    .io_pixelVal_out_4(KernelConvolution_2_io_pixelVal_out_4),
    .io_pixelVal_out_5(KernelConvolution_2_io_pixelVal_out_5),
    .io_pixelVal_out_6(KernelConvolution_2_io_pixelVal_out_6),
    .io_pixelVal_out_7(KernelConvolution_2_io_pixelVal_out_7),
    .io_valid_out(KernelConvolution_2_io_valid_out)
  );
  assign io_pixelVal_out_0_0 = _GEN_27877[3:0]; // @[Filter.scala 213:35 Filter.scala 215:37 Filter.scala 218:35 Filter.scala 220:35 Filter.scala 222:35 Filter.scala 224:35]
  assign io_pixelVal_out_0_1 = _GEN_27882[3:0]; // @[Filter.scala 213:35 Filter.scala 215:37 Filter.scala 218:35 Filter.scala 220:35 Filter.scala 222:35 Filter.scala 224:35]
  assign io_pixelVal_out_0_2 = _GEN_27887[3:0]; // @[Filter.scala 213:35 Filter.scala 215:37 Filter.scala 218:35 Filter.scala 220:35 Filter.scala 222:35 Filter.scala 224:35]
  assign io_pixelVal_out_0_3 = _GEN_27892[3:0]; // @[Filter.scala 213:35 Filter.scala 215:37 Filter.scala 218:35 Filter.scala 220:35 Filter.scala 222:35 Filter.scala 224:35]
  assign io_pixelVal_out_0_4 = _GEN_27897[3:0]; // @[Filter.scala 213:35 Filter.scala 215:37 Filter.scala 218:35 Filter.scala 220:35 Filter.scala 222:35 Filter.scala 224:35]
  assign io_pixelVal_out_0_5 = _GEN_27902[3:0]; // @[Filter.scala 213:35 Filter.scala 215:37 Filter.scala 218:35 Filter.scala 220:35 Filter.scala 222:35 Filter.scala 224:35]
  assign io_pixelVal_out_0_6 = _GEN_27907[3:0]; // @[Filter.scala 213:35 Filter.scala 215:37 Filter.scala 218:35 Filter.scala 220:35 Filter.scala 222:35 Filter.scala 224:35]
  assign io_pixelVal_out_0_7 = _GEN_27912[3:0]; // @[Filter.scala 213:35 Filter.scala 215:37 Filter.scala 218:35 Filter.scala 220:35 Filter.scala 222:35 Filter.scala 224:35]
  assign io_pixelVal_out_1_0 = _GEN_27917[3:0]; // @[Filter.scala 213:35 Filter.scala 215:37 Filter.scala 218:35 Filter.scala 220:35 Filter.scala 222:35 Filter.scala 224:35]
  assign io_pixelVal_out_1_1 = _GEN_27922[3:0]; // @[Filter.scala 213:35 Filter.scala 215:37 Filter.scala 218:35 Filter.scala 220:35 Filter.scala 222:35 Filter.scala 224:35]
  assign io_pixelVal_out_1_2 = _GEN_27927[3:0]; // @[Filter.scala 213:35 Filter.scala 215:37 Filter.scala 218:35 Filter.scala 220:35 Filter.scala 222:35 Filter.scala 224:35]
  assign io_pixelVal_out_1_3 = _GEN_27932[3:0]; // @[Filter.scala 213:35 Filter.scala 215:37 Filter.scala 218:35 Filter.scala 220:35 Filter.scala 222:35 Filter.scala 224:35]
  assign io_pixelVal_out_1_4 = _GEN_27937[3:0]; // @[Filter.scala 213:35 Filter.scala 215:37 Filter.scala 218:35 Filter.scala 220:35 Filter.scala 222:35 Filter.scala 224:35]
  assign io_pixelVal_out_1_5 = _GEN_27942[3:0]; // @[Filter.scala 213:35 Filter.scala 215:37 Filter.scala 218:35 Filter.scala 220:35 Filter.scala 222:35 Filter.scala 224:35]
  assign io_pixelVal_out_1_6 = _GEN_27947[3:0]; // @[Filter.scala 213:35 Filter.scala 215:37 Filter.scala 218:35 Filter.scala 220:35 Filter.scala 222:35 Filter.scala 224:35]
  assign io_pixelVal_out_1_7 = _GEN_27952[3:0]; // @[Filter.scala 213:35 Filter.scala 215:37 Filter.scala 218:35 Filter.scala 220:35 Filter.scala 222:35 Filter.scala 224:35]
  assign io_pixelVal_out_2_0 = _GEN_27957[3:0]; // @[Filter.scala 213:35 Filter.scala 215:37 Filter.scala 218:35 Filter.scala 220:35 Filter.scala 222:35 Filter.scala 224:35]
  assign io_pixelVal_out_2_1 = _GEN_27962[3:0]; // @[Filter.scala 213:35 Filter.scala 215:37 Filter.scala 218:35 Filter.scala 220:35 Filter.scala 222:35 Filter.scala 224:35]
  assign io_pixelVal_out_2_2 = _GEN_27967[3:0]; // @[Filter.scala 213:35 Filter.scala 215:37 Filter.scala 218:35 Filter.scala 220:35 Filter.scala 222:35 Filter.scala 224:35]
  assign io_pixelVal_out_2_3 = _GEN_27972[3:0]; // @[Filter.scala 213:35 Filter.scala 215:37 Filter.scala 218:35 Filter.scala 220:35 Filter.scala 222:35 Filter.scala 224:35]
  assign io_pixelVal_out_2_4 = _GEN_27977[3:0]; // @[Filter.scala 213:35 Filter.scala 215:37 Filter.scala 218:35 Filter.scala 220:35 Filter.scala 222:35 Filter.scala 224:35]
  assign io_pixelVal_out_2_5 = _GEN_27982[3:0]; // @[Filter.scala 213:35 Filter.scala 215:37 Filter.scala 218:35 Filter.scala 220:35 Filter.scala 222:35 Filter.scala 224:35]
  assign io_pixelVal_out_2_6 = _GEN_27987[3:0]; // @[Filter.scala 213:35 Filter.scala 215:37 Filter.scala 218:35 Filter.scala 220:35 Filter.scala 222:35 Filter.scala 224:35]
  assign io_pixelVal_out_2_7 = _GEN_27992[3:0]; // @[Filter.scala 213:35 Filter.scala 215:37 Filter.scala 218:35 Filter.scala 220:35 Filter.scala 222:35 Filter.scala 224:35]
  assign io_valid_out = validOut; // @[Filter.scala 231:18]
  assign KernelConvolution_clock = clock;
  assign KernelConvolution_reset = reset;
  assign KernelConvolution_io_kernelVal_in = _GEN_28077 & _GEN_28004 ? $signed(5'sh0) : $signed(_GEN_55); // @[Filter.scala 181:41]
  assign KernelConvolution_io_pixelVal_in_0 = _GEN_2476[3:0]; // @[Filter.scala 195:53 Filter.scala 197:51 Filter.scala 199:51]
  assign KernelConvolution_io_pixelVal_in_1 = _GEN_5938[3:0]; // @[Filter.scala 195:53 Filter.scala 197:51 Filter.scala 199:51]
  assign KernelConvolution_io_pixelVal_in_2 = _GEN_9400[3:0]; // @[Filter.scala 195:53 Filter.scala 197:51 Filter.scala 199:51]
  assign KernelConvolution_io_pixelVal_in_3 = _GEN_12862[3:0]; // @[Filter.scala 195:53 Filter.scala 197:51 Filter.scala 199:51]
  assign KernelConvolution_io_pixelVal_in_4 = _GEN_16324[3:0]; // @[Filter.scala 195:53 Filter.scala 197:51 Filter.scala 199:51]
  assign KernelConvolution_io_pixelVal_in_5 = _GEN_19786[3:0]; // @[Filter.scala 195:53 Filter.scala 197:51 Filter.scala 199:51]
  assign KernelConvolution_io_pixelVal_in_6 = _GEN_23248[3:0]; // @[Filter.scala 195:53 Filter.scala 197:51 Filter.scala 199:51]
  assign KernelConvolution_io_pixelVal_in_7 = _GEN_26710[3:0]; // @[Filter.scala 195:53 Filter.scala 197:51 Filter.scala 199:51]
  assign KernelConvolution_1_clock = clock;
  assign KernelConvolution_1_reset = reset;
  assign KernelConvolution_1_io_kernelVal_in = _GEN_28077 & _GEN_28004 ? $signed(5'sh0) : $signed(_GEN_55); // @[Filter.scala 181:41]
  assign KernelConvolution_1_io_pixelVal_in_0 = _GEN_3054[3:0]; // @[Filter.scala 195:53 Filter.scala 197:51 Filter.scala 199:51]
  assign KernelConvolution_1_io_pixelVal_in_1 = _GEN_6516[3:0]; // @[Filter.scala 195:53 Filter.scala 197:51 Filter.scala 199:51]
  assign KernelConvolution_1_io_pixelVal_in_2 = _GEN_9978[3:0]; // @[Filter.scala 195:53 Filter.scala 197:51 Filter.scala 199:51]
  assign KernelConvolution_1_io_pixelVal_in_3 = _GEN_13440[3:0]; // @[Filter.scala 195:53 Filter.scala 197:51 Filter.scala 199:51]
  assign KernelConvolution_1_io_pixelVal_in_4 = _GEN_16902[3:0]; // @[Filter.scala 195:53 Filter.scala 197:51 Filter.scala 199:51]
  assign KernelConvolution_1_io_pixelVal_in_5 = _GEN_20364[3:0]; // @[Filter.scala 195:53 Filter.scala 197:51 Filter.scala 199:51]
  assign KernelConvolution_1_io_pixelVal_in_6 = _GEN_23826[3:0]; // @[Filter.scala 195:53 Filter.scala 197:51 Filter.scala 199:51]
  assign KernelConvolution_1_io_pixelVal_in_7 = _GEN_27288[3:0]; // @[Filter.scala 195:53 Filter.scala 197:51 Filter.scala 199:51]
  assign KernelConvolution_2_clock = clock;
  assign KernelConvolution_2_reset = reset;
  assign KernelConvolution_2_io_kernelVal_in = _GEN_28077 & _GEN_28004 ? $signed(5'sh0) : $signed(_GEN_55); // @[Filter.scala 181:41]
  assign KernelConvolution_2_io_pixelVal_in_0 = _GEN_3632[3:0]; // @[Filter.scala 195:53 Filter.scala 197:51 Filter.scala 199:51]
  assign KernelConvolution_2_io_pixelVal_in_1 = _GEN_7094[3:0]; // @[Filter.scala 195:53 Filter.scala 197:51 Filter.scala 199:51]
  assign KernelConvolution_2_io_pixelVal_in_2 = _GEN_10556[3:0]; // @[Filter.scala 195:53 Filter.scala 197:51 Filter.scala 199:51]
  assign KernelConvolution_2_io_pixelVal_in_3 = _GEN_14018[3:0]; // @[Filter.scala 195:53 Filter.scala 197:51 Filter.scala 199:51]
  assign KernelConvolution_2_io_pixelVal_in_4 = _GEN_17480[3:0]; // @[Filter.scala 195:53 Filter.scala 197:51 Filter.scala 199:51]
  assign KernelConvolution_2_io_pixelVal_in_5 = _GEN_20942[3:0]; // @[Filter.scala 195:53 Filter.scala 197:51 Filter.scala 199:51]
  assign KernelConvolution_2_io_pixelVal_in_6 = _GEN_24404[3:0]; // @[Filter.scala 195:53 Filter.scala 197:51 Filter.scala 199:51]
  assign KernelConvolution_2_io_pixelVal_in_7 = _GEN_27866[3:0]; // @[Filter.scala 195:53 Filter.scala 197:51 Filter.scala 199:51]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  kernelCounter = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  imageCounterX = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  imageCounterY = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  pixelIndex = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  pixOut_0_0 = _RAND_4[8:0];
  _RAND_5 = {1{`RANDOM}};
  pixOut_0_1 = _RAND_5[8:0];
  _RAND_6 = {1{`RANDOM}};
  pixOut_0_2 = _RAND_6[8:0];
  _RAND_7 = {1{`RANDOM}};
  pixOut_0_3 = _RAND_7[8:0];
  _RAND_8 = {1{`RANDOM}};
  pixOut_0_4 = _RAND_8[8:0];
  _RAND_9 = {1{`RANDOM}};
  pixOut_0_5 = _RAND_9[8:0];
  _RAND_10 = {1{`RANDOM}};
  pixOut_0_6 = _RAND_10[8:0];
  _RAND_11 = {1{`RANDOM}};
  pixOut_0_7 = _RAND_11[8:0];
  _RAND_12 = {1{`RANDOM}};
  pixOut_1_0 = _RAND_12[8:0];
  _RAND_13 = {1{`RANDOM}};
  pixOut_1_1 = _RAND_13[8:0];
  _RAND_14 = {1{`RANDOM}};
  pixOut_1_2 = _RAND_14[8:0];
  _RAND_15 = {1{`RANDOM}};
  pixOut_1_3 = _RAND_15[8:0];
  _RAND_16 = {1{`RANDOM}};
  pixOut_1_4 = _RAND_16[8:0];
  _RAND_17 = {1{`RANDOM}};
  pixOut_1_5 = _RAND_17[8:0];
  _RAND_18 = {1{`RANDOM}};
  pixOut_1_6 = _RAND_18[8:0];
  _RAND_19 = {1{`RANDOM}};
  pixOut_1_7 = _RAND_19[8:0];
  _RAND_20 = {1{`RANDOM}};
  pixOut_2_0 = _RAND_20[8:0];
  _RAND_21 = {1{`RANDOM}};
  pixOut_2_1 = _RAND_21[8:0];
  _RAND_22 = {1{`RANDOM}};
  pixOut_2_2 = _RAND_22[8:0];
  _RAND_23 = {1{`RANDOM}};
  pixOut_2_3 = _RAND_23[8:0];
  _RAND_24 = {1{`RANDOM}};
  pixOut_2_4 = _RAND_24[8:0];
  _RAND_25 = {1{`RANDOM}};
  pixOut_2_5 = _RAND_25[8:0];
  _RAND_26 = {1{`RANDOM}};
  pixOut_2_6 = _RAND_26[8:0];
  _RAND_27 = {1{`RANDOM}};
  pixOut_2_7 = _RAND_27[8:0];
  _RAND_28 = {1{`RANDOM}};
  validOut = _RAND_28[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      kernelCounter <= 4'h0;
    end else if (kernelCountReset) begin
      kernelCounter <= 4'h0;
    end else begin
      kernelCounter <= _T_17;
    end
    if (reset) begin
      imageCounterX <= 2'h0;
    end else if (imageCounterXReset) begin
      imageCounterX <= 2'h0;
    end else begin
      imageCounterX <= _T_23;
    end
    if (reset) begin
      imageCounterY <= 2'h0;
    end else if (imageCounterXReset) begin
      if (_T_24) begin
        imageCounterY <= 2'h0;
      end else begin
        imageCounterY <= _T_26;
      end
    end
    if (reset) begin
      pixelIndex <= 32'h0;
    end else if (kernelCountReset) begin
      if (_T_834) begin
        pixelIndex <= 32'h0;
      end else begin
        pixelIndex <= _T_832;
      end
    end
    if (reset) begin
      pixOut_0_0 <= 9'sh0;
    end else begin
      pixOut_0_0 <= _T_567[8:0];
    end
    if (reset) begin
      pixOut_0_1 <= 9'sh0;
    end else begin
      pixOut_0_1 <= _T_578[8:0];
    end
    if (reset) begin
      pixOut_0_2 <= 9'sh0;
    end else begin
      pixOut_0_2 <= _T_589[8:0];
    end
    if (reset) begin
      pixOut_0_3 <= 9'sh0;
    end else begin
      pixOut_0_3 <= _T_600[8:0];
    end
    if (reset) begin
      pixOut_0_4 <= 9'sh0;
    end else begin
      pixOut_0_4 <= _T_611[8:0];
    end
    if (reset) begin
      pixOut_0_5 <= 9'sh0;
    end else begin
      pixOut_0_5 <= _T_622[8:0];
    end
    if (reset) begin
      pixOut_0_6 <= 9'sh0;
    end else begin
      pixOut_0_6 <= _T_633[8:0];
    end
    if (reset) begin
      pixOut_0_7 <= 9'sh0;
    end else begin
      pixOut_0_7 <= _T_644[8:0];
    end
    if (reset) begin
      pixOut_1_0 <= 9'sh0;
    end else begin
      pixOut_1_0 <= _T_655[8:0];
    end
    if (reset) begin
      pixOut_1_1 <= 9'sh0;
    end else begin
      pixOut_1_1 <= _T_666[8:0];
    end
    if (reset) begin
      pixOut_1_2 <= 9'sh0;
    end else begin
      pixOut_1_2 <= _T_677[8:0];
    end
    if (reset) begin
      pixOut_1_3 <= 9'sh0;
    end else begin
      pixOut_1_3 <= _T_688[8:0];
    end
    if (reset) begin
      pixOut_1_4 <= 9'sh0;
    end else begin
      pixOut_1_4 <= _T_699[8:0];
    end
    if (reset) begin
      pixOut_1_5 <= 9'sh0;
    end else begin
      pixOut_1_5 <= _T_710[8:0];
    end
    if (reset) begin
      pixOut_1_6 <= 9'sh0;
    end else begin
      pixOut_1_6 <= _T_721[8:0];
    end
    if (reset) begin
      pixOut_1_7 <= 9'sh0;
    end else begin
      pixOut_1_7 <= _T_732[8:0];
    end
    if (reset) begin
      pixOut_2_0 <= 9'sh0;
    end else begin
      pixOut_2_0 <= _T_743[8:0];
    end
    if (reset) begin
      pixOut_2_1 <= 9'sh0;
    end else begin
      pixOut_2_1 <= _T_754[8:0];
    end
    if (reset) begin
      pixOut_2_2 <= 9'sh0;
    end else begin
      pixOut_2_2 <= _T_765[8:0];
    end
    if (reset) begin
      pixOut_2_3 <= 9'sh0;
    end else begin
      pixOut_2_3 <= _T_776[8:0];
    end
    if (reset) begin
      pixOut_2_4 <= 9'sh0;
    end else begin
      pixOut_2_4 <= _T_787[8:0];
    end
    if (reset) begin
      pixOut_2_5 <= 9'sh0;
    end else begin
      pixOut_2_5 <= _T_798[8:0];
    end
    if (reset) begin
      pixOut_2_6 <= 9'sh0;
    end else begin
      pixOut_2_6 <= _T_809[8:0];
    end
    if (reset) begin
      pixOut_2_7 <= 9'sh0;
    end else begin
      pixOut_2_7 <= _T_820[8:0];
    end
    if (reset) begin
      validOut <= 1'h0;
    end else begin
      validOut <= KernelConvolution_io_valid_out;
    end
  end
endmodule
module VideoBuffer(
  input         clock,
  input         reset,
  input  [3:0]  io_pixelVal_in_0_0,
  input  [3:0]  io_pixelVal_in_0_1,
  input  [3:0]  io_pixelVal_in_0_2,
  input  [3:0]  io_pixelVal_in_0_3,
  input  [3:0]  io_pixelVal_in_0_4,
  input  [3:0]  io_pixelVal_in_0_5,
  input  [3:0]  io_pixelVal_in_0_6,
  input  [3:0]  io_pixelVal_in_0_7,
  input  [3:0]  io_pixelVal_in_1_0,
  input  [3:0]  io_pixelVal_in_1_1,
  input  [3:0]  io_pixelVal_in_1_2,
  input  [3:0]  io_pixelVal_in_1_3,
  input  [3:0]  io_pixelVal_in_1_4,
  input  [3:0]  io_pixelVal_in_1_5,
  input  [3:0]  io_pixelVal_in_1_6,
  input  [3:0]  io_pixelVal_in_1_7,
  input  [3:0]  io_pixelVal_in_2_0,
  input  [3:0]  io_pixelVal_in_2_1,
  input  [3:0]  io_pixelVal_in_2_2,
  input  [3:0]  io_pixelVal_in_2_3,
  input  [3:0]  io_pixelVal_in_2_4,
  input  [3:0]  io_pixelVal_in_2_5,
  input  [3:0]  io_pixelVal_in_2_6,
  input  [3:0]  io_pixelVal_in_2_7,
  input         io_valid_in,
  input  [10:0] io_rowIndex,
  input  [10:0] io_colIndex,
  output [3:0]  io_pixelVal_out_0,
  output [3:0]  io_pixelVal_out_1,
  output [3:0]  io_pixelVal_out_2
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1041;
  reg [31:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1045;
  reg [31:0] _RAND_1046;
  reg [31:0] _RAND_1047;
  reg [31:0] _RAND_1048;
  reg [31:0] _RAND_1049;
  reg [31:0] _RAND_1050;
  reg [31:0] _RAND_1051;
  reg [31:0] _RAND_1052;
  reg [31:0] _RAND_1053;
  reg [31:0] _RAND_1054;
  reg [31:0] _RAND_1055;
  reg [31:0] _RAND_1056;
  reg [31:0] _RAND_1057;
  reg [31:0] _RAND_1058;
  reg [31:0] _RAND_1059;
  reg [31:0] _RAND_1060;
  reg [31:0] _RAND_1061;
  reg [31:0] _RAND_1062;
  reg [31:0] _RAND_1063;
  reg [31:0] _RAND_1064;
  reg [31:0] _RAND_1065;
  reg [31:0] _RAND_1066;
  reg [31:0] _RAND_1067;
  reg [31:0] _RAND_1068;
  reg [31:0] _RAND_1069;
  reg [31:0] _RAND_1070;
  reg [31:0] _RAND_1071;
  reg [31:0] _RAND_1072;
  reg [31:0] _RAND_1073;
  reg [31:0] _RAND_1074;
  reg [31:0] _RAND_1075;
  reg [31:0] _RAND_1076;
  reg [31:0] _RAND_1077;
  reg [31:0] _RAND_1078;
  reg [31:0] _RAND_1079;
  reg [31:0] _RAND_1080;
  reg [31:0] _RAND_1081;
  reg [31:0] _RAND_1082;
  reg [31:0] _RAND_1083;
  reg [31:0] _RAND_1084;
  reg [31:0] _RAND_1085;
  reg [31:0] _RAND_1086;
  reg [31:0] _RAND_1087;
  reg [31:0] _RAND_1088;
  reg [31:0] _RAND_1089;
  reg [31:0] _RAND_1090;
  reg [31:0] _RAND_1091;
  reg [31:0] _RAND_1092;
  reg [31:0] _RAND_1093;
  reg [31:0] _RAND_1094;
  reg [31:0] _RAND_1095;
  reg [31:0] _RAND_1096;
  reg [31:0] _RAND_1097;
  reg [31:0] _RAND_1098;
  reg [31:0] _RAND_1099;
  reg [31:0] _RAND_1100;
  reg [31:0] _RAND_1101;
  reg [31:0] _RAND_1102;
  reg [31:0] _RAND_1103;
  reg [31:0] _RAND_1104;
  reg [31:0] _RAND_1105;
  reg [31:0] _RAND_1106;
  reg [31:0] _RAND_1107;
  reg [31:0] _RAND_1108;
  reg [31:0] _RAND_1109;
  reg [31:0] _RAND_1110;
  reg [31:0] _RAND_1111;
  reg [31:0] _RAND_1112;
  reg [31:0] _RAND_1113;
  reg [31:0] _RAND_1114;
  reg [31:0] _RAND_1115;
  reg [31:0] _RAND_1116;
  reg [31:0] _RAND_1117;
  reg [31:0] _RAND_1118;
  reg [31:0] _RAND_1119;
  reg [31:0] _RAND_1120;
  reg [31:0] _RAND_1121;
  reg [31:0] _RAND_1122;
  reg [31:0] _RAND_1123;
  reg [31:0] _RAND_1124;
  reg [31:0] _RAND_1125;
  reg [31:0] _RAND_1126;
  reg [31:0] _RAND_1127;
  reg [31:0] _RAND_1128;
  reg [31:0] _RAND_1129;
  reg [31:0] _RAND_1130;
  reg [31:0] _RAND_1131;
  reg [31:0] _RAND_1132;
  reg [31:0] _RAND_1133;
  reg [31:0] _RAND_1134;
  reg [31:0] _RAND_1135;
  reg [31:0] _RAND_1136;
  reg [31:0] _RAND_1137;
  reg [31:0] _RAND_1138;
  reg [31:0] _RAND_1139;
  reg [31:0] _RAND_1140;
  reg [31:0] _RAND_1141;
  reg [31:0] _RAND_1142;
  reg [31:0] _RAND_1143;
  reg [31:0] _RAND_1144;
  reg [31:0] _RAND_1145;
  reg [31:0] _RAND_1146;
  reg [31:0] _RAND_1147;
  reg [31:0] _RAND_1148;
  reg [31:0] _RAND_1149;
  reg [31:0] _RAND_1150;
  reg [31:0] _RAND_1151;
  reg [31:0] _RAND_1152;
  reg [31:0] _RAND_1153;
  reg [31:0] _RAND_1154;
  reg [31:0] _RAND_1155;
  reg [31:0] _RAND_1156;
  reg [31:0] _RAND_1157;
  reg [31:0] _RAND_1158;
  reg [31:0] _RAND_1159;
  reg [31:0] _RAND_1160;
  reg [31:0] _RAND_1161;
  reg [31:0] _RAND_1162;
  reg [31:0] _RAND_1163;
  reg [31:0] _RAND_1164;
  reg [31:0] _RAND_1165;
  reg [31:0] _RAND_1166;
  reg [31:0] _RAND_1167;
  reg [31:0] _RAND_1168;
  reg [31:0] _RAND_1169;
  reg [31:0] _RAND_1170;
  reg [31:0] _RAND_1171;
  reg [31:0] _RAND_1172;
  reg [31:0] _RAND_1173;
  reg [31:0] _RAND_1174;
  reg [31:0] _RAND_1175;
  reg [31:0] _RAND_1176;
  reg [31:0] _RAND_1177;
  reg [31:0] _RAND_1178;
  reg [31:0] _RAND_1179;
  reg [31:0] _RAND_1180;
  reg [31:0] _RAND_1181;
  reg [31:0] _RAND_1182;
  reg [31:0] _RAND_1183;
  reg [31:0] _RAND_1184;
  reg [31:0] _RAND_1185;
  reg [31:0] _RAND_1186;
  reg [31:0] _RAND_1187;
  reg [31:0] _RAND_1188;
  reg [31:0] _RAND_1189;
  reg [31:0] _RAND_1190;
  reg [31:0] _RAND_1191;
  reg [31:0] _RAND_1192;
  reg [31:0] _RAND_1193;
  reg [31:0] _RAND_1194;
  reg [31:0] _RAND_1195;
  reg [31:0] _RAND_1196;
  reg [31:0] _RAND_1197;
  reg [31:0] _RAND_1198;
  reg [31:0] _RAND_1199;
  reg [31:0] _RAND_1200;
  reg [31:0] _RAND_1201;
  reg [31:0] _RAND_1202;
  reg [31:0] _RAND_1203;
  reg [31:0] _RAND_1204;
  reg [31:0] _RAND_1205;
  reg [31:0] _RAND_1206;
  reg [31:0] _RAND_1207;
  reg [31:0] _RAND_1208;
  reg [31:0] _RAND_1209;
  reg [31:0] _RAND_1210;
  reg [31:0] _RAND_1211;
  reg [31:0] _RAND_1212;
  reg [31:0] _RAND_1213;
  reg [31:0] _RAND_1214;
  reg [31:0] _RAND_1215;
  reg [31:0] _RAND_1216;
  reg [31:0] _RAND_1217;
  reg [31:0] _RAND_1218;
  reg [31:0] _RAND_1219;
  reg [31:0] _RAND_1220;
  reg [31:0] _RAND_1221;
  reg [31:0] _RAND_1222;
  reg [31:0] _RAND_1223;
  reg [31:0] _RAND_1224;
  reg [31:0] _RAND_1225;
  reg [31:0] _RAND_1226;
  reg [31:0] _RAND_1227;
  reg [31:0] _RAND_1228;
  reg [31:0] _RAND_1229;
  reg [31:0] _RAND_1230;
  reg [31:0] _RAND_1231;
  reg [31:0] _RAND_1232;
  reg [31:0] _RAND_1233;
  reg [31:0] _RAND_1234;
  reg [31:0] _RAND_1235;
  reg [31:0] _RAND_1236;
  reg [31:0] _RAND_1237;
  reg [31:0] _RAND_1238;
  reg [31:0] _RAND_1239;
  reg [31:0] _RAND_1240;
  reg [31:0] _RAND_1241;
  reg [31:0] _RAND_1242;
  reg [31:0] _RAND_1243;
  reg [31:0] _RAND_1244;
  reg [31:0] _RAND_1245;
  reg [31:0] _RAND_1246;
  reg [31:0] _RAND_1247;
  reg [31:0] _RAND_1248;
  reg [31:0] _RAND_1249;
  reg [31:0] _RAND_1250;
  reg [31:0] _RAND_1251;
  reg [31:0] _RAND_1252;
  reg [31:0] _RAND_1253;
  reg [31:0] _RAND_1254;
  reg [31:0] _RAND_1255;
  reg [31:0] _RAND_1256;
  reg [31:0] _RAND_1257;
  reg [31:0] _RAND_1258;
  reg [31:0] _RAND_1259;
  reg [31:0] _RAND_1260;
  reg [31:0] _RAND_1261;
  reg [31:0] _RAND_1262;
  reg [31:0] _RAND_1263;
  reg [31:0] _RAND_1264;
  reg [31:0] _RAND_1265;
  reg [31:0] _RAND_1266;
  reg [31:0] _RAND_1267;
  reg [31:0] _RAND_1268;
  reg [31:0] _RAND_1269;
  reg [31:0] _RAND_1270;
  reg [31:0] _RAND_1271;
  reg [31:0] _RAND_1272;
  reg [31:0] _RAND_1273;
  reg [31:0] _RAND_1274;
  reg [31:0] _RAND_1275;
  reg [31:0] _RAND_1276;
  reg [31:0] _RAND_1277;
  reg [31:0] _RAND_1278;
  reg [31:0] _RAND_1279;
  reg [31:0] _RAND_1280;
  reg [31:0] _RAND_1281;
  reg [31:0] _RAND_1282;
  reg [31:0] _RAND_1283;
  reg [31:0] _RAND_1284;
  reg [31:0] _RAND_1285;
  reg [31:0] _RAND_1286;
  reg [31:0] _RAND_1287;
  reg [31:0] _RAND_1288;
  reg [31:0] _RAND_1289;
  reg [31:0] _RAND_1290;
  reg [31:0] _RAND_1291;
  reg [31:0] _RAND_1292;
  reg [31:0] _RAND_1293;
  reg [31:0] _RAND_1294;
  reg [31:0] _RAND_1295;
  reg [31:0] _RAND_1296;
  reg [31:0] _RAND_1297;
  reg [31:0] _RAND_1298;
  reg [31:0] _RAND_1299;
  reg [31:0] _RAND_1300;
  reg [31:0] _RAND_1301;
  reg [31:0] _RAND_1302;
  reg [31:0] _RAND_1303;
  reg [31:0] _RAND_1304;
  reg [31:0] _RAND_1305;
  reg [31:0] _RAND_1306;
  reg [31:0] _RAND_1307;
  reg [31:0] _RAND_1308;
  reg [31:0] _RAND_1309;
  reg [31:0] _RAND_1310;
  reg [31:0] _RAND_1311;
  reg [31:0] _RAND_1312;
  reg [31:0] _RAND_1313;
  reg [31:0] _RAND_1314;
  reg [31:0] _RAND_1315;
  reg [31:0] _RAND_1316;
  reg [31:0] _RAND_1317;
  reg [31:0] _RAND_1318;
  reg [31:0] _RAND_1319;
  reg [31:0] _RAND_1320;
  reg [31:0] _RAND_1321;
  reg [31:0] _RAND_1322;
  reg [31:0] _RAND_1323;
  reg [31:0] _RAND_1324;
  reg [31:0] _RAND_1325;
  reg [31:0] _RAND_1326;
  reg [31:0] _RAND_1327;
  reg [31:0] _RAND_1328;
  reg [31:0] _RAND_1329;
  reg [31:0] _RAND_1330;
  reg [31:0] _RAND_1331;
  reg [31:0] _RAND_1332;
  reg [31:0] _RAND_1333;
  reg [31:0] _RAND_1334;
  reg [31:0] _RAND_1335;
  reg [31:0] _RAND_1336;
  reg [31:0] _RAND_1337;
  reg [31:0] _RAND_1338;
  reg [31:0] _RAND_1339;
  reg [31:0] _RAND_1340;
  reg [31:0] _RAND_1341;
  reg [31:0] _RAND_1342;
  reg [31:0] _RAND_1343;
  reg [31:0] _RAND_1344;
  reg [31:0] _RAND_1345;
  reg [31:0] _RAND_1346;
  reg [31:0] _RAND_1347;
  reg [31:0] _RAND_1348;
  reg [31:0] _RAND_1349;
  reg [31:0] _RAND_1350;
  reg [31:0] _RAND_1351;
  reg [31:0] _RAND_1352;
  reg [31:0] _RAND_1353;
  reg [31:0] _RAND_1354;
  reg [31:0] _RAND_1355;
  reg [31:0] _RAND_1356;
  reg [31:0] _RAND_1357;
  reg [31:0] _RAND_1358;
  reg [31:0] _RAND_1359;
  reg [31:0] _RAND_1360;
  reg [31:0] _RAND_1361;
  reg [31:0] _RAND_1362;
  reg [31:0] _RAND_1363;
  reg [31:0] _RAND_1364;
  reg [31:0] _RAND_1365;
  reg [31:0] _RAND_1366;
  reg [31:0] _RAND_1367;
  reg [31:0] _RAND_1368;
  reg [31:0] _RAND_1369;
  reg [31:0] _RAND_1370;
  reg [31:0] _RAND_1371;
  reg [31:0] _RAND_1372;
  reg [31:0] _RAND_1373;
  reg [31:0] _RAND_1374;
  reg [31:0] _RAND_1375;
  reg [31:0] _RAND_1376;
  reg [31:0] _RAND_1377;
  reg [31:0] _RAND_1378;
  reg [31:0] _RAND_1379;
  reg [31:0] _RAND_1380;
  reg [31:0] _RAND_1381;
  reg [31:0] _RAND_1382;
  reg [31:0] _RAND_1383;
  reg [31:0] _RAND_1384;
  reg [31:0] _RAND_1385;
  reg [31:0] _RAND_1386;
  reg [31:0] _RAND_1387;
  reg [31:0] _RAND_1388;
  reg [31:0] _RAND_1389;
  reg [31:0] _RAND_1390;
  reg [31:0] _RAND_1391;
  reg [31:0] _RAND_1392;
  reg [31:0] _RAND_1393;
  reg [31:0] _RAND_1394;
  reg [31:0] _RAND_1395;
  reg [31:0] _RAND_1396;
  reg [31:0] _RAND_1397;
  reg [31:0] _RAND_1398;
  reg [31:0] _RAND_1399;
  reg [31:0] _RAND_1400;
  reg [31:0] _RAND_1401;
  reg [31:0] _RAND_1402;
  reg [31:0] _RAND_1403;
  reg [31:0] _RAND_1404;
  reg [31:0] _RAND_1405;
  reg [31:0] _RAND_1406;
  reg [31:0] _RAND_1407;
  reg [31:0] _RAND_1408;
  reg [31:0] _RAND_1409;
  reg [31:0] _RAND_1410;
  reg [31:0] _RAND_1411;
  reg [31:0] _RAND_1412;
  reg [31:0] _RAND_1413;
  reg [31:0] _RAND_1414;
  reg [31:0] _RAND_1415;
  reg [31:0] _RAND_1416;
  reg [31:0] _RAND_1417;
  reg [31:0] _RAND_1418;
  reg [31:0] _RAND_1419;
  reg [31:0] _RAND_1420;
  reg [31:0] _RAND_1421;
  reg [31:0] _RAND_1422;
  reg [31:0] _RAND_1423;
  reg [31:0] _RAND_1424;
  reg [31:0] _RAND_1425;
  reg [31:0] _RAND_1426;
  reg [31:0] _RAND_1427;
  reg [31:0] _RAND_1428;
  reg [31:0] _RAND_1429;
  reg [31:0] _RAND_1430;
  reg [31:0] _RAND_1431;
  reg [31:0] _RAND_1432;
  reg [31:0] _RAND_1433;
  reg [31:0] _RAND_1434;
  reg [31:0] _RAND_1435;
  reg [31:0] _RAND_1436;
  reg [31:0] _RAND_1437;
  reg [31:0] _RAND_1438;
  reg [31:0] _RAND_1439;
  reg [31:0] _RAND_1440;
  reg [31:0] _RAND_1441;
  reg [31:0] _RAND_1442;
  reg [31:0] _RAND_1443;
  reg [31:0] _RAND_1444;
  reg [31:0] _RAND_1445;
  reg [31:0] _RAND_1446;
  reg [31:0] _RAND_1447;
  reg [31:0] _RAND_1448;
  reg [31:0] _RAND_1449;
  reg [31:0] _RAND_1450;
  reg [31:0] _RAND_1451;
  reg [31:0] _RAND_1452;
  reg [31:0] _RAND_1453;
  reg [31:0] _RAND_1454;
  reg [31:0] _RAND_1455;
  reg [31:0] _RAND_1456;
  reg [31:0] _RAND_1457;
  reg [31:0] _RAND_1458;
  reg [31:0] _RAND_1459;
  reg [31:0] _RAND_1460;
  reg [31:0] _RAND_1461;
  reg [31:0] _RAND_1462;
  reg [31:0] _RAND_1463;
  reg [31:0] _RAND_1464;
  reg [31:0] _RAND_1465;
  reg [31:0] _RAND_1466;
  reg [31:0] _RAND_1467;
  reg [31:0] _RAND_1468;
  reg [31:0] _RAND_1469;
  reg [31:0] _RAND_1470;
  reg [31:0] _RAND_1471;
  reg [31:0] _RAND_1472;
  reg [31:0] _RAND_1473;
  reg [31:0] _RAND_1474;
  reg [31:0] _RAND_1475;
  reg [31:0] _RAND_1476;
  reg [31:0] _RAND_1477;
  reg [31:0] _RAND_1478;
  reg [31:0] _RAND_1479;
  reg [31:0] _RAND_1480;
  reg [31:0] _RAND_1481;
  reg [31:0] _RAND_1482;
  reg [31:0] _RAND_1483;
  reg [31:0] _RAND_1484;
  reg [31:0] _RAND_1485;
  reg [31:0] _RAND_1486;
  reg [31:0] _RAND_1487;
  reg [31:0] _RAND_1488;
  reg [31:0] _RAND_1489;
  reg [31:0] _RAND_1490;
  reg [31:0] _RAND_1491;
  reg [31:0] _RAND_1492;
  reg [31:0] _RAND_1493;
  reg [31:0] _RAND_1494;
  reg [31:0] _RAND_1495;
  reg [31:0] _RAND_1496;
  reg [31:0] _RAND_1497;
  reg [31:0] _RAND_1498;
  reg [31:0] _RAND_1499;
  reg [31:0] _RAND_1500;
  reg [31:0] _RAND_1501;
  reg [31:0] _RAND_1502;
  reg [31:0] _RAND_1503;
  reg [31:0] _RAND_1504;
  reg [31:0] _RAND_1505;
  reg [31:0] _RAND_1506;
  reg [31:0] _RAND_1507;
  reg [31:0] _RAND_1508;
  reg [31:0] _RAND_1509;
  reg [31:0] _RAND_1510;
  reg [31:0] _RAND_1511;
  reg [31:0] _RAND_1512;
  reg [31:0] _RAND_1513;
  reg [31:0] _RAND_1514;
  reg [31:0] _RAND_1515;
  reg [31:0] _RAND_1516;
  reg [31:0] _RAND_1517;
  reg [31:0] _RAND_1518;
  reg [31:0] _RAND_1519;
  reg [31:0] _RAND_1520;
  reg [31:0] _RAND_1521;
  reg [31:0] _RAND_1522;
  reg [31:0] _RAND_1523;
  reg [31:0] _RAND_1524;
  reg [31:0] _RAND_1525;
  reg [31:0] _RAND_1526;
  reg [31:0] _RAND_1527;
  reg [31:0] _RAND_1528;
  reg [31:0] _RAND_1529;
  reg [31:0] _RAND_1530;
  reg [31:0] _RAND_1531;
  reg [31:0] _RAND_1532;
  reg [31:0] _RAND_1533;
  reg [31:0] _RAND_1534;
  reg [31:0] _RAND_1535;
  reg [31:0] _RAND_1536;
  reg [31:0] _RAND_1537;
  reg [31:0] _RAND_1538;
  reg [31:0] _RAND_1539;
  reg [31:0] _RAND_1540;
  reg [31:0] _RAND_1541;
  reg [31:0] _RAND_1542;
  reg [31:0] _RAND_1543;
  reg [31:0] _RAND_1544;
  reg [31:0] _RAND_1545;
  reg [31:0] _RAND_1546;
  reg [31:0] _RAND_1547;
  reg [31:0] _RAND_1548;
  reg [31:0] _RAND_1549;
  reg [31:0] _RAND_1550;
  reg [31:0] _RAND_1551;
  reg [31:0] _RAND_1552;
  reg [31:0] _RAND_1553;
  reg [31:0] _RAND_1554;
  reg [31:0] _RAND_1555;
  reg [31:0] _RAND_1556;
  reg [31:0] _RAND_1557;
  reg [31:0] _RAND_1558;
  reg [31:0] _RAND_1559;
  reg [31:0] _RAND_1560;
  reg [31:0] _RAND_1561;
  reg [31:0] _RAND_1562;
  reg [31:0] _RAND_1563;
  reg [31:0] _RAND_1564;
  reg [31:0] _RAND_1565;
  reg [31:0] _RAND_1566;
  reg [31:0] _RAND_1567;
  reg [31:0] _RAND_1568;
  reg [31:0] _RAND_1569;
  reg [31:0] _RAND_1570;
  reg [31:0] _RAND_1571;
  reg [31:0] _RAND_1572;
  reg [31:0] _RAND_1573;
  reg [31:0] _RAND_1574;
  reg [31:0] _RAND_1575;
  reg [31:0] _RAND_1576;
  reg [31:0] _RAND_1577;
  reg [31:0] _RAND_1578;
  reg [31:0] _RAND_1579;
  reg [31:0] _RAND_1580;
  reg [31:0] _RAND_1581;
  reg [31:0] _RAND_1582;
  reg [31:0] _RAND_1583;
  reg [31:0] _RAND_1584;
  reg [31:0] _RAND_1585;
  reg [31:0] _RAND_1586;
  reg [31:0] _RAND_1587;
  reg [31:0] _RAND_1588;
  reg [31:0] _RAND_1589;
  reg [31:0] _RAND_1590;
  reg [31:0] _RAND_1591;
  reg [31:0] _RAND_1592;
  reg [31:0] _RAND_1593;
  reg [31:0] _RAND_1594;
  reg [31:0] _RAND_1595;
  reg [31:0] _RAND_1596;
  reg [31:0] _RAND_1597;
  reg [31:0] _RAND_1598;
  reg [31:0] _RAND_1599;
  reg [31:0] _RAND_1600;
  reg [31:0] _RAND_1601;
  reg [31:0] _RAND_1602;
  reg [31:0] _RAND_1603;
  reg [31:0] _RAND_1604;
  reg [31:0] _RAND_1605;
  reg [31:0] _RAND_1606;
  reg [31:0] _RAND_1607;
  reg [31:0] _RAND_1608;
  reg [31:0] _RAND_1609;
  reg [31:0] _RAND_1610;
  reg [31:0] _RAND_1611;
  reg [31:0] _RAND_1612;
  reg [31:0] _RAND_1613;
  reg [31:0] _RAND_1614;
  reg [31:0] _RAND_1615;
  reg [31:0] _RAND_1616;
  reg [31:0] _RAND_1617;
  reg [31:0] _RAND_1618;
  reg [31:0] _RAND_1619;
  reg [31:0] _RAND_1620;
  reg [31:0] _RAND_1621;
  reg [31:0] _RAND_1622;
  reg [31:0] _RAND_1623;
  reg [31:0] _RAND_1624;
  reg [31:0] _RAND_1625;
  reg [31:0] _RAND_1626;
  reg [31:0] _RAND_1627;
  reg [31:0] _RAND_1628;
  reg [31:0] _RAND_1629;
  reg [31:0] _RAND_1630;
  reg [31:0] _RAND_1631;
  reg [31:0] _RAND_1632;
  reg [31:0] _RAND_1633;
  reg [31:0] _RAND_1634;
  reg [31:0] _RAND_1635;
  reg [31:0] _RAND_1636;
  reg [31:0] _RAND_1637;
  reg [31:0] _RAND_1638;
  reg [31:0] _RAND_1639;
  reg [31:0] _RAND_1640;
  reg [31:0] _RAND_1641;
  reg [31:0] _RAND_1642;
  reg [31:0] _RAND_1643;
  reg [31:0] _RAND_1644;
  reg [31:0] _RAND_1645;
  reg [31:0] _RAND_1646;
  reg [31:0] _RAND_1647;
  reg [31:0] _RAND_1648;
  reg [31:0] _RAND_1649;
  reg [31:0] _RAND_1650;
  reg [31:0] _RAND_1651;
  reg [31:0] _RAND_1652;
  reg [31:0] _RAND_1653;
  reg [31:0] _RAND_1654;
  reg [31:0] _RAND_1655;
  reg [31:0] _RAND_1656;
  reg [31:0] _RAND_1657;
  reg [31:0] _RAND_1658;
  reg [31:0] _RAND_1659;
  reg [31:0] _RAND_1660;
  reg [31:0] _RAND_1661;
  reg [31:0] _RAND_1662;
  reg [31:0] _RAND_1663;
  reg [31:0] _RAND_1664;
  reg [31:0] _RAND_1665;
  reg [31:0] _RAND_1666;
  reg [31:0] _RAND_1667;
  reg [31:0] _RAND_1668;
  reg [31:0] _RAND_1669;
  reg [31:0] _RAND_1670;
  reg [31:0] _RAND_1671;
  reg [31:0] _RAND_1672;
  reg [31:0] _RAND_1673;
  reg [31:0] _RAND_1674;
  reg [31:0] _RAND_1675;
  reg [31:0] _RAND_1676;
  reg [31:0] _RAND_1677;
  reg [31:0] _RAND_1678;
  reg [31:0] _RAND_1679;
  reg [31:0] _RAND_1680;
  reg [31:0] _RAND_1681;
  reg [31:0] _RAND_1682;
  reg [31:0] _RAND_1683;
  reg [31:0] _RAND_1684;
  reg [31:0] _RAND_1685;
  reg [31:0] _RAND_1686;
  reg [31:0] _RAND_1687;
  reg [31:0] _RAND_1688;
  reg [31:0] _RAND_1689;
  reg [31:0] _RAND_1690;
  reg [31:0] _RAND_1691;
  reg [31:0] _RAND_1692;
  reg [31:0] _RAND_1693;
  reg [31:0] _RAND_1694;
  reg [31:0] _RAND_1695;
  reg [31:0] _RAND_1696;
  reg [31:0] _RAND_1697;
  reg [31:0] _RAND_1698;
  reg [31:0] _RAND_1699;
  reg [31:0] _RAND_1700;
  reg [31:0] _RAND_1701;
  reg [31:0] _RAND_1702;
  reg [31:0] _RAND_1703;
  reg [31:0] _RAND_1704;
  reg [31:0] _RAND_1705;
  reg [31:0] _RAND_1706;
  reg [31:0] _RAND_1707;
  reg [31:0] _RAND_1708;
  reg [31:0] _RAND_1709;
  reg [31:0] _RAND_1710;
  reg [31:0] _RAND_1711;
  reg [31:0] _RAND_1712;
  reg [31:0] _RAND_1713;
  reg [31:0] _RAND_1714;
  reg [31:0] _RAND_1715;
  reg [31:0] _RAND_1716;
  reg [31:0] _RAND_1717;
  reg [31:0] _RAND_1718;
  reg [31:0] _RAND_1719;
  reg [31:0] _RAND_1720;
  reg [31:0] _RAND_1721;
  reg [31:0] _RAND_1722;
  reg [31:0] _RAND_1723;
  reg [31:0] _RAND_1724;
  reg [31:0] _RAND_1725;
  reg [31:0] _RAND_1726;
  reg [31:0] _RAND_1727;
  reg [31:0] _RAND_1728;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] image_0_0; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_1; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_2; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_3; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_4; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_5; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_6; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_7; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_8; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_9; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_10; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_11; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_12; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_13; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_14; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_15; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_16; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_17; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_18; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_19; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_20; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_21; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_22; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_23; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_24; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_25; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_26; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_27; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_28; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_29; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_30; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_31; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_32; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_33; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_34; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_35; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_36; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_37; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_38; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_39; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_40; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_41; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_42; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_43; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_44; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_45; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_46; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_47; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_48; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_49; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_50; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_51; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_52; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_53; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_54; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_55; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_56; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_57; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_58; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_59; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_60; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_61; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_62; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_63; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_64; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_65; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_66; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_67; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_68; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_69; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_70; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_71; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_72; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_73; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_74; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_75; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_76; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_77; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_78; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_79; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_80; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_81; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_82; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_83; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_84; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_85; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_86; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_87; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_88; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_89; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_90; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_91; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_92; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_93; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_94; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_95; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_96; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_97; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_98; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_99; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_100; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_101; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_102; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_103; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_104; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_105; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_106; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_107; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_108; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_109; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_110; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_111; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_112; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_113; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_114; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_115; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_116; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_117; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_118; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_119; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_120; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_121; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_122; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_123; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_124; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_125; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_126; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_127; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_128; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_129; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_130; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_131; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_132; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_133; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_134; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_135; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_136; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_137; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_138; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_139; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_140; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_141; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_142; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_143; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_144; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_145; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_146; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_147; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_148; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_149; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_150; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_151; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_152; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_153; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_154; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_155; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_156; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_157; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_158; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_159; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_160; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_161; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_162; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_163; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_164; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_165; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_166; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_167; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_168; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_169; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_170; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_171; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_172; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_173; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_174; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_175; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_176; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_177; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_178; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_179; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_180; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_181; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_182; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_183; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_184; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_185; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_186; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_187; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_188; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_189; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_190; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_191; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_192; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_193; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_194; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_195; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_196; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_197; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_198; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_199; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_200; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_201; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_202; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_203; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_204; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_205; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_206; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_207; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_208; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_209; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_210; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_211; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_212; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_213; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_214; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_215; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_216; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_217; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_218; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_219; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_220; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_221; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_222; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_223; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_224; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_225; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_226; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_227; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_228; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_229; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_230; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_231; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_232; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_233; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_234; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_235; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_236; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_237; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_238; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_239; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_240; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_241; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_242; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_243; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_244; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_245; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_246; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_247; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_248; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_249; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_250; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_251; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_252; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_253; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_254; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_255; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_256; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_257; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_258; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_259; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_260; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_261; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_262; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_263; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_264; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_265; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_266; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_267; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_268; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_269; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_270; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_271; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_272; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_273; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_274; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_275; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_276; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_277; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_278; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_279; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_280; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_281; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_282; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_283; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_284; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_285; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_286; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_287; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_288; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_289; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_290; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_291; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_292; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_293; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_294; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_295; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_296; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_297; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_298; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_299; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_300; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_301; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_302; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_303; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_304; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_305; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_306; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_307; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_308; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_309; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_310; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_311; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_312; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_313; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_314; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_315; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_316; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_317; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_318; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_319; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_320; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_321; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_322; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_323; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_324; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_325; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_326; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_327; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_328; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_329; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_330; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_331; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_332; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_333; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_334; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_335; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_336; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_337; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_338; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_339; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_340; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_341; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_342; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_343; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_344; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_345; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_346; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_347; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_348; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_349; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_350; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_351; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_352; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_353; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_354; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_355; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_356; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_357; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_358; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_359; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_360; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_361; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_362; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_363; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_364; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_365; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_366; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_367; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_368; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_369; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_370; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_371; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_372; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_373; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_374; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_375; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_376; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_377; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_378; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_379; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_380; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_381; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_382; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_383; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_384; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_385; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_386; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_387; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_388; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_389; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_390; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_391; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_392; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_393; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_394; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_395; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_396; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_397; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_398; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_399; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_400; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_401; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_402; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_403; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_404; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_405; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_406; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_407; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_408; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_409; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_410; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_411; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_412; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_413; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_414; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_415; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_416; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_417; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_418; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_419; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_420; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_421; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_422; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_423; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_424; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_425; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_426; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_427; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_428; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_429; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_430; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_431; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_432; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_433; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_434; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_435; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_436; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_437; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_438; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_439; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_440; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_441; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_442; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_443; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_444; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_445; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_446; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_447; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_448; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_449; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_450; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_451; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_452; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_453; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_454; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_455; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_456; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_457; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_458; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_459; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_460; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_461; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_462; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_463; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_464; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_465; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_466; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_467; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_468; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_469; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_470; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_471; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_472; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_473; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_474; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_475; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_476; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_477; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_478; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_479; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_480; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_481; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_482; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_483; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_484; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_485; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_486; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_487; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_488; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_489; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_490; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_491; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_492; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_493; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_494; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_495; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_496; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_497; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_498; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_499; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_500; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_501; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_502; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_503; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_504; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_505; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_506; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_507; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_508; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_509; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_510; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_511; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_512; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_513; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_514; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_515; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_516; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_517; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_518; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_519; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_520; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_521; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_522; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_523; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_524; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_525; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_526; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_527; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_528; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_529; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_530; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_531; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_532; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_533; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_534; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_535; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_536; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_537; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_538; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_539; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_540; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_541; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_542; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_543; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_544; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_545; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_546; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_547; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_548; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_549; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_550; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_551; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_552; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_553; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_554; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_555; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_556; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_557; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_558; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_559; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_560; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_561; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_562; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_563; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_564; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_565; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_566; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_567; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_568; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_569; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_570; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_571; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_572; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_573; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_574; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_0_575; // @[VideoBuffer.scala 19:25]
  reg [3:0] image_1_0; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_1; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_2; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_3; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_4; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_5; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_6; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_7; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_8; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_9; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_10; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_11; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_12; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_13; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_14; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_15; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_16; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_17; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_18; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_19; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_20; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_21; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_22; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_23; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_24; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_25; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_26; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_27; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_28; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_29; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_30; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_31; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_32; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_33; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_34; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_35; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_36; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_37; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_38; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_39; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_40; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_41; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_42; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_43; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_44; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_45; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_46; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_47; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_48; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_49; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_50; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_51; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_52; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_53; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_54; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_55; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_56; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_57; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_58; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_59; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_60; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_61; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_62; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_63; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_64; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_65; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_66; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_67; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_68; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_69; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_70; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_71; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_72; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_73; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_74; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_75; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_76; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_77; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_78; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_79; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_80; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_81; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_82; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_83; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_84; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_85; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_86; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_87; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_88; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_89; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_90; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_91; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_92; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_93; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_94; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_95; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_96; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_97; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_98; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_99; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_100; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_101; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_102; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_103; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_104; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_105; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_106; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_107; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_108; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_109; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_110; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_111; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_112; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_113; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_114; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_115; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_116; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_117; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_118; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_119; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_120; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_121; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_122; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_123; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_124; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_125; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_126; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_127; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_128; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_129; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_130; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_131; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_132; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_133; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_134; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_135; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_136; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_137; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_138; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_139; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_140; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_141; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_142; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_143; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_144; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_145; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_146; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_147; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_148; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_149; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_150; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_151; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_152; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_153; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_154; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_155; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_156; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_157; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_158; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_159; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_160; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_161; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_162; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_163; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_164; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_165; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_166; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_167; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_168; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_169; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_170; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_171; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_172; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_173; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_174; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_175; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_176; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_177; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_178; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_179; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_180; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_181; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_182; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_183; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_184; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_185; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_186; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_187; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_188; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_189; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_190; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_191; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_192; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_193; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_194; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_195; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_196; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_197; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_198; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_199; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_200; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_201; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_202; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_203; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_204; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_205; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_206; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_207; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_208; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_209; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_210; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_211; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_212; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_213; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_214; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_215; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_216; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_217; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_218; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_219; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_220; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_221; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_222; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_223; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_224; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_225; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_226; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_227; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_228; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_229; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_230; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_231; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_232; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_233; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_234; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_235; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_236; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_237; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_238; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_239; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_240; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_241; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_242; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_243; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_244; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_245; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_246; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_247; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_248; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_249; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_250; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_251; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_252; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_253; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_254; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_255; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_256; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_257; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_258; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_259; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_260; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_261; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_262; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_263; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_264; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_265; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_266; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_267; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_268; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_269; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_270; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_271; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_272; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_273; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_274; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_275; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_276; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_277; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_278; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_279; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_280; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_281; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_282; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_283; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_284; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_285; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_286; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_287; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_288; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_289; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_290; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_291; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_292; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_293; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_294; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_295; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_296; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_297; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_298; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_299; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_300; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_301; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_302; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_303; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_304; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_305; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_306; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_307; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_308; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_309; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_310; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_311; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_312; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_313; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_314; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_315; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_316; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_317; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_318; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_319; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_320; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_321; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_322; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_323; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_324; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_325; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_326; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_327; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_328; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_329; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_330; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_331; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_332; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_333; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_334; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_335; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_336; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_337; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_338; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_339; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_340; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_341; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_342; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_343; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_344; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_345; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_346; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_347; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_348; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_349; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_350; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_351; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_352; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_353; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_354; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_355; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_356; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_357; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_358; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_359; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_360; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_361; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_362; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_363; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_364; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_365; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_366; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_367; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_368; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_369; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_370; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_371; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_372; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_373; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_374; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_375; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_376; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_377; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_378; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_379; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_380; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_381; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_382; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_383; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_384; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_385; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_386; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_387; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_388; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_389; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_390; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_391; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_392; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_393; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_394; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_395; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_396; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_397; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_398; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_399; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_400; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_401; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_402; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_403; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_404; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_405; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_406; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_407; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_408; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_409; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_410; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_411; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_412; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_413; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_414; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_415; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_416; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_417; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_418; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_419; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_420; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_421; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_422; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_423; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_424; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_425; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_426; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_427; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_428; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_429; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_430; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_431; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_432; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_433; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_434; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_435; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_436; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_437; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_438; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_439; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_440; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_441; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_442; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_443; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_444; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_445; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_446; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_447; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_448; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_449; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_450; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_451; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_452; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_453; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_454; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_455; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_456; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_457; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_458; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_459; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_460; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_461; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_462; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_463; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_464; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_465; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_466; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_467; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_468; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_469; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_470; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_471; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_472; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_473; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_474; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_475; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_476; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_477; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_478; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_479; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_480; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_481; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_482; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_483; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_484; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_485; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_486; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_487; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_488; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_489; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_490; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_491; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_492; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_493; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_494; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_495; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_496; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_497; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_498; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_499; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_500; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_501; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_502; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_503; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_504; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_505; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_506; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_507; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_508; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_509; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_510; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_511; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_512; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_513; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_514; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_515; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_516; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_517; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_518; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_519; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_520; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_521; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_522; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_523; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_524; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_525; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_526; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_527; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_528; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_529; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_530; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_531; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_532; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_533; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_534; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_535; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_536; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_537; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_538; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_539; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_540; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_541; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_542; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_543; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_544; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_545; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_546; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_547; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_548; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_549; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_550; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_551; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_552; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_553; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_554; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_555; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_556; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_557; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_558; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_559; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_560; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_561; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_562; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_563; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_564; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_565; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_566; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_567; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_568; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_569; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_570; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_571; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_572; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_573; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_574; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_1_575; // @[VideoBuffer.scala 20:25]
  reg [3:0] image_2_0; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_1; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_2; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_3; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_4; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_5; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_6; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_7; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_8; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_9; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_10; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_11; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_12; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_13; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_14; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_15; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_16; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_17; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_18; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_19; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_20; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_21; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_22; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_23; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_24; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_25; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_26; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_27; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_28; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_29; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_30; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_31; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_32; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_33; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_34; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_35; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_36; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_37; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_38; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_39; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_40; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_41; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_42; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_43; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_44; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_45; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_46; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_47; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_48; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_49; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_50; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_51; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_52; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_53; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_54; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_55; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_56; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_57; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_58; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_59; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_60; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_61; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_62; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_63; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_64; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_65; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_66; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_67; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_68; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_69; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_70; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_71; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_72; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_73; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_74; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_75; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_76; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_77; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_78; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_79; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_80; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_81; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_82; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_83; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_84; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_85; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_86; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_87; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_88; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_89; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_90; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_91; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_92; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_93; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_94; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_95; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_96; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_97; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_98; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_99; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_100; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_101; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_102; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_103; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_104; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_105; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_106; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_107; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_108; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_109; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_110; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_111; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_112; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_113; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_114; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_115; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_116; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_117; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_118; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_119; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_120; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_121; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_122; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_123; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_124; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_125; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_126; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_127; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_128; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_129; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_130; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_131; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_132; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_133; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_134; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_135; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_136; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_137; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_138; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_139; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_140; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_141; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_142; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_143; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_144; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_145; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_146; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_147; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_148; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_149; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_150; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_151; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_152; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_153; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_154; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_155; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_156; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_157; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_158; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_159; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_160; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_161; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_162; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_163; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_164; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_165; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_166; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_167; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_168; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_169; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_170; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_171; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_172; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_173; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_174; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_175; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_176; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_177; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_178; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_179; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_180; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_181; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_182; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_183; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_184; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_185; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_186; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_187; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_188; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_189; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_190; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_191; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_192; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_193; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_194; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_195; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_196; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_197; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_198; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_199; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_200; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_201; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_202; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_203; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_204; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_205; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_206; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_207; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_208; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_209; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_210; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_211; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_212; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_213; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_214; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_215; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_216; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_217; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_218; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_219; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_220; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_221; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_222; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_223; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_224; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_225; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_226; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_227; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_228; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_229; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_230; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_231; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_232; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_233; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_234; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_235; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_236; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_237; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_238; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_239; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_240; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_241; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_242; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_243; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_244; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_245; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_246; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_247; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_248; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_249; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_250; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_251; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_252; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_253; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_254; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_255; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_256; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_257; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_258; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_259; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_260; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_261; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_262; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_263; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_264; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_265; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_266; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_267; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_268; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_269; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_270; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_271; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_272; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_273; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_274; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_275; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_276; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_277; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_278; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_279; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_280; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_281; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_282; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_283; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_284; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_285; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_286; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_287; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_288; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_289; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_290; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_291; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_292; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_293; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_294; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_295; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_296; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_297; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_298; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_299; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_300; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_301; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_302; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_303; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_304; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_305; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_306; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_307; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_308; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_309; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_310; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_311; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_312; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_313; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_314; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_315; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_316; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_317; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_318; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_319; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_320; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_321; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_322; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_323; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_324; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_325; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_326; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_327; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_328; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_329; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_330; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_331; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_332; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_333; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_334; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_335; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_336; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_337; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_338; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_339; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_340; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_341; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_342; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_343; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_344; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_345; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_346; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_347; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_348; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_349; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_350; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_351; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_352; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_353; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_354; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_355; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_356; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_357; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_358; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_359; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_360; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_361; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_362; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_363; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_364; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_365; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_366; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_367; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_368; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_369; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_370; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_371; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_372; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_373; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_374; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_375; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_376; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_377; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_378; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_379; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_380; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_381; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_382; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_383; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_384; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_385; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_386; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_387; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_388; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_389; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_390; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_391; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_392; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_393; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_394; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_395; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_396; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_397; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_398; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_399; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_400; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_401; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_402; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_403; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_404; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_405; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_406; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_407; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_408; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_409; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_410; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_411; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_412; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_413; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_414; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_415; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_416; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_417; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_418; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_419; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_420; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_421; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_422; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_423; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_424; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_425; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_426; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_427; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_428; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_429; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_430; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_431; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_432; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_433; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_434; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_435; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_436; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_437; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_438; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_439; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_440; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_441; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_442; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_443; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_444; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_445; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_446; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_447; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_448; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_449; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_450; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_451; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_452; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_453; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_454; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_455; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_456; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_457; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_458; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_459; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_460; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_461; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_462; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_463; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_464; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_465; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_466; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_467; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_468; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_469; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_470; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_471; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_472; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_473; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_474; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_475; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_476; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_477; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_478; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_479; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_480; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_481; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_482; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_483; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_484; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_485; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_486; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_487; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_488; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_489; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_490; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_491; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_492; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_493; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_494; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_495; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_496; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_497; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_498; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_499; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_500; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_501; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_502; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_503; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_504; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_505; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_506; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_507; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_508; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_509; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_510; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_511; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_512; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_513; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_514; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_515; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_516; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_517; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_518; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_519; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_520; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_521; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_522; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_523; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_524; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_525; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_526; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_527; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_528; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_529; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_530; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_531; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_532; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_533; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_534; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_535; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_536; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_537; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_538; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_539; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_540; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_541; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_542; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_543; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_544; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_545; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_546; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_547; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_548; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_549; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_550; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_551; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_552; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_553; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_554; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_555; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_556; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_557; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_558; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_559; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_560; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_561; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_562; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_563; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_564; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_565; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_566; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_567; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_568; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_569; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_570; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_571; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_572; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_573; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_574; // @[VideoBuffer.scala 21:25]
  reg [3:0] image_2_575; // @[VideoBuffer.scala 21:25]
  reg [31:0] pixelIndex; // @[VideoBuffer.scala 24:33]
  wire [16:0] _T_3 = io_rowIndex * 11'h20; // @[VideoBuffer.scala 27:54]
  wire [16:0] _GEN_17282 = {{6'd0}, io_colIndex}; // @[VideoBuffer.scala 27:69]
  wire [16:0] _T_5 = _T_3 + _GEN_17282; // @[VideoBuffer.scala 27:69]
  wire [3:0] _GEN_1 = 10'h1 == _T_5[9:0] ? image_0_1 : image_0_0; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_2 = 10'h2 == _T_5[9:0] ? image_0_2 : _GEN_1; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_3 = 10'h3 == _T_5[9:0] ? image_0_3 : _GEN_2; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_4 = 10'h4 == _T_5[9:0] ? image_0_4 : _GEN_3; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_5 = 10'h5 == _T_5[9:0] ? image_0_5 : _GEN_4; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_6 = 10'h6 == _T_5[9:0] ? image_0_6 : _GEN_5; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_7 = 10'h7 == _T_5[9:0] ? image_0_7 : _GEN_6; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_8 = 10'h8 == _T_5[9:0] ? image_0_8 : _GEN_7; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_9 = 10'h9 == _T_5[9:0] ? image_0_9 : _GEN_8; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_10 = 10'ha == _T_5[9:0] ? image_0_10 : _GEN_9; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_11 = 10'hb == _T_5[9:0] ? image_0_11 : _GEN_10; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_12 = 10'hc == _T_5[9:0] ? image_0_12 : _GEN_11; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_13 = 10'hd == _T_5[9:0] ? image_0_13 : _GEN_12; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_14 = 10'he == _T_5[9:0] ? image_0_14 : _GEN_13; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_15 = 10'hf == _T_5[9:0] ? image_0_15 : _GEN_14; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_16 = 10'h10 == _T_5[9:0] ? image_0_16 : _GEN_15; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_17 = 10'h11 == _T_5[9:0] ? image_0_17 : _GEN_16; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_18 = 10'h12 == _T_5[9:0] ? image_0_18 : _GEN_17; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_19 = 10'h13 == _T_5[9:0] ? image_0_19 : _GEN_18; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_20 = 10'h14 == _T_5[9:0] ? image_0_20 : _GEN_19; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_21 = 10'h15 == _T_5[9:0] ? image_0_21 : _GEN_20; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_22 = 10'h16 == _T_5[9:0] ? image_0_22 : _GEN_21; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_23 = 10'h17 == _T_5[9:0] ? image_0_23 : _GEN_22; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_24 = 10'h18 == _T_5[9:0] ? image_0_24 : _GEN_23; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_25 = 10'h19 == _T_5[9:0] ? image_0_25 : _GEN_24; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_26 = 10'h1a == _T_5[9:0] ? image_0_26 : _GEN_25; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_27 = 10'h1b == _T_5[9:0] ? image_0_27 : _GEN_26; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_28 = 10'h1c == _T_5[9:0] ? image_0_28 : _GEN_27; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_29 = 10'h1d == _T_5[9:0] ? image_0_29 : _GEN_28; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_30 = 10'h1e == _T_5[9:0] ? image_0_30 : _GEN_29; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_31 = 10'h1f == _T_5[9:0] ? image_0_31 : _GEN_30; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_32 = 10'h20 == _T_5[9:0] ? image_0_32 : _GEN_31; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_33 = 10'h21 == _T_5[9:0] ? image_0_33 : _GEN_32; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_34 = 10'h22 == _T_5[9:0] ? image_0_34 : _GEN_33; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_35 = 10'h23 == _T_5[9:0] ? image_0_35 : _GEN_34; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_36 = 10'h24 == _T_5[9:0] ? image_0_36 : _GEN_35; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_37 = 10'h25 == _T_5[9:0] ? image_0_37 : _GEN_36; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_38 = 10'h26 == _T_5[9:0] ? image_0_38 : _GEN_37; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_39 = 10'h27 == _T_5[9:0] ? image_0_39 : _GEN_38; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_40 = 10'h28 == _T_5[9:0] ? image_0_40 : _GEN_39; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_41 = 10'h29 == _T_5[9:0] ? image_0_41 : _GEN_40; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_42 = 10'h2a == _T_5[9:0] ? image_0_42 : _GEN_41; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_43 = 10'h2b == _T_5[9:0] ? image_0_43 : _GEN_42; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_44 = 10'h2c == _T_5[9:0] ? image_0_44 : _GEN_43; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_45 = 10'h2d == _T_5[9:0] ? image_0_45 : _GEN_44; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_46 = 10'h2e == _T_5[9:0] ? image_0_46 : _GEN_45; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_47 = 10'h2f == _T_5[9:0] ? image_0_47 : _GEN_46; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_48 = 10'h30 == _T_5[9:0] ? image_0_48 : _GEN_47; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_49 = 10'h31 == _T_5[9:0] ? image_0_49 : _GEN_48; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_50 = 10'h32 == _T_5[9:0] ? image_0_50 : _GEN_49; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_51 = 10'h33 == _T_5[9:0] ? image_0_51 : _GEN_50; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_52 = 10'h34 == _T_5[9:0] ? image_0_52 : _GEN_51; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_53 = 10'h35 == _T_5[9:0] ? image_0_53 : _GEN_52; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_54 = 10'h36 == _T_5[9:0] ? image_0_54 : _GEN_53; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_55 = 10'h37 == _T_5[9:0] ? image_0_55 : _GEN_54; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_56 = 10'h38 == _T_5[9:0] ? image_0_56 : _GEN_55; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_57 = 10'h39 == _T_5[9:0] ? image_0_57 : _GEN_56; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_58 = 10'h3a == _T_5[9:0] ? image_0_58 : _GEN_57; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_59 = 10'h3b == _T_5[9:0] ? image_0_59 : _GEN_58; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_60 = 10'h3c == _T_5[9:0] ? image_0_60 : _GEN_59; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_61 = 10'h3d == _T_5[9:0] ? image_0_61 : _GEN_60; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_62 = 10'h3e == _T_5[9:0] ? image_0_62 : _GEN_61; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_63 = 10'h3f == _T_5[9:0] ? image_0_63 : _GEN_62; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_64 = 10'h40 == _T_5[9:0] ? image_0_64 : _GEN_63; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_65 = 10'h41 == _T_5[9:0] ? image_0_65 : _GEN_64; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_66 = 10'h42 == _T_5[9:0] ? image_0_66 : _GEN_65; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_67 = 10'h43 == _T_5[9:0] ? image_0_67 : _GEN_66; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_68 = 10'h44 == _T_5[9:0] ? image_0_68 : _GEN_67; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_69 = 10'h45 == _T_5[9:0] ? image_0_69 : _GEN_68; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_70 = 10'h46 == _T_5[9:0] ? image_0_70 : _GEN_69; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_71 = 10'h47 == _T_5[9:0] ? image_0_71 : _GEN_70; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_72 = 10'h48 == _T_5[9:0] ? image_0_72 : _GEN_71; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_73 = 10'h49 == _T_5[9:0] ? image_0_73 : _GEN_72; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_74 = 10'h4a == _T_5[9:0] ? image_0_74 : _GEN_73; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_75 = 10'h4b == _T_5[9:0] ? image_0_75 : _GEN_74; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_76 = 10'h4c == _T_5[9:0] ? image_0_76 : _GEN_75; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_77 = 10'h4d == _T_5[9:0] ? image_0_77 : _GEN_76; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_78 = 10'h4e == _T_5[9:0] ? image_0_78 : _GEN_77; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_79 = 10'h4f == _T_5[9:0] ? image_0_79 : _GEN_78; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_80 = 10'h50 == _T_5[9:0] ? image_0_80 : _GEN_79; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_81 = 10'h51 == _T_5[9:0] ? image_0_81 : _GEN_80; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_82 = 10'h52 == _T_5[9:0] ? image_0_82 : _GEN_81; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_83 = 10'h53 == _T_5[9:0] ? image_0_83 : _GEN_82; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_84 = 10'h54 == _T_5[9:0] ? image_0_84 : _GEN_83; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_85 = 10'h55 == _T_5[9:0] ? image_0_85 : _GEN_84; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_86 = 10'h56 == _T_5[9:0] ? image_0_86 : _GEN_85; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_87 = 10'h57 == _T_5[9:0] ? image_0_87 : _GEN_86; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_88 = 10'h58 == _T_5[9:0] ? image_0_88 : _GEN_87; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_89 = 10'h59 == _T_5[9:0] ? image_0_89 : _GEN_88; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_90 = 10'h5a == _T_5[9:0] ? image_0_90 : _GEN_89; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_91 = 10'h5b == _T_5[9:0] ? image_0_91 : _GEN_90; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_92 = 10'h5c == _T_5[9:0] ? image_0_92 : _GEN_91; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_93 = 10'h5d == _T_5[9:0] ? image_0_93 : _GEN_92; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_94 = 10'h5e == _T_5[9:0] ? image_0_94 : _GEN_93; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_95 = 10'h5f == _T_5[9:0] ? image_0_95 : _GEN_94; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_96 = 10'h60 == _T_5[9:0] ? image_0_96 : _GEN_95; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_97 = 10'h61 == _T_5[9:0] ? image_0_97 : _GEN_96; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_98 = 10'h62 == _T_5[9:0] ? image_0_98 : _GEN_97; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_99 = 10'h63 == _T_5[9:0] ? image_0_99 : _GEN_98; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_100 = 10'h64 == _T_5[9:0] ? image_0_100 : _GEN_99; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_101 = 10'h65 == _T_5[9:0] ? image_0_101 : _GEN_100; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_102 = 10'h66 == _T_5[9:0] ? image_0_102 : _GEN_101; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_103 = 10'h67 == _T_5[9:0] ? image_0_103 : _GEN_102; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_104 = 10'h68 == _T_5[9:0] ? image_0_104 : _GEN_103; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_105 = 10'h69 == _T_5[9:0] ? image_0_105 : _GEN_104; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_106 = 10'h6a == _T_5[9:0] ? image_0_106 : _GEN_105; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_107 = 10'h6b == _T_5[9:0] ? image_0_107 : _GEN_106; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_108 = 10'h6c == _T_5[9:0] ? image_0_108 : _GEN_107; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_109 = 10'h6d == _T_5[9:0] ? image_0_109 : _GEN_108; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_110 = 10'h6e == _T_5[9:0] ? image_0_110 : _GEN_109; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_111 = 10'h6f == _T_5[9:0] ? image_0_111 : _GEN_110; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_112 = 10'h70 == _T_5[9:0] ? image_0_112 : _GEN_111; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_113 = 10'h71 == _T_5[9:0] ? image_0_113 : _GEN_112; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_114 = 10'h72 == _T_5[9:0] ? image_0_114 : _GEN_113; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_115 = 10'h73 == _T_5[9:0] ? image_0_115 : _GEN_114; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_116 = 10'h74 == _T_5[9:0] ? image_0_116 : _GEN_115; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_117 = 10'h75 == _T_5[9:0] ? image_0_117 : _GEN_116; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_118 = 10'h76 == _T_5[9:0] ? image_0_118 : _GEN_117; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_119 = 10'h77 == _T_5[9:0] ? image_0_119 : _GEN_118; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_120 = 10'h78 == _T_5[9:0] ? image_0_120 : _GEN_119; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_121 = 10'h79 == _T_5[9:0] ? image_0_121 : _GEN_120; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_122 = 10'h7a == _T_5[9:0] ? image_0_122 : _GEN_121; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_123 = 10'h7b == _T_5[9:0] ? image_0_123 : _GEN_122; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_124 = 10'h7c == _T_5[9:0] ? image_0_124 : _GEN_123; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_125 = 10'h7d == _T_5[9:0] ? image_0_125 : _GEN_124; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_126 = 10'h7e == _T_5[9:0] ? image_0_126 : _GEN_125; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_127 = 10'h7f == _T_5[9:0] ? image_0_127 : _GEN_126; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_128 = 10'h80 == _T_5[9:0] ? image_0_128 : _GEN_127; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_129 = 10'h81 == _T_5[9:0] ? image_0_129 : _GEN_128; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_130 = 10'h82 == _T_5[9:0] ? image_0_130 : _GEN_129; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_131 = 10'h83 == _T_5[9:0] ? image_0_131 : _GEN_130; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_132 = 10'h84 == _T_5[9:0] ? image_0_132 : _GEN_131; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_133 = 10'h85 == _T_5[9:0] ? image_0_133 : _GEN_132; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_134 = 10'h86 == _T_5[9:0] ? image_0_134 : _GEN_133; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_135 = 10'h87 == _T_5[9:0] ? image_0_135 : _GEN_134; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_136 = 10'h88 == _T_5[9:0] ? image_0_136 : _GEN_135; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_137 = 10'h89 == _T_5[9:0] ? image_0_137 : _GEN_136; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_138 = 10'h8a == _T_5[9:0] ? image_0_138 : _GEN_137; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_139 = 10'h8b == _T_5[9:0] ? image_0_139 : _GEN_138; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_140 = 10'h8c == _T_5[9:0] ? image_0_140 : _GEN_139; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_141 = 10'h8d == _T_5[9:0] ? image_0_141 : _GEN_140; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_142 = 10'h8e == _T_5[9:0] ? image_0_142 : _GEN_141; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_143 = 10'h8f == _T_5[9:0] ? image_0_143 : _GEN_142; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_144 = 10'h90 == _T_5[9:0] ? image_0_144 : _GEN_143; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_145 = 10'h91 == _T_5[9:0] ? image_0_145 : _GEN_144; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_146 = 10'h92 == _T_5[9:0] ? image_0_146 : _GEN_145; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_147 = 10'h93 == _T_5[9:0] ? image_0_147 : _GEN_146; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_148 = 10'h94 == _T_5[9:0] ? image_0_148 : _GEN_147; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_149 = 10'h95 == _T_5[9:0] ? image_0_149 : _GEN_148; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_150 = 10'h96 == _T_5[9:0] ? image_0_150 : _GEN_149; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_151 = 10'h97 == _T_5[9:0] ? image_0_151 : _GEN_150; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_152 = 10'h98 == _T_5[9:0] ? image_0_152 : _GEN_151; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_153 = 10'h99 == _T_5[9:0] ? image_0_153 : _GEN_152; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_154 = 10'h9a == _T_5[9:0] ? image_0_154 : _GEN_153; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_155 = 10'h9b == _T_5[9:0] ? image_0_155 : _GEN_154; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_156 = 10'h9c == _T_5[9:0] ? image_0_156 : _GEN_155; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_157 = 10'h9d == _T_5[9:0] ? image_0_157 : _GEN_156; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_158 = 10'h9e == _T_5[9:0] ? image_0_158 : _GEN_157; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_159 = 10'h9f == _T_5[9:0] ? image_0_159 : _GEN_158; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_160 = 10'ha0 == _T_5[9:0] ? image_0_160 : _GEN_159; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_161 = 10'ha1 == _T_5[9:0] ? image_0_161 : _GEN_160; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_162 = 10'ha2 == _T_5[9:0] ? image_0_162 : _GEN_161; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_163 = 10'ha3 == _T_5[9:0] ? image_0_163 : _GEN_162; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_164 = 10'ha4 == _T_5[9:0] ? image_0_164 : _GEN_163; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_165 = 10'ha5 == _T_5[9:0] ? image_0_165 : _GEN_164; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_166 = 10'ha6 == _T_5[9:0] ? image_0_166 : _GEN_165; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_167 = 10'ha7 == _T_5[9:0] ? image_0_167 : _GEN_166; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_168 = 10'ha8 == _T_5[9:0] ? image_0_168 : _GEN_167; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_169 = 10'ha9 == _T_5[9:0] ? image_0_169 : _GEN_168; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_170 = 10'haa == _T_5[9:0] ? image_0_170 : _GEN_169; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_171 = 10'hab == _T_5[9:0] ? image_0_171 : _GEN_170; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_172 = 10'hac == _T_5[9:0] ? image_0_172 : _GEN_171; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_173 = 10'had == _T_5[9:0] ? image_0_173 : _GEN_172; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_174 = 10'hae == _T_5[9:0] ? image_0_174 : _GEN_173; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_175 = 10'haf == _T_5[9:0] ? image_0_175 : _GEN_174; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_176 = 10'hb0 == _T_5[9:0] ? image_0_176 : _GEN_175; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_177 = 10'hb1 == _T_5[9:0] ? image_0_177 : _GEN_176; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_178 = 10'hb2 == _T_5[9:0] ? image_0_178 : _GEN_177; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_179 = 10'hb3 == _T_5[9:0] ? image_0_179 : _GEN_178; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_180 = 10'hb4 == _T_5[9:0] ? image_0_180 : _GEN_179; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_181 = 10'hb5 == _T_5[9:0] ? image_0_181 : _GEN_180; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_182 = 10'hb6 == _T_5[9:0] ? image_0_182 : _GEN_181; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_183 = 10'hb7 == _T_5[9:0] ? image_0_183 : _GEN_182; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_184 = 10'hb8 == _T_5[9:0] ? image_0_184 : _GEN_183; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_185 = 10'hb9 == _T_5[9:0] ? image_0_185 : _GEN_184; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_186 = 10'hba == _T_5[9:0] ? image_0_186 : _GEN_185; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_187 = 10'hbb == _T_5[9:0] ? image_0_187 : _GEN_186; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_188 = 10'hbc == _T_5[9:0] ? image_0_188 : _GEN_187; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_189 = 10'hbd == _T_5[9:0] ? image_0_189 : _GEN_188; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_190 = 10'hbe == _T_5[9:0] ? image_0_190 : _GEN_189; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_191 = 10'hbf == _T_5[9:0] ? image_0_191 : _GEN_190; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_192 = 10'hc0 == _T_5[9:0] ? image_0_192 : _GEN_191; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_193 = 10'hc1 == _T_5[9:0] ? image_0_193 : _GEN_192; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_194 = 10'hc2 == _T_5[9:0] ? image_0_194 : _GEN_193; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_195 = 10'hc3 == _T_5[9:0] ? image_0_195 : _GEN_194; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_196 = 10'hc4 == _T_5[9:0] ? image_0_196 : _GEN_195; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_197 = 10'hc5 == _T_5[9:0] ? image_0_197 : _GEN_196; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_198 = 10'hc6 == _T_5[9:0] ? image_0_198 : _GEN_197; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_199 = 10'hc7 == _T_5[9:0] ? image_0_199 : _GEN_198; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_200 = 10'hc8 == _T_5[9:0] ? image_0_200 : _GEN_199; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_201 = 10'hc9 == _T_5[9:0] ? image_0_201 : _GEN_200; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_202 = 10'hca == _T_5[9:0] ? image_0_202 : _GEN_201; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_203 = 10'hcb == _T_5[9:0] ? image_0_203 : _GEN_202; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_204 = 10'hcc == _T_5[9:0] ? image_0_204 : _GEN_203; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_205 = 10'hcd == _T_5[9:0] ? image_0_205 : _GEN_204; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_206 = 10'hce == _T_5[9:0] ? image_0_206 : _GEN_205; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_207 = 10'hcf == _T_5[9:0] ? image_0_207 : _GEN_206; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_208 = 10'hd0 == _T_5[9:0] ? image_0_208 : _GEN_207; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_209 = 10'hd1 == _T_5[9:0] ? image_0_209 : _GEN_208; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_210 = 10'hd2 == _T_5[9:0] ? image_0_210 : _GEN_209; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_211 = 10'hd3 == _T_5[9:0] ? image_0_211 : _GEN_210; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_212 = 10'hd4 == _T_5[9:0] ? image_0_212 : _GEN_211; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_213 = 10'hd5 == _T_5[9:0] ? image_0_213 : _GEN_212; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_214 = 10'hd6 == _T_5[9:0] ? image_0_214 : _GEN_213; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_215 = 10'hd7 == _T_5[9:0] ? image_0_215 : _GEN_214; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_216 = 10'hd8 == _T_5[9:0] ? image_0_216 : _GEN_215; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_217 = 10'hd9 == _T_5[9:0] ? image_0_217 : _GEN_216; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_218 = 10'hda == _T_5[9:0] ? image_0_218 : _GEN_217; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_219 = 10'hdb == _T_5[9:0] ? image_0_219 : _GEN_218; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_220 = 10'hdc == _T_5[9:0] ? image_0_220 : _GEN_219; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_221 = 10'hdd == _T_5[9:0] ? image_0_221 : _GEN_220; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_222 = 10'hde == _T_5[9:0] ? image_0_222 : _GEN_221; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_223 = 10'hdf == _T_5[9:0] ? image_0_223 : _GEN_222; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_224 = 10'he0 == _T_5[9:0] ? image_0_224 : _GEN_223; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_225 = 10'he1 == _T_5[9:0] ? image_0_225 : _GEN_224; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_226 = 10'he2 == _T_5[9:0] ? image_0_226 : _GEN_225; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_227 = 10'he3 == _T_5[9:0] ? image_0_227 : _GEN_226; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_228 = 10'he4 == _T_5[9:0] ? image_0_228 : _GEN_227; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_229 = 10'he5 == _T_5[9:0] ? image_0_229 : _GEN_228; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_230 = 10'he6 == _T_5[9:0] ? image_0_230 : _GEN_229; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_231 = 10'he7 == _T_5[9:0] ? image_0_231 : _GEN_230; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_232 = 10'he8 == _T_5[9:0] ? image_0_232 : _GEN_231; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_233 = 10'he9 == _T_5[9:0] ? image_0_233 : _GEN_232; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_234 = 10'hea == _T_5[9:0] ? image_0_234 : _GEN_233; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_235 = 10'heb == _T_5[9:0] ? image_0_235 : _GEN_234; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_236 = 10'hec == _T_5[9:0] ? image_0_236 : _GEN_235; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_237 = 10'hed == _T_5[9:0] ? image_0_237 : _GEN_236; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_238 = 10'hee == _T_5[9:0] ? image_0_238 : _GEN_237; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_239 = 10'hef == _T_5[9:0] ? image_0_239 : _GEN_238; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_240 = 10'hf0 == _T_5[9:0] ? image_0_240 : _GEN_239; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_241 = 10'hf1 == _T_5[9:0] ? image_0_241 : _GEN_240; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_242 = 10'hf2 == _T_5[9:0] ? image_0_242 : _GEN_241; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_243 = 10'hf3 == _T_5[9:0] ? image_0_243 : _GEN_242; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_244 = 10'hf4 == _T_5[9:0] ? image_0_244 : _GEN_243; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_245 = 10'hf5 == _T_5[9:0] ? image_0_245 : _GEN_244; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_246 = 10'hf6 == _T_5[9:0] ? image_0_246 : _GEN_245; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_247 = 10'hf7 == _T_5[9:0] ? image_0_247 : _GEN_246; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_248 = 10'hf8 == _T_5[9:0] ? image_0_248 : _GEN_247; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_249 = 10'hf9 == _T_5[9:0] ? image_0_249 : _GEN_248; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_250 = 10'hfa == _T_5[9:0] ? image_0_250 : _GEN_249; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_251 = 10'hfb == _T_5[9:0] ? image_0_251 : _GEN_250; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_252 = 10'hfc == _T_5[9:0] ? image_0_252 : _GEN_251; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_253 = 10'hfd == _T_5[9:0] ? image_0_253 : _GEN_252; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_254 = 10'hfe == _T_5[9:0] ? image_0_254 : _GEN_253; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_255 = 10'hff == _T_5[9:0] ? image_0_255 : _GEN_254; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_256 = 10'h100 == _T_5[9:0] ? image_0_256 : _GEN_255; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_257 = 10'h101 == _T_5[9:0] ? image_0_257 : _GEN_256; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_258 = 10'h102 == _T_5[9:0] ? image_0_258 : _GEN_257; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_259 = 10'h103 == _T_5[9:0] ? image_0_259 : _GEN_258; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_260 = 10'h104 == _T_5[9:0] ? image_0_260 : _GEN_259; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_261 = 10'h105 == _T_5[9:0] ? image_0_261 : _GEN_260; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_262 = 10'h106 == _T_5[9:0] ? image_0_262 : _GEN_261; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_263 = 10'h107 == _T_5[9:0] ? image_0_263 : _GEN_262; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_264 = 10'h108 == _T_5[9:0] ? image_0_264 : _GEN_263; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_265 = 10'h109 == _T_5[9:0] ? image_0_265 : _GEN_264; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_266 = 10'h10a == _T_5[9:0] ? image_0_266 : _GEN_265; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_267 = 10'h10b == _T_5[9:0] ? image_0_267 : _GEN_266; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_268 = 10'h10c == _T_5[9:0] ? image_0_268 : _GEN_267; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_269 = 10'h10d == _T_5[9:0] ? image_0_269 : _GEN_268; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_270 = 10'h10e == _T_5[9:0] ? image_0_270 : _GEN_269; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_271 = 10'h10f == _T_5[9:0] ? image_0_271 : _GEN_270; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_272 = 10'h110 == _T_5[9:0] ? image_0_272 : _GEN_271; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_273 = 10'h111 == _T_5[9:0] ? image_0_273 : _GEN_272; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_274 = 10'h112 == _T_5[9:0] ? image_0_274 : _GEN_273; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_275 = 10'h113 == _T_5[9:0] ? image_0_275 : _GEN_274; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_276 = 10'h114 == _T_5[9:0] ? image_0_276 : _GEN_275; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_277 = 10'h115 == _T_5[9:0] ? image_0_277 : _GEN_276; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_278 = 10'h116 == _T_5[9:0] ? image_0_278 : _GEN_277; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_279 = 10'h117 == _T_5[9:0] ? image_0_279 : _GEN_278; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_280 = 10'h118 == _T_5[9:0] ? image_0_280 : _GEN_279; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_281 = 10'h119 == _T_5[9:0] ? image_0_281 : _GEN_280; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_282 = 10'h11a == _T_5[9:0] ? image_0_282 : _GEN_281; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_283 = 10'h11b == _T_5[9:0] ? image_0_283 : _GEN_282; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_284 = 10'h11c == _T_5[9:0] ? image_0_284 : _GEN_283; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_285 = 10'h11d == _T_5[9:0] ? image_0_285 : _GEN_284; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_286 = 10'h11e == _T_5[9:0] ? image_0_286 : _GEN_285; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_287 = 10'h11f == _T_5[9:0] ? image_0_287 : _GEN_286; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_288 = 10'h120 == _T_5[9:0] ? image_0_288 : _GEN_287; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_289 = 10'h121 == _T_5[9:0] ? image_0_289 : _GEN_288; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_290 = 10'h122 == _T_5[9:0] ? image_0_290 : _GEN_289; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_291 = 10'h123 == _T_5[9:0] ? image_0_291 : _GEN_290; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_292 = 10'h124 == _T_5[9:0] ? image_0_292 : _GEN_291; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_293 = 10'h125 == _T_5[9:0] ? image_0_293 : _GEN_292; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_294 = 10'h126 == _T_5[9:0] ? image_0_294 : _GEN_293; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_295 = 10'h127 == _T_5[9:0] ? image_0_295 : _GEN_294; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_296 = 10'h128 == _T_5[9:0] ? image_0_296 : _GEN_295; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_297 = 10'h129 == _T_5[9:0] ? image_0_297 : _GEN_296; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_298 = 10'h12a == _T_5[9:0] ? image_0_298 : _GEN_297; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_299 = 10'h12b == _T_5[9:0] ? image_0_299 : _GEN_298; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_300 = 10'h12c == _T_5[9:0] ? image_0_300 : _GEN_299; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_301 = 10'h12d == _T_5[9:0] ? image_0_301 : _GEN_300; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_302 = 10'h12e == _T_5[9:0] ? image_0_302 : _GEN_301; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_303 = 10'h12f == _T_5[9:0] ? image_0_303 : _GEN_302; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_304 = 10'h130 == _T_5[9:0] ? image_0_304 : _GEN_303; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_305 = 10'h131 == _T_5[9:0] ? image_0_305 : _GEN_304; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_306 = 10'h132 == _T_5[9:0] ? image_0_306 : _GEN_305; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_307 = 10'h133 == _T_5[9:0] ? image_0_307 : _GEN_306; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_308 = 10'h134 == _T_5[9:0] ? image_0_308 : _GEN_307; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_309 = 10'h135 == _T_5[9:0] ? image_0_309 : _GEN_308; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_310 = 10'h136 == _T_5[9:0] ? image_0_310 : _GEN_309; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_311 = 10'h137 == _T_5[9:0] ? image_0_311 : _GEN_310; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_312 = 10'h138 == _T_5[9:0] ? image_0_312 : _GEN_311; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_313 = 10'h139 == _T_5[9:0] ? image_0_313 : _GEN_312; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_314 = 10'h13a == _T_5[9:0] ? image_0_314 : _GEN_313; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_315 = 10'h13b == _T_5[9:0] ? image_0_315 : _GEN_314; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_316 = 10'h13c == _T_5[9:0] ? image_0_316 : _GEN_315; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_317 = 10'h13d == _T_5[9:0] ? image_0_317 : _GEN_316; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_318 = 10'h13e == _T_5[9:0] ? image_0_318 : _GEN_317; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_319 = 10'h13f == _T_5[9:0] ? image_0_319 : _GEN_318; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_320 = 10'h140 == _T_5[9:0] ? image_0_320 : _GEN_319; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_321 = 10'h141 == _T_5[9:0] ? image_0_321 : _GEN_320; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_322 = 10'h142 == _T_5[9:0] ? image_0_322 : _GEN_321; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_323 = 10'h143 == _T_5[9:0] ? image_0_323 : _GEN_322; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_324 = 10'h144 == _T_5[9:0] ? image_0_324 : _GEN_323; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_325 = 10'h145 == _T_5[9:0] ? image_0_325 : _GEN_324; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_326 = 10'h146 == _T_5[9:0] ? image_0_326 : _GEN_325; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_327 = 10'h147 == _T_5[9:0] ? image_0_327 : _GEN_326; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_328 = 10'h148 == _T_5[9:0] ? image_0_328 : _GEN_327; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_329 = 10'h149 == _T_5[9:0] ? image_0_329 : _GEN_328; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_330 = 10'h14a == _T_5[9:0] ? image_0_330 : _GEN_329; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_331 = 10'h14b == _T_5[9:0] ? image_0_331 : _GEN_330; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_332 = 10'h14c == _T_5[9:0] ? image_0_332 : _GEN_331; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_333 = 10'h14d == _T_5[9:0] ? image_0_333 : _GEN_332; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_334 = 10'h14e == _T_5[9:0] ? image_0_334 : _GEN_333; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_335 = 10'h14f == _T_5[9:0] ? image_0_335 : _GEN_334; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_336 = 10'h150 == _T_5[9:0] ? image_0_336 : _GEN_335; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_337 = 10'h151 == _T_5[9:0] ? image_0_337 : _GEN_336; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_338 = 10'h152 == _T_5[9:0] ? image_0_338 : _GEN_337; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_339 = 10'h153 == _T_5[9:0] ? image_0_339 : _GEN_338; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_340 = 10'h154 == _T_5[9:0] ? image_0_340 : _GEN_339; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_341 = 10'h155 == _T_5[9:0] ? image_0_341 : _GEN_340; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_342 = 10'h156 == _T_5[9:0] ? image_0_342 : _GEN_341; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_343 = 10'h157 == _T_5[9:0] ? image_0_343 : _GEN_342; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_344 = 10'h158 == _T_5[9:0] ? image_0_344 : _GEN_343; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_345 = 10'h159 == _T_5[9:0] ? image_0_345 : _GEN_344; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_346 = 10'h15a == _T_5[9:0] ? image_0_346 : _GEN_345; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_347 = 10'h15b == _T_5[9:0] ? image_0_347 : _GEN_346; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_348 = 10'h15c == _T_5[9:0] ? image_0_348 : _GEN_347; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_349 = 10'h15d == _T_5[9:0] ? image_0_349 : _GEN_348; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_350 = 10'h15e == _T_5[9:0] ? image_0_350 : _GEN_349; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_351 = 10'h15f == _T_5[9:0] ? image_0_351 : _GEN_350; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_352 = 10'h160 == _T_5[9:0] ? image_0_352 : _GEN_351; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_353 = 10'h161 == _T_5[9:0] ? image_0_353 : _GEN_352; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_354 = 10'h162 == _T_5[9:0] ? image_0_354 : _GEN_353; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_355 = 10'h163 == _T_5[9:0] ? image_0_355 : _GEN_354; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_356 = 10'h164 == _T_5[9:0] ? image_0_356 : _GEN_355; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_357 = 10'h165 == _T_5[9:0] ? image_0_357 : _GEN_356; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_358 = 10'h166 == _T_5[9:0] ? image_0_358 : _GEN_357; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_359 = 10'h167 == _T_5[9:0] ? image_0_359 : _GEN_358; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_360 = 10'h168 == _T_5[9:0] ? image_0_360 : _GEN_359; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_361 = 10'h169 == _T_5[9:0] ? image_0_361 : _GEN_360; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_362 = 10'h16a == _T_5[9:0] ? image_0_362 : _GEN_361; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_363 = 10'h16b == _T_5[9:0] ? image_0_363 : _GEN_362; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_364 = 10'h16c == _T_5[9:0] ? image_0_364 : _GEN_363; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_365 = 10'h16d == _T_5[9:0] ? image_0_365 : _GEN_364; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_366 = 10'h16e == _T_5[9:0] ? image_0_366 : _GEN_365; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_367 = 10'h16f == _T_5[9:0] ? image_0_367 : _GEN_366; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_368 = 10'h170 == _T_5[9:0] ? image_0_368 : _GEN_367; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_369 = 10'h171 == _T_5[9:0] ? image_0_369 : _GEN_368; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_370 = 10'h172 == _T_5[9:0] ? image_0_370 : _GEN_369; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_371 = 10'h173 == _T_5[9:0] ? image_0_371 : _GEN_370; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_372 = 10'h174 == _T_5[9:0] ? image_0_372 : _GEN_371; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_373 = 10'h175 == _T_5[9:0] ? image_0_373 : _GEN_372; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_374 = 10'h176 == _T_5[9:0] ? image_0_374 : _GEN_373; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_375 = 10'h177 == _T_5[9:0] ? image_0_375 : _GEN_374; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_376 = 10'h178 == _T_5[9:0] ? image_0_376 : _GEN_375; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_377 = 10'h179 == _T_5[9:0] ? image_0_377 : _GEN_376; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_378 = 10'h17a == _T_5[9:0] ? image_0_378 : _GEN_377; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_379 = 10'h17b == _T_5[9:0] ? image_0_379 : _GEN_378; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_380 = 10'h17c == _T_5[9:0] ? image_0_380 : _GEN_379; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_381 = 10'h17d == _T_5[9:0] ? image_0_381 : _GEN_380; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_382 = 10'h17e == _T_5[9:0] ? image_0_382 : _GEN_381; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_383 = 10'h17f == _T_5[9:0] ? image_0_383 : _GEN_382; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_384 = 10'h180 == _T_5[9:0] ? image_0_384 : _GEN_383; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_385 = 10'h181 == _T_5[9:0] ? image_0_385 : _GEN_384; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_386 = 10'h182 == _T_5[9:0] ? image_0_386 : _GEN_385; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_387 = 10'h183 == _T_5[9:0] ? image_0_387 : _GEN_386; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_388 = 10'h184 == _T_5[9:0] ? image_0_388 : _GEN_387; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_389 = 10'h185 == _T_5[9:0] ? image_0_389 : _GEN_388; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_390 = 10'h186 == _T_5[9:0] ? image_0_390 : _GEN_389; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_391 = 10'h187 == _T_5[9:0] ? image_0_391 : _GEN_390; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_392 = 10'h188 == _T_5[9:0] ? image_0_392 : _GEN_391; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_393 = 10'h189 == _T_5[9:0] ? image_0_393 : _GEN_392; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_394 = 10'h18a == _T_5[9:0] ? image_0_394 : _GEN_393; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_395 = 10'h18b == _T_5[9:0] ? image_0_395 : _GEN_394; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_396 = 10'h18c == _T_5[9:0] ? image_0_396 : _GEN_395; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_397 = 10'h18d == _T_5[9:0] ? image_0_397 : _GEN_396; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_398 = 10'h18e == _T_5[9:0] ? image_0_398 : _GEN_397; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_399 = 10'h18f == _T_5[9:0] ? image_0_399 : _GEN_398; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_400 = 10'h190 == _T_5[9:0] ? image_0_400 : _GEN_399; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_401 = 10'h191 == _T_5[9:0] ? image_0_401 : _GEN_400; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_402 = 10'h192 == _T_5[9:0] ? image_0_402 : _GEN_401; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_403 = 10'h193 == _T_5[9:0] ? image_0_403 : _GEN_402; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_404 = 10'h194 == _T_5[9:0] ? image_0_404 : _GEN_403; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_405 = 10'h195 == _T_5[9:0] ? image_0_405 : _GEN_404; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_406 = 10'h196 == _T_5[9:0] ? image_0_406 : _GEN_405; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_407 = 10'h197 == _T_5[9:0] ? image_0_407 : _GEN_406; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_408 = 10'h198 == _T_5[9:0] ? image_0_408 : _GEN_407; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_409 = 10'h199 == _T_5[9:0] ? image_0_409 : _GEN_408; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_410 = 10'h19a == _T_5[9:0] ? image_0_410 : _GEN_409; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_411 = 10'h19b == _T_5[9:0] ? image_0_411 : _GEN_410; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_412 = 10'h19c == _T_5[9:0] ? image_0_412 : _GEN_411; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_413 = 10'h19d == _T_5[9:0] ? image_0_413 : _GEN_412; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_414 = 10'h19e == _T_5[9:0] ? image_0_414 : _GEN_413; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_415 = 10'h19f == _T_5[9:0] ? image_0_415 : _GEN_414; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_416 = 10'h1a0 == _T_5[9:0] ? image_0_416 : _GEN_415; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_417 = 10'h1a1 == _T_5[9:0] ? image_0_417 : _GEN_416; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_418 = 10'h1a2 == _T_5[9:0] ? image_0_418 : _GEN_417; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_419 = 10'h1a3 == _T_5[9:0] ? image_0_419 : _GEN_418; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_420 = 10'h1a4 == _T_5[9:0] ? image_0_420 : _GEN_419; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_421 = 10'h1a5 == _T_5[9:0] ? image_0_421 : _GEN_420; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_422 = 10'h1a6 == _T_5[9:0] ? image_0_422 : _GEN_421; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_423 = 10'h1a7 == _T_5[9:0] ? image_0_423 : _GEN_422; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_424 = 10'h1a8 == _T_5[9:0] ? image_0_424 : _GEN_423; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_425 = 10'h1a9 == _T_5[9:0] ? image_0_425 : _GEN_424; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_426 = 10'h1aa == _T_5[9:0] ? image_0_426 : _GEN_425; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_427 = 10'h1ab == _T_5[9:0] ? image_0_427 : _GEN_426; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_428 = 10'h1ac == _T_5[9:0] ? image_0_428 : _GEN_427; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_429 = 10'h1ad == _T_5[9:0] ? image_0_429 : _GEN_428; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_430 = 10'h1ae == _T_5[9:0] ? image_0_430 : _GEN_429; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_431 = 10'h1af == _T_5[9:0] ? image_0_431 : _GEN_430; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_432 = 10'h1b0 == _T_5[9:0] ? image_0_432 : _GEN_431; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_433 = 10'h1b1 == _T_5[9:0] ? image_0_433 : _GEN_432; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_434 = 10'h1b2 == _T_5[9:0] ? image_0_434 : _GEN_433; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_435 = 10'h1b3 == _T_5[9:0] ? image_0_435 : _GEN_434; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_436 = 10'h1b4 == _T_5[9:0] ? image_0_436 : _GEN_435; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_437 = 10'h1b5 == _T_5[9:0] ? image_0_437 : _GEN_436; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_438 = 10'h1b6 == _T_5[9:0] ? image_0_438 : _GEN_437; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_439 = 10'h1b7 == _T_5[9:0] ? image_0_439 : _GEN_438; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_440 = 10'h1b8 == _T_5[9:0] ? image_0_440 : _GEN_439; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_441 = 10'h1b9 == _T_5[9:0] ? image_0_441 : _GEN_440; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_442 = 10'h1ba == _T_5[9:0] ? image_0_442 : _GEN_441; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_443 = 10'h1bb == _T_5[9:0] ? image_0_443 : _GEN_442; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_444 = 10'h1bc == _T_5[9:0] ? image_0_444 : _GEN_443; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_445 = 10'h1bd == _T_5[9:0] ? image_0_445 : _GEN_444; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_446 = 10'h1be == _T_5[9:0] ? image_0_446 : _GEN_445; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_447 = 10'h1bf == _T_5[9:0] ? image_0_447 : _GEN_446; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_448 = 10'h1c0 == _T_5[9:0] ? image_0_448 : _GEN_447; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_449 = 10'h1c1 == _T_5[9:0] ? image_0_449 : _GEN_448; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_450 = 10'h1c2 == _T_5[9:0] ? image_0_450 : _GEN_449; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_451 = 10'h1c3 == _T_5[9:0] ? image_0_451 : _GEN_450; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_452 = 10'h1c4 == _T_5[9:0] ? image_0_452 : _GEN_451; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_453 = 10'h1c5 == _T_5[9:0] ? image_0_453 : _GEN_452; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_454 = 10'h1c6 == _T_5[9:0] ? image_0_454 : _GEN_453; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_455 = 10'h1c7 == _T_5[9:0] ? image_0_455 : _GEN_454; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_456 = 10'h1c8 == _T_5[9:0] ? image_0_456 : _GEN_455; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_457 = 10'h1c9 == _T_5[9:0] ? image_0_457 : _GEN_456; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_458 = 10'h1ca == _T_5[9:0] ? image_0_458 : _GEN_457; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_459 = 10'h1cb == _T_5[9:0] ? image_0_459 : _GEN_458; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_460 = 10'h1cc == _T_5[9:0] ? image_0_460 : _GEN_459; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_461 = 10'h1cd == _T_5[9:0] ? image_0_461 : _GEN_460; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_462 = 10'h1ce == _T_5[9:0] ? image_0_462 : _GEN_461; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_463 = 10'h1cf == _T_5[9:0] ? image_0_463 : _GEN_462; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_464 = 10'h1d0 == _T_5[9:0] ? image_0_464 : _GEN_463; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_465 = 10'h1d1 == _T_5[9:0] ? image_0_465 : _GEN_464; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_466 = 10'h1d2 == _T_5[9:0] ? image_0_466 : _GEN_465; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_467 = 10'h1d3 == _T_5[9:0] ? image_0_467 : _GEN_466; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_468 = 10'h1d4 == _T_5[9:0] ? image_0_468 : _GEN_467; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_469 = 10'h1d5 == _T_5[9:0] ? image_0_469 : _GEN_468; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_470 = 10'h1d6 == _T_5[9:0] ? image_0_470 : _GEN_469; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_471 = 10'h1d7 == _T_5[9:0] ? image_0_471 : _GEN_470; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_472 = 10'h1d8 == _T_5[9:0] ? image_0_472 : _GEN_471; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_473 = 10'h1d9 == _T_5[9:0] ? image_0_473 : _GEN_472; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_474 = 10'h1da == _T_5[9:0] ? image_0_474 : _GEN_473; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_475 = 10'h1db == _T_5[9:0] ? image_0_475 : _GEN_474; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_476 = 10'h1dc == _T_5[9:0] ? image_0_476 : _GEN_475; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_477 = 10'h1dd == _T_5[9:0] ? image_0_477 : _GEN_476; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_478 = 10'h1de == _T_5[9:0] ? image_0_478 : _GEN_477; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_479 = 10'h1df == _T_5[9:0] ? image_0_479 : _GEN_478; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_480 = 10'h1e0 == _T_5[9:0] ? image_0_480 : _GEN_479; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_481 = 10'h1e1 == _T_5[9:0] ? image_0_481 : _GEN_480; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_482 = 10'h1e2 == _T_5[9:0] ? image_0_482 : _GEN_481; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_483 = 10'h1e3 == _T_5[9:0] ? image_0_483 : _GEN_482; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_484 = 10'h1e4 == _T_5[9:0] ? image_0_484 : _GEN_483; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_485 = 10'h1e5 == _T_5[9:0] ? image_0_485 : _GEN_484; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_486 = 10'h1e6 == _T_5[9:0] ? image_0_486 : _GEN_485; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_487 = 10'h1e7 == _T_5[9:0] ? image_0_487 : _GEN_486; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_488 = 10'h1e8 == _T_5[9:0] ? image_0_488 : _GEN_487; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_489 = 10'h1e9 == _T_5[9:0] ? image_0_489 : _GEN_488; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_490 = 10'h1ea == _T_5[9:0] ? image_0_490 : _GEN_489; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_491 = 10'h1eb == _T_5[9:0] ? image_0_491 : _GEN_490; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_492 = 10'h1ec == _T_5[9:0] ? image_0_492 : _GEN_491; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_493 = 10'h1ed == _T_5[9:0] ? image_0_493 : _GEN_492; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_494 = 10'h1ee == _T_5[9:0] ? image_0_494 : _GEN_493; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_495 = 10'h1ef == _T_5[9:0] ? image_0_495 : _GEN_494; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_496 = 10'h1f0 == _T_5[9:0] ? image_0_496 : _GEN_495; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_497 = 10'h1f1 == _T_5[9:0] ? image_0_497 : _GEN_496; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_498 = 10'h1f2 == _T_5[9:0] ? image_0_498 : _GEN_497; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_499 = 10'h1f3 == _T_5[9:0] ? image_0_499 : _GEN_498; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_500 = 10'h1f4 == _T_5[9:0] ? image_0_500 : _GEN_499; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_501 = 10'h1f5 == _T_5[9:0] ? image_0_501 : _GEN_500; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_502 = 10'h1f6 == _T_5[9:0] ? image_0_502 : _GEN_501; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_503 = 10'h1f7 == _T_5[9:0] ? image_0_503 : _GEN_502; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_504 = 10'h1f8 == _T_5[9:0] ? image_0_504 : _GEN_503; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_505 = 10'h1f9 == _T_5[9:0] ? image_0_505 : _GEN_504; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_506 = 10'h1fa == _T_5[9:0] ? image_0_506 : _GEN_505; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_507 = 10'h1fb == _T_5[9:0] ? image_0_507 : _GEN_506; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_508 = 10'h1fc == _T_5[9:0] ? image_0_508 : _GEN_507; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_509 = 10'h1fd == _T_5[9:0] ? image_0_509 : _GEN_508; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_510 = 10'h1fe == _T_5[9:0] ? image_0_510 : _GEN_509; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_511 = 10'h1ff == _T_5[9:0] ? image_0_511 : _GEN_510; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_512 = 10'h200 == _T_5[9:0] ? image_0_512 : _GEN_511; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_513 = 10'h201 == _T_5[9:0] ? image_0_513 : _GEN_512; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_514 = 10'h202 == _T_5[9:0] ? image_0_514 : _GEN_513; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_515 = 10'h203 == _T_5[9:0] ? image_0_515 : _GEN_514; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_516 = 10'h204 == _T_5[9:0] ? image_0_516 : _GEN_515; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_517 = 10'h205 == _T_5[9:0] ? image_0_517 : _GEN_516; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_518 = 10'h206 == _T_5[9:0] ? image_0_518 : _GEN_517; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_519 = 10'h207 == _T_5[9:0] ? image_0_519 : _GEN_518; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_520 = 10'h208 == _T_5[9:0] ? image_0_520 : _GEN_519; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_521 = 10'h209 == _T_5[9:0] ? image_0_521 : _GEN_520; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_522 = 10'h20a == _T_5[9:0] ? image_0_522 : _GEN_521; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_523 = 10'h20b == _T_5[9:0] ? image_0_523 : _GEN_522; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_524 = 10'h20c == _T_5[9:0] ? image_0_524 : _GEN_523; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_525 = 10'h20d == _T_5[9:0] ? image_0_525 : _GEN_524; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_526 = 10'h20e == _T_5[9:0] ? image_0_526 : _GEN_525; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_527 = 10'h20f == _T_5[9:0] ? image_0_527 : _GEN_526; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_528 = 10'h210 == _T_5[9:0] ? image_0_528 : _GEN_527; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_529 = 10'h211 == _T_5[9:0] ? image_0_529 : _GEN_528; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_530 = 10'h212 == _T_5[9:0] ? image_0_530 : _GEN_529; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_531 = 10'h213 == _T_5[9:0] ? image_0_531 : _GEN_530; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_532 = 10'h214 == _T_5[9:0] ? image_0_532 : _GEN_531; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_533 = 10'h215 == _T_5[9:0] ? image_0_533 : _GEN_532; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_534 = 10'h216 == _T_5[9:0] ? image_0_534 : _GEN_533; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_535 = 10'h217 == _T_5[9:0] ? image_0_535 : _GEN_534; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_536 = 10'h218 == _T_5[9:0] ? image_0_536 : _GEN_535; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_537 = 10'h219 == _T_5[9:0] ? image_0_537 : _GEN_536; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_538 = 10'h21a == _T_5[9:0] ? image_0_538 : _GEN_537; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_539 = 10'h21b == _T_5[9:0] ? image_0_539 : _GEN_538; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_540 = 10'h21c == _T_5[9:0] ? image_0_540 : _GEN_539; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_541 = 10'h21d == _T_5[9:0] ? image_0_541 : _GEN_540; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_542 = 10'h21e == _T_5[9:0] ? image_0_542 : _GEN_541; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_543 = 10'h21f == _T_5[9:0] ? image_0_543 : _GEN_542; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_544 = 10'h220 == _T_5[9:0] ? image_0_544 : _GEN_543; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_545 = 10'h221 == _T_5[9:0] ? image_0_545 : _GEN_544; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_546 = 10'h222 == _T_5[9:0] ? image_0_546 : _GEN_545; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_547 = 10'h223 == _T_5[9:0] ? image_0_547 : _GEN_546; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_548 = 10'h224 == _T_5[9:0] ? image_0_548 : _GEN_547; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_549 = 10'h225 == _T_5[9:0] ? image_0_549 : _GEN_548; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_550 = 10'h226 == _T_5[9:0] ? image_0_550 : _GEN_549; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_551 = 10'h227 == _T_5[9:0] ? image_0_551 : _GEN_550; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_552 = 10'h228 == _T_5[9:0] ? image_0_552 : _GEN_551; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_553 = 10'h229 == _T_5[9:0] ? image_0_553 : _GEN_552; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_554 = 10'h22a == _T_5[9:0] ? image_0_554 : _GEN_553; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_555 = 10'h22b == _T_5[9:0] ? image_0_555 : _GEN_554; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_556 = 10'h22c == _T_5[9:0] ? image_0_556 : _GEN_555; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_557 = 10'h22d == _T_5[9:0] ? image_0_557 : _GEN_556; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_558 = 10'h22e == _T_5[9:0] ? image_0_558 : _GEN_557; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_559 = 10'h22f == _T_5[9:0] ? image_0_559 : _GEN_558; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_560 = 10'h230 == _T_5[9:0] ? image_0_560 : _GEN_559; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_561 = 10'h231 == _T_5[9:0] ? image_0_561 : _GEN_560; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_562 = 10'h232 == _T_5[9:0] ? image_0_562 : _GEN_561; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_563 = 10'h233 == _T_5[9:0] ? image_0_563 : _GEN_562; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_564 = 10'h234 == _T_5[9:0] ? image_0_564 : _GEN_563; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_565 = 10'h235 == _T_5[9:0] ? image_0_565 : _GEN_564; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_566 = 10'h236 == _T_5[9:0] ? image_0_566 : _GEN_565; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_567 = 10'h237 == _T_5[9:0] ? image_0_567 : _GEN_566; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_568 = 10'h238 == _T_5[9:0] ? image_0_568 : _GEN_567; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_569 = 10'h239 == _T_5[9:0] ? image_0_569 : _GEN_568; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_570 = 10'h23a == _T_5[9:0] ? image_0_570 : _GEN_569; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_571 = 10'h23b == _T_5[9:0] ? image_0_571 : _GEN_570; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_572 = 10'h23c == _T_5[9:0] ? image_0_572 : _GEN_571; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_573 = 10'h23d == _T_5[9:0] ? image_0_573 : _GEN_572; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_574 = 10'h23e == _T_5[9:0] ? image_0_574 : _GEN_573; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_577 = 10'h1 == _T_5[9:0] ? image_1_1 : image_1_0; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_578 = 10'h2 == _T_5[9:0] ? image_1_2 : _GEN_577; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_579 = 10'h3 == _T_5[9:0] ? image_1_3 : _GEN_578; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_580 = 10'h4 == _T_5[9:0] ? image_1_4 : _GEN_579; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_581 = 10'h5 == _T_5[9:0] ? image_1_5 : _GEN_580; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_582 = 10'h6 == _T_5[9:0] ? image_1_6 : _GEN_581; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_583 = 10'h7 == _T_5[9:0] ? image_1_7 : _GEN_582; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_584 = 10'h8 == _T_5[9:0] ? image_1_8 : _GEN_583; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_585 = 10'h9 == _T_5[9:0] ? image_1_9 : _GEN_584; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_586 = 10'ha == _T_5[9:0] ? image_1_10 : _GEN_585; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_587 = 10'hb == _T_5[9:0] ? image_1_11 : _GEN_586; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_588 = 10'hc == _T_5[9:0] ? image_1_12 : _GEN_587; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_589 = 10'hd == _T_5[9:0] ? image_1_13 : _GEN_588; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_590 = 10'he == _T_5[9:0] ? image_1_14 : _GEN_589; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_591 = 10'hf == _T_5[9:0] ? image_1_15 : _GEN_590; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_592 = 10'h10 == _T_5[9:0] ? image_1_16 : _GEN_591; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_593 = 10'h11 == _T_5[9:0] ? image_1_17 : _GEN_592; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_594 = 10'h12 == _T_5[9:0] ? image_1_18 : _GEN_593; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_595 = 10'h13 == _T_5[9:0] ? image_1_19 : _GEN_594; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_596 = 10'h14 == _T_5[9:0] ? image_1_20 : _GEN_595; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_597 = 10'h15 == _T_5[9:0] ? image_1_21 : _GEN_596; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_598 = 10'h16 == _T_5[9:0] ? image_1_22 : _GEN_597; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_599 = 10'h17 == _T_5[9:0] ? image_1_23 : _GEN_598; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_600 = 10'h18 == _T_5[9:0] ? image_1_24 : _GEN_599; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_601 = 10'h19 == _T_5[9:0] ? image_1_25 : _GEN_600; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_602 = 10'h1a == _T_5[9:0] ? image_1_26 : _GEN_601; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_603 = 10'h1b == _T_5[9:0] ? image_1_27 : _GEN_602; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_604 = 10'h1c == _T_5[9:0] ? image_1_28 : _GEN_603; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_605 = 10'h1d == _T_5[9:0] ? image_1_29 : _GEN_604; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_606 = 10'h1e == _T_5[9:0] ? image_1_30 : _GEN_605; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_607 = 10'h1f == _T_5[9:0] ? image_1_31 : _GEN_606; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_608 = 10'h20 == _T_5[9:0] ? image_1_32 : _GEN_607; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_609 = 10'h21 == _T_5[9:0] ? image_1_33 : _GEN_608; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_610 = 10'h22 == _T_5[9:0] ? image_1_34 : _GEN_609; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_611 = 10'h23 == _T_5[9:0] ? image_1_35 : _GEN_610; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_612 = 10'h24 == _T_5[9:0] ? image_1_36 : _GEN_611; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_613 = 10'h25 == _T_5[9:0] ? image_1_37 : _GEN_612; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_614 = 10'h26 == _T_5[9:0] ? image_1_38 : _GEN_613; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_615 = 10'h27 == _T_5[9:0] ? image_1_39 : _GEN_614; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_616 = 10'h28 == _T_5[9:0] ? image_1_40 : _GEN_615; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_617 = 10'h29 == _T_5[9:0] ? image_1_41 : _GEN_616; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_618 = 10'h2a == _T_5[9:0] ? image_1_42 : _GEN_617; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_619 = 10'h2b == _T_5[9:0] ? image_1_43 : _GEN_618; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_620 = 10'h2c == _T_5[9:0] ? image_1_44 : _GEN_619; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_621 = 10'h2d == _T_5[9:0] ? image_1_45 : _GEN_620; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_622 = 10'h2e == _T_5[9:0] ? image_1_46 : _GEN_621; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_623 = 10'h2f == _T_5[9:0] ? image_1_47 : _GEN_622; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_624 = 10'h30 == _T_5[9:0] ? image_1_48 : _GEN_623; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_625 = 10'h31 == _T_5[9:0] ? image_1_49 : _GEN_624; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_626 = 10'h32 == _T_5[9:0] ? image_1_50 : _GEN_625; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_627 = 10'h33 == _T_5[9:0] ? image_1_51 : _GEN_626; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_628 = 10'h34 == _T_5[9:0] ? image_1_52 : _GEN_627; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_629 = 10'h35 == _T_5[9:0] ? image_1_53 : _GEN_628; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_630 = 10'h36 == _T_5[9:0] ? image_1_54 : _GEN_629; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_631 = 10'h37 == _T_5[9:0] ? image_1_55 : _GEN_630; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_632 = 10'h38 == _T_5[9:0] ? image_1_56 : _GEN_631; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_633 = 10'h39 == _T_5[9:0] ? image_1_57 : _GEN_632; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_634 = 10'h3a == _T_5[9:0] ? image_1_58 : _GEN_633; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_635 = 10'h3b == _T_5[9:0] ? image_1_59 : _GEN_634; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_636 = 10'h3c == _T_5[9:0] ? image_1_60 : _GEN_635; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_637 = 10'h3d == _T_5[9:0] ? image_1_61 : _GEN_636; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_638 = 10'h3e == _T_5[9:0] ? image_1_62 : _GEN_637; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_639 = 10'h3f == _T_5[9:0] ? image_1_63 : _GEN_638; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_640 = 10'h40 == _T_5[9:0] ? image_1_64 : _GEN_639; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_641 = 10'h41 == _T_5[9:0] ? image_1_65 : _GEN_640; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_642 = 10'h42 == _T_5[9:0] ? image_1_66 : _GEN_641; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_643 = 10'h43 == _T_5[9:0] ? image_1_67 : _GEN_642; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_644 = 10'h44 == _T_5[9:0] ? image_1_68 : _GEN_643; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_645 = 10'h45 == _T_5[9:0] ? image_1_69 : _GEN_644; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_646 = 10'h46 == _T_5[9:0] ? image_1_70 : _GEN_645; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_647 = 10'h47 == _T_5[9:0] ? image_1_71 : _GEN_646; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_648 = 10'h48 == _T_5[9:0] ? image_1_72 : _GEN_647; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_649 = 10'h49 == _T_5[9:0] ? image_1_73 : _GEN_648; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_650 = 10'h4a == _T_5[9:0] ? image_1_74 : _GEN_649; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_651 = 10'h4b == _T_5[9:0] ? image_1_75 : _GEN_650; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_652 = 10'h4c == _T_5[9:0] ? image_1_76 : _GEN_651; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_653 = 10'h4d == _T_5[9:0] ? image_1_77 : _GEN_652; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_654 = 10'h4e == _T_5[9:0] ? image_1_78 : _GEN_653; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_655 = 10'h4f == _T_5[9:0] ? image_1_79 : _GEN_654; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_656 = 10'h50 == _T_5[9:0] ? image_1_80 : _GEN_655; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_657 = 10'h51 == _T_5[9:0] ? image_1_81 : _GEN_656; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_658 = 10'h52 == _T_5[9:0] ? image_1_82 : _GEN_657; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_659 = 10'h53 == _T_5[9:0] ? image_1_83 : _GEN_658; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_660 = 10'h54 == _T_5[9:0] ? image_1_84 : _GEN_659; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_661 = 10'h55 == _T_5[9:0] ? image_1_85 : _GEN_660; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_662 = 10'h56 == _T_5[9:0] ? image_1_86 : _GEN_661; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_663 = 10'h57 == _T_5[9:0] ? image_1_87 : _GEN_662; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_664 = 10'h58 == _T_5[9:0] ? image_1_88 : _GEN_663; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_665 = 10'h59 == _T_5[9:0] ? image_1_89 : _GEN_664; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_666 = 10'h5a == _T_5[9:0] ? image_1_90 : _GEN_665; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_667 = 10'h5b == _T_5[9:0] ? image_1_91 : _GEN_666; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_668 = 10'h5c == _T_5[9:0] ? image_1_92 : _GEN_667; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_669 = 10'h5d == _T_5[9:0] ? image_1_93 : _GEN_668; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_670 = 10'h5e == _T_5[9:0] ? image_1_94 : _GEN_669; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_671 = 10'h5f == _T_5[9:0] ? image_1_95 : _GEN_670; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_672 = 10'h60 == _T_5[9:0] ? image_1_96 : _GEN_671; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_673 = 10'h61 == _T_5[9:0] ? image_1_97 : _GEN_672; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_674 = 10'h62 == _T_5[9:0] ? image_1_98 : _GEN_673; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_675 = 10'h63 == _T_5[9:0] ? image_1_99 : _GEN_674; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_676 = 10'h64 == _T_5[9:0] ? image_1_100 : _GEN_675; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_677 = 10'h65 == _T_5[9:0] ? image_1_101 : _GEN_676; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_678 = 10'h66 == _T_5[9:0] ? image_1_102 : _GEN_677; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_679 = 10'h67 == _T_5[9:0] ? image_1_103 : _GEN_678; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_680 = 10'h68 == _T_5[9:0] ? image_1_104 : _GEN_679; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_681 = 10'h69 == _T_5[9:0] ? image_1_105 : _GEN_680; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_682 = 10'h6a == _T_5[9:0] ? image_1_106 : _GEN_681; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_683 = 10'h6b == _T_5[9:0] ? image_1_107 : _GEN_682; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_684 = 10'h6c == _T_5[9:0] ? image_1_108 : _GEN_683; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_685 = 10'h6d == _T_5[9:0] ? image_1_109 : _GEN_684; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_686 = 10'h6e == _T_5[9:0] ? image_1_110 : _GEN_685; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_687 = 10'h6f == _T_5[9:0] ? image_1_111 : _GEN_686; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_688 = 10'h70 == _T_5[9:0] ? image_1_112 : _GEN_687; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_689 = 10'h71 == _T_5[9:0] ? image_1_113 : _GEN_688; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_690 = 10'h72 == _T_5[9:0] ? image_1_114 : _GEN_689; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_691 = 10'h73 == _T_5[9:0] ? image_1_115 : _GEN_690; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_692 = 10'h74 == _T_5[9:0] ? image_1_116 : _GEN_691; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_693 = 10'h75 == _T_5[9:0] ? image_1_117 : _GEN_692; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_694 = 10'h76 == _T_5[9:0] ? image_1_118 : _GEN_693; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_695 = 10'h77 == _T_5[9:0] ? image_1_119 : _GEN_694; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_696 = 10'h78 == _T_5[9:0] ? image_1_120 : _GEN_695; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_697 = 10'h79 == _T_5[9:0] ? image_1_121 : _GEN_696; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_698 = 10'h7a == _T_5[9:0] ? image_1_122 : _GEN_697; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_699 = 10'h7b == _T_5[9:0] ? image_1_123 : _GEN_698; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_700 = 10'h7c == _T_5[9:0] ? image_1_124 : _GEN_699; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_701 = 10'h7d == _T_5[9:0] ? image_1_125 : _GEN_700; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_702 = 10'h7e == _T_5[9:0] ? image_1_126 : _GEN_701; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_703 = 10'h7f == _T_5[9:0] ? image_1_127 : _GEN_702; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_704 = 10'h80 == _T_5[9:0] ? image_1_128 : _GEN_703; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_705 = 10'h81 == _T_5[9:0] ? image_1_129 : _GEN_704; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_706 = 10'h82 == _T_5[9:0] ? image_1_130 : _GEN_705; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_707 = 10'h83 == _T_5[9:0] ? image_1_131 : _GEN_706; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_708 = 10'h84 == _T_5[9:0] ? image_1_132 : _GEN_707; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_709 = 10'h85 == _T_5[9:0] ? image_1_133 : _GEN_708; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_710 = 10'h86 == _T_5[9:0] ? image_1_134 : _GEN_709; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_711 = 10'h87 == _T_5[9:0] ? image_1_135 : _GEN_710; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_712 = 10'h88 == _T_5[9:0] ? image_1_136 : _GEN_711; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_713 = 10'h89 == _T_5[9:0] ? image_1_137 : _GEN_712; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_714 = 10'h8a == _T_5[9:0] ? image_1_138 : _GEN_713; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_715 = 10'h8b == _T_5[9:0] ? image_1_139 : _GEN_714; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_716 = 10'h8c == _T_5[9:0] ? image_1_140 : _GEN_715; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_717 = 10'h8d == _T_5[9:0] ? image_1_141 : _GEN_716; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_718 = 10'h8e == _T_5[9:0] ? image_1_142 : _GEN_717; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_719 = 10'h8f == _T_5[9:0] ? image_1_143 : _GEN_718; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_720 = 10'h90 == _T_5[9:0] ? image_1_144 : _GEN_719; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_721 = 10'h91 == _T_5[9:0] ? image_1_145 : _GEN_720; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_722 = 10'h92 == _T_5[9:0] ? image_1_146 : _GEN_721; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_723 = 10'h93 == _T_5[9:0] ? image_1_147 : _GEN_722; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_724 = 10'h94 == _T_5[9:0] ? image_1_148 : _GEN_723; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_725 = 10'h95 == _T_5[9:0] ? image_1_149 : _GEN_724; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_726 = 10'h96 == _T_5[9:0] ? image_1_150 : _GEN_725; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_727 = 10'h97 == _T_5[9:0] ? image_1_151 : _GEN_726; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_728 = 10'h98 == _T_5[9:0] ? image_1_152 : _GEN_727; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_729 = 10'h99 == _T_5[9:0] ? image_1_153 : _GEN_728; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_730 = 10'h9a == _T_5[9:0] ? image_1_154 : _GEN_729; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_731 = 10'h9b == _T_5[9:0] ? image_1_155 : _GEN_730; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_732 = 10'h9c == _T_5[9:0] ? image_1_156 : _GEN_731; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_733 = 10'h9d == _T_5[9:0] ? image_1_157 : _GEN_732; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_734 = 10'h9e == _T_5[9:0] ? image_1_158 : _GEN_733; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_735 = 10'h9f == _T_5[9:0] ? image_1_159 : _GEN_734; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_736 = 10'ha0 == _T_5[9:0] ? image_1_160 : _GEN_735; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_737 = 10'ha1 == _T_5[9:0] ? image_1_161 : _GEN_736; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_738 = 10'ha2 == _T_5[9:0] ? image_1_162 : _GEN_737; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_739 = 10'ha3 == _T_5[9:0] ? image_1_163 : _GEN_738; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_740 = 10'ha4 == _T_5[9:0] ? image_1_164 : _GEN_739; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_741 = 10'ha5 == _T_5[9:0] ? image_1_165 : _GEN_740; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_742 = 10'ha6 == _T_5[9:0] ? image_1_166 : _GEN_741; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_743 = 10'ha7 == _T_5[9:0] ? image_1_167 : _GEN_742; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_744 = 10'ha8 == _T_5[9:0] ? image_1_168 : _GEN_743; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_745 = 10'ha9 == _T_5[9:0] ? image_1_169 : _GEN_744; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_746 = 10'haa == _T_5[9:0] ? image_1_170 : _GEN_745; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_747 = 10'hab == _T_5[9:0] ? image_1_171 : _GEN_746; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_748 = 10'hac == _T_5[9:0] ? image_1_172 : _GEN_747; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_749 = 10'had == _T_5[9:0] ? image_1_173 : _GEN_748; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_750 = 10'hae == _T_5[9:0] ? image_1_174 : _GEN_749; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_751 = 10'haf == _T_5[9:0] ? image_1_175 : _GEN_750; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_752 = 10'hb0 == _T_5[9:0] ? image_1_176 : _GEN_751; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_753 = 10'hb1 == _T_5[9:0] ? image_1_177 : _GEN_752; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_754 = 10'hb2 == _T_5[9:0] ? image_1_178 : _GEN_753; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_755 = 10'hb3 == _T_5[9:0] ? image_1_179 : _GEN_754; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_756 = 10'hb4 == _T_5[9:0] ? image_1_180 : _GEN_755; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_757 = 10'hb5 == _T_5[9:0] ? image_1_181 : _GEN_756; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_758 = 10'hb6 == _T_5[9:0] ? image_1_182 : _GEN_757; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_759 = 10'hb7 == _T_5[9:0] ? image_1_183 : _GEN_758; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_760 = 10'hb8 == _T_5[9:0] ? image_1_184 : _GEN_759; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_761 = 10'hb9 == _T_5[9:0] ? image_1_185 : _GEN_760; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_762 = 10'hba == _T_5[9:0] ? image_1_186 : _GEN_761; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_763 = 10'hbb == _T_5[9:0] ? image_1_187 : _GEN_762; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_764 = 10'hbc == _T_5[9:0] ? image_1_188 : _GEN_763; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_765 = 10'hbd == _T_5[9:0] ? image_1_189 : _GEN_764; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_766 = 10'hbe == _T_5[9:0] ? image_1_190 : _GEN_765; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_767 = 10'hbf == _T_5[9:0] ? image_1_191 : _GEN_766; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_768 = 10'hc0 == _T_5[9:0] ? image_1_192 : _GEN_767; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_769 = 10'hc1 == _T_5[9:0] ? image_1_193 : _GEN_768; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_770 = 10'hc2 == _T_5[9:0] ? image_1_194 : _GEN_769; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_771 = 10'hc3 == _T_5[9:0] ? image_1_195 : _GEN_770; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_772 = 10'hc4 == _T_5[9:0] ? image_1_196 : _GEN_771; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_773 = 10'hc5 == _T_5[9:0] ? image_1_197 : _GEN_772; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_774 = 10'hc6 == _T_5[9:0] ? image_1_198 : _GEN_773; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_775 = 10'hc7 == _T_5[9:0] ? image_1_199 : _GEN_774; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_776 = 10'hc8 == _T_5[9:0] ? image_1_200 : _GEN_775; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_777 = 10'hc9 == _T_5[9:0] ? image_1_201 : _GEN_776; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_778 = 10'hca == _T_5[9:0] ? image_1_202 : _GEN_777; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_779 = 10'hcb == _T_5[9:0] ? image_1_203 : _GEN_778; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_780 = 10'hcc == _T_5[9:0] ? image_1_204 : _GEN_779; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_781 = 10'hcd == _T_5[9:0] ? image_1_205 : _GEN_780; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_782 = 10'hce == _T_5[9:0] ? image_1_206 : _GEN_781; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_783 = 10'hcf == _T_5[9:0] ? image_1_207 : _GEN_782; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_784 = 10'hd0 == _T_5[9:0] ? image_1_208 : _GEN_783; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_785 = 10'hd1 == _T_5[9:0] ? image_1_209 : _GEN_784; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_786 = 10'hd2 == _T_5[9:0] ? image_1_210 : _GEN_785; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_787 = 10'hd3 == _T_5[9:0] ? image_1_211 : _GEN_786; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_788 = 10'hd4 == _T_5[9:0] ? image_1_212 : _GEN_787; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_789 = 10'hd5 == _T_5[9:0] ? image_1_213 : _GEN_788; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_790 = 10'hd6 == _T_5[9:0] ? image_1_214 : _GEN_789; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_791 = 10'hd7 == _T_5[9:0] ? image_1_215 : _GEN_790; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_792 = 10'hd8 == _T_5[9:0] ? image_1_216 : _GEN_791; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_793 = 10'hd9 == _T_5[9:0] ? image_1_217 : _GEN_792; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_794 = 10'hda == _T_5[9:0] ? image_1_218 : _GEN_793; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_795 = 10'hdb == _T_5[9:0] ? image_1_219 : _GEN_794; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_796 = 10'hdc == _T_5[9:0] ? image_1_220 : _GEN_795; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_797 = 10'hdd == _T_5[9:0] ? image_1_221 : _GEN_796; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_798 = 10'hde == _T_5[9:0] ? image_1_222 : _GEN_797; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_799 = 10'hdf == _T_5[9:0] ? image_1_223 : _GEN_798; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_800 = 10'he0 == _T_5[9:0] ? image_1_224 : _GEN_799; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_801 = 10'he1 == _T_5[9:0] ? image_1_225 : _GEN_800; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_802 = 10'he2 == _T_5[9:0] ? image_1_226 : _GEN_801; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_803 = 10'he3 == _T_5[9:0] ? image_1_227 : _GEN_802; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_804 = 10'he4 == _T_5[9:0] ? image_1_228 : _GEN_803; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_805 = 10'he5 == _T_5[9:0] ? image_1_229 : _GEN_804; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_806 = 10'he6 == _T_5[9:0] ? image_1_230 : _GEN_805; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_807 = 10'he7 == _T_5[9:0] ? image_1_231 : _GEN_806; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_808 = 10'he8 == _T_5[9:0] ? image_1_232 : _GEN_807; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_809 = 10'he9 == _T_5[9:0] ? image_1_233 : _GEN_808; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_810 = 10'hea == _T_5[9:0] ? image_1_234 : _GEN_809; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_811 = 10'heb == _T_5[9:0] ? image_1_235 : _GEN_810; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_812 = 10'hec == _T_5[9:0] ? image_1_236 : _GEN_811; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_813 = 10'hed == _T_5[9:0] ? image_1_237 : _GEN_812; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_814 = 10'hee == _T_5[9:0] ? image_1_238 : _GEN_813; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_815 = 10'hef == _T_5[9:0] ? image_1_239 : _GEN_814; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_816 = 10'hf0 == _T_5[9:0] ? image_1_240 : _GEN_815; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_817 = 10'hf1 == _T_5[9:0] ? image_1_241 : _GEN_816; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_818 = 10'hf2 == _T_5[9:0] ? image_1_242 : _GEN_817; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_819 = 10'hf3 == _T_5[9:0] ? image_1_243 : _GEN_818; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_820 = 10'hf4 == _T_5[9:0] ? image_1_244 : _GEN_819; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_821 = 10'hf5 == _T_5[9:0] ? image_1_245 : _GEN_820; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_822 = 10'hf6 == _T_5[9:0] ? image_1_246 : _GEN_821; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_823 = 10'hf7 == _T_5[9:0] ? image_1_247 : _GEN_822; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_824 = 10'hf8 == _T_5[9:0] ? image_1_248 : _GEN_823; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_825 = 10'hf9 == _T_5[9:0] ? image_1_249 : _GEN_824; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_826 = 10'hfa == _T_5[9:0] ? image_1_250 : _GEN_825; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_827 = 10'hfb == _T_5[9:0] ? image_1_251 : _GEN_826; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_828 = 10'hfc == _T_5[9:0] ? image_1_252 : _GEN_827; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_829 = 10'hfd == _T_5[9:0] ? image_1_253 : _GEN_828; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_830 = 10'hfe == _T_5[9:0] ? image_1_254 : _GEN_829; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_831 = 10'hff == _T_5[9:0] ? image_1_255 : _GEN_830; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_832 = 10'h100 == _T_5[9:0] ? image_1_256 : _GEN_831; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_833 = 10'h101 == _T_5[9:0] ? image_1_257 : _GEN_832; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_834 = 10'h102 == _T_5[9:0] ? image_1_258 : _GEN_833; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_835 = 10'h103 == _T_5[9:0] ? image_1_259 : _GEN_834; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_836 = 10'h104 == _T_5[9:0] ? image_1_260 : _GEN_835; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_837 = 10'h105 == _T_5[9:0] ? image_1_261 : _GEN_836; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_838 = 10'h106 == _T_5[9:0] ? image_1_262 : _GEN_837; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_839 = 10'h107 == _T_5[9:0] ? image_1_263 : _GEN_838; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_840 = 10'h108 == _T_5[9:0] ? image_1_264 : _GEN_839; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_841 = 10'h109 == _T_5[9:0] ? image_1_265 : _GEN_840; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_842 = 10'h10a == _T_5[9:0] ? image_1_266 : _GEN_841; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_843 = 10'h10b == _T_5[9:0] ? image_1_267 : _GEN_842; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_844 = 10'h10c == _T_5[9:0] ? image_1_268 : _GEN_843; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_845 = 10'h10d == _T_5[9:0] ? image_1_269 : _GEN_844; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_846 = 10'h10e == _T_5[9:0] ? image_1_270 : _GEN_845; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_847 = 10'h10f == _T_5[9:0] ? image_1_271 : _GEN_846; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_848 = 10'h110 == _T_5[9:0] ? image_1_272 : _GEN_847; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_849 = 10'h111 == _T_5[9:0] ? image_1_273 : _GEN_848; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_850 = 10'h112 == _T_5[9:0] ? image_1_274 : _GEN_849; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_851 = 10'h113 == _T_5[9:0] ? image_1_275 : _GEN_850; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_852 = 10'h114 == _T_5[9:0] ? image_1_276 : _GEN_851; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_853 = 10'h115 == _T_5[9:0] ? image_1_277 : _GEN_852; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_854 = 10'h116 == _T_5[9:0] ? image_1_278 : _GEN_853; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_855 = 10'h117 == _T_5[9:0] ? image_1_279 : _GEN_854; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_856 = 10'h118 == _T_5[9:0] ? image_1_280 : _GEN_855; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_857 = 10'h119 == _T_5[9:0] ? image_1_281 : _GEN_856; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_858 = 10'h11a == _T_5[9:0] ? image_1_282 : _GEN_857; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_859 = 10'h11b == _T_5[9:0] ? image_1_283 : _GEN_858; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_860 = 10'h11c == _T_5[9:0] ? image_1_284 : _GEN_859; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_861 = 10'h11d == _T_5[9:0] ? image_1_285 : _GEN_860; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_862 = 10'h11e == _T_5[9:0] ? image_1_286 : _GEN_861; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_863 = 10'h11f == _T_5[9:0] ? image_1_287 : _GEN_862; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_864 = 10'h120 == _T_5[9:0] ? image_1_288 : _GEN_863; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_865 = 10'h121 == _T_5[9:0] ? image_1_289 : _GEN_864; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_866 = 10'h122 == _T_5[9:0] ? image_1_290 : _GEN_865; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_867 = 10'h123 == _T_5[9:0] ? image_1_291 : _GEN_866; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_868 = 10'h124 == _T_5[9:0] ? image_1_292 : _GEN_867; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_869 = 10'h125 == _T_5[9:0] ? image_1_293 : _GEN_868; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_870 = 10'h126 == _T_5[9:0] ? image_1_294 : _GEN_869; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_871 = 10'h127 == _T_5[9:0] ? image_1_295 : _GEN_870; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_872 = 10'h128 == _T_5[9:0] ? image_1_296 : _GEN_871; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_873 = 10'h129 == _T_5[9:0] ? image_1_297 : _GEN_872; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_874 = 10'h12a == _T_5[9:0] ? image_1_298 : _GEN_873; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_875 = 10'h12b == _T_5[9:0] ? image_1_299 : _GEN_874; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_876 = 10'h12c == _T_5[9:0] ? image_1_300 : _GEN_875; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_877 = 10'h12d == _T_5[9:0] ? image_1_301 : _GEN_876; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_878 = 10'h12e == _T_5[9:0] ? image_1_302 : _GEN_877; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_879 = 10'h12f == _T_5[9:0] ? image_1_303 : _GEN_878; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_880 = 10'h130 == _T_5[9:0] ? image_1_304 : _GEN_879; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_881 = 10'h131 == _T_5[9:0] ? image_1_305 : _GEN_880; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_882 = 10'h132 == _T_5[9:0] ? image_1_306 : _GEN_881; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_883 = 10'h133 == _T_5[9:0] ? image_1_307 : _GEN_882; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_884 = 10'h134 == _T_5[9:0] ? image_1_308 : _GEN_883; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_885 = 10'h135 == _T_5[9:0] ? image_1_309 : _GEN_884; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_886 = 10'h136 == _T_5[9:0] ? image_1_310 : _GEN_885; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_887 = 10'h137 == _T_5[9:0] ? image_1_311 : _GEN_886; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_888 = 10'h138 == _T_5[9:0] ? image_1_312 : _GEN_887; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_889 = 10'h139 == _T_5[9:0] ? image_1_313 : _GEN_888; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_890 = 10'h13a == _T_5[9:0] ? image_1_314 : _GEN_889; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_891 = 10'h13b == _T_5[9:0] ? image_1_315 : _GEN_890; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_892 = 10'h13c == _T_5[9:0] ? image_1_316 : _GEN_891; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_893 = 10'h13d == _T_5[9:0] ? image_1_317 : _GEN_892; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_894 = 10'h13e == _T_5[9:0] ? image_1_318 : _GEN_893; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_895 = 10'h13f == _T_5[9:0] ? image_1_319 : _GEN_894; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_896 = 10'h140 == _T_5[9:0] ? image_1_320 : _GEN_895; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_897 = 10'h141 == _T_5[9:0] ? image_1_321 : _GEN_896; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_898 = 10'h142 == _T_5[9:0] ? image_1_322 : _GEN_897; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_899 = 10'h143 == _T_5[9:0] ? image_1_323 : _GEN_898; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_900 = 10'h144 == _T_5[9:0] ? image_1_324 : _GEN_899; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_901 = 10'h145 == _T_5[9:0] ? image_1_325 : _GEN_900; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_902 = 10'h146 == _T_5[9:0] ? image_1_326 : _GEN_901; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_903 = 10'h147 == _T_5[9:0] ? image_1_327 : _GEN_902; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_904 = 10'h148 == _T_5[9:0] ? image_1_328 : _GEN_903; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_905 = 10'h149 == _T_5[9:0] ? image_1_329 : _GEN_904; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_906 = 10'h14a == _T_5[9:0] ? image_1_330 : _GEN_905; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_907 = 10'h14b == _T_5[9:0] ? image_1_331 : _GEN_906; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_908 = 10'h14c == _T_5[9:0] ? image_1_332 : _GEN_907; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_909 = 10'h14d == _T_5[9:0] ? image_1_333 : _GEN_908; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_910 = 10'h14e == _T_5[9:0] ? image_1_334 : _GEN_909; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_911 = 10'h14f == _T_5[9:0] ? image_1_335 : _GEN_910; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_912 = 10'h150 == _T_5[9:0] ? image_1_336 : _GEN_911; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_913 = 10'h151 == _T_5[9:0] ? image_1_337 : _GEN_912; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_914 = 10'h152 == _T_5[9:0] ? image_1_338 : _GEN_913; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_915 = 10'h153 == _T_5[9:0] ? image_1_339 : _GEN_914; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_916 = 10'h154 == _T_5[9:0] ? image_1_340 : _GEN_915; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_917 = 10'h155 == _T_5[9:0] ? image_1_341 : _GEN_916; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_918 = 10'h156 == _T_5[9:0] ? image_1_342 : _GEN_917; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_919 = 10'h157 == _T_5[9:0] ? image_1_343 : _GEN_918; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_920 = 10'h158 == _T_5[9:0] ? image_1_344 : _GEN_919; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_921 = 10'h159 == _T_5[9:0] ? image_1_345 : _GEN_920; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_922 = 10'h15a == _T_5[9:0] ? image_1_346 : _GEN_921; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_923 = 10'h15b == _T_5[9:0] ? image_1_347 : _GEN_922; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_924 = 10'h15c == _T_5[9:0] ? image_1_348 : _GEN_923; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_925 = 10'h15d == _T_5[9:0] ? image_1_349 : _GEN_924; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_926 = 10'h15e == _T_5[9:0] ? image_1_350 : _GEN_925; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_927 = 10'h15f == _T_5[9:0] ? image_1_351 : _GEN_926; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_928 = 10'h160 == _T_5[9:0] ? image_1_352 : _GEN_927; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_929 = 10'h161 == _T_5[9:0] ? image_1_353 : _GEN_928; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_930 = 10'h162 == _T_5[9:0] ? image_1_354 : _GEN_929; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_931 = 10'h163 == _T_5[9:0] ? image_1_355 : _GEN_930; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_932 = 10'h164 == _T_5[9:0] ? image_1_356 : _GEN_931; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_933 = 10'h165 == _T_5[9:0] ? image_1_357 : _GEN_932; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_934 = 10'h166 == _T_5[9:0] ? image_1_358 : _GEN_933; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_935 = 10'h167 == _T_5[9:0] ? image_1_359 : _GEN_934; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_936 = 10'h168 == _T_5[9:0] ? image_1_360 : _GEN_935; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_937 = 10'h169 == _T_5[9:0] ? image_1_361 : _GEN_936; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_938 = 10'h16a == _T_5[9:0] ? image_1_362 : _GEN_937; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_939 = 10'h16b == _T_5[9:0] ? image_1_363 : _GEN_938; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_940 = 10'h16c == _T_5[9:0] ? image_1_364 : _GEN_939; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_941 = 10'h16d == _T_5[9:0] ? image_1_365 : _GEN_940; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_942 = 10'h16e == _T_5[9:0] ? image_1_366 : _GEN_941; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_943 = 10'h16f == _T_5[9:0] ? image_1_367 : _GEN_942; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_944 = 10'h170 == _T_5[9:0] ? image_1_368 : _GEN_943; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_945 = 10'h171 == _T_5[9:0] ? image_1_369 : _GEN_944; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_946 = 10'h172 == _T_5[9:0] ? image_1_370 : _GEN_945; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_947 = 10'h173 == _T_5[9:0] ? image_1_371 : _GEN_946; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_948 = 10'h174 == _T_5[9:0] ? image_1_372 : _GEN_947; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_949 = 10'h175 == _T_5[9:0] ? image_1_373 : _GEN_948; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_950 = 10'h176 == _T_5[9:0] ? image_1_374 : _GEN_949; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_951 = 10'h177 == _T_5[9:0] ? image_1_375 : _GEN_950; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_952 = 10'h178 == _T_5[9:0] ? image_1_376 : _GEN_951; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_953 = 10'h179 == _T_5[9:0] ? image_1_377 : _GEN_952; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_954 = 10'h17a == _T_5[9:0] ? image_1_378 : _GEN_953; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_955 = 10'h17b == _T_5[9:0] ? image_1_379 : _GEN_954; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_956 = 10'h17c == _T_5[9:0] ? image_1_380 : _GEN_955; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_957 = 10'h17d == _T_5[9:0] ? image_1_381 : _GEN_956; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_958 = 10'h17e == _T_5[9:0] ? image_1_382 : _GEN_957; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_959 = 10'h17f == _T_5[9:0] ? image_1_383 : _GEN_958; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_960 = 10'h180 == _T_5[9:0] ? image_1_384 : _GEN_959; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_961 = 10'h181 == _T_5[9:0] ? image_1_385 : _GEN_960; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_962 = 10'h182 == _T_5[9:0] ? image_1_386 : _GEN_961; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_963 = 10'h183 == _T_5[9:0] ? image_1_387 : _GEN_962; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_964 = 10'h184 == _T_5[9:0] ? image_1_388 : _GEN_963; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_965 = 10'h185 == _T_5[9:0] ? image_1_389 : _GEN_964; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_966 = 10'h186 == _T_5[9:0] ? image_1_390 : _GEN_965; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_967 = 10'h187 == _T_5[9:0] ? image_1_391 : _GEN_966; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_968 = 10'h188 == _T_5[9:0] ? image_1_392 : _GEN_967; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_969 = 10'h189 == _T_5[9:0] ? image_1_393 : _GEN_968; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_970 = 10'h18a == _T_5[9:0] ? image_1_394 : _GEN_969; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_971 = 10'h18b == _T_5[9:0] ? image_1_395 : _GEN_970; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_972 = 10'h18c == _T_5[9:0] ? image_1_396 : _GEN_971; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_973 = 10'h18d == _T_5[9:0] ? image_1_397 : _GEN_972; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_974 = 10'h18e == _T_5[9:0] ? image_1_398 : _GEN_973; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_975 = 10'h18f == _T_5[9:0] ? image_1_399 : _GEN_974; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_976 = 10'h190 == _T_5[9:0] ? image_1_400 : _GEN_975; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_977 = 10'h191 == _T_5[9:0] ? image_1_401 : _GEN_976; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_978 = 10'h192 == _T_5[9:0] ? image_1_402 : _GEN_977; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_979 = 10'h193 == _T_5[9:0] ? image_1_403 : _GEN_978; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_980 = 10'h194 == _T_5[9:0] ? image_1_404 : _GEN_979; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_981 = 10'h195 == _T_5[9:0] ? image_1_405 : _GEN_980; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_982 = 10'h196 == _T_5[9:0] ? image_1_406 : _GEN_981; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_983 = 10'h197 == _T_5[9:0] ? image_1_407 : _GEN_982; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_984 = 10'h198 == _T_5[9:0] ? image_1_408 : _GEN_983; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_985 = 10'h199 == _T_5[9:0] ? image_1_409 : _GEN_984; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_986 = 10'h19a == _T_5[9:0] ? image_1_410 : _GEN_985; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_987 = 10'h19b == _T_5[9:0] ? image_1_411 : _GEN_986; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_988 = 10'h19c == _T_5[9:0] ? image_1_412 : _GEN_987; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_989 = 10'h19d == _T_5[9:0] ? image_1_413 : _GEN_988; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_990 = 10'h19e == _T_5[9:0] ? image_1_414 : _GEN_989; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_991 = 10'h19f == _T_5[9:0] ? image_1_415 : _GEN_990; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_992 = 10'h1a0 == _T_5[9:0] ? image_1_416 : _GEN_991; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_993 = 10'h1a1 == _T_5[9:0] ? image_1_417 : _GEN_992; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_994 = 10'h1a2 == _T_5[9:0] ? image_1_418 : _GEN_993; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_995 = 10'h1a3 == _T_5[9:0] ? image_1_419 : _GEN_994; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_996 = 10'h1a4 == _T_5[9:0] ? image_1_420 : _GEN_995; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_997 = 10'h1a5 == _T_5[9:0] ? image_1_421 : _GEN_996; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_998 = 10'h1a6 == _T_5[9:0] ? image_1_422 : _GEN_997; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_999 = 10'h1a7 == _T_5[9:0] ? image_1_423 : _GEN_998; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1000 = 10'h1a8 == _T_5[9:0] ? image_1_424 : _GEN_999; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1001 = 10'h1a9 == _T_5[9:0] ? image_1_425 : _GEN_1000; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1002 = 10'h1aa == _T_5[9:0] ? image_1_426 : _GEN_1001; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1003 = 10'h1ab == _T_5[9:0] ? image_1_427 : _GEN_1002; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1004 = 10'h1ac == _T_5[9:0] ? image_1_428 : _GEN_1003; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1005 = 10'h1ad == _T_5[9:0] ? image_1_429 : _GEN_1004; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1006 = 10'h1ae == _T_5[9:0] ? image_1_430 : _GEN_1005; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1007 = 10'h1af == _T_5[9:0] ? image_1_431 : _GEN_1006; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1008 = 10'h1b0 == _T_5[9:0] ? image_1_432 : _GEN_1007; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1009 = 10'h1b1 == _T_5[9:0] ? image_1_433 : _GEN_1008; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1010 = 10'h1b2 == _T_5[9:0] ? image_1_434 : _GEN_1009; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1011 = 10'h1b3 == _T_5[9:0] ? image_1_435 : _GEN_1010; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1012 = 10'h1b4 == _T_5[9:0] ? image_1_436 : _GEN_1011; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1013 = 10'h1b5 == _T_5[9:0] ? image_1_437 : _GEN_1012; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1014 = 10'h1b6 == _T_5[9:0] ? image_1_438 : _GEN_1013; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1015 = 10'h1b7 == _T_5[9:0] ? image_1_439 : _GEN_1014; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1016 = 10'h1b8 == _T_5[9:0] ? image_1_440 : _GEN_1015; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1017 = 10'h1b9 == _T_5[9:0] ? image_1_441 : _GEN_1016; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1018 = 10'h1ba == _T_5[9:0] ? image_1_442 : _GEN_1017; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1019 = 10'h1bb == _T_5[9:0] ? image_1_443 : _GEN_1018; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1020 = 10'h1bc == _T_5[9:0] ? image_1_444 : _GEN_1019; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1021 = 10'h1bd == _T_5[9:0] ? image_1_445 : _GEN_1020; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1022 = 10'h1be == _T_5[9:0] ? image_1_446 : _GEN_1021; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1023 = 10'h1bf == _T_5[9:0] ? image_1_447 : _GEN_1022; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1024 = 10'h1c0 == _T_5[9:0] ? image_1_448 : _GEN_1023; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1025 = 10'h1c1 == _T_5[9:0] ? image_1_449 : _GEN_1024; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1026 = 10'h1c2 == _T_5[9:0] ? image_1_450 : _GEN_1025; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1027 = 10'h1c3 == _T_5[9:0] ? image_1_451 : _GEN_1026; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1028 = 10'h1c4 == _T_5[9:0] ? image_1_452 : _GEN_1027; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1029 = 10'h1c5 == _T_5[9:0] ? image_1_453 : _GEN_1028; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1030 = 10'h1c6 == _T_5[9:0] ? image_1_454 : _GEN_1029; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1031 = 10'h1c7 == _T_5[9:0] ? image_1_455 : _GEN_1030; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1032 = 10'h1c8 == _T_5[9:0] ? image_1_456 : _GEN_1031; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1033 = 10'h1c9 == _T_5[9:0] ? image_1_457 : _GEN_1032; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1034 = 10'h1ca == _T_5[9:0] ? image_1_458 : _GEN_1033; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1035 = 10'h1cb == _T_5[9:0] ? image_1_459 : _GEN_1034; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1036 = 10'h1cc == _T_5[9:0] ? image_1_460 : _GEN_1035; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1037 = 10'h1cd == _T_5[9:0] ? image_1_461 : _GEN_1036; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1038 = 10'h1ce == _T_5[9:0] ? image_1_462 : _GEN_1037; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1039 = 10'h1cf == _T_5[9:0] ? image_1_463 : _GEN_1038; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1040 = 10'h1d0 == _T_5[9:0] ? image_1_464 : _GEN_1039; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1041 = 10'h1d1 == _T_5[9:0] ? image_1_465 : _GEN_1040; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1042 = 10'h1d2 == _T_5[9:0] ? image_1_466 : _GEN_1041; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1043 = 10'h1d3 == _T_5[9:0] ? image_1_467 : _GEN_1042; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1044 = 10'h1d4 == _T_5[9:0] ? image_1_468 : _GEN_1043; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1045 = 10'h1d5 == _T_5[9:0] ? image_1_469 : _GEN_1044; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1046 = 10'h1d6 == _T_5[9:0] ? image_1_470 : _GEN_1045; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1047 = 10'h1d7 == _T_5[9:0] ? image_1_471 : _GEN_1046; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1048 = 10'h1d8 == _T_5[9:0] ? image_1_472 : _GEN_1047; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1049 = 10'h1d9 == _T_5[9:0] ? image_1_473 : _GEN_1048; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1050 = 10'h1da == _T_5[9:0] ? image_1_474 : _GEN_1049; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1051 = 10'h1db == _T_5[9:0] ? image_1_475 : _GEN_1050; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1052 = 10'h1dc == _T_5[9:0] ? image_1_476 : _GEN_1051; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1053 = 10'h1dd == _T_5[9:0] ? image_1_477 : _GEN_1052; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1054 = 10'h1de == _T_5[9:0] ? image_1_478 : _GEN_1053; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1055 = 10'h1df == _T_5[9:0] ? image_1_479 : _GEN_1054; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1056 = 10'h1e0 == _T_5[9:0] ? image_1_480 : _GEN_1055; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1057 = 10'h1e1 == _T_5[9:0] ? image_1_481 : _GEN_1056; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1058 = 10'h1e2 == _T_5[9:0] ? image_1_482 : _GEN_1057; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1059 = 10'h1e3 == _T_5[9:0] ? image_1_483 : _GEN_1058; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1060 = 10'h1e4 == _T_5[9:0] ? image_1_484 : _GEN_1059; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1061 = 10'h1e5 == _T_5[9:0] ? image_1_485 : _GEN_1060; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1062 = 10'h1e6 == _T_5[9:0] ? image_1_486 : _GEN_1061; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1063 = 10'h1e7 == _T_5[9:0] ? image_1_487 : _GEN_1062; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1064 = 10'h1e8 == _T_5[9:0] ? image_1_488 : _GEN_1063; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1065 = 10'h1e9 == _T_5[9:0] ? image_1_489 : _GEN_1064; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1066 = 10'h1ea == _T_5[9:0] ? image_1_490 : _GEN_1065; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1067 = 10'h1eb == _T_5[9:0] ? image_1_491 : _GEN_1066; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1068 = 10'h1ec == _T_5[9:0] ? image_1_492 : _GEN_1067; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1069 = 10'h1ed == _T_5[9:0] ? image_1_493 : _GEN_1068; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1070 = 10'h1ee == _T_5[9:0] ? image_1_494 : _GEN_1069; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1071 = 10'h1ef == _T_5[9:0] ? image_1_495 : _GEN_1070; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1072 = 10'h1f0 == _T_5[9:0] ? image_1_496 : _GEN_1071; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1073 = 10'h1f1 == _T_5[9:0] ? image_1_497 : _GEN_1072; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1074 = 10'h1f2 == _T_5[9:0] ? image_1_498 : _GEN_1073; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1075 = 10'h1f3 == _T_5[9:0] ? image_1_499 : _GEN_1074; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1076 = 10'h1f4 == _T_5[9:0] ? image_1_500 : _GEN_1075; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1077 = 10'h1f5 == _T_5[9:0] ? image_1_501 : _GEN_1076; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1078 = 10'h1f6 == _T_5[9:0] ? image_1_502 : _GEN_1077; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1079 = 10'h1f7 == _T_5[9:0] ? image_1_503 : _GEN_1078; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1080 = 10'h1f8 == _T_5[9:0] ? image_1_504 : _GEN_1079; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1081 = 10'h1f9 == _T_5[9:0] ? image_1_505 : _GEN_1080; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1082 = 10'h1fa == _T_5[9:0] ? image_1_506 : _GEN_1081; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1083 = 10'h1fb == _T_5[9:0] ? image_1_507 : _GEN_1082; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1084 = 10'h1fc == _T_5[9:0] ? image_1_508 : _GEN_1083; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1085 = 10'h1fd == _T_5[9:0] ? image_1_509 : _GEN_1084; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1086 = 10'h1fe == _T_5[9:0] ? image_1_510 : _GEN_1085; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1087 = 10'h1ff == _T_5[9:0] ? image_1_511 : _GEN_1086; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1088 = 10'h200 == _T_5[9:0] ? image_1_512 : _GEN_1087; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1089 = 10'h201 == _T_5[9:0] ? image_1_513 : _GEN_1088; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1090 = 10'h202 == _T_5[9:0] ? image_1_514 : _GEN_1089; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1091 = 10'h203 == _T_5[9:0] ? image_1_515 : _GEN_1090; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1092 = 10'h204 == _T_5[9:0] ? image_1_516 : _GEN_1091; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1093 = 10'h205 == _T_5[9:0] ? image_1_517 : _GEN_1092; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1094 = 10'h206 == _T_5[9:0] ? image_1_518 : _GEN_1093; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1095 = 10'h207 == _T_5[9:0] ? image_1_519 : _GEN_1094; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1096 = 10'h208 == _T_5[9:0] ? image_1_520 : _GEN_1095; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1097 = 10'h209 == _T_5[9:0] ? image_1_521 : _GEN_1096; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1098 = 10'h20a == _T_5[9:0] ? image_1_522 : _GEN_1097; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1099 = 10'h20b == _T_5[9:0] ? image_1_523 : _GEN_1098; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1100 = 10'h20c == _T_5[9:0] ? image_1_524 : _GEN_1099; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1101 = 10'h20d == _T_5[9:0] ? image_1_525 : _GEN_1100; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1102 = 10'h20e == _T_5[9:0] ? image_1_526 : _GEN_1101; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1103 = 10'h20f == _T_5[9:0] ? image_1_527 : _GEN_1102; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1104 = 10'h210 == _T_5[9:0] ? image_1_528 : _GEN_1103; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1105 = 10'h211 == _T_5[9:0] ? image_1_529 : _GEN_1104; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1106 = 10'h212 == _T_5[9:0] ? image_1_530 : _GEN_1105; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1107 = 10'h213 == _T_5[9:0] ? image_1_531 : _GEN_1106; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1108 = 10'h214 == _T_5[9:0] ? image_1_532 : _GEN_1107; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1109 = 10'h215 == _T_5[9:0] ? image_1_533 : _GEN_1108; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1110 = 10'h216 == _T_5[9:0] ? image_1_534 : _GEN_1109; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1111 = 10'h217 == _T_5[9:0] ? image_1_535 : _GEN_1110; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1112 = 10'h218 == _T_5[9:0] ? image_1_536 : _GEN_1111; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1113 = 10'h219 == _T_5[9:0] ? image_1_537 : _GEN_1112; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1114 = 10'h21a == _T_5[9:0] ? image_1_538 : _GEN_1113; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1115 = 10'h21b == _T_5[9:0] ? image_1_539 : _GEN_1114; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1116 = 10'h21c == _T_5[9:0] ? image_1_540 : _GEN_1115; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1117 = 10'h21d == _T_5[9:0] ? image_1_541 : _GEN_1116; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1118 = 10'h21e == _T_5[9:0] ? image_1_542 : _GEN_1117; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1119 = 10'h21f == _T_5[9:0] ? image_1_543 : _GEN_1118; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1120 = 10'h220 == _T_5[9:0] ? image_1_544 : _GEN_1119; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1121 = 10'h221 == _T_5[9:0] ? image_1_545 : _GEN_1120; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1122 = 10'h222 == _T_5[9:0] ? image_1_546 : _GEN_1121; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1123 = 10'h223 == _T_5[9:0] ? image_1_547 : _GEN_1122; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1124 = 10'h224 == _T_5[9:0] ? image_1_548 : _GEN_1123; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1125 = 10'h225 == _T_5[9:0] ? image_1_549 : _GEN_1124; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1126 = 10'h226 == _T_5[9:0] ? image_1_550 : _GEN_1125; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1127 = 10'h227 == _T_5[9:0] ? image_1_551 : _GEN_1126; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1128 = 10'h228 == _T_5[9:0] ? image_1_552 : _GEN_1127; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1129 = 10'h229 == _T_5[9:0] ? image_1_553 : _GEN_1128; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1130 = 10'h22a == _T_5[9:0] ? image_1_554 : _GEN_1129; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1131 = 10'h22b == _T_5[9:0] ? image_1_555 : _GEN_1130; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1132 = 10'h22c == _T_5[9:0] ? image_1_556 : _GEN_1131; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1133 = 10'h22d == _T_5[9:0] ? image_1_557 : _GEN_1132; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1134 = 10'h22e == _T_5[9:0] ? image_1_558 : _GEN_1133; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1135 = 10'h22f == _T_5[9:0] ? image_1_559 : _GEN_1134; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1136 = 10'h230 == _T_5[9:0] ? image_1_560 : _GEN_1135; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1137 = 10'h231 == _T_5[9:0] ? image_1_561 : _GEN_1136; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1138 = 10'h232 == _T_5[9:0] ? image_1_562 : _GEN_1137; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1139 = 10'h233 == _T_5[9:0] ? image_1_563 : _GEN_1138; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1140 = 10'h234 == _T_5[9:0] ? image_1_564 : _GEN_1139; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1141 = 10'h235 == _T_5[9:0] ? image_1_565 : _GEN_1140; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1142 = 10'h236 == _T_5[9:0] ? image_1_566 : _GEN_1141; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1143 = 10'h237 == _T_5[9:0] ? image_1_567 : _GEN_1142; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1144 = 10'h238 == _T_5[9:0] ? image_1_568 : _GEN_1143; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1145 = 10'h239 == _T_5[9:0] ? image_1_569 : _GEN_1144; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1146 = 10'h23a == _T_5[9:0] ? image_1_570 : _GEN_1145; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1147 = 10'h23b == _T_5[9:0] ? image_1_571 : _GEN_1146; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1148 = 10'h23c == _T_5[9:0] ? image_1_572 : _GEN_1147; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1149 = 10'h23d == _T_5[9:0] ? image_1_573 : _GEN_1148; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1150 = 10'h23e == _T_5[9:0] ? image_1_574 : _GEN_1149; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1153 = 10'h1 == _T_5[9:0] ? image_2_1 : image_2_0; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1154 = 10'h2 == _T_5[9:0] ? image_2_2 : _GEN_1153; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1155 = 10'h3 == _T_5[9:0] ? image_2_3 : _GEN_1154; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1156 = 10'h4 == _T_5[9:0] ? image_2_4 : _GEN_1155; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1157 = 10'h5 == _T_5[9:0] ? image_2_5 : _GEN_1156; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1158 = 10'h6 == _T_5[9:0] ? image_2_6 : _GEN_1157; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1159 = 10'h7 == _T_5[9:0] ? image_2_7 : _GEN_1158; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1160 = 10'h8 == _T_5[9:0] ? image_2_8 : _GEN_1159; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1161 = 10'h9 == _T_5[9:0] ? image_2_9 : _GEN_1160; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1162 = 10'ha == _T_5[9:0] ? image_2_10 : _GEN_1161; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1163 = 10'hb == _T_5[9:0] ? image_2_11 : _GEN_1162; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1164 = 10'hc == _T_5[9:0] ? image_2_12 : _GEN_1163; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1165 = 10'hd == _T_5[9:0] ? image_2_13 : _GEN_1164; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1166 = 10'he == _T_5[9:0] ? image_2_14 : _GEN_1165; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1167 = 10'hf == _T_5[9:0] ? image_2_15 : _GEN_1166; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1168 = 10'h10 == _T_5[9:0] ? image_2_16 : _GEN_1167; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1169 = 10'h11 == _T_5[9:0] ? image_2_17 : _GEN_1168; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1170 = 10'h12 == _T_5[9:0] ? image_2_18 : _GEN_1169; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1171 = 10'h13 == _T_5[9:0] ? image_2_19 : _GEN_1170; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1172 = 10'h14 == _T_5[9:0] ? image_2_20 : _GEN_1171; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1173 = 10'h15 == _T_5[9:0] ? image_2_21 : _GEN_1172; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1174 = 10'h16 == _T_5[9:0] ? image_2_22 : _GEN_1173; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1175 = 10'h17 == _T_5[9:0] ? image_2_23 : _GEN_1174; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1176 = 10'h18 == _T_5[9:0] ? image_2_24 : _GEN_1175; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1177 = 10'h19 == _T_5[9:0] ? image_2_25 : _GEN_1176; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1178 = 10'h1a == _T_5[9:0] ? image_2_26 : _GEN_1177; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1179 = 10'h1b == _T_5[9:0] ? image_2_27 : _GEN_1178; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1180 = 10'h1c == _T_5[9:0] ? image_2_28 : _GEN_1179; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1181 = 10'h1d == _T_5[9:0] ? image_2_29 : _GEN_1180; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1182 = 10'h1e == _T_5[9:0] ? image_2_30 : _GEN_1181; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1183 = 10'h1f == _T_5[9:0] ? image_2_31 : _GEN_1182; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1184 = 10'h20 == _T_5[9:0] ? image_2_32 : _GEN_1183; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1185 = 10'h21 == _T_5[9:0] ? image_2_33 : _GEN_1184; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1186 = 10'h22 == _T_5[9:0] ? image_2_34 : _GEN_1185; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1187 = 10'h23 == _T_5[9:0] ? image_2_35 : _GEN_1186; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1188 = 10'h24 == _T_5[9:0] ? image_2_36 : _GEN_1187; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1189 = 10'h25 == _T_5[9:0] ? image_2_37 : _GEN_1188; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1190 = 10'h26 == _T_5[9:0] ? image_2_38 : _GEN_1189; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1191 = 10'h27 == _T_5[9:0] ? image_2_39 : _GEN_1190; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1192 = 10'h28 == _T_5[9:0] ? image_2_40 : _GEN_1191; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1193 = 10'h29 == _T_5[9:0] ? image_2_41 : _GEN_1192; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1194 = 10'h2a == _T_5[9:0] ? image_2_42 : _GEN_1193; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1195 = 10'h2b == _T_5[9:0] ? image_2_43 : _GEN_1194; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1196 = 10'h2c == _T_5[9:0] ? image_2_44 : _GEN_1195; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1197 = 10'h2d == _T_5[9:0] ? image_2_45 : _GEN_1196; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1198 = 10'h2e == _T_5[9:0] ? image_2_46 : _GEN_1197; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1199 = 10'h2f == _T_5[9:0] ? image_2_47 : _GEN_1198; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1200 = 10'h30 == _T_5[9:0] ? image_2_48 : _GEN_1199; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1201 = 10'h31 == _T_5[9:0] ? image_2_49 : _GEN_1200; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1202 = 10'h32 == _T_5[9:0] ? image_2_50 : _GEN_1201; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1203 = 10'h33 == _T_5[9:0] ? image_2_51 : _GEN_1202; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1204 = 10'h34 == _T_5[9:0] ? image_2_52 : _GEN_1203; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1205 = 10'h35 == _T_5[9:0] ? image_2_53 : _GEN_1204; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1206 = 10'h36 == _T_5[9:0] ? image_2_54 : _GEN_1205; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1207 = 10'h37 == _T_5[9:0] ? image_2_55 : _GEN_1206; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1208 = 10'h38 == _T_5[9:0] ? image_2_56 : _GEN_1207; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1209 = 10'h39 == _T_5[9:0] ? image_2_57 : _GEN_1208; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1210 = 10'h3a == _T_5[9:0] ? image_2_58 : _GEN_1209; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1211 = 10'h3b == _T_5[9:0] ? image_2_59 : _GEN_1210; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1212 = 10'h3c == _T_5[9:0] ? image_2_60 : _GEN_1211; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1213 = 10'h3d == _T_5[9:0] ? image_2_61 : _GEN_1212; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1214 = 10'h3e == _T_5[9:0] ? image_2_62 : _GEN_1213; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1215 = 10'h3f == _T_5[9:0] ? image_2_63 : _GEN_1214; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1216 = 10'h40 == _T_5[9:0] ? image_2_64 : _GEN_1215; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1217 = 10'h41 == _T_5[9:0] ? image_2_65 : _GEN_1216; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1218 = 10'h42 == _T_5[9:0] ? image_2_66 : _GEN_1217; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1219 = 10'h43 == _T_5[9:0] ? image_2_67 : _GEN_1218; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1220 = 10'h44 == _T_5[9:0] ? image_2_68 : _GEN_1219; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1221 = 10'h45 == _T_5[9:0] ? image_2_69 : _GEN_1220; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1222 = 10'h46 == _T_5[9:0] ? image_2_70 : _GEN_1221; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1223 = 10'h47 == _T_5[9:0] ? image_2_71 : _GEN_1222; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1224 = 10'h48 == _T_5[9:0] ? image_2_72 : _GEN_1223; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1225 = 10'h49 == _T_5[9:0] ? image_2_73 : _GEN_1224; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1226 = 10'h4a == _T_5[9:0] ? image_2_74 : _GEN_1225; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1227 = 10'h4b == _T_5[9:0] ? image_2_75 : _GEN_1226; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1228 = 10'h4c == _T_5[9:0] ? image_2_76 : _GEN_1227; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1229 = 10'h4d == _T_5[9:0] ? image_2_77 : _GEN_1228; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1230 = 10'h4e == _T_5[9:0] ? image_2_78 : _GEN_1229; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1231 = 10'h4f == _T_5[9:0] ? image_2_79 : _GEN_1230; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1232 = 10'h50 == _T_5[9:0] ? image_2_80 : _GEN_1231; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1233 = 10'h51 == _T_5[9:0] ? image_2_81 : _GEN_1232; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1234 = 10'h52 == _T_5[9:0] ? image_2_82 : _GEN_1233; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1235 = 10'h53 == _T_5[9:0] ? image_2_83 : _GEN_1234; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1236 = 10'h54 == _T_5[9:0] ? image_2_84 : _GEN_1235; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1237 = 10'h55 == _T_5[9:0] ? image_2_85 : _GEN_1236; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1238 = 10'h56 == _T_5[9:0] ? image_2_86 : _GEN_1237; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1239 = 10'h57 == _T_5[9:0] ? image_2_87 : _GEN_1238; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1240 = 10'h58 == _T_5[9:0] ? image_2_88 : _GEN_1239; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1241 = 10'h59 == _T_5[9:0] ? image_2_89 : _GEN_1240; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1242 = 10'h5a == _T_5[9:0] ? image_2_90 : _GEN_1241; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1243 = 10'h5b == _T_5[9:0] ? image_2_91 : _GEN_1242; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1244 = 10'h5c == _T_5[9:0] ? image_2_92 : _GEN_1243; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1245 = 10'h5d == _T_5[9:0] ? image_2_93 : _GEN_1244; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1246 = 10'h5e == _T_5[9:0] ? image_2_94 : _GEN_1245; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1247 = 10'h5f == _T_5[9:0] ? image_2_95 : _GEN_1246; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1248 = 10'h60 == _T_5[9:0] ? image_2_96 : _GEN_1247; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1249 = 10'h61 == _T_5[9:0] ? image_2_97 : _GEN_1248; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1250 = 10'h62 == _T_5[9:0] ? image_2_98 : _GEN_1249; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1251 = 10'h63 == _T_5[9:0] ? image_2_99 : _GEN_1250; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1252 = 10'h64 == _T_5[9:0] ? image_2_100 : _GEN_1251; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1253 = 10'h65 == _T_5[9:0] ? image_2_101 : _GEN_1252; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1254 = 10'h66 == _T_5[9:0] ? image_2_102 : _GEN_1253; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1255 = 10'h67 == _T_5[9:0] ? image_2_103 : _GEN_1254; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1256 = 10'h68 == _T_5[9:0] ? image_2_104 : _GEN_1255; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1257 = 10'h69 == _T_5[9:0] ? image_2_105 : _GEN_1256; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1258 = 10'h6a == _T_5[9:0] ? image_2_106 : _GEN_1257; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1259 = 10'h6b == _T_5[9:0] ? image_2_107 : _GEN_1258; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1260 = 10'h6c == _T_5[9:0] ? image_2_108 : _GEN_1259; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1261 = 10'h6d == _T_5[9:0] ? image_2_109 : _GEN_1260; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1262 = 10'h6e == _T_5[9:0] ? image_2_110 : _GEN_1261; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1263 = 10'h6f == _T_5[9:0] ? image_2_111 : _GEN_1262; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1264 = 10'h70 == _T_5[9:0] ? image_2_112 : _GEN_1263; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1265 = 10'h71 == _T_5[9:0] ? image_2_113 : _GEN_1264; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1266 = 10'h72 == _T_5[9:0] ? image_2_114 : _GEN_1265; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1267 = 10'h73 == _T_5[9:0] ? image_2_115 : _GEN_1266; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1268 = 10'h74 == _T_5[9:0] ? image_2_116 : _GEN_1267; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1269 = 10'h75 == _T_5[9:0] ? image_2_117 : _GEN_1268; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1270 = 10'h76 == _T_5[9:0] ? image_2_118 : _GEN_1269; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1271 = 10'h77 == _T_5[9:0] ? image_2_119 : _GEN_1270; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1272 = 10'h78 == _T_5[9:0] ? image_2_120 : _GEN_1271; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1273 = 10'h79 == _T_5[9:0] ? image_2_121 : _GEN_1272; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1274 = 10'h7a == _T_5[9:0] ? image_2_122 : _GEN_1273; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1275 = 10'h7b == _T_5[9:0] ? image_2_123 : _GEN_1274; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1276 = 10'h7c == _T_5[9:0] ? image_2_124 : _GEN_1275; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1277 = 10'h7d == _T_5[9:0] ? image_2_125 : _GEN_1276; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1278 = 10'h7e == _T_5[9:0] ? image_2_126 : _GEN_1277; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1279 = 10'h7f == _T_5[9:0] ? image_2_127 : _GEN_1278; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1280 = 10'h80 == _T_5[9:0] ? image_2_128 : _GEN_1279; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1281 = 10'h81 == _T_5[9:0] ? image_2_129 : _GEN_1280; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1282 = 10'h82 == _T_5[9:0] ? image_2_130 : _GEN_1281; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1283 = 10'h83 == _T_5[9:0] ? image_2_131 : _GEN_1282; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1284 = 10'h84 == _T_5[9:0] ? image_2_132 : _GEN_1283; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1285 = 10'h85 == _T_5[9:0] ? image_2_133 : _GEN_1284; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1286 = 10'h86 == _T_5[9:0] ? image_2_134 : _GEN_1285; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1287 = 10'h87 == _T_5[9:0] ? image_2_135 : _GEN_1286; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1288 = 10'h88 == _T_5[9:0] ? image_2_136 : _GEN_1287; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1289 = 10'h89 == _T_5[9:0] ? image_2_137 : _GEN_1288; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1290 = 10'h8a == _T_5[9:0] ? image_2_138 : _GEN_1289; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1291 = 10'h8b == _T_5[9:0] ? image_2_139 : _GEN_1290; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1292 = 10'h8c == _T_5[9:0] ? image_2_140 : _GEN_1291; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1293 = 10'h8d == _T_5[9:0] ? image_2_141 : _GEN_1292; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1294 = 10'h8e == _T_5[9:0] ? image_2_142 : _GEN_1293; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1295 = 10'h8f == _T_5[9:0] ? image_2_143 : _GEN_1294; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1296 = 10'h90 == _T_5[9:0] ? image_2_144 : _GEN_1295; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1297 = 10'h91 == _T_5[9:0] ? image_2_145 : _GEN_1296; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1298 = 10'h92 == _T_5[9:0] ? image_2_146 : _GEN_1297; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1299 = 10'h93 == _T_5[9:0] ? image_2_147 : _GEN_1298; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1300 = 10'h94 == _T_5[9:0] ? image_2_148 : _GEN_1299; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1301 = 10'h95 == _T_5[9:0] ? image_2_149 : _GEN_1300; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1302 = 10'h96 == _T_5[9:0] ? image_2_150 : _GEN_1301; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1303 = 10'h97 == _T_5[9:0] ? image_2_151 : _GEN_1302; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1304 = 10'h98 == _T_5[9:0] ? image_2_152 : _GEN_1303; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1305 = 10'h99 == _T_5[9:0] ? image_2_153 : _GEN_1304; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1306 = 10'h9a == _T_5[9:0] ? image_2_154 : _GEN_1305; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1307 = 10'h9b == _T_5[9:0] ? image_2_155 : _GEN_1306; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1308 = 10'h9c == _T_5[9:0] ? image_2_156 : _GEN_1307; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1309 = 10'h9d == _T_5[9:0] ? image_2_157 : _GEN_1308; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1310 = 10'h9e == _T_5[9:0] ? image_2_158 : _GEN_1309; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1311 = 10'h9f == _T_5[9:0] ? image_2_159 : _GEN_1310; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1312 = 10'ha0 == _T_5[9:0] ? image_2_160 : _GEN_1311; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1313 = 10'ha1 == _T_5[9:0] ? image_2_161 : _GEN_1312; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1314 = 10'ha2 == _T_5[9:0] ? image_2_162 : _GEN_1313; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1315 = 10'ha3 == _T_5[9:0] ? image_2_163 : _GEN_1314; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1316 = 10'ha4 == _T_5[9:0] ? image_2_164 : _GEN_1315; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1317 = 10'ha5 == _T_5[9:0] ? image_2_165 : _GEN_1316; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1318 = 10'ha6 == _T_5[9:0] ? image_2_166 : _GEN_1317; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1319 = 10'ha7 == _T_5[9:0] ? image_2_167 : _GEN_1318; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1320 = 10'ha8 == _T_5[9:0] ? image_2_168 : _GEN_1319; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1321 = 10'ha9 == _T_5[9:0] ? image_2_169 : _GEN_1320; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1322 = 10'haa == _T_5[9:0] ? image_2_170 : _GEN_1321; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1323 = 10'hab == _T_5[9:0] ? image_2_171 : _GEN_1322; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1324 = 10'hac == _T_5[9:0] ? image_2_172 : _GEN_1323; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1325 = 10'had == _T_5[9:0] ? image_2_173 : _GEN_1324; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1326 = 10'hae == _T_5[9:0] ? image_2_174 : _GEN_1325; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1327 = 10'haf == _T_5[9:0] ? image_2_175 : _GEN_1326; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1328 = 10'hb0 == _T_5[9:0] ? image_2_176 : _GEN_1327; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1329 = 10'hb1 == _T_5[9:0] ? image_2_177 : _GEN_1328; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1330 = 10'hb2 == _T_5[9:0] ? image_2_178 : _GEN_1329; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1331 = 10'hb3 == _T_5[9:0] ? image_2_179 : _GEN_1330; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1332 = 10'hb4 == _T_5[9:0] ? image_2_180 : _GEN_1331; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1333 = 10'hb5 == _T_5[9:0] ? image_2_181 : _GEN_1332; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1334 = 10'hb6 == _T_5[9:0] ? image_2_182 : _GEN_1333; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1335 = 10'hb7 == _T_5[9:0] ? image_2_183 : _GEN_1334; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1336 = 10'hb8 == _T_5[9:0] ? image_2_184 : _GEN_1335; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1337 = 10'hb9 == _T_5[9:0] ? image_2_185 : _GEN_1336; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1338 = 10'hba == _T_5[9:0] ? image_2_186 : _GEN_1337; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1339 = 10'hbb == _T_5[9:0] ? image_2_187 : _GEN_1338; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1340 = 10'hbc == _T_5[9:0] ? image_2_188 : _GEN_1339; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1341 = 10'hbd == _T_5[9:0] ? image_2_189 : _GEN_1340; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1342 = 10'hbe == _T_5[9:0] ? image_2_190 : _GEN_1341; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1343 = 10'hbf == _T_5[9:0] ? image_2_191 : _GEN_1342; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1344 = 10'hc0 == _T_5[9:0] ? image_2_192 : _GEN_1343; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1345 = 10'hc1 == _T_5[9:0] ? image_2_193 : _GEN_1344; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1346 = 10'hc2 == _T_5[9:0] ? image_2_194 : _GEN_1345; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1347 = 10'hc3 == _T_5[9:0] ? image_2_195 : _GEN_1346; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1348 = 10'hc4 == _T_5[9:0] ? image_2_196 : _GEN_1347; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1349 = 10'hc5 == _T_5[9:0] ? image_2_197 : _GEN_1348; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1350 = 10'hc6 == _T_5[9:0] ? image_2_198 : _GEN_1349; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1351 = 10'hc7 == _T_5[9:0] ? image_2_199 : _GEN_1350; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1352 = 10'hc8 == _T_5[9:0] ? image_2_200 : _GEN_1351; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1353 = 10'hc9 == _T_5[9:0] ? image_2_201 : _GEN_1352; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1354 = 10'hca == _T_5[9:0] ? image_2_202 : _GEN_1353; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1355 = 10'hcb == _T_5[9:0] ? image_2_203 : _GEN_1354; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1356 = 10'hcc == _T_5[9:0] ? image_2_204 : _GEN_1355; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1357 = 10'hcd == _T_5[9:0] ? image_2_205 : _GEN_1356; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1358 = 10'hce == _T_5[9:0] ? image_2_206 : _GEN_1357; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1359 = 10'hcf == _T_5[9:0] ? image_2_207 : _GEN_1358; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1360 = 10'hd0 == _T_5[9:0] ? image_2_208 : _GEN_1359; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1361 = 10'hd1 == _T_5[9:0] ? image_2_209 : _GEN_1360; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1362 = 10'hd2 == _T_5[9:0] ? image_2_210 : _GEN_1361; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1363 = 10'hd3 == _T_5[9:0] ? image_2_211 : _GEN_1362; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1364 = 10'hd4 == _T_5[9:0] ? image_2_212 : _GEN_1363; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1365 = 10'hd5 == _T_5[9:0] ? image_2_213 : _GEN_1364; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1366 = 10'hd6 == _T_5[9:0] ? image_2_214 : _GEN_1365; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1367 = 10'hd7 == _T_5[9:0] ? image_2_215 : _GEN_1366; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1368 = 10'hd8 == _T_5[9:0] ? image_2_216 : _GEN_1367; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1369 = 10'hd9 == _T_5[9:0] ? image_2_217 : _GEN_1368; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1370 = 10'hda == _T_5[9:0] ? image_2_218 : _GEN_1369; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1371 = 10'hdb == _T_5[9:0] ? image_2_219 : _GEN_1370; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1372 = 10'hdc == _T_5[9:0] ? image_2_220 : _GEN_1371; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1373 = 10'hdd == _T_5[9:0] ? image_2_221 : _GEN_1372; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1374 = 10'hde == _T_5[9:0] ? image_2_222 : _GEN_1373; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1375 = 10'hdf == _T_5[9:0] ? image_2_223 : _GEN_1374; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1376 = 10'he0 == _T_5[9:0] ? image_2_224 : _GEN_1375; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1377 = 10'he1 == _T_5[9:0] ? image_2_225 : _GEN_1376; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1378 = 10'he2 == _T_5[9:0] ? image_2_226 : _GEN_1377; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1379 = 10'he3 == _T_5[9:0] ? image_2_227 : _GEN_1378; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1380 = 10'he4 == _T_5[9:0] ? image_2_228 : _GEN_1379; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1381 = 10'he5 == _T_5[9:0] ? image_2_229 : _GEN_1380; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1382 = 10'he6 == _T_5[9:0] ? image_2_230 : _GEN_1381; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1383 = 10'he7 == _T_5[9:0] ? image_2_231 : _GEN_1382; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1384 = 10'he8 == _T_5[9:0] ? image_2_232 : _GEN_1383; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1385 = 10'he9 == _T_5[9:0] ? image_2_233 : _GEN_1384; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1386 = 10'hea == _T_5[9:0] ? image_2_234 : _GEN_1385; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1387 = 10'heb == _T_5[9:0] ? image_2_235 : _GEN_1386; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1388 = 10'hec == _T_5[9:0] ? image_2_236 : _GEN_1387; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1389 = 10'hed == _T_5[9:0] ? image_2_237 : _GEN_1388; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1390 = 10'hee == _T_5[9:0] ? image_2_238 : _GEN_1389; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1391 = 10'hef == _T_5[9:0] ? image_2_239 : _GEN_1390; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1392 = 10'hf0 == _T_5[9:0] ? image_2_240 : _GEN_1391; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1393 = 10'hf1 == _T_5[9:0] ? image_2_241 : _GEN_1392; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1394 = 10'hf2 == _T_5[9:0] ? image_2_242 : _GEN_1393; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1395 = 10'hf3 == _T_5[9:0] ? image_2_243 : _GEN_1394; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1396 = 10'hf4 == _T_5[9:0] ? image_2_244 : _GEN_1395; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1397 = 10'hf5 == _T_5[9:0] ? image_2_245 : _GEN_1396; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1398 = 10'hf6 == _T_5[9:0] ? image_2_246 : _GEN_1397; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1399 = 10'hf7 == _T_5[9:0] ? image_2_247 : _GEN_1398; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1400 = 10'hf8 == _T_5[9:0] ? image_2_248 : _GEN_1399; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1401 = 10'hf9 == _T_5[9:0] ? image_2_249 : _GEN_1400; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1402 = 10'hfa == _T_5[9:0] ? image_2_250 : _GEN_1401; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1403 = 10'hfb == _T_5[9:0] ? image_2_251 : _GEN_1402; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1404 = 10'hfc == _T_5[9:0] ? image_2_252 : _GEN_1403; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1405 = 10'hfd == _T_5[9:0] ? image_2_253 : _GEN_1404; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1406 = 10'hfe == _T_5[9:0] ? image_2_254 : _GEN_1405; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1407 = 10'hff == _T_5[9:0] ? image_2_255 : _GEN_1406; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1408 = 10'h100 == _T_5[9:0] ? image_2_256 : _GEN_1407; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1409 = 10'h101 == _T_5[9:0] ? image_2_257 : _GEN_1408; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1410 = 10'h102 == _T_5[9:0] ? image_2_258 : _GEN_1409; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1411 = 10'h103 == _T_5[9:0] ? image_2_259 : _GEN_1410; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1412 = 10'h104 == _T_5[9:0] ? image_2_260 : _GEN_1411; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1413 = 10'h105 == _T_5[9:0] ? image_2_261 : _GEN_1412; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1414 = 10'h106 == _T_5[9:0] ? image_2_262 : _GEN_1413; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1415 = 10'h107 == _T_5[9:0] ? image_2_263 : _GEN_1414; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1416 = 10'h108 == _T_5[9:0] ? image_2_264 : _GEN_1415; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1417 = 10'h109 == _T_5[9:0] ? image_2_265 : _GEN_1416; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1418 = 10'h10a == _T_5[9:0] ? image_2_266 : _GEN_1417; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1419 = 10'h10b == _T_5[9:0] ? image_2_267 : _GEN_1418; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1420 = 10'h10c == _T_5[9:0] ? image_2_268 : _GEN_1419; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1421 = 10'h10d == _T_5[9:0] ? image_2_269 : _GEN_1420; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1422 = 10'h10e == _T_5[9:0] ? image_2_270 : _GEN_1421; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1423 = 10'h10f == _T_5[9:0] ? image_2_271 : _GEN_1422; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1424 = 10'h110 == _T_5[9:0] ? image_2_272 : _GEN_1423; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1425 = 10'h111 == _T_5[9:0] ? image_2_273 : _GEN_1424; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1426 = 10'h112 == _T_5[9:0] ? image_2_274 : _GEN_1425; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1427 = 10'h113 == _T_5[9:0] ? image_2_275 : _GEN_1426; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1428 = 10'h114 == _T_5[9:0] ? image_2_276 : _GEN_1427; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1429 = 10'h115 == _T_5[9:0] ? image_2_277 : _GEN_1428; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1430 = 10'h116 == _T_5[9:0] ? image_2_278 : _GEN_1429; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1431 = 10'h117 == _T_5[9:0] ? image_2_279 : _GEN_1430; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1432 = 10'h118 == _T_5[9:0] ? image_2_280 : _GEN_1431; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1433 = 10'h119 == _T_5[9:0] ? image_2_281 : _GEN_1432; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1434 = 10'h11a == _T_5[9:0] ? image_2_282 : _GEN_1433; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1435 = 10'h11b == _T_5[9:0] ? image_2_283 : _GEN_1434; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1436 = 10'h11c == _T_5[9:0] ? image_2_284 : _GEN_1435; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1437 = 10'h11d == _T_5[9:0] ? image_2_285 : _GEN_1436; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1438 = 10'h11e == _T_5[9:0] ? image_2_286 : _GEN_1437; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1439 = 10'h11f == _T_5[9:0] ? image_2_287 : _GEN_1438; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1440 = 10'h120 == _T_5[9:0] ? image_2_288 : _GEN_1439; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1441 = 10'h121 == _T_5[9:0] ? image_2_289 : _GEN_1440; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1442 = 10'h122 == _T_5[9:0] ? image_2_290 : _GEN_1441; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1443 = 10'h123 == _T_5[9:0] ? image_2_291 : _GEN_1442; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1444 = 10'h124 == _T_5[9:0] ? image_2_292 : _GEN_1443; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1445 = 10'h125 == _T_5[9:0] ? image_2_293 : _GEN_1444; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1446 = 10'h126 == _T_5[9:0] ? image_2_294 : _GEN_1445; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1447 = 10'h127 == _T_5[9:0] ? image_2_295 : _GEN_1446; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1448 = 10'h128 == _T_5[9:0] ? image_2_296 : _GEN_1447; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1449 = 10'h129 == _T_5[9:0] ? image_2_297 : _GEN_1448; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1450 = 10'h12a == _T_5[9:0] ? image_2_298 : _GEN_1449; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1451 = 10'h12b == _T_5[9:0] ? image_2_299 : _GEN_1450; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1452 = 10'h12c == _T_5[9:0] ? image_2_300 : _GEN_1451; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1453 = 10'h12d == _T_5[9:0] ? image_2_301 : _GEN_1452; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1454 = 10'h12e == _T_5[9:0] ? image_2_302 : _GEN_1453; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1455 = 10'h12f == _T_5[9:0] ? image_2_303 : _GEN_1454; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1456 = 10'h130 == _T_5[9:0] ? image_2_304 : _GEN_1455; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1457 = 10'h131 == _T_5[9:0] ? image_2_305 : _GEN_1456; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1458 = 10'h132 == _T_5[9:0] ? image_2_306 : _GEN_1457; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1459 = 10'h133 == _T_5[9:0] ? image_2_307 : _GEN_1458; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1460 = 10'h134 == _T_5[9:0] ? image_2_308 : _GEN_1459; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1461 = 10'h135 == _T_5[9:0] ? image_2_309 : _GEN_1460; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1462 = 10'h136 == _T_5[9:0] ? image_2_310 : _GEN_1461; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1463 = 10'h137 == _T_5[9:0] ? image_2_311 : _GEN_1462; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1464 = 10'h138 == _T_5[9:0] ? image_2_312 : _GEN_1463; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1465 = 10'h139 == _T_5[9:0] ? image_2_313 : _GEN_1464; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1466 = 10'h13a == _T_5[9:0] ? image_2_314 : _GEN_1465; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1467 = 10'h13b == _T_5[9:0] ? image_2_315 : _GEN_1466; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1468 = 10'h13c == _T_5[9:0] ? image_2_316 : _GEN_1467; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1469 = 10'h13d == _T_5[9:0] ? image_2_317 : _GEN_1468; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1470 = 10'h13e == _T_5[9:0] ? image_2_318 : _GEN_1469; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1471 = 10'h13f == _T_5[9:0] ? image_2_319 : _GEN_1470; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1472 = 10'h140 == _T_5[9:0] ? image_2_320 : _GEN_1471; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1473 = 10'h141 == _T_5[9:0] ? image_2_321 : _GEN_1472; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1474 = 10'h142 == _T_5[9:0] ? image_2_322 : _GEN_1473; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1475 = 10'h143 == _T_5[9:0] ? image_2_323 : _GEN_1474; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1476 = 10'h144 == _T_5[9:0] ? image_2_324 : _GEN_1475; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1477 = 10'h145 == _T_5[9:0] ? image_2_325 : _GEN_1476; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1478 = 10'h146 == _T_5[9:0] ? image_2_326 : _GEN_1477; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1479 = 10'h147 == _T_5[9:0] ? image_2_327 : _GEN_1478; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1480 = 10'h148 == _T_5[9:0] ? image_2_328 : _GEN_1479; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1481 = 10'h149 == _T_5[9:0] ? image_2_329 : _GEN_1480; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1482 = 10'h14a == _T_5[9:0] ? image_2_330 : _GEN_1481; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1483 = 10'h14b == _T_5[9:0] ? image_2_331 : _GEN_1482; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1484 = 10'h14c == _T_5[9:0] ? image_2_332 : _GEN_1483; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1485 = 10'h14d == _T_5[9:0] ? image_2_333 : _GEN_1484; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1486 = 10'h14e == _T_5[9:0] ? image_2_334 : _GEN_1485; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1487 = 10'h14f == _T_5[9:0] ? image_2_335 : _GEN_1486; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1488 = 10'h150 == _T_5[9:0] ? image_2_336 : _GEN_1487; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1489 = 10'h151 == _T_5[9:0] ? image_2_337 : _GEN_1488; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1490 = 10'h152 == _T_5[9:0] ? image_2_338 : _GEN_1489; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1491 = 10'h153 == _T_5[9:0] ? image_2_339 : _GEN_1490; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1492 = 10'h154 == _T_5[9:0] ? image_2_340 : _GEN_1491; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1493 = 10'h155 == _T_5[9:0] ? image_2_341 : _GEN_1492; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1494 = 10'h156 == _T_5[9:0] ? image_2_342 : _GEN_1493; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1495 = 10'h157 == _T_5[9:0] ? image_2_343 : _GEN_1494; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1496 = 10'h158 == _T_5[9:0] ? image_2_344 : _GEN_1495; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1497 = 10'h159 == _T_5[9:0] ? image_2_345 : _GEN_1496; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1498 = 10'h15a == _T_5[9:0] ? image_2_346 : _GEN_1497; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1499 = 10'h15b == _T_5[9:0] ? image_2_347 : _GEN_1498; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1500 = 10'h15c == _T_5[9:0] ? image_2_348 : _GEN_1499; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1501 = 10'h15d == _T_5[9:0] ? image_2_349 : _GEN_1500; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1502 = 10'h15e == _T_5[9:0] ? image_2_350 : _GEN_1501; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1503 = 10'h15f == _T_5[9:0] ? image_2_351 : _GEN_1502; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1504 = 10'h160 == _T_5[9:0] ? image_2_352 : _GEN_1503; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1505 = 10'h161 == _T_5[9:0] ? image_2_353 : _GEN_1504; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1506 = 10'h162 == _T_5[9:0] ? image_2_354 : _GEN_1505; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1507 = 10'h163 == _T_5[9:0] ? image_2_355 : _GEN_1506; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1508 = 10'h164 == _T_5[9:0] ? image_2_356 : _GEN_1507; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1509 = 10'h165 == _T_5[9:0] ? image_2_357 : _GEN_1508; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1510 = 10'h166 == _T_5[9:0] ? image_2_358 : _GEN_1509; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1511 = 10'h167 == _T_5[9:0] ? image_2_359 : _GEN_1510; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1512 = 10'h168 == _T_5[9:0] ? image_2_360 : _GEN_1511; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1513 = 10'h169 == _T_5[9:0] ? image_2_361 : _GEN_1512; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1514 = 10'h16a == _T_5[9:0] ? image_2_362 : _GEN_1513; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1515 = 10'h16b == _T_5[9:0] ? image_2_363 : _GEN_1514; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1516 = 10'h16c == _T_5[9:0] ? image_2_364 : _GEN_1515; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1517 = 10'h16d == _T_5[9:0] ? image_2_365 : _GEN_1516; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1518 = 10'h16e == _T_5[9:0] ? image_2_366 : _GEN_1517; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1519 = 10'h16f == _T_5[9:0] ? image_2_367 : _GEN_1518; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1520 = 10'h170 == _T_5[9:0] ? image_2_368 : _GEN_1519; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1521 = 10'h171 == _T_5[9:0] ? image_2_369 : _GEN_1520; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1522 = 10'h172 == _T_5[9:0] ? image_2_370 : _GEN_1521; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1523 = 10'h173 == _T_5[9:0] ? image_2_371 : _GEN_1522; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1524 = 10'h174 == _T_5[9:0] ? image_2_372 : _GEN_1523; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1525 = 10'h175 == _T_5[9:0] ? image_2_373 : _GEN_1524; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1526 = 10'h176 == _T_5[9:0] ? image_2_374 : _GEN_1525; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1527 = 10'h177 == _T_5[9:0] ? image_2_375 : _GEN_1526; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1528 = 10'h178 == _T_5[9:0] ? image_2_376 : _GEN_1527; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1529 = 10'h179 == _T_5[9:0] ? image_2_377 : _GEN_1528; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1530 = 10'h17a == _T_5[9:0] ? image_2_378 : _GEN_1529; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1531 = 10'h17b == _T_5[9:0] ? image_2_379 : _GEN_1530; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1532 = 10'h17c == _T_5[9:0] ? image_2_380 : _GEN_1531; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1533 = 10'h17d == _T_5[9:0] ? image_2_381 : _GEN_1532; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1534 = 10'h17e == _T_5[9:0] ? image_2_382 : _GEN_1533; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1535 = 10'h17f == _T_5[9:0] ? image_2_383 : _GEN_1534; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1536 = 10'h180 == _T_5[9:0] ? image_2_384 : _GEN_1535; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1537 = 10'h181 == _T_5[9:0] ? image_2_385 : _GEN_1536; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1538 = 10'h182 == _T_5[9:0] ? image_2_386 : _GEN_1537; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1539 = 10'h183 == _T_5[9:0] ? image_2_387 : _GEN_1538; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1540 = 10'h184 == _T_5[9:0] ? image_2_388 : _GEN_1539; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1541 = 10'h185 == _T_5[9:0] ? image_2_389 : _GEN_1540; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1542 = 10'h186 == _T_5[9:0] ? image_2_390 : _GEN_1541; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1543 = 10'h187 == _T_5[9:0] ? image_2_391 : _GEN_1542; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1544 = 10'h188 == _T_5[9:0] ? image_2_392 : _GEN_1543; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1545 = 10'h189 == _T_5[9:0] ? image_2_393 : _GEN_1544; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1546 = 10'h18a == _T_5[9:0] ? image_2_394 : _GEN_1545; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1547 = 10'h18b == _T_5[9:0] ? image_2_395 : _GEN_1546; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1548 = 10'h18c == _T_5[9:0] ? image_2_396 : _GEN_1547; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1549 = 10'h18d == _T_5[9:0] ? image_2_397 : _GEN_1548; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1550 = 10'h18e == _T_5[9:0] ? image_2_398 : _GEN_1549; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1551 = 10'h18f == _T_5[9:0] ? image_2_399 : _GEN_1550; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1552 = 10'h190 == _T_5[9:0] ? image_2_400 : _GEN_1551; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1553 = 10'h191 == _T_5[9:0] ? image_2_401 : _GEN_1552; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1554 = 10'h192 == _T_5[9:0] ? image_2_402 : _GEN_1553; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1555 = 10'h193 == _T_5[9:0] ? image_2_403 : _GEN_1554; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1556 = 10'h194 == _T_5[9:0] ? image_2_404 : _GEN_1555; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1557 = 10'h195 == _T_5[9:0] ? image_2_405 : _GEN_1556; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1558 = 10'h196 == _T_5[9:0] ? image_2_406 : _GEN_1557; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1559 = 10'h197 == _T_5[9:0] ? image_2_407 : _GEN_1558; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1560 = 10'h198 == _T_5[9:0] ? image_2_408 : _GEN_1559; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1561 = 10'h199 == _T_5[9:0] ? image_2_409 : _GEN_1560; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1562 = 10'h19a == _T_5[9:0] ? image_2_410 : _GEN_1561; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1563 = 10'h19b == _T_5[9:0] ? image_2_411 : _GEN_1562; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1564 = 10'h19c == _T_5[9:0] ? image_2_412 : _GEN_1563; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1565 = 10'h19d == _T_5[9:0] ? image_2_413 : _GEN_1564; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1566 = 10'h19e == _T_5[9:0] ? image_2_414 : _GEN_1565; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1567 = 10'h19f == _T_5[9:0] ? image_2_415 : _GEN_1566; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1568 = 10'h1a0 == _T_5[9:0] ? image_2_416 : _GEN_1567; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1569 = 10'h1a1 == _T_5[9:0] ? image_2_417 : _GEN_1568; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1570 = 10'h1a2 == _T_5[9:0] ? image_2_418 : _GEN_1569; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1571 = 10'h1a3 == _T_5[9:0] ? image_2_419 : _GEN_1570; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1572 = 10'h1a4 == _T_5[9:0] ? image_2_420 : _GEN_1571; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1573 = 10'h1a5 == _T_5[9:0] ? image_2_421 : _GEN_1572; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1574 = 10'h1a6 == _T_5[9:0] ? image_2_422 : _GEN_1573; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1575 = 10'h1a7 == _T_5[9:0] ? image_2_423 : _GEN_1574; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1576 = 10'h1a8 == _T_5[9:0] ? image_2_424 : _GEN_1575; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1577 = 10'h1a9 == _T_5[9:0] ? image_2_425 : _GEN_1576; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1578 = 10'h1aa == _T_5[9:0] ? image_2_426 : _GEN_1577; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1579 = 10'h1ab == _T_5[9:0] ? image_2_427 : _GEN_1578; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1580 = 10'h1ac == _T_5[9:0] ? image_2_428 : _GEN_1579; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1581 = 10'h1ad == _T_5[9:0] ? image_2_429 : _GEN_1580; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1582 = 10'h1ae == _T_5[9:0] ? image_2_430 : _GEN_1581; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1583 = 10'h1af == _T_5[9:0] ? image_2_431 : _GEN_1582; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1584 = 10'h1b0 == _T_5[9:0] ? image_2_432 : _GEN_1583; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1585 = 10'h1b1 == _T_5[9:0] ? image_2_433 : _GEN_1584; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1586 = 10'h1b2 == _T_5[9:0] ? image_2_434 : _GEN_1585; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1587 = 10'h1b3 == _T_5[9:0] ? image_2_435 : _GEN_1586; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1588 = 10'h1b4 == _T_5[9:0] ? image_2_436 : _GEN_1587; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1589 = 10'h1b5 == _T_5[9:0] ? image_2_437 : _GEN_1588; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1590 = 10'h1b6 == _T_5[9:0] ? image_2_438 : _GEN_1589; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1591 = 10'h1b7 == _T_5[9:0] ? image_2_439 : _GEN_1590; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1592 = 10'h1b8 == _T_5[9:0] ? image_2_440 : _GEN_1591; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1593 = 10'h1b9 == _T_5[9:0] ? image_2_441 : _GEN_1592; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1594 = 10'h1ba == _T_5[9:0] ? image_2_442 : _GEN_1593; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1595 = 10'h1bb == _T_5[9:0] ? image_2_443 : _GEN_1594; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1596 = 10'h1bc == _T_5[9:0] ? image_2_444 : _GEN_1595; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1597 = 10'h1bd == _T_5[9:0] ? image_2_445 : _GEN_1596; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1598 = 10'h1be == _T_5[9:0] ? image_2_446 : _GEN_1597; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1599 = 10'h1bf == _T_5[9:0] ? image_2_447 : _GEN_1598; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1600 = 10'h1c0 == _T_5[9:0] ? image_2_448 : _GEN_1599; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1601 = 10'h1c1 == _T_5[9:0] ? image_2_449 : _GEN_1600; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1602 = 10'h1c2 == _T_5[9:0] ? image_2_450 : _GEN_1601; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1603 = 10'h1c3 == _T_5[9:0] ? image_2_451 : _GEN_1602; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1604 = 10'h1c4 == _T_5[9:0] ? image_2_452 : _GEN_1603; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1605 = 10'h1c5 == _T_5[9:0] ? image_2_453 : _GEN_1604; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1606 = 10'h1c6 == _T_5[9:0] ? image_2_454 : _GEN_1605; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1607 = 10'h1c7 == _T_5[9:0] ? image_2_455 : _GEN_1606; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1608 = 10'h1c8 == _T_5[9:0] ? image_2_456 : _GEN_1607; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1609 = 10'h1c9 == _T_5[9:0] ? image_2_457 : _GEN_1608; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1610 = 10'h1ca == _T_5[9:0] ? image_2_458 : _GEN_1609; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1611 = 10'h1cb == _T_5[9:0] ? image_2_459 : _GEN_1610; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1612 = 10'h1cc == _T_5[9:0] ? image_2_460 : _GEN_1611; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1613 = 10'h1cd == _T_5[9:0] ? image_2_461 : _GEN_1612; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1614 = 10'h1ce == _T_5[9:0] ? image_2_462 : _GEN_1613; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1615 = 10'h1cf == _T_5[9:0] ? image_2_463 : _GEN_1614; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1616 = 10'h1d0 == _T_5[9:0] ? image_2_464 : _GEN_1615; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1617 = 10'h1d1 == _T_5[9:0] ? image_2_465 : _GEN_1616; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1618 = 10'h1d2 == _T_5[9:0] ? image_2_466 : _GEN_1617; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1619 = 10'h1d3 == _T_5[9:0] ? image_2_467 : _GEN_1618; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1620 = 10'h1d4 == _T_5[9:0] ? image_2_468 : _GEN_1619; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1621 = 10'h1d5 == _T_5[9:0] ? image_2_469 : _GEN_1620; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1622 = 10'h1d6 == _T_5[9:0] ? image_2_470 : _GEN_1621; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1623 = 10'h1d7 == _T_5[9:0] ? image_2_471 : _GEN_1622; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1624 = 10'h1d8 == _T_5[9:0] ? image_2_472 : _GEN_1623; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1625 = 10'h1d9 == _T_5[9:0] ? image_2_473 : _GEN_1624; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1626 = 10'h1da == _T_5[9:0] ? image_2_474 : _GEN_1625; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1627 = 10'h1db == _T_5[9:0] ? image_2_475 : _GEN_1626; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1628 = 10'h1dc == _T_5[9:0] ? image_2_476 : _GEN_1627; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1629 = 10'h1dd == _T_5[9:0] ? image_2_477 : _GEN_1628; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1630 = 10'h1de == _T_5[9:0] ? image_2_478 : _GEN_1629; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1631 = 10'h1df == _T_5[9:0] ? image_2_479 : _GEN_1630; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1632 = 10'h1e0 == _T_5[9:0] ? image_2_480 : _GEN_1631; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1633 = 10'h1e1 == _T_5[9:0] ? image_2_481 : _GEN_1632; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1634 = 10'h1e2 == _T_5[9:0] ? image_2_482 : _GEN_1633; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1635 = 10'h1e3 == _T_5[9:0] ? image_2_483 : _GEN_1634; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1636 = 10'h1e4 == _T_5[9:0] ? image_2_484 : _GEN_1635; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1637 = 10'h1e5 == _T_5[9:0] ? image_2_485 : _GEN_1636; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1638 = 10'h1e6 == _T_5[9:0] ? image_2_486 : _GEN_1637; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1639 = 10'h1e7 == _T_5[9:0] ? image_2_487 : _GEN_1638; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1640 = 10'h1e8 == _T_5[9:0] ? image_2_488 : _GEN_1639; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1641 = 10'h1e9 == _T_5[9:0] ? image_2_489 : _GEN_1640; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1642 = 10'h1ea == _T_5[9:0] ? image_2_490 : _GEN_1641; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1643 = 10'h1eb == _T_5[9:0] ? image_2_491 : _GEN_1642; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1644 = 10'h1ec == _T_5[9:0] ? image_2_492 : _GEN_1643; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1645 = 10'h1ed == _T_5[9:0] ? image_2_493 : _GEN_1644; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1646 = 10'h1ee == _T_5[9:0] ? image_2_494 : _GEN_1645; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1647 = 10'h1ef == _T_5[9:0] ? image_2_495 : _GEN_1646; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1648 = 10'h1f0 == _T_5[9:0] ? image_2_496 : _GEN_1647; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1649 = 10'h1f1 == _T_5[9:0] ? image_2_497 : _GEN_1648; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1650 = 10'h1f2 == _T_5[9:0] ? image_2_498 : _GEN_1649; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1651 = 10'h1f3 == _T_5[9:0] ? image_2_499 : _GEN_1650; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1652 = 10'h1f4 == _T_5[9:0] ? image_2_500 : _GEN_1651; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1653 = 10'h1f5 == _T_5[9:0] ? image_2_501 : _GEN_1652; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1654 = 10'h1f6 == _T_5[9:0] ? image_2_502 : _GEN_1653; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1655 = 10'h1f7 == _T_5[9:0] ? image_2_503 : _GEN_1654; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1656 = 10'h1f8 == _T_5[9:0] ? image_2_504 : _GEN_1655; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1657 = 10'h1f9 == _T_5[9:0] ? image_2_505 : _GEN_1656; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1658 = 10'h1fa == _T_5[9:0] ? image_2_506 : _GEN_1657; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1659 = 10'h1fb == _T_5[9:0] ? image_2_507 : _GEN_1658; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1660 = 10'h1fc == _T_5[9:0] ? image_2_508 : _GEN_1659; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1661 = 10'h1fd == _T_5[9:0] ? image_2_509 : _GEN_1660; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1662 = 10'h1fe == _T_5[9:0] ? image_2_510 : _GEN_1661; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1663 = 10'h1ff == _T_5[9:0] ? image_2_511 : _GEN_1662; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1664 = 10'h200 == _T_5[9:0] ? image_2_512 : _GEN_1663; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1665 = 10'h201 == _T_5[9:0] ? image_2_513 : _GEN_1664; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1666 = 10'h202 == _T_5[9:0] ? image_2_514 : _GEN_1665; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1667 = 10'h203 == _T_5[9:0] ? image_2_515 : _GEN_1666; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1668 = 10'h204 == _T_5[9:0] ? image_2_516 : _GEN_1667; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1669 = 10'h205 == _T_5[9:0] ? image_2_517 : _GEN_1668; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1670 = 10'h206 == _T_5[9:0] ? image_2_518 : _GEN_1669; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1671 = 10'h207 == _T_5[9:0] ? image_2_519 : _GEN_1670; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1672 = 10'h208 == _T_5[9:0] ? image_2_520 : _GEN_1671; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1673 = 10'h209 == _T_5[9:0] ? image_2_521 : _GEN_1672; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1674 = 10'h20a == _T_5[9:0] ? image_2_522 : _GEN_1673; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1675 = 10'h20b == _T_5[9:0] ? image_2_523 : _GEN_1674; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1676 = 10'h20c == _T_5[9:0] ? image_2_524 : _GEN_1675; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1677 = 10'h20d == _T_5[9:0] ? image_2_525 : _GEN_1676; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1678 = 10'h20e == _T_5[9:0] ? image_2_526 : _GEN_1677; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1679 = 10'h20f == _T_5[9:0] ? image_2_527 : _GEN_1678; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1680 = 10'h210 == _T_5[9:0] ? image_2_528 : _GEN_1679; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1681 = 10'h211 == _T_5[9:0] ? image_2_529 : _GEN_1680; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1682 = 10'h212 == _T_5[9:0] ? image_2_530 : _GEN_1681; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1683 = 10'h213 == _T_5[9:0] ? image_2_531 : _GEN_1682; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1684 = 10'h214 == _T_5[9:0] ? image_2_532 : _GEN_1683; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1685 = 10'h215 == _T_5[9:0] ? image_2_533 : _GEN_1684; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1686 = 10'h216 == _T_5[9:0] ? image_2_534 : _GEN_1685; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1687 = 10'h217 == _T_5[9:0] ? image_2_535 : _GEN_1686; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1688 = 10'h218 == _T_5[9:0] ? image_2_536 : _GEN_1687; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1689 = 10'h219 == _T_5[9:0] ? image_2_537 : _GEN_1688; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1690 = 10'h21a == _T_5[9:0] ? image_2_538 : _GEN_1689; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1691 = 10'h21b == _T_5[9:0] ? image_2_539 : _GEN_1690; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1692 = 10'h21c == _T_5[9:0] ? image_2_540 : _GEN_1691; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1693 = 10'h21d == _T_5[9:0] ? image_2_541 : _GEN_1692; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1694 = 10'h21e == _T_5[9:0] ? image_2_542 : _GEN_1693; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1695 = 10'h21f == _T_5[9:0] ? image_2_543 : _GEN_1694; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1696 = 10'h220 == _T_5[9:0] ? image_2_544 : _GEN_1695; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1697 = 10'h221 == _T_5[9:0] ? image_2_545 : _GEN_1696; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1698 = 10'h222 == _T_5[9:0] ? image_2_546 : _GEN_1697; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1699 = 10'h223 == _T_5[9:0] ? image_2_547 : _GEN_1698; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1700 = 10'h224 == _T_5[9:0] ? image_2_548 : _GEN_1699; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1701 = 10'h225 == _T_5[9:0] ? image_2_549 : _GEN_1700; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1702 = 10'h226 == _T_5[9:0] ? image_2_550 : _GEN_1701; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1703 = 10'h227 == _T_5[9:0] ? image_2_551 : _GEN_1702; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1704 = 10'h228 == _T_5[9:0] ? image_2_552 : _GEN_1703; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1705 = 10'h229 == _T_5[9:0] ? image_2_553 : _GEN_1704; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1706 = 10'h22a == _T_5[9:0] ? image_2_554 : _GEN_1705; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1707 = 10'h22b == _T_5[9:0] ? image_2_555 : _GEN_1706; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1708 = 10'h22c == _T_5[9:0] ? image_2_556 : _GEN_1707; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1709 = 10'h22d == _T_5[9:0] ? image_2_557 : _GEN_1708; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1710 = 10'h22e == _T_5[9:0] ? image_2_558 : _GEN_1709; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1711 = 10'h22f == _T_5[9:0] ? image_2_559 : _GEN_1710; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1712 = 10'h230 == _T_5[9:0] ? image_2_560 : _GEN_1711; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1713 = 10'h231 == _T_5[9:0] ? image_2_561 : _GEN_1712; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1714 = 10'h232 == _T_5[9:0] ? image_2_562 : _GEN_1713; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1715 = 10'h233 == _T_5[9:0] ? image_2_563 : _GEN_1714; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1716 = 10'h234 == _T_5[9:0] ? image_2_564 : _GEN_1715; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1717 = 10'h235 == _T_5[9:0] ? image_2_565 : _GEN_1716; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1718 = 10'h236 == _T_5[9:0] ? image_2_566 : _GEN_1717; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1719 = 10'h237 == _T_5[9:0] ? image_2_567 : _GEN_1718; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1720 = 10'h238 == _T_5[9:0] ? image_2_568 : _GEN_1719; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1721 = 10'h239 == _T_5[9:0] ? image_2_569 : _GEN_1720; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1722 = 10'h23a == _T_5[9:0] ? image_2_570 : _GEN_1721; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1723 = 10'h23b == _T_5[9:0] ? image_2_571 : _GEN_1722; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1724 = 10'h23c == _T_5[9:0] ? image_2_572 : _GEN_1723; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1725 = 10'h23d == _T_5[9:0] ? image_2_573 : _GEN_1724; // @[VideoBuffer.scala 27:30]
  wire [3:0] _GEN_1726 = 10'h23e == _T_5[9:0] ? image_2_574 : _GEN_1725; // @[VideoBuffer.scala 27:30]
  wire [32:0] _T_15 = {{1'd0}, pixelIndex}; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_19 = pixelIndex + 32'h1; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_22 = pixelIndex + 32'h2; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_25 = pixelIndex + 32'h3; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_28 = pixelIndex + 32'h4; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_31 = pixelIndex + 32'h5; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_34 = pixelIndex + 32'h6; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_37 = pixelIndex + 32'h7; // @[VideoBuffer.scala 33:35]
  wire [31:0] _T_88 = pixelIndex + 32'h8; // @[VideoBuffer.scala 36:34]
  wire [10:0] _T_89 = 6'h20 * 6'h12; // @[VideoBuffer.scala 37:42]
  wire [31:0] _GEN_17285 = {{21'd0}, _T_89}; // @[VideoBuffer.scala 37:25]
  wire  _T_90 = pixelIndex == _GEN_17285; // @[VideoBuffer.scala 37:25]
  assign io_pixelVal_out_0 = 10'h23f == _T_5[9:0] ? image_0_575 : _GEN_574; // @[VideoBuffer.scala 27:30]
  assign io_pixelVal_out_1 = 10'h23f == _T_5[9:0] ? image_1_575 : _GEN_1150; // @[VideoBuffer.scala 27:30]
  assign io_pixelVal_out_2 = 10'h23f == _T_5[9:0] ? image_2_575 : _GEN_1726; // @[VideoBuffer.scala 27:30]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  image_0_0 = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  image_0_1 = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  image_0_2 = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  image_0_3 = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  image_0_4 = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  image_0_5 = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  image_0_6 = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  image_0_7 = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  image_0_8 = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  image_0_9 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  image_0_10 = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  image_0_11 = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  image_0_12 = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  image_0_13 = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  image_0_14 = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  image_0_15 = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  image_0_16 = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  image_0_17 = _RAND_17[3:0];
  _RAND_18 = {1{`RANDOM}};
  image_0_18 = _RAND_18[3:0];
  _RAND_19 = {1{`RANDOM}};
  image_0_19 = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  image_0_20 = _RAND_20[3:0];
  _RAND_21 = {1{`RANDOM}};
  image_0_21 = _RAND_21[3:0];
  _RAND_22 = {1{`RANDOM}};
  image_0_22 = _RAND_22[3:0];
  _RAND_23 = {1{`RANDOM}};
  image_0_23 = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
  image_0_24 = _RAND_24[3:0];
  _RAND_25 = {1{`RANDOM}};
  image_0_25 = _RAND_25[3:0];
  _RAND_26 = {1{`RANDOM}};
  image_0_26 = _RAND_26[3:0];
  _RAND_27 = {1{`RANDOM}};
  image_0_27 = _RAND_27[3:0];
  _RAND_28 = {1{`RANDOM}};
  image_0_28 = _RAND_28[3:0];
  _RAND_29 = {1{`RANDOM}};
  image_0_29 = _RAND_29[3:0];
  _RAND_30 = {1{`RANDOM}};
  image_0_30 = _RAND_30[3:0];
  _RAND_31 = {1{`RANDOM}};
  image_0_31 = _RAND_31[3:0];
  _RAND_32 = {1{`RANDOM}};
  image_0_32 = _RAND_32[3:0];
  _RAND_33 = {1{`RANDOM}};
  image_0_33 = _RAND_33[3:0];
  _RAND_34 = {1{`RANDOM}};
  image_0_34 = _RAND_34[3:0];
  _RAND_35 = {1{`RANDOM}};
  image_0_35 = _RAND_35[3:0];
  _RAND_36 = {1{`RANDOM}};
  image_0_36 = _RAND_36[3:0];
  _RAND_37 = {1{`RANDOM}};
  image_0_37 = _RAND_37[3:0];
  _RAND_38 = {1{`RANDOM}};
  image_0_38 = _RAND_38[3:0];
  _RAND_39 = {1{`RANDOM}};
  image_0_39 = _RAND_39[3:0];
  _RAND_40 = {1{`RANDOM}};
  image_0_40 = _RAND_40[3:0];
  _RAND_41 = {1{`RANDOM}};
  image_0_41 = _RAND_41[3:0];
  _RAND_42 = {1{`RANDOM}};
  image_0_42 = _RAND_42[3:0];
  _RAND_43 = {1{`RANDOM}};
  image_0_43 = _RAND_43[3:0];
  _RAND_44 = {1{`RANDOM}};
  image_0_44 = _RAND_44[3:0];
  _RAND_45 = {1{`RANDOM}};
  image_0_45 = _RAND_45[3:0];
  _RAND_46 = {1{`RANDOM}};
  image_0_46 = _RAND_46[3:0];
  _RAND_47 = {1{`RANDOM}};
  image_0_47 = _RAND_47[3:0];
  _RAND_48 = {1{`RANDOM}};
  image_0_48 = _RAND_48[3:0];
  _RAND_49 = {1{`RANDOM}};
  image_0_49 = _RAND_49[3:0];
  _RAND_50 = {1{`RANDOM}};
  image_0_50 = _RAND_50[3:0];
  _RAND_51 = {1{`RANDOM}};
  image_0_51 = _RAND_51[3:0];
  _RAND_52 = {1{`RANDOM}};
  image_0_52 = _RAND_52[3:0];
  _RAND_53 = {1{`RANDOM}};
  image_0_53 = _RAND_53[3:0];
  _RAND_54 = {1{`RANDOM}};
  image_0_54 = _RAND_54[3:0];
  _RAND_55 = {1{`RANDOM}};
  image_0_55 = _RAND_55[3:0];
  _RAND_56 = {1{`RANDOM}};
  image_0_56 = _RAND_56[3:0];
  _RAND_57 = {1{`RANDOM}};
  image_0_57 = _RAND_57[3:0];
  _RAND_58 = {1{`RANDOM}};
  image_0_58 = _RAND_58[3:0];
  _RAND_59 = {1{`RANDOM}};
  image_0_59 = _RAND_59[3:0];
  _RAND_60 = {1{`RANDOM}};
  image_0_60 = _RAND_60[3:0];
  _RAND_61 = {1{`RANDOM}};
  image_0_61 = _RAND_61[3:0];
  _RAND_62 = {1{`RANDOM}};
  image_0_62 = _RAND_62[3:0];
  _RAND_63 = {1{`RANDOM}};
  image_0_63 = _RAND_63[3:0];
  _RAND_64 = {1{`RANDOM}};
  image_0_64 = _RAND_64[3:0];
  _RAND_65 = {1{`RANDOM}};
  image_0_65 = _RAND_65[3:0];
  _RAND_66 = {1{`RANDOM}};
  image_0_66 = _RAND_66[3:0];
  _RAND_67 = {1{`RANDOM}};
  image_0_67 = _RAND_67[3:0];
  _RAND_68 = {1{`RANDOM}};
  image_0_68 = _RAND_68[3:0];
  _RAND_69 = {1{`RANDOM}};
  image_0_69 = _RAND_69[3:0];
  _RAND_70 = {1{`RANDOM}};
  image_0_70 = _RAND_70[3:0];
  _RAND_71 = {1{`RANDOM}};
  image_0_71 = _RAND_71[3:0];
  _RAND_72 = {1{`RANDOM}};
  image_0_72 = _RAND_72[3:0];
  _RAND_73 = {1{`RANDOM}};
  image_0_73 = _RAND_73[3:0];
  _RAND_74 = {1{`RANDOM}};
  image_0_74 = _RAND_74[3:0];
  _RAND_75 = {1{`RANDOM}};
  image_0_75 = _RAND_75[3:0];
  _RAND_76 = {1{`RANDOM}};
  image_0_76 = _RAND_76[3:0];
  _RAND_77 = {1{`RANDOM}};
  image_0_77 = _RAND_77[3:0];
  _RAND_78 = {1{`RANDOM}};
  image_0_78 = _RAND_78[3:0];
  _RAND_79 = {1{`RANDOM}};
  image_0_79 = _RAND_79[3:0];
  _RAND_80 = {1{`RANDOM}};
  image_0_80 = _RAND_80[3:0];
  _RAND_81 = {1{`RANDOM}};
  image_0_81 = _RAND_81[3:0];
  _RAND_82 = {1{`RANDOM}};
  image_0_82 = _RAND_82[3:0];
  _RAND_83 = {1{`RANDOM}};
  image_0_83 = _RAND_83[3:0];
  _RAND_84 = {1{`RANDOM}};
  image_0_84 = _RAND_84[3:0];
  _RAND_85 = {1{`RANDOM}};
  image_0_85 = _RAND_85[3:0];
  _RAND_86 = {1{`RANDOM}};
  image_0_86 = _RAND_86[3:0];
  _RAND_87 = {1{`RANDOM}};
  image_0_87 = _RAND_87[3:0];
  _RAND_88 = {1{`RANDOM}};
  image_0_88 = _RAND_88[3:0];
  _RAND_89 = {1{`RANDOM}};
  image_0_89 = _RAND_89[3:0];
  _RAND_90 = {1{`RANDOM}};
  image_0_90 = _RAND_90[3:0];
  _RAND_91 = {1{`RANDOM}};
  image_0_91 = _RAND_91[3:0];
  _RAND_92 = {1{`RANDOM}};
  image_0_92 = _RAND_92[3:0];
  _RAND_93 = {1{`RANDOM}};
  image_0_93 = _RAND_93[3:0];
  _RAND_94 = {1{`RANDOM}};
  image_0_94 = _RAND_94[3:0];
  _RAND_95 = {1{`RANDOM}};
  image_0_95 = _RAND_95[3:0];
  _RAND_96 = {1{`RANDOM}};
  image_0_96 = _RAND_96[3:0];
  _RAND_97 = {1{`RANDOM}};
  image_0_97 = _RAND_97[3:0];
  _RAND_98 = {1{`RANDOM}};
  image_0_98 = _RAND_98[3:0];
  _RAND_99 = {1{`RANDOM}};
  image_0_99 = _RAND_99[3:0];
  _RAND_100 = {1{`RANDOM}};
  image_0_100 = _RAND_100[3:0];
  _RAND_101 = {1{`RANDOM}};
  image_0_101 = _RAND_101[3:0];
  _RAND_102 = {1{`RANDOM}};
  image_0_102 = _RAND_102[3:0];
  _RAND_103 = {1{`RANDOM}};
  image_0_103 = _RAND_103[3:0];
  _RAND_104 = {1{`RANDOM}};
  image_0_104 = _RAND_104[3:0];
  _RAND_105 = {1{`RANDOM}};
  image_0_105 = _RAND_105[3:0];
  _RAND_106 = {1{`RANDOM}};
  image_0_106 = _RAND_106[3:0];
  _RAND_107 = {1{`RANDOM}};
  image_0_107 = _RAND_107[3:0];
  _RAND_108 = {1{`RANDOM}};
  image_0_108 = _RAND_108[3:0];
  _RAND_109 = {1{`RANDOM}};
  image_0_109 = _RAND_109[3:0];
  _RAND_110 = {1{`RANDOM}};
  image_0_110 = _RAND_110[3:0];
  _RAND_111 = {1{`RANDOM}};
  image_0_111 = _RAND_111[3:0];
  _RAND_112 = {1{`RANDOM}};
  image_0_112 = _RAND_112[3:0];
  _RAND_113 = {1{`RANDOM}};
  image_0_113 = _RAND_113[3:0];
  _RAND_114 = {1{`RANDOM}};
  image_0_114 = _RAND_114[3:0];
  _RAND_115 = {1{`RANDOM}};
  image_0_115 = _RAND_115[3:0];
  _RAND_116 = {1{`RANDOM}};
  image_0_116 = _RAND_116[3:0];
  _RAND_117 = {1{`RANDOM}};
  image_0_117 = _RAND_117[3:0];
  _RAND_118 = {1{`RANDOM}};
  image_0_118 = _RAND_118[3:0];
  _RAND_119 = {1{`RANDOM}};
  image_0_119 = _RAND_119[3:0];
  _RAND_120 = {1{`RANDOM}};
  image_0_120 = _RAND_120[3:0];
  _RAND_121 = {1{`RANDOM}};
  image_0_121 = _RAND_121[3:0];
  _RAND_122 = {1{`RANDOM}};
  image_0_122 = _RAND_122[3:0];
  _RAND_123 = {1{`RANDOM}};
  image_0_123 = _RAND_123[3:0];
  _RAND_124 = {1{`RANDOM}};
  image_0_124 = _RAND_124[3:0];
  _RAND_125 = {1{`RANDOM}};
  image_0_125 = _RAND_125[3:0];
  _RAND_126 = {1{`RANDOM}};
  image_0_126 = _RAND_126[3:0];
  _RAND_127 = {1{`RANDOM}};
  image_0_127 = _RAND_127[3:0];
  _RAND_128 = {1{`RANDOM}};
  image_0_128 = _RAND_128[3:0];
  _RAND_129 = {1{`RANDOM}};
  image_0_129 = _RAND_129[3:0];
  _RAND_130 = {1{`RANDOM}};
  image_0_130 = _RAND_130[3:0];
  _RAND_131 = {1{`RANDOM}};
  image_0_131 = _RAND_131[3:0];
  _RAND_132 = {1{`RANDOM}};
  image_0_132 = _RAND_132[3:0];
  _RAND_133 = {1{`RANDOM}};
  image_0_133 = _RAND_133[3:0];
  _RAND_134 = {1{`RANDOM}};
  image_0_134 = _RAND_134[3:0];
  _RAND_135 = {1{`RANDOM}};
  image_0_135 = _RAND_135[3:0];
  _RAND_136 = {1{`RANDOM}};
  image_0_136 = _RAND_136[3:0];
  _RAND_137 = {1{`RANDOM}};
  image_0_137 = _RAND_137[3:0];
  _RAND_138 = {1{`RANDOM}};
  image_0_138 = _RAND_138[3:0];
  _RAND_139 = {1{`RANDOM}};
  image_0_139 = _RAND_139[3:0];
  _RAND_140 = {1{`RANDOM}};
  image_0_140 = _RAND_140[3:0];
  _RAND_141 = {1{`RANDOM}};
  image_0_141 = _RAND_141[3:0];
  _RAND_142 = {1{`RANDOM}};
  image_0_142 = _RAND_142[3:0];
  _RAND_143 = {1{`RANDOM}};
  image_0_143 = _RAND_143[3:0];
  _RAND_144 = {1{`RANDOM}};
  image_0_144 = _RAND_144[3:0];
  _RAND_145 = {1{`RANDOM}};
  image_0_145 = _RAND_145[3:0];
  _RAND_146 = {1{`RANDOM}};
  image_0_146 = _RAND_146[3:0];
  _RAND_147 = {1{`RANDOM}};
  image_0_147 = _RAND_147[3:0];
  _RAND_148 = {1{`RANDOM}};
  image_0_148 = _RAND_148[3:0];
  _RAND_149 = {1{`RANDOM}};
  image_0_149 = _RAND_149[3:0];
  _RAND_150 = {1{`RANDOM}};
  image_0_150 = _RAND_150[3:0];
  _RAND_151 = {1{`RANDOM}};
  image_0_151 = _RAND_151[3:0];
  _RAND_152 = {1{`RANDOM}};
  image_0_152 = _RAND_152[3:0];
  _RAND_153 = {1{`RANDOM}};
  image_0_153 = _RAND_153[3:0];
  _RAND_154 = {1{`RANDOM}};
  image_0_154 = _RAND_154[3:0];
  _RAND_155 = {1{`RANDOM}};
  image_0_155 = _RAND_155[3:0];
  _RAND_156 = {1{`RANDOM}};
  image_0_156 = _RAND_156[3:0];
  _RAND_157 = {1{`RANDOM}};
  image_0_157 = _RAND_157[3:0];
  _RAND_158 = {1{`RANDOM}};
  image_0_158 = _RAND_158[3:0];
  _RAND_159 = {1{`RANDOM}};
  image_0_159 = _RAND_159[3:0];
  _RAND_160 = {1{`RANDOM}};
  image_0_160 = _RAND_160[3:0];
  _RAND_161 = {1{`RANDOM}};
  image_0_161 = _RAND_161[3:0];
  _RAND_162 = {1{`RANDOM}};
  image_0_162 = _RAND_162[3:0];
  _RAND_163 = {1{`RANDOM}};
  image_0_163 = _RAND_163[3:0];
  _RAND_164 = {1{`RANDOM}};
  image_0_164 = _RAND_164[3:0];
  _RAND_165 = {1{`RANDOM}};
  image_0_165 = _RAND_165[3:0];
  _RAND_166 = {1{`RANDOM}};
  image_0_166 = _RAND_166[3:0];
  _RAND_167 = {1{`RANDOM}};
  image_0_167 = _RAND_167[3:0];
  _RAND_168 = {1{`RANDOM}};
  image_0_168 = _RAND_168[3:0];
  _RAND_169 = {1{`RANDOM}};
  image_0_169 = _RAND_169[3:0];
  _RAND_170 = {1{`RANDOM}};
  image_0_170 = _RAND_170[3:0];
  _RAND_171 = {1{`RANDOM}};
  image_0_171 = _RAND_171[3:0];
  _RAND_172 = {1{`RANDOM}};
  image_0_172 = _RAND_172[3:0];
  _RAND_173 = {1{`RANDOM}};
  image_0_173 = _RAND_173[3:0];
  _RAND_174 = {1{`RANDOM}};
  image_0_174 = _RAND_174[3:0];
  _RAND_175 = {1{`RANDOM}};
  image_0_175 = _RAND_175[3:0];
  _RAND_176 = {1{`RANDOM}};
  image_0_176 = _RAND_176[3:0];
  _RAND_177 = {1{`RANDOM}};
  image_0_177 = _RAND_177[3:0];
  _RAND_178 = {1{`RANDOM}};
  image_0_178 = _RAND_178[3:0];
  _RAND_179 = {1{`RANDOM}};
  image_0_179 = _RAND_179[3:0];
  _RAND_180 = {1{`RANDOM}};
  image_0_180 = _RAND_180[3:0];
  _RAND_181 = {1{`RANDOM}};
  image_0_181 = _RAND_181[3:0];
  _RAND_182 = {1{`RANDOM}};
  image_0_182 = _RAND_182[3:0];
  _RAND_183 = {1{`RANDOM}};
  image_0_183 = _RAND_183[3:0];
  _RAND_184 = {1{`RANDOM}};
  image_0_184 = _RAND_184[3:0];
  _RAND_185 = {1{`RANDOM}};
  image_0_185 = _RAND_185[3:0];
  _RAND_186 = {1{`RANDOM}};
  image_0_186 = _RAND_186[3:0];
  _RAND_187 = {1{`RANDOM}};
  image_0_187 = _RAND_187[3:0];
  _RAND_188 = {1{`RANDOM}};
  image_0_188 = _RAND_188[3:0];
  _RAND_189 = {1{`RANDOM}};
  image_0_189 = _RAND_189[3:0];
  _RAND_190 = {1{`RANDOM}};
  image_0_190 = _RAND_190[3:0];
  _RAND_191 = {1{`RANDOM}};
  image_0_191 = _RAND_191[3:0];
  _RAND_192 = {1{`RANDOM}};
  image_0_192 = _RAND_192[3:0];
  _RAND_193 = {1{`RANDOM}};
  image_0_193 = _RAND_193[3:0];
  _RAND_194 = {1{`RANDOM}};
  image_0_194 = _RAND_194[3:0];
  _RAND_195 = {1{`RANDOM}};
  image_0_195 = _RAND_195[3:0];
  _RAND_196 = {1{`RANDOM}};
  image_0_196 = _RAND_196[3:0];
  _RAND_197 = {1{`RANDOM}};
  image_0_197 = _RAND_197[3:0];
  _RAND_198 = {1{`RANDOM}};
  image_0_198 = _RAND_198[3:0];
  _RAND_199 = {1{`RANDOM}};
  image_0_199 = _RAND_199[3:0];
  _RAND_200 = {1{`RANDOM}};
  image_0_200 = _RAND_200[3:0];
  _RAND_201 = {1{`RANDOM}};
  image_0_201 = _RAND_201[3:0];
  _RAND_202 = {1{`RANDOM}};
  image_0_202 = _RAND_202[3:0];
  _RAND_203 = {1{`RANDOM}};
  image_0_203 = _RAND_203[3:0];
  _RAND_204 = {1{`RANDOM}};
  image_0_204 = _RAND_204[3:0];
  _RAND_205 = {1{`RANDOM}};
  image_0_205 = _RAND_205[3:0];
  _RAND_206 = {1{`RANDOM}};
  image_0_206 = _RAND_206[3:0];
  _RAND_207 = {1{`RANDOM}};
  image_0_207 = _RAND_207[3:0];
  _RAND_208 = {1{`RANDOM}};
  image_0_208 = _RAND_208[3:0];
  _RAND_209 = {1{`RANDOM}};
  image_0_209 = _RAND_209[3:0];
  _RAND_210 = {1{`RANDOM}};
  image_0_210 = _RAND_210[3:0];
  _RAND_211 = {1{`RANDOM}};
  image_0_211 = _RAND_211[3:0];
  _RAND_212 = {1{`RANDOM}};
  image_0_212 = _RAND_212[3:0];
  _RAND_213 = {1{`RANDOM}};
  image_0_213 = _RAND_213[3:0];
  _RAND_214 = {1{`RANDOM}};
  image_0_214 = _RAND_214[3:0];
  _RAND_215 = {1{`RANDOM}};
  image_0_215 = _RAND_215[3:0];
  _RAND_216 = {1{`RANDOM}};
  image_0_216 = _RAND_216[3:0];
  _RAND_217 = {1{`RANDOM}};
  image_0_217 = _RAND_217[3:0];
  _RAND_218 = {1{`RANDOM}};
  image_0_218 = _RAND_218[3:0];
  _RAND_219 = {1{`RANDOM}};
  image_0_219 = _RAND_219[3:0];
  _RAND_220 = {1{`RANDOM}};
  image_0_220 = _RAND_220[3:0];
  _RAND_221 = {1{`RANDOM}};
  image_0_221 = _RAND_221[3:0];
  _RAND_222 = {1{`RANDOM}};
  image_0_222 = _RAND_222[3:0];
  _RAND_223 = {1{`RANDOM}};
  image_0_223 = _RAND_223[3:0];
  _RAND_224 = {1{`RANDOM}};
  image_0_224 = _RAND_224[3:0];
  _RAND_225 = {1{`RANDOM}};
  image_0_225 = _RAND_225[3:0];
  _RAND_226 = {1{`RANDOM}};
  image_0_226 = _RAND_226[3:0];
  _RAND_227 = {1{`RANDOM}};
  image_0_227 = _RAND_227[3:0];
  _RAND_228 = {1{`RANDOM}};
  image_0_228 = _RAND_228[3:0];
  _RAND_229 = {1{`RANDOM}};
  image_0_229 = _RAND_229[3:0];
  _RAND_230 = {1{`RANDOM}};
  image_0_230 = _RAND_230[3:0];
  _RAND_231 = {1{`RANDOM}};
  image_0_231 = _RAND_231[3:0];
  _RAND_232 = {1{`RANDOM}};
  image_0_232 = _RAND_232[3:0];
  _RAND_233 = {1{`RANDOM}};
  image_0_233 = _RAND_233[3:0];
  _RAND_234 = {1{`RANDOM}};
  image_0_234 = _RAND_234[3:0];
  _RAND_235 = {1{`RANDOM}};
  image_0_235 = _RAND_235[3:0];
  _RAND_236 = {1{`RANDOM}};
  image_0_236 = _RAND_236[3:0];
  _RAND_237 = {1{`RANDOM}};
  image_0_237 = _RAND_237[3:0];
  _RAND_238 = {1{`RANDOM}};
  image_0_238 = _RAND_238[3:0];
  _RAND_239 = {1{`RANDOM}};
  image_0_239 = _RAND_239[3:0];
  _RAND_240 = {1{`RANDOM}};
  image_0_240 = _RAND_240[3:0];
  _RAND_241 = {1{`RANDOM}};
  image_0_241 = _RAND_241[3:0];
  _RAND_242 = {1{`RANDOM}};
  image_0_242 = _RAND_242[3:0];
  _RAND_243 = {1{`RANDOM}};
  image_0_243 = _RAND_243[3:0];
  _RAND_244 = {1{`RANDOM}};
  image_0_244 = _RAND_244[3:0];
  _RAND_245 = {1{`RANDOM}};
  image_0_245 = _RAND_245[3:0];
  _RAND_246 = {1{`RANDOM}};
  image_0_246 = _RAND_246[3:0];
  _RAND_247 = {1{`RANDOM}};
  image_0_247 = _RAND_247[3:0];
  _RAND_248 = {1{`RANDOM}};
  image_0_248 = _RAND_248[3:0];
  _RAND_249 = {1{`RANDOM}};
  image_0_249 = _RAND_249[3:0];
  _RAND_250 = {1{`RANDOM}};
  image_0_250 = _RAND_250[3:0];
  _RAND_251 = {1{`RANDOM}};
  image_0_251 = _RAND_251[3:0];
  _RAND_252 = {1{`RANDOM}};
  image_0_252 = _RAND_252[3:0];
  _RAND_253 = {1{`RANDOM}};
  image_0_253 = _RAND_253[3:0];
  _RAND_254 = {1{`RANDOM}};
  image_0_254 = _RAND_254[3:0];
  _RAND_255 = {1{`RANDOM}};
  image_0_255 = _RAND_255[3:0];
  _RAND_256 = {1{`RANDOM}};
  image_0_256 = _RAND_256[3:0];
  _RAND_257 = {1{`RANDOM}};
  image_0_257 = _RAND_257[3:0];
  _RAND_258 = {1{`RANDOM}};
  image_0_258 = _RAND_258[3:0];
  _RAND_259 = {1{`RANDOM}};
  image_0_259 = _RAND_259[3:0];
  _RAND_260 = {1{`RANDOM}};
  image_0_260 = _RAND_260[3:0];
  _RAND_261 = {1{`RANDOM}};
  image_0_261 = _RAND_261[3:0];
  _RAND_262 = {1{`RANDOM}};
  image_0_262 = _RAND_262[3:0];
  _RAND_263 = {1{`RANDOM}};
  image_0_263 = _RAND_263[3:0];
  _RAND_264 = {1{`RANDOM}};
  image_0_264 = _RAND_264[3:0];
  _RAND_265 = {1{`RANDOM}};
  image_0_265 = _RAND_265[3:0];
  _RAND_266 = {1{`RANDOM}};
  image_0_266 = _RAND_266[3:0];
  _RAND_267 = {1{`RANDOM}};
  image_0_267 = _RAND_267[3:0];
  _RAND_268 = {1{`RANDOM}};
  image_0_268 = _RAND_268[3:0];
  _RAND_269 = {1{`RANDOM}};
  image_0_269 = _RAND_269[3:0];
  _RAND_270 = {1{`RANDOM}};
  image_0_270 = _RAND_270[3:0];
  _RAND_271 = {1{`RANDOM}};
  image_0_271 = _RAND_271[3:0];
  _RAND_272 = {1{`RANDOM}};
  image_0_272 = _RAND_272[3:0];
  _RAND_273 = {1{`RANDOM}};
  image_0_273 = _RAND_273[3:0];
  _RAND_274 = {1{`RANDOM}};
  image_0_274 = _RAND_274[3:0];
  _RAND_275 = {1{`RANDOM}};
  image_0_275 = _RAND_275[3:0];
  _RAND_276 = {1{`RANDOM}};
  image_0_276 = _RAND_276[3:0];
  _RAND_277 = {1{`RANDOM}};
  image_0_277 = _RAND_277[3:0];
  _RAND_278 = {1{`RANDOM}};
  image_0_278 = _RAND_278[3:0];
  _RAND_279 = {1{`RANDOM}};
  image_0_279 = _RAND_279[3:0];
  _RAND_280 = {1{`RANDOM}};
  image_0_280 = _RAND_280[3:0];
  _RAND_281 = {1{`RANDOM}};
  image_0_281 = _RAND_281[3:0];
  _RAND_282 = {1{`RANDOM}};
  image_0_282 = _RAND_282[3:0];
  _RAND_283 = {1{`RANDOM}};
  image_0_283 = _RAND_283[3:0];
  _RAND_284 = {1{`RANDOM}};
  image_0_284 = _RAND_284[3:0];
  _RAND_285 = {1{`RANDOM}};
  image_0_285 = _RAND_285[3:0];
  _RAND_286 = {1{`RANDOM}};
  image_0_286 = _RAND_286[3:0];
  _RAND_287 = {1{`RANDOM}};
  image_0_287 = _RAND_287[3:0];
  _RAND_288 = {1{`RANDOM}};
  image_0_288 = _RAND_288[3:0];
  _RAND_289 = {1{`RANDOM}};
  image_0_289 = _RAND_289[3:0];
  _RAND_290 = {1{`RANDOM}};
  image_0_290 = _RAND_290[3:0];
  _RAND_291 = {1{`RANDOM}};
  image_0_291 = _RAND_291[3:0];
  _RAND_292 = {1{`RANDOM}};
  image_0_292 = _RAND_292[3:0];
  _RAND_293 = {1{`RANDOM}};
  image_0_293 = _RAND_293[3:0];
  _RAND_294 = {1{`RANDOM}};
  image_0_294 = _RAND_294[3:0];
  _RAND_295 = {1{`RANDOM}};
  image_0_295 = _RAND_295[3:0];
  _RAND_296 = {1{`RANDOM}};
  image_0_296 = _RAND_296[3:0];
  _RAND_297 = {1{`RANDOM}};
  image_0_297 = _RAND_297[3:0];
  _RAND_298 = {1{`RANDOM}};
  image_0_298 = _RAND_298[3:0];
  _RAND_299 = {1{`RANDOM}};
  image_0_299 = _RAND_299[3:0];
  _RAND_300 = {1{`RANDOM}};
  image_0_300 = _RAND_300[3:0];
  _RAND_301 = {1{`RANDOM}};
  image_0_301 = _RAND_301[3:0];
  _RAND_302 = {1{`RANDOM}};
  image_0_302 = _RAND_302[3:0];
  _RAND_303 = {1{`RANDOM}};
  image_0_303 = _RAND_303[3:0];
  _RAND_304 = {1{`RANDOM}};
  image_0_304 = _RAND_304[3:0];
  _RAND_305 = {1{`RANDOM}};
  image_0_305 = _RAND_305[3:0];
  _RAND_306 = {1{`RANDOM}};
  image_0_306 = _RAND_306[3:0];
  _RAND_307 = {1{`RANDOM}};
  image_0_307 = _RAND_307[3:0];
  _RAND_308 = {1{`RANDOM}};
  image_0_308 = _RAND_308[3:0];
  _RAND_309 = {1{`RANDOM}};
  image_0_309 = _RAND_309[3:0];
  _RAND_310 = {1{`RANDOM}};
  image_0_310 = _RAND_310[3:0];
  _RAND_311 = {1{`RANDOM}};
  image_0_311 = _RAND_311[3:0];
  _RAND_312 = {1{`RANDOM}};
  image_0_312 = _RAND_312[3:0];
  _RAND_313 = {1{`RANDOM}};
  image_0_313 = _RAND_313[3:0];
  _RAND_314 = {1{`RANDOM}};
  image_0_314 = _RAND_314[3:0];
  _RAND_315 = {1{`RANDOM}};
  image_0_315 = _RAND_315[3:0];
  _RAND_316 = {1{`RANDOM}};
  image_0_316 = _RAND_316[3:0];
  _RAND_317 = {1{`RANDOM}};
  image_0_317 = _RAND_317[3:0];
  _RAND_318 = {1{`RANDOM}};
  image_0_318 = _RAND_318[3:0];
  _RAND_319 = {1{`RANDOM}};
  image_0_319 = _RAND_319[3:0];
  _RAND_320 = {1{`RANDOM}};
  image_0_320 = _RAND_320[3:0];
  _RAND_321 = {1{`RANDOM}};
  image_0_321 = _RAND_321[3:0];
  _RAND_322 = {1{`RANDOM}};
  image_0_322 = _RAND_322[3:0];
  _RAND_323 = {1{`RANDOM}};
  image_0_323 = _RAND_323[3:0];
  _RAND_324 = {1{`RANDOM}};
  image_0_324 = _RAND_324[3:0];
  _RAND_325 = {1{`RANDOM}};
  image_0_325 = _RAND_325[3:0];
  _RAND_326 = {1{`RANDOM}};
  image_0_326 = _RAND_326[3:0];
  _RAND_327 = {1{`RANDOM}};
  image_0_327 = _RAND_327[3:0];
  _RAND_328 = {1{`RANDOM}};
  image_0_328 = _RAND_328[3:0];
  _RAND_329 = {1{`RANDOM}};
  image_0_329 = _RAND_329[3:0];
  _RAND_330 = {1{`RANDOM}};
  image_0_330 = _RAND_330[3:0];
  _RAND_331 = {1{`RANDOM}};
  image_0_331 = _RAND_331[3:0];
  _RAND_332 = {1{`RANDOM}};
  image_0_332 = _RAND_332[3:0];
  _RAND_333 = {1{`RANDOM}};
  image_0_333 = _RAND_333[3:0];
  _RAND_334 = {1{`RANDOM}};
  image_0_334 = _RAND_334[3:0];
  _RAND_335 = {1{`RANDOM}};
  image_0_335 = _RAND_335[3:0];
  _RAND_336 = {1{`RANDOM}};
  image_0_336 = _RAND_336[3:0];
  _RAND_337 = {1{`RANDOM}};
  image_0_337 = _RAND_337[3:0];
  _RAND_338 = {1{`RANDOM}};
  image_0_338 = _RAND_338[3:0];
  _RAND_339 = {1{`RANDOM}};
  image_0_339 = _RAND_339[3:0];
  _RAND_340 = {1{`RANDOM}};
  image_0_340 = _RAND_340[3:0];
  _RAND_341 = {1{`RANDOM}};
  image_0_341 = _RAND_341[3:0];
  _RAND_342 = {1{`RANDOM}};
  image_0_342 = _RAND_342[3:0];
  _RAND_343 = {1{`RANDOM}};
  image_0_343 = _RAND_343[3:0];
  _RAND_344 = {1{`RANDOM}};
  image_0_344 = _RAND_344[3:0];
  _RAND_345 = {1{`RANDOM}};
  image_0_345 = _RAND_345[3:0];
  _RAND_346 = {1{`RANDOM}};
  image_0_346 = _RAND_346[3:0];
  _RAND_347 = {1{`RANDOM}};
  image_0_347 = _RAND_347[3:0];
  _RAND_348 = {1{`RANDOM}};
  image_0_348 = _RAND_348[3:0];
  _RAND_349 = {1{`RANDOM}};
  image_0_349 = _RAND_349[3:0];
  _RAND_350 = {1{`RANDOM}};
  image_0_350 = _RAND_350[3:0];
  _RAND_351 = {1{`RANDOM}};
  image_0_351 = _RAND_351[3:0];
  _RAND_352 = {1{`RANDOM}};
  image_0_352 = _RAND_352[3:0];
  _RAND_353 = {1{`RANDOM}};
  image_0_353 = _RAND_353[3:0];
  _RAND_354 = {1{`RANDOM}};
  image_0_354 = _RAND_354[3:0];
  _RAND_355 = {1{`RANDOM}};
  image_0_355 = _RAND_355[3:0];
  _RAND_356 = {1{`RANDOM}};
  image_0_356 = _RAND_356[3:0];
  _RAND_357 = {1{`RANDOM}};
  image_0_357 = _RAND_357[3:0];
  _RAND_358 = {1{`RANDOM}};
  image_0_358 = _RAND_358[3:0];
  _RAND_359 = {1{`RANDOM}};
  image_0_359 = _RAND_359[3:0];
  _RAND_360 = {1{`RANDOM}};
  image_0_360 = _RAND_360[3:0];
  _RAND_361 = {1{`RANDOM}};
  image_0_361 = _RAND_361[3:0];
  _RAND_362 = {1{`RANDOM}};
  image_0_362 = _RAND_362[3:0];
  _RAND_363 = {1{`RANDOM}};
  image_0_363 = _RAND_363[3:0];
  _RAND_364 = {1{`RANDOM}};
  image_0_364 = _RAND_364[3:0];
  _RAND_365 = {1{`RANDOM}};
  image_0_365 = _RAND_365[3:0];
  _RAND_366 = {1{`RANDOM}};
  image_0_366 = _RAND_366[3:0];
  _RAND_367 = {1{`RANDOM}};
  image_0_367 = _RAND_367[3:0];
  _RAND_368 = {1{`RANDOM}};
  image_0_368 = _RAND_368[3:0];
  _RAND_369 = {1{`RANDOM}};
  image_0_369 = _RAND_369[3:0];
  _RAND_370 = {1{`RANDOM}};
  image_0_370 = _RAND_370[3:0];
  _RAND_371 = {1{`RANDOM}};
  image_0_371 = _RAND_371[3:0];
  _RAND_372 = {1{`RANDOM}};
  image_0_372 = _RAND_372[3:0];
  _RAND_373 = {1{`RANDOM}};
  image_0_373 = _RAND_373[3:0];
  _RAND_374 = {1{`RANDOM}};
  image_0_374 = _RAND_374[3:0];
  _RAND_375 = {1{`RANDOM}};
  image_0_375 = _RAND_375[3:0];
  _RAND_376 = {1{`RANDOM}};
  image_0_376 = _RAND_376[3:0];
  _RAND_377 = {1{`RANDOM}};
  image_0_377 = _RAND_377[3:0];
  _RAND_378 = {1{`RANDOM}};
  image_0_378 = _RAND_378[3:0];
  _RAND_379 = {1{`RANDOM}};
  image_0_379 = _RAND_379[3:0];
  _RAND_380 = {1{`RANDOM}};
  image_0_380 = _RAND_380[3:0];
  _RAND_381 = {1{`RANDOM}};
  image_0_381 = _RAND_381[3:0];
  _RAND_382 = {1{`RANDOM}};
  image_0_382 = _RAND_382[3:0];
  _RAND_383 = {1{`RANDOM}};
  image_0_383 = _RAND_383[3:0];
  _RAND_384 = {1{`RANDOM}};
  image_0_384 = _RAND_384[3:0];
  _RAND_385 = {1{`RANDOM}};
  image_0_385 = _RAND_385[3:0];
  _RAND_386 = {1{`RANDOM}};
  image_0_386 = _RAND_386[3:0];
  _RAND_387 = {1{`RANDOM}};
  image_0_387 = _RAND_387[3:0];
  _RAND_388 = {1{`RANDOM}};
  image_0_388 = _RAND_388[3:0];
  _RAND_389 = {1{`RANDOM}};
  image_0_389 = _RAND_389[3:0];
  _RAND_390 = {1{`RANDOM}};
  image_0_390 = _RAND_390[3:0];
  _RAND_391 = {1{`RANDOM}};
  image_0_391 = _RAND_391[3:0];
  _RAND_392 = {1{`RANDOM}};
  image_0_392 = _RAND_392[3:0];
  _RAND_393 = {1{`RANDOM}};
  image_0_393 = _RAND_393[3:0];
  _RAND_394 = {1{`RANDOM}};
  image_0_394 = _RAND_394[3:0];
  _RAND_395 = {1{`RANDOM}};
  image_0_395 = _RAND_395[3:0];
  _RAND_396 = {1{`RANDOM}};
  image_0_396 = _RAND_396[3:0];
  _RAND_397 = {1{`RANDOM}};
  image_0_397 = _RAND_397[3:0];
  _RAND_398 = {1{`RANDOM}};
  image_0_398 = _RAND_398[3:0];
  _RAND_399 = {1{`RANDOM}};
  image_0_399 = _RAND_399[3:0];
  _RAND_400 = {1{`RANDOM}};
  image_0_400 = _RAND_400[3:0];
  _RAND_401 = {1{`RANDOM}};
  image_0_401 = _RAND_401[3:0];
  _RAND_402 = {1{`RANDOM}};
  image_0_402 = _RAND_402[3:0];
  _RAND_403 = {1{`RANDOM}};
  image_0_403 = _RAND_403[3:0];
  _RAND_404 = {1{`RANDOM}};
  image_0_404 = _RAND_404[3:0];
  _RAND_405 = {1{`RANDOM}};
  image_0_405 = _RAND_405[3:0];
  _RAND_406 = {1{`RANDOM}};
  image_0_406 = _RAND_406[3:0];
  _RAND_407 = {1{`RANDOM}};
  image_0_407 = _RAND_407[3:0];
  _RAND_408 = {1{`RANDOM}};
  image_0_408 = _RAND_408[3:0];
  _RAND_409 = {1{`RANDOM}};
  image_0_409 = _RAND_409[3:0];
  _RAND_410 = {1{`RANDOM}};
  image_0_410 = _RAND_410[3:0];
  _RAND_411 = {1{`RANDOM}};
  image_0_411 = _RAND_411[3:0];
  _RAND_412 = {1{`RANDOM}};
  image_0_412 = _RAND_412[3:0];
  _RAND_413 = {1{`RANDOM}};
  image_0_413 = _RAND_413[3:0];
  _RAND_414 = {1{`RANDOM}};
  image_0_414 = _RAND_414[3:0];
  _RAND_415 = {1{`RANDOM}};
  image_0_415 = _RAND_415[3:0];
  _RAND_416 = {1{`RANDOM}};
  image_0_416 = _RAND_416[3:0];
  _RAND_417 = {1{`RANDOM}};
  image_0_417 = _RAND_417[3:0];
  _RAND_418 = {1{`RANDOM}};
  image_0_418 = _RAND_418[3:0];
  _RAND_419 = {1{`RANDOM}};
  image_0_419 = _RAND_419[3:0];
  _RAND_420 = {1{`RANDOM}};
  image_0_420 = _RAND_420[3:0];
  _RAND_421 = {1{`RANDOM}};
  image_0_421 = _RAND_421[3:0];
  _RAND_422 = {1{`RANDOM}};
  image_0_422 = _RAND_422[3:0];
  _RAND_423 = {1{`RANDOM}};
  image_0_423 = _RAND_423[3:0];
  _RAND_424 = {1{`RANDOM}};
  image_0_424 = _RAND_424[3:0];
  _RAND_425 = {1{`RANDOM}};
  image_0_425 = _RAND_425[3:0];
  _RAND_426 = {1{`RANDOM}};
  image_0_426 = _RAND_426[3:0];
  _RAND_427 = {1{`RANDOM}};
  image_0_427 = _RAND_427[3:0];
  _RAND_428 = {1{`RANDOM}};
  image_0_428 = _RAND_428[3:0];
  _RAND_429 = {1{`RANDOM}};
  image_0_429 = _RAND_429[3:0];
  _RAND_430 = {1{`RANDOM}};
  image_0_430 = _RAND_430[3:0];
  _RAND_431 = {1{`RANDOM}};
  image_0_431 = _RAND_431[3:0];
  _RAND_432 = {1{`RANDOM}};
  image_0_432 = _RAND_432[3:0];
  _RAND_433 = {1{`RANDOM}};
  image_0_433 = _RAND_433[3:0];
  _RAND_434 = {1{`RANDOM}};
  image_0_434 = _RAND_434[3:0];
  _RAND_435 = {1{`RANDOM}};
  image_0_435 = _RAND_435[3:0];
  _RAND_436 = {1{`RANDOM}};
  image_0_436 = _RAND_436[3:0];
  _RAND_437 = {1{`RANDOM}};
  image_0_437 = _RAND_437[3:0];
  _RAND_438 = {1{`RANDOM}};
  image_0_438 = _RAND_438[3:0];
  _RAND_439 = {1{`RANDOM}};
  image_0_439 = _RAND_439[3:0];
  _RAND_440 = {1{`RANDOM}};
  image_0_440 = _RAND_440[3:0];
  _RAND_441 = {1{`RANDOM}};
  image_0_441 = _RAND_441[3:0];
  _RAND_442 = {1{`RANDOM}};
  image_0_442 = _RAND_442[3:0];
  _RAND_443 = {1{`RANDOM}};
  image_0_443 = _RAND_443[3:0];
  _RAND_444 = {1{`RANDOM}};
  image_0_444 = _RAND_444[3:0];
  _RAND_445 = {1{`RANDOM}};
  image_0_445 = _RAND_445[3:0];
  _RAND_446 = {1{`RANDOM}};
  image_0_446 = _RAND_446[3:0];
  _RAND_447 = {1{`RANDOM}};
  image_0_447 = _RAND_447[3:0];
  _RAND_448 = {1{`RANDOM}};
  image_0_448 = _RAND_448[3:0];
  _RAND_449 = {1{`RANDOM}};
  image_0_449 = _RAND_449[3:0];
  _RAND_450 = {1{`RANDOM}};
  image_0_450 = _RAND_450[3:0];
  _RAND_451 = {1{`RANDOM}};
  image_0_451 = _RAND_451[3:0];
  _RAND_452 = {1{`RANDOM}};
  image_0_452 = _RAND_452[3:0];
  _RAND_453 = {1{`RANDOM}};
  image_0_453 = _RAND_453[3:0];
  _RAND_454 = {1{`RANDOM}};
  image_0_454 = _RAND_454[3:0];
  _RAND_455 = {1{`RANDOM}};
  image_0_455 = _RAND_455[3:0];
  _RAND_456 = {1{`RANDOM}};
  image_0_456 = _RAND_456[3:0];
  _RAND_457 = {1{`RANDOM}};
  image_0_457 = _RAND_457[3:0];
  _RAND_458 = {1{`RANDOM}};
  image_0_458 = _RAND_458[3:0];
  _RAND_459 = {1{`RANDOM}};
  image_0_459 = _RAND_459[3:0];
  _RAND_460 = {1{`RANDOM}};
  image_0_460 = _RAND_460[3:0];
  _RAND_461 = {1{`RANDOM}};
  image_0_461 = _RAND_461[3:0];
  _RAND_462 = {1{`RANDOM}};
  image_0_462 = _RAND_462[3:0];
  _RAND_463 = {1{`RANDOM}};
  image_0_463 = _RAND_463[3:0];
  _RAND_464 = {1{`RANDOM}};
  image_0_464 = _RAND_464[3:0];
  _RAND_465 = {1{`RANDOM}};
  image_0_465 = _RAND_465[3:0];
  _RAND_466 = {1{`RANDOM}};
  image_0_466 = _RAND_466[3:0];
  _RAND_467 = {1{`RANDOM}};
  image_0_467 = _RAND_467[3:0];
  _RAND_468 = {1{`RANDOM}};
  image_0_468 = _RAND_468[3:0];
  _RAND_469 = {1{`RANDOM}};
  image_0_469 = _RAND_469[3:0];
  _RAND_470 = {1{`RANDOM}};
  image_0_470 = _RAND_470[3:0];
  _RAND_471 = {1{`RANDOM}};
  image_0_471 = _RAND_471[3:0];
  _RAND_472 = {1{`RANDOM}};
  image_0_472 = _RAND_472[3:0];
  _RAND_473 = {1{`RANDOM}};
  image_0_473 = _RAND_473[3:0];
  _RAND_474 = {1{`RANDOM}};
  image_0_474 = _RAND_474[3:0];
  _RAND_475 = {1{`RANDOM}};
  image_0_475 = _RAND_475[3:0];
  _RAND_476 = {1{`RANDOM}};
  image_0_476 = _RAND_476[3:0];
  _RAND_477 = {1{`RANDOM}};
  image_0_477 = _RAND_477[3:0];
  _RAND_478 = {1{`RANDOM}};
  image_0_478 = _RAND_478[3:0];
  _RAND_479 = {1{`RANDOM}};
  image_0_479 = _RAND_479[3:0];
  _RAND_480 = {1{`RANDOM}};
  image_0_480 = _RAND_480[3:0];
  _RAND_481 = {1{`RANDOM}};
  image_0_481 = _RAND_481[3:0];
  _RAND_482 = {1{`RANDOM}};
  image_0_482 = _RAND_482[3:0];
  _RAND_483 = {1{`RANDOM}};
  image_0_483 = _RAND_483[3:0];
  _RAND_484 = {1{`RANDOM}};
  image_0_484 = _RAND_484[3:0];
  _RAND_485 = {1{`RANDOM}};
  image_0_485 = _RAND_485[3:0];
  _RAND_486 = {1{`RANDOM}};
  image_0_486 = _RAND_486[3:0];
  _RAND_487 = {1{`RANDOM}};
  image_0_487 = _RAND_487[3:0];
  _RAND_488 = {1{`RANDOM}};
  image_0_488 = _RAND_488[3:0];
  _RAND_489 = {1{`RANDOM}};
  image_0_489 = _RAND_489[3:0];
  _RAND_490 = {1{`RANDOM}};
  image_0_490 = _RAND_490[3:0];
  _RAND_491 = {1{`RANDOM}};
  image_0_491 = _RAND_491[3:0];
  _RAND_492 = {1{`RANDOM}};
  image_0_492 = _RAND_492[3:0];
  _RAND_493 = {1{`RANDOM}};
  image_0_493 = _RAND_493[3:0];
  _RAND_494 = {1{`RANDOM}};
  image_0_494 = _RAND_494[3:0];
  _RAND_495 = {1{`RANDOM}};
  image_0_495 = _RAND_495[3:0];
  _RAND_496 = {1{`RANDOM}};
  image_0_496 = _RAND_496[3:0];
  _RAND_497 = {1{`RANDOM}};
  image_0_497 = _RAND_497[3:0];
  _RAND_498 = {1{`RANDOM}};
  image_0_498 = _RAND_498[3:0];
  _RAND_499 = {1{`RANDOM}};
  image_0_499 = _RAND_499[3:0];
  _RAND_500 = {1{`RANDOM}};
  image_0_500 = _RAND_500[3:0];
  _RAND_501 = {1{`RANDOM}};
  image_0_501 = _RAND_501[3:0];
  _RAND_502 = {1{`RANDOM}};
  image_0_502 = _RAND_502[3:0];
  _RAND_503 = {1{`RANDOM}};
  image_0_503 = _RAND_503[3:0];
  _RAND_504 = {1{`RANDOM}};
  image_0_504 = _RAND_504[3:0];
  _RAND_505 = {1{`RANDOM}};
  image_0_505 = _RAND_505[3:0];
  _RAND_506 = {1{`RANDOM}};
  image_0_506 = _RAND_506[3:0];
  _RAND_507 = {1{`RANDOM}};
  image_0_507 = _RAND_507[3:0];
  _RAND_508 = {1{`RANDOM}};
  image_0_508 = _RAND_508[3:0];
  _RAND_509 = {1{`RANDOM}};
  image_0_509 = _RAND_509[3:0];
  _RAND_510 = {1{`RANDOM}};
  image_0_510 = _RAND_510[3:0];
  _RAND_511 = {1{`RANDOM}};
  image_0_511 = _RAND_511[3:0];
  _RAND_512 = {1{`RANDOM}};
  image_0_512 = _RAND_512[3:0];
  _RAND_513 = {1{`RANDOM}};
  image_0_513 = _RAND_513[3:0];
  _RAND_514 = {1{`RANDOM}};
  image_0_514 = _RAND_514[3:0];
  _RAND_515 = {1{`RANDOM}};
  image_0_515 = _RAND_515[3:0];
  _RAND_516 = {1{`RANDOM}};
  image_0_516 = _RAND_516[3:0];
  _RAND_517 = {1{`RANDOM}};
  image_0_517 = _RAND_517[3:0];
  _RAND_518 = {1{`RANDOM}};
  image_0_518 = _RAND_518[3:0];
  _RAND_519 = {1{`RANDOM}};
  image_0_519 = _RAND_519[3:0];
  _RAND_520 = {1{`RANDOM}};
  image_0_520 = _RAND_520[3:0];
  _RAND_521 = {1{`RANDOM}};
  image_0_521 = _RAND_521[3:0];
  _RAND_522 = {1{`RANDOM}};
  image_0_522 = _RAND_522[3:0];
  _RAND_523 = {1{`RANDOM}};
  image_0_523 = _RAND_523[3:0];
  _RAND_524 = {1{`RANDOM}};
  image_0_524 = _RAND_524[3:0];
  _RAND_525 = {1{`RANDOM}};
  image_0_525 = _RAND_525[3:0];
  _RAND_526 = {1{`RANDOM}};
  image_0_526 = _RAND_526[3:0];
  _RAND_527 = {1{`RANDOM}};
  image_0_527 = _RAND_527[3:0];
  _RAND_528 = {1{`RANDOM}};
  image_0_528 = _RAND_528[3:0];
  _RAND_529 = {1{`RANDOM}};
  image_0_529 = _RAND_529[3:0];
  _RAND_530 = {1{`RANDOM}};
  image_0_530 = _RAND_530[3:0];
  _RAND_531 = {1{`RANDOM}};
  image_0_531 = _RAND_531[3:0];
  _RAND_532 = {1{`RANDOM}};
  image_0_532 = _RAND_532[3:0];
  _RAND_533 = {1{`RANDOM}};
  image_0_533 = _RAND_533[3:0];
  _RAND_534 = {1{`RANDOM}};
  image_0_534 = _RAND_534[3:0];
  _RAND_535 = {1{`RANDOM}};
  image_0_535 = _RAND_535[3:0];
  _RAND_536 = {1{`RANDOM}};
  image_0_536 = _RAND_536[3:0];
  _RAND_537 = {1{`RANDOM}};
  image_0_537 = _RAND_537[3:0];
  _RAND_538 = {1{`RANDOM}};
  image_0_538 = _RAND_538[3:0];
  _RAND_539 = {1{`RANDOM}};
  image_0_539 = _RAND_539[3:0];
  _RAND_540 = {1{`RANDOM}};
  image_0_540 = _RAND_540[3:0];
  _RAND_541 = {1{`RANDOM}};
  image_0_541 = _RAND_541[3:0];
  _RAND_542 = {1{`RANDOM}};
  image_0_542 = _RAND_542[3:0];
  _RAND_543 = {1{`RANDOM}};
  image_0_543 = _RAND_543[3:0];
  _RAND_544 = {1{`RANDOM}};
  image_0_544 = _RAND_544[3:0];
  _RAND_545 = {1{`RANDOM}};
  image_0_545 = _RAND_545[3:0];
  _RAND_546 = {1{`RANDOM}};
  image_0_546 = _RAND_546[3:0];
  _RAND_547 = {1{`RANDOM}};
  image_0_547 = _RAND_547[3:0];
  _RAND_548 = {1{`RANDOM}};
  image_0_548 = _RAND_548[3:0];
  _RAND_549 = {1{`RANDOM}};
  image_0_549 = _RAND_549[3:0];
  _RAND_550 = {1{`RANDOM}};
  image_0_550 = _RAND_550[3:0];
  _RAND_551 = {1{`RANDOM}};
  image_0_551 = _RAND_551[3:0];
  _RAND_552 = {1{`RANDOM}};
  image_0_552 = _RAND_552[3:0];
  _RAND_553 = {1{`RANDOM}};
  image_0_553 = _RAND_553[3:0];
  _RAND_554 = {1{`RANDOM}};
  image_0_554 = _RAND_554[3:0];
  _RAND_555 = {1{`RANDOM}};
  image_0_555 = _RAND_555[3:0];
  _RAND_556 = {1{`RANDOM}};
  image_0_556 = _RAND_556[3:0];
  _RAND_557 = {1{`RANDOM}};
  image_0_557 = _RAND_557[3:0];
  _RAND_558 = {1{`RANDOM}};
  image_0_558 = _RAND_558[3:0];
  _RAND_559 = {1{`RANDOM}};
  image_0_559 = _RAND_559[3:0];
  _RAND_560 = {1{`RANDOM}};
  image_0_560 = _RAND_560[3:0];
  _RAND_561 = {1{`RANDOM}};
  image_0_561 = _RAND_561[3:0];
  _RAND_562 = {1{`RANDOM}};
  image_0_562 = _RAND_562[3:0];
  _RAND_563 = {1{`RANDOM}};
  image_0_563 = _RAND_563[3:0];
  _RAND_564 = {1{`RANDOM}};
  image_0_564 = _RAND_564[3:0];
  _RAND_565 = {1{`RANDOM}};
  image_0_565 = _RAND_565[3:0];
  _RAND_566 = {1{`RANDOM}};
  image_0_566 = _RAND_566[3:0];
  _RAND_567 = {1{`RANDOM}};
  image_0_567 = _RAND_567[3:0];
  _RAND_568 = {1{`RANDOM}};
  image_0_568 = _RAND_568[3:0];
  _RAND_569 = {1{`RANDOM}};
  image_0_569 = _RAND_569[3:0];
  _RAND_570 = {1{`RANDOM}};
  image_0_570 = _RAND_570[3:0];
  _RAND_571 = {1{`RANDOM}};
  image_0_571 = _RAND_571[3:0];
  _RAND_572 = {1{`RANDOM}};
  image_0_572 = _RAND_572[3:0];
  _RAND_573 = {1{`RANDOM}};
  image_0_573 = _RAND_573[3:0];
  _RAND_574 = {1{`RANDOM}};
  image_0_574 = _RAND_574[3:0];
  _RAND_575 = {1{`RANDOM}};
  image_0_575 = _RAND_575[3:0];
  _RAND_576 = {1{`RANDOM}};
  image_1_0 = _RAND_576[3:0];
  _RAND_577 = {1{`RANDOM}};
  image_1_1 = _RAND_577[3:0];
  _RAND_578 = {1{`RANDOM}};
  image_1_2 = _RAND_578[3:0];
  _RAND_579 = {1{`RANDOM}};
  image_1_3 = _RAND_579[3:0];
  _RAND_580 = {1{`RANDOM}};
  image_1_4 = _RAND_580[3:0];
  _RAND_581 = {1{`RANDOM}};
  image_1_5 = _RAND_581[3:0];
  _RAND_582 = {1{`RANDOM}};
  image_1_6 = _RAND_582[3:0];
  _RAND_583 = {1{`RANDOM}};
  image_1_7 = _RAND_583[3:0];
  _RAND_584 = {1{`RANDOM}};
  image_1_8 = _RAND_584[3:0];
  _RAND_585 = {1{`RANDOM}};
  image_1_9 = _RAND_585[3:0];
  _RAND_586 = {1{`RANDOM}};
  image_1_10 = _RAND_586[3:0];
  _RAND_587 = {1{`RANDOM}};
  image_1_11 = _RAND_587[3:0];
  _RAND_588 = {1{`RANDOM}};
  image_1_12 = _RAND_588[3:0];
  _RAND_589 = {1{`RANDOM}};
  image_1_13 = _RAND_589[3:0];
  _RAND_590 = {1{`RANDOM}};
  image_1_14 = _RAND_590[3:0];
  _RAND_591 = {1{`RANDOM}};
  image_1_15 = _RAND_591[3:0];
  _RAND_592 = {1{`RANDOM}};
  image_1_16 = _RAND_592[3:0];
  _RAND_593 = {1{`RANDOM}};
  image_1_17 = _RAND_593[3:0];
  _RAND_594 = {1{`RANDOM}};
  image_1_18 = _RAND_594[3:0];
  _RAND_595 = {1{`RANDOM}};
  image_1_19 = _RAND_595[3:0];
  _RAND_596 = {1{`RANDOM}};
  image_1_20 = _RAND_596[3:0];
  _RAND_597 = {1{`RANDOM}};
  image_1_21 = _RAND_597[3:0];
  _RAND_598 = {1{`RANDOM}};
  image_1_22 = _RAND_598[3:0];
  _RAND_599 = {1{`RANDOM}};
  image_1_23 = _RAND_599[3:0];
  _RAND_600 = {1{`RANDOM}};
  image_1_24 = _RAND_600[3:0];
  _RAND_601 = {1{`RANDOM}};
  image_1_25 = _RAND_601[3:0];
  _RAND_602 = {1{`RANDOM}};
  image_1_26 = _RAND_602[3:0];
  _RAND_603 = {1{`RANDOM}};
  image_1_27 = _RAND_603[3:0];
  _RAND_604 = {1{`RANDOM}};
  image_1_28 = _RAND_604[3:0];
  _RAND_605 = {1{`RANDOM}};
  image_1_29 = _RAND_605[3:0];
  _RAND_606 = {1{`RANDOM}};
  image_1_30 = _RAND_606[3:0];
  _RAND_607 = {1{`RANDOM}};
  image_1_31 = _RAND_607[3:0];
  _RAND_608 = {1{`RANDOM}};
  image_1_32 = _RAND_608[3:0];
  _RAND_609 = {1{`RANDOM}};
  image_1_33 = _RAND_609[3:0];
  _RAND_610 = {1{`RANDOM}};
  image_1_34 = _RAND_610[3:0];
  _RAND_611 = {1{`RANDOM}};
  image_1_35 = _RAND_611[3:0];
  _RAND_612 = {1{`RANDOM}};
  image_1_36 = _RAND_612[3:0];
  _RAND_613 = {1{`RANDOM}};
  image_1_37 = _RAND_613[3:0];
  _RAND_614 = {1{`RANDOM}};
  image_1_38 = _RAND_614[3:0];
  _RAND_615 = {1{`RANDOM}};
  image_1_39 = _RAND_615[3:0];
  _RAND_616 = {1{`RANDOM}};
  image_1_40 = _RAND_616[3:0];
  _RAND_617 = {1{`RANDOM}};
  image_1_41 = _RAND_617[3:0];
  _RAND_618 = {1{`RANDOM}};
  image_1_42 = _RAND_618[3:0];
  _RAND_619 = {1{`RANDOM}};
  image_1_43 = _RAND_619[3:0];
  _RAND_620 = {1{`RANDOM}};
  image_1_44 = _RAND_620[3:0];
  _RAND_621 = {1{`RANDOM}};
  image_1_45 = _RAND_621[3:0];
  _RAND_622 = {1{`RANDOM}};
  image_1_46 = _RAND_622[3:0];
  _RAND_623 = {1{`RANDOM}};
  image_1_47 = _RAND_623[3:0];
  _RAND_624 = {1{`RANDOM}};
  image_1_48 = _RAND_624[3:0];
  _RAND_625 = {1{`RANDOM}};
  image_1_49 = _RAND_625[3:0];
  _RAND_626 = {1{`RANDOM}};
  image_1_50 = _RAND_626[3:0];
  _RAND_627 = {1{`RANDOM}};
  image_1_51 = _RAND_627[3:0];
  _RAND_628 = {1{`RANDOM}};
  image_1_52 = _RAND_628[3:0];
  _RAND_629 = {1{`RANDOM}};
  image_1_53 = _RAND_629[3:0];
  _RAND_630 = {1{`RANDOM}};
  image_1_54 = _RAND_630[3:0];
  _RAND_631 = {1{`RANDOM}};
  image_1_55 = _RAND_631[3:0];
  _RAND_632 = {1{`RANDOM}};
  image_1_56 = _RAND_632[3:0];
  _RAND_633 = {1{`RANDOM}};
  image_1_57 = _RAND_633[3:0];
  _RAND_634 = {1{`RANDOM}};
  image_1_58 = _RAND_634[3:0];
  _RAND_635 = {1{`RANDOM}};
  image_1_59 = _RAND_635[3:0];
  _RAND_636 = {1{`RANDOM}};
  image_1_60 = _RAND_636[3:0];
  _RAND_637 = {1{`RANDOM}};
  image_1_61 = _RAND_637[3:0];
  _RAND_638 = {1{`RANDOM}};
  image_1_62 = _RAND_638[3:0];
  _RAND_639 = {1{`RANDOM}};
  image_1_63 = _RAND_639[3:0];
  _RAND_640 = {1{`RANDOM}};
  image_1_64 = _RAND_640[3:0];
  _RAND_641 = {1{`RANDOM}};
  image_1_65 = _RAND_641[3:0];
  _RAND_642 = {1{`RANDOM}};
  image_1_66 = _RAND_642[3:0];
  _RAND_643 = {1{`RANDOM}};
  image_1_67 = _RAND_643[3:0];
  _RAND_644 = {1{`RANDOM}};
  image_1_68 = _RAND_644[3:0];
  _RAND_645 = {1{`RANDOM}};
  image_1_69 = _RAND_645[3:0];
  _RAND_646 = {1{`RANDOM}};
  image_1_70 = _RAND_646[3:0];
  _RAND_647 = {1{`RANDOM}};
  image_1_71 = _RAND_647[3:0];
  _RAND_648 = {1{`RANDOM}};
  image_1_72 = _RAND_648[3:0];
  _RAND_649 = {1{`RANDOM}};
  image_1_73 = _RAND_649[3:0];
  _RAND_650 = {1{`RANDOM}};
  image_1_74 = _RAND_650[3:0];
  _RAND_651 = {1{`RANDOM}};
  image_1_75 = _RAND_651[3:0];
  _RAND_652 = {1{`RANDOM}};
  image_1_76 = _RAND_652[3:0];
  _RAND_653 = {1{`RANDOM}};
  image_1_77 = _RAND_653[3:0];
  _RAND_654 = {1{`RANDOM}};
  image_1_78 = _RAND_654[3:0];
  _RAND_655 = {1{`RANDOM}};
  image_1_79 = _RAND_655[3:0];
  _RAND_656 = {1{`RANDOM}};
  image_1_80 = _RAND_656[3:0];
  _RAND_657 = {1{`RANDOM}};
  image_1_81 = _RAND_657[3:0];
  _RAND_658 = {1{`RANDOM}};
  image_1_82 = _RAND_658[3:0];
  _RAND_659 = {1{`RANDOM}};
  image_1_83 = _RAND_659[3:0];
  _RAND_660 = {1{`RANDOM}};
  image_1_84 = _RAND_660[3:0];
  _RAND_661 = {1{`RANDOM}};
  image_1_85 = _RAND_661[3:0];
  _RAND_662 = {1{`RANDOM}};
  image_1_86 = _RAND_662[3:0];
  _RAND_663 = {1{`RANDOM}};
  image_1_87 = _RAND_663[3:0];
  _RAND_664 = {1{`RANDOM}};
  image_1_88 = _RAND_664[3:0];
  _RAND_665 = {1{`RANDOM}};
  image_1_89 = _RAND_665[3:0];
  _RAND_666 = {1{`RANDOM}};
  image_1_90 = _RAND_666[3:0];
  _RAND_667 = {1{`RANDOM}};
  image_1_91 = _RAND_667[3:0];
  _RAND_668 = {1{`RANDOM}};
  image_1_92 = _RAND_668[3:0];
  _RAND_669 = {1{`RANDOM}};
  image_1_93 = _RAND_669[3:0];
  _RAND_670 = {1{`RANDOM}};
  image_1_94 = _RAND_670[3:0];
  _RAND_671 = {1{`RANDOM}};
  image_1_95 = _RAND_671[3:0];
  _RAND_672 = {1{`RANDOM}};
  image_1_96 = _RAND_672[3:0];
  _RAND_673 = {1{`RANDOM}};
  image_1_97 = _RAND_673[3:0];
  _RAND_674 = {1{`RANDOM}};
  image_1_98 = _RAND_674[3:0];
  _RAND_675 = {1{`RANDOM}};
  image_1_99 = _RAND_675[3:0];
  _RAND_676 = {1{`RANDOM}};
  image_1_100 = _RAND_676[3:0];
  _RAND_677 = {1{`RANDOM}};
  image_1_101 = _RAND_677[3:0];
  _RAND_678 = {1{`RANDOM}};
  image_1_102 = _RAND_678[3:0];
  _RAND_679 = {1{`RANDOM}};
  image_1_103 = _RAND_679[3:0];
  _RAND_680 = {1{`RANDOM}};
  image_1_104 = _RAND_680[3:0];
  _RAND_681 = {1{`RANDOM}};
  image_1_105 = _RAND_681[3:0];
  _RAND_682 = {1{`RANDOM}};
  image_1_106 = _RAND_682[3:0];
  _RAND_683 = {1{`RANDOM}};
  image_1_107 = _RAND_683[3:0];
  _RAND_684 = {1{`RANDOM}};
  image_1_108 = _RAND_684[3:0];
  _RAND_685 = {1{`RANDOM}};
  image_1_109 = _RAND_685[3:0];
  _RAND_686 = {1{`RANDOM}};
  image_1_110 = _RAND_686[3:0];
  _RAND_687 = {1{`RANDOM}};
  image_1_111 = _RAND_687[3:0];
  _RAND_688 = {1{`RANDOM}};
  image_1_112 = _RAND_688[3:0];
  _RAND_689 = {1{`RANDOM}};
  image_1_113 = _RAND_689[3:0];
  _RAND_690 = {1{`RANDOM}};
  image_1_114 = _RAND_690[3:0];
  _RAND_691 = {1{`RANDOM}};
  image_1_115 = _RAND_691[3:0];
  _RAND_692 = {1{`RANDOM}};
  image_1_116 = _RAND_692[3:0];
  _RAND_693 = {1{`RANDOM}};
  image_1_117 = _RAND_693[3:0];
  _RAND_694 = {1{`RANDOM}};
  image_1_118 = _RAND_694[3:0];
  _RAND_695 = {1{`RANDOM}};
  image_1_119 = _RAND_695[3:0];
  _RAND_696 = {1{`RANDOM}};
  image_1_120 = _RAND_696[3:0];
  _RAND_697 = {1{`RANDOM}};
  image_1_121 = _RAND_697[3:0];
  _RAND_698 = {1{`RANDOM}};
  image_1_122 = _RAND_698[3:0];
  _RAND_699 = {1{`RANDOM}};
  image_1_123 = _RAND_699[3:0];
  _RAND_700 = {1{`RANDOM}};
  image_1_124 = _RAND_700[3:0];
  _RAND_701 = {1{`RANDOM}};
  image_1_125 = _RAND_701[3:0];
  _RAND_702 = {1{`RANDOM}};
  image_1_126 = _RAND_702[3:0];
  _RAND_703 = {1{`RANDOM}};
  image_1_127 = _RAND_703[3:0];
  _RAND_704 = {1{`RANDOM}};
  image_1_128 = _RAND_704[3:0];
  _RAND_705 = {1{`RANDOM}};
  image_1_129 = _RAND_705[3:0];
  _RAND_706 = {1{`RANDOM}};
  image_1_130 = _RAND_706[3:0];
  _RAND_707 = {1{`RANDOM}};
  image_1_131 = _RAND_707[3:0];
  _RAND_708 = {1{`RANDOM}};
  image_1_132 = _RAND_708[3:0];
  _RAND_709 = {1{`RANDOM}};
  image_1_133 = _RAND_709[3:0];
  _RAND_710 = {1{`RANDOM}};
  image_1_134 = _RAND_710[3:0];
  _RAND_711 = {1{`RANDOM}};
  image_1_135 = _RAND_711[3:0];
  _RAND_712 = {1{`RANDOM}};
  image_1_136 = _RAND_712[3:0];
  _RAND_713 = {1{`RANDOM}};
  image_1_137 = _RAND_713[3:0];
  _RAND_714 = {1{`RANDOM}};
  image_1_138 = _RAND_714[3:0];
  _RAND_715 = {1{`RANDOM}};
  image_1_139 = _RAND_715[3:0];
  _RAND_716 = {1{`RANDOM}};
  image_1_140 = _RAND_716[3:0];
  _RAND_717 = {1{`RANDOM}};
  image_1_141 = _RAND_717[3:0];
  _RAND_718 = {1{`RANDOM}};
  image_1_142 = _RAND_718[3:0];
  _RAND_719 = {1{`RANDOM}};
  image_1_143 = _RAND_719[3:0];
  _RAND_720 = {1{`RANDOM}};
  image_1_144 = _RAND_720[3:0];
  _RAND_721 = {1{`RANDOM}};
  image_1_145 = _RAND_721[3:0];
  _RAND_722 = {1{`RANDOM}};
  image_1_146 = _RAND_722[3:0];
  _RAND_723 = {1{`RANDOM}};
  image_1_147 = _RAND_723[3:0];
  _RAND_724 = {1{`RANDOM}};
  image_1_148 = _RAND_724[3:0];
  _RAND_725 = {1{`RANDOM}};
  image_1_149 = _RAND_725[3:0];
  _RAND_726 = {1{`RANDOM}};
  image_1_150 = _RAND_726[3:0];
  _RAND_727 = {1{`RANDOM}};
  image_1_151 = _RAND_727[3:0];
  _RAND_728 = {1{`RANDOM}};
  image_1_152 = _RAND_728[3:0];
  _RAND_729 = {1{`RANDOM}};
  image_1_153 = _RAND_729[3:0];
  _RAND_730 = {1{`RANDOM}};
  image_1_154 = _RAND_730[3:0];
  _RAND_731 = {1{`RANDOM}};
  image_1_155 = _RAND_731[3:0];
  _RAND_732 = {1{`RANDOM}};
  image_1_156 = _RAND_732[3:0];
  _RAND_733 = {1{`RANDOM}};
  image_1_157 = _RAND_733[3:0];
  _RAND_734 = {1{`RANDOM}};
  image_1_158 = _RAND_734[3:0];
  _RAND_735 = {1{`RANDOM}};
  image_1_159 = _RAND_735[3:0];
  _RAND_736 = {1{`RANDOM}};
  image_1_160 = _RAND_736[3:0];
  _RAND_737 = {1{`RANDOM}};
  image_1_161 = _RAND_737[3:0];
  _RAND_738 = {1{`RANDOM}};
  image_1_162 = _RAND_738[3:0];
  _RAND_739 = {1{`RANDOM}};
  image_1_163 = _RAND_739[3:0];
  _RAND_740 = {1{`RANDOM}};
  image_1_164 = _RAND_740[3:0];
  _RAND_741 = {1{`RANDOM}};
  image_1_165 = _RAND_741[3:0];
  _RAND_742 = {1{`RANDOM}};
  image_1_166 = _RAND_742[3:0];
  _RAND_743 = {1{`RANDOM}};
  image_1_167 = _RAND_743[3:0];
  _RAND_744 = {1{`RANDOM}};
  image_1_168 = _RAND_744[3:0];
  _RAND_745 = {1{`RANDOM}};
  image_1_169 = _RAND_745[3:0];
  _RAND_746 = {1{`RANDOM}};
  image_1_170 = _RAND_746[3:0];
  _RAND_747 = {1{`RANDOM}};
  image_1_171 = _RAND_747[3:0];
  _RAND_748 = {1{`RANDOM}};
  image_1_172 = _RAND_748[3:0];
  _RAND_749 = {1{`RANDOM}};
  image_1_173 = _RAND_749[3:0];
  _RAND_750 = {1{`RANDOM}};
  image_1_174 = _RAND_750[3:0];
  _RAND_751 = {1{`RANDOM}};
  image_1_175 = _RAND_751[3:0];
  _RAND_752 = {1{`RANDOM}};
  image_1_176 = _RAND_752[3:0];
  _RAND_753 = {1{`RANDOM}};
  image_1_177 = _RAND_753[3:0];
  _RAND_754 = {1{`RANDOM}};
  image_1_178 = _RAND_754[3:0];
  _RAND_755 = {1{`RANDOM}};
  image_1_179 = _RAND_755[3:0];
  _RAND_756 = {1{`RANDOM}};
  image_1_180 = _RAND_756[3:0];
  _RAND_757 = {1{`RANDOM}};
  image_1_181 = _RAND_757[3:0];
  _RAND_758 = {1{`RANDOM}};
  image_1_182 = _RAND_758[3:0];
  _RAND_759 = {1{`RANDOM}};
  image_1_183 = _RAND_759[3:0];
  _RAND_760 = {1{`RANDOM}};
  image_1_184 = _RAND_760[3:0];
  _RAND_761 = {1{`RANDOM}};
  image_1_185 = _RAND_761[3:0];
  _RAND_762 = {1{`RANDOM}};
  image_1_186 = _RAND_762[3:0];
  _RAND_763 = {1{`RANDOM}};
  image_1_187 = _RAND_763[3:0];
  _RAND_764 = {1{`RANDOM}};
  image_1_188 = _RAND_764[3:0];
  _RAND_765 = {1{`RANDOM}};
  image_1_189 = _RAND_765[3:0];
  _RAND_766 = {1{`RANDOM}};
  image_1_190 = _RAND_766[3:0];
  _RAND_767 = {1{`RANDOM}};
  image_1_191 = _RAND_767[3:0];
  _RAND_768 = {1{`RANDOM}};
  image_1_192 = _RAND_768[3:0];
  _RAND_769 = {1{`RANDOM}};
  image_1_193 = _RAND_769[3:0];
  _RAND_770 = {1{`RANDOM}};
  image_1_194 = _RAND_770[3:0];
  _RAND_771 = {1{`RANDOM}};
  image_1_195 = _RAND_771[3:0];
  _RAND_772 = {1{`RANDOM}};
  image_1_196 = _RAND_772[3:0];
  _RAND_773 = {1{`RANDOM}};
  image_1_197 = _RAND_773[3:0];
  _RAND_774 = {1{`RANDOM}};
  image_1_198 = _RAND_774[3:0];
  _RAND_775 = {1{`RANDOM}};
  image_1_199 = _RAND_775[3:0];
  _RAND_776 = {1{`RANDOM}};
  image_1_200 = _RAND_776[3:0];
  _RAND_777 = {1{`RANDOM}};
  image_1_201 = _RAND_777[3:0];
  _RAND_778 = {1{`RANDOM}};
  image_1_202 = _RAND_778[3:0];
  _RAND_779 = {1{`RANDOM}};
  image_1_203 = _RAND_779[3:0];
  _RAND_780 = {1{`RANDOM}};
  image_1_204 = _RAND_780[3:0];
  _RAND_781 = {1{`RANDOM}};
  image_1_205 = _RAND_781[3:0];
  _RAND_782 = {1{`RANDOM}};
  image_1_206 = _RAND_782[3:0];
  _RAND_783 = {1{`RANDOM}};
  image_1_207 = _RAND_783[3:0];
  _RAND_784 = {1{`RANDOM}};
  image_1_208 = _RAND_784[3:0];
  _RAND_785 = {1{`RANDOM}};
  image_1_209 = _RAND_785[3:0];
  _RAND_786 = {1{`RANDOM}};
  image_1_210 = _RAND_786[3:0];
  _RAND_787 = {1{`RANDOM}};
  image_1_211 = _RAND_787[3:0];
  _RAND_788 = {1{`RANDOM}};
  image_1_212 = _RAND_788[3:0];
  _RAND_789 = {1{`RANDOM}};
  image_1_213 = _RAND_789[3:0];
  _RAND_790 = {1{`RANDOM}};
  image_1_214 = _RAND_790[3:0];
  _RAND_791 = {1{`RANDOM}};
  image_1_215 = _RAND_791[3:0];
  _RAND_792 = {1{`RANDOM}};
  image_1_216 = _RAND_792[3:0];
  _RAND_793 = {1{`RANDOM}};
  image_1_217 = _RAND_793[3:0];
  _RAND_794 = {1{`RANDOM}};
  image_1_218 = _RAND_794[3:0];
  _RAND_795 = {1{`RANDOM}};
  image_1_219 = _RAND_795[3:0];
  _RAND_796 = {1{`RANDOM}};
  image_1_220 = _RAND_796[3:0];
  _RAND_797 = {1{`RANDOM}};
  image_1_221 = _RAND_797[3:0];
  _RAND_798 = {1{`RANDOM}};
  image_1_222 = _RAND_798[3:0];
  _RAND_799 = {1{`RANDOM}};
  image_1_223 = _RAND_799[3:0];
  _RAND_800 = {1{`RANDOM}};
  image_1_224 = _RAND_800[3:0];
  _RAND_801 = {1{`RANDOM}};
  image_1_225 = _RAND_801[3:0];
  _RAND_802 = {1{`RANDOM}};
  image_1_226 = _RAND_802[3:0];
  _RAND_803 = {1{`RANDOM}};
  image_1_227 = _RAND_803[3:0];
  _RAND_804 = {1{`RANDOM}};
  image_1_228 = _RAND_804[3:0];
  _RAND_805 = {1{`RANDOM}};
  image_1_229 = _RAND_805[3:0];
  _RAND_806 = {1{`RANDOM}};
  image_1_230 = _RAND_806[3:0];
  _RAND_807 = {1{`RANDOM}};
  image_1_231 = _RAND_807[3:0];
  _RAND_808 = {1{`RANDOM}};
  image_1_232 = _RAND_808[3:0];
  _RAND_809 = {1{`RANDOM}};
  image_1_233 = _RAND_809[3:0];
  _RAND_810 = {1{`RANDOM}};
  image_1_234 = _RAND_810[3:0];
  _RAND_811 = {1{`RANDOM}};
  image_1_235 = _RAND_811[3:0];
  _RAND_812 = {1{`RANDOM}};
  image_1_236 = _RAND_812[3:0];
  _RAND_813 = {1{`RANDOM}};
  image_1_237 = _RAND_813[3:0];
  _RAND_814 = {1{`RANDOM}};
  image_1_238 = _RAND_814[3:0];
  _RAND_815 = {1{`RANDOM}};
  image_1_239 = _RAND_815[3:0];
  _RAND_816 = {1{`RANDOM}};
  image_1_240 = _RAND_816[3:0];
  _RAND_817 = {1{`RANDOM}};
  image_1_241 = _RAND_817[3:0];
  _RAND_818 = {1{`RANDOM}};
  image_1_242 = _RAND_818[3:0];
  _RAND_819 = {1{`RANDOM}};
  image_1_243 = _RAND_819[3:0];
  _RAND_820 = {1{`RANDOM}};
  image_1_244 = _RAND_820[3:0];
  _RAND_821 = {1{`RANDOM}};
  image_1_245 = _RAND_821[3:0];
  _RAND_822 = {1{`RANDOM}};
  image_1_246 = _RAND_822[3:0];
  _RAND_823 = {1{`RANDOM}};
  image_1_247 = _RAND_823[3:0];
  _RAND_824 = {1{`RANDOM}};
  image_1_248 = _RAND_824[3:0];
  _RAND_825 = {1{`RANDOM}};
  image_1_249 = _RAND_825[3:0];
  _RAND_826 = {1{`RANDOM}};
  image_1_250 = _RAND_826[3:0];
  _RAND_827 = {1{`RANDOM}};
  image_1_251 = _RAND_827[3:0];
  _RAND_828 = {1{`RANDOM}};
  image_1_252 = _RAND_828[3:0];
  _RAND_829 = {1{`RANDOM}};
  image_1_253 = _RAND_829[3:0];
  _RAND_830 = {1{`RANDOM}};
  image_1_254 = _RAND_830[3:0];
  _RAND_831 = {1{`RANDOM}};
  image_1_255 = _RAND_831[3:0];
  _RAND_832 = {1{`RANDOM}};
  image_1_256 = _RAND_832[3:0];
  _RAND_833 = {1{`RANDOM}};
  image_1_257 = _RAND_833[3:0];
  _RAND_834 = {1{`RANDOM}};
  image_1_258 = _RAND_834[3:0];
  _RAND_835 = {1{`RANDOM}};
  image_1_259 = _RAND_835[3:0];
  _RAND_836 = {1{`RANDOM}};
  image_1_260 = _RAND_836[3:0];
  _RAND_837 = {1{`RANDOM}};
  image_1_261 = _RAND_837[3:0];
  _RAND_838 = {1{`RANDOM}};
  image_1_262 = _RAND_838[3:0];
  _RAND_839 = {1{`RANDOM}};
  image_1_263 = _RAND_839[3:0];
  _RAND_840 = {1{`RANDOM}};
  image_1_264 = _RAND_840[3:0];
  _RAND_841 = {1{`RANDOM}};
  image_1_265 = _RAND_841[3:0];
  _RAND_842 = {1{`RANDOM}};
  image_1_266 = _RAND_842[3:0];
  _RAND_843 = {1{`RANDOM}};
  image_1_267 = _RAND_843[3:0];
  _RAND_844 = {1{`RANDOM}};
  image_1_268 = _RAND_844[3:0];
  _RAND_845 = {1{`RANDOM}};
  image_1_269 = _RAND_845[3:0];
  _RAND_846 = {1{`RANDOM}};
  image_1_270 = _RAND_846[3:0];
  _RAND_847 = {1{`RANDOM}};
  image_1_271 = _RAND_847[3:0];
  _RAND_848 = {1{`RANDOM}};
  image_1_272 = _RAND_848[3:0];
  _RAND_849 = {1{`RANDOM}};
  image_1_273 = _RAND_849[3:0];
  _RAND_850 = {1{`RANDOM}};
  image_1_274 = _RAND_850[3:0];
  _RAND_851 = {1{`RANDOM}};
  image_1_275 = _RAND_851[3:0];
  _RAND_852 = {1{`RANDOM}};
  image_1_276 = _RAND_852[3:0];
  _RAND_853 = {1{`RANDOM}};
  image_1_277 = _RAND_853[3:0];
  _RAND_854 = {1{`RANDOM}};
  image_1_278 = _RAND_854[3:0];
  _RAND_855 = {1{`RANDOM}};
  image_1_279 = _RAND_855[3:0];
  _RAND_856 = {1{`RANDOM}};
  image_1_280 = _RAND_856[3:0];
  _RAND_857 = {1{`RANDOM}};
  image_1_281 = _RAND_857[3:0];
  _RAND_858 = {1{`RANDOM}};
  image_1_282 = _RAND_858[3:0];
  _RAND_859 = {1{`RANDOM}};
  image_1_283 = _RAND_859[3:0];
  _RAND_860 = {1{`RANDOM}};
  image_1_284 = _RAND_860[3:0];
  _RAND_861 = {1{`RANDOM}};
  image_1_285 = _RAND_861[3:0];
  _RAND_862 = {1{`RANDOM}};
  image_1_286 = _RAND_862[3:0];
  _RAND_863 = {1{`RANDOM}};
  image_1_287 = _RAND_863[3:0];
  _RAND_864 = {1{`RANDOM}};
  image_1_288 = _RAND_864[3:0];
  _RAND_865 = {1{`RANDOM}};
  image_1_289 = _RAND_865[3:0];
  _RAND_866 = {1{`RANDOM}};
  image_1_290 = _RAND_866[3:0];
  _RAND_867 = {1{`RANDOM}};
  image_1_291 = _RAND_867[3:0];
  _RAND_868 = {1{`RANDOM}};
  image_1_292 = _RAND_868[3:0];
  _RAND_869 = {1{`RANDOM}};
  image_1_293 = _RAND_869[3:0];
  _RAND_870 = {1{`RANDOM}};
  image_1_294 = _RAND_870[3:0];
  _RAND_871 = {1{`RANDOM}};
  image_1_295 = _RAND_871[3:0];
  _RAND_872 = {1{`RANDOM}};
  image_1_296 = _RAND_872[3:0];
  _RAND_873 = {1{`RANDOM}};
  image_1_297 = _RAND_873[3:0];
  _RAND_874 = {1{`RANDOM}};
  image_1_298 = _RAND_874[3:0];
  _RAND_875 = {1{`RANDOM}};
  image_1_299 = _RAND_875[3:0];
  _RAND_876 = {1{`RANDOM}};
  image_1_300 = _RAND_876[3:0];
  _RAND_877 = {1{`RANDOM}};
  image_1_301 = _RAND_877[3:0];
  _RAND_878 = {1{`RANDOM}};
  image_1_302 = _RAND_878[3:0];
  _RAND_879 = {1{`RANDOM}};
  image_1_303 = _RAND_879[3:0];
  _RAND_880 = {1{`RANDOM}};
  image_1_304 = _RAND_880[3:0];
  _RAND_881 = {1{`RANDOM}};
  image_1_305 = _RAND_881[3:0];
  _RAND_882 = {1{`RANDOM}};
  image_1_306 = _RAND_882[3:0];
  _RAND_883 = {1{`RANDOM}};
  image_1_307 = _RAND_883[3:0];
  _RAND_884 = {1{`RANDOM}};
  image_1_308 = _RAND_884[3:0];
  _RAND_885 = {1{`RANDOM}};
  image_1_309 = _RAND_885[3:0];
  _RAND_886 = {1{`RANDOM}};
  image_1_310 = _RAND_886[3:0];
  _RAND_887 = {1{`RANDOM}};
  image_1_311 = _RAND_887[3:0];
  _RAND_888 = {1{`RANDOM}};
  image_1_312 = _RAND_888[3:0];
  _RAND_889 = {1{`RANDOM}};
  image_1_313 = _RAND_889[3:0];
  _RAND_890 = {1{`RANDOM}};
  image_1_314 = _RAND_890[3:0];
  _RAND_891 = {1{`RANDOM}};
  image_1_315 = _RAND_891[3:0];
  _RAND_892 = {1{`RANDOM}};
  image_1_316 = _RAND_892[3:0];
  _RAND_893 = {1{`RANDOM}};
  image_1_317 = _RAND_893[3:0];
  _RAND_894 = {1{`RANDOM}};
  image_1_318 = _RAND_894[3:0];
  _RAND_895 = {1{`RANDOM}};
  image_1_319 = _RAND_895[3:0];
  _RAND_896 = {1{`RANDOM}};
  image_1_320 = _RAND_896[3:0];
  _RAND_897 = {1{`RANDOM}};
  image_1_321 = _RAND_897[3:0];
  _RAND_898 = {1{`RANDOM}};
  image_1_322 = _RAND_898[3:0];
  _RAND_899 = {1{`RANDOM}};
  image_1_323 = _RAND_899[3:0];
  _RAND_900 = {1{`RANDOM}};
  image_1_324 = _RAND_900[3:0];
  _RAND_901 = {1{`RANDOM}};
  image_1_325 = _RAND_901[3:0];
  _RAND_902 = {1{`RANDOM}};
  image_1_326 = _RAND_902[3:0];
  _RAND_903 = {1{`RANDOM}};
  image_1_327 = _RAND_903[3:0];
  _RAND_904 = {1{`RANDOM}};
  image_1_328 = _RAND_904[3:0];
  _RAND_905 = {1{`RANDOM}};
  image_1_329 = _RAND_905[3:0];
  _RAND_906 = {1{`RANDOM}};
  image_1_330 = _RAND_906[3:0];
  _RAND_907 = {1{`RANDOM}};
  image_1_331 = _RAND_907[3:0];
  _RAND_908 = {1{`RANDOM}};
  image_1_332 = _RAND_908[3:0];
  _RAND_909 = {1{`RANDOM}};
  image_1_333 = _RAND_909[3:0];
  _RAND_910 = {1{`RANDOM}};
  image_1_334 = _RAND_910[3:0];
  _RAND_911 = {1{`RANDOM}};
  image_1_335 = _RAND_911[3:0];
  _RAND_912 = {1{`RANDOM}};
  image_1_336 = _RAND_912[3:0];
  _RAND_913 = {1{`RANDOM}};
  image_1_337 = _RAND_913[3:0];
  _RAND_914 = {1{`RANDOM}};
  image_1_338 = _RAND_914[3:0];
  _RAND_915 = {1{`RANDOM}};
  image_1_339 = _RAND_915[3:0];
  _RAND_916 = {1{`RANDOM}};
  image_1_340 = _RAND_916[3:0];
  _RAND_917 = {1{`RANDOM}};
  image_1_341 = _RAND_917[3:0];
  _RAND_918 = {1{`RANDOM}};
  image_1_342 = _RAND_918[3:0];
  _RAND_919 = {1{`RANDOM}};
  image_1_343 = _RAND_919[3:0];
  _RAND_920 = {1{`RANDOM}};
  image_1_344 = _RAND_920[3:0];
  _RAND_921 = {1{`RANDOM}};
  image_1_345 = _RAND_921[3:0];
  _RAND_922 = {1{`RANDOM}};
  image_1_346 = _RAND_922[3:0];
  _RAND_923 = {1{`RANDOM}};
  image_1_347 = _RAND_923[3:0];
  _RAND_924 = {1{`RANDOM}};
  image_1_348 = _RAND_924[3:0];
  _RAND_925 = {1{`RANDOM}};
  image_1_349 = _RAND_925[3:0];
  _RAND_926 = {1{`RANDOM}};
  image_1_350 = _RAND_926[3:0];
  _RAND_927 = {1{`RANDOM}};
  image_1_351 = _RAND_927[3:0];
  _RAND_928 = {1{`RANDOM}};
  image_1_352 = _RAND_928[3:0];
  _RAND_929 = {1{`RANDOM}};
  image_1_353 = _RAND_929[3:0];
  _RAND_930 = {1{`RANDOM}};
  image_1_354 = _RAND_930[3:0];
  _RAND_931 = {1{`RANDOM}};
  image_1_355 = _RAND_931[3:0];
  _RAND_932 = {1{`RANDOM}};
  image_1_356 = _RAND_932[3:0];
  _RAND_933 = {1{`RANDOM}};
  image_1_357 = _RAND_933[3:0];
  _RAND_934 = {1{`RANDOM}};
  image_1_358 = _RAND_934[3:0];
  _RAND_935 = {1{`RANDOM}};
  image_1_359 = _RAND_935[3:0];
  _RAND_936 = {1{`RANDOM}};
  image_1_360 = _RAND_936[3:0];
  _RAND_937 = {1{`RANDOM}};
  image_1_361 = _RAND_937[3:0];
  _RAND_938 = {1{`RANDOM}};
  image_1_362 = _RAND_938[3:0];
  _RAND_939 = {1{`RANDOM}};
  image_1_363 = _RAND_939[3:0];
  _RAND_940 = {1{`RANDOM}};
  image_1_364 = _RAND_940[3:0];
  _RAND_941 = {1{`RANDOM}};
  image_1_365 = _RAND_941[3:0];
  _RAND_942 = {1{`RANDOM}};
  image_1_366 = _RAND_942[3:0];
  _RAND_943 = {1{`RANDOM}};
  image_1_367 = _RAND_943[3:0];
  _RAND_944 = {1{`RANDOM}};
  image_1_368 = _RAND_944[3:0];
  _RAND_945 = {1{`RANDOM}};
  image_1_369 = _RAND_945[3:0];
  _RAND_946 = {1{`RANDOM}};
  image_1_370 = _RAND_946[3:0];
  _RAND_947 = {1{`RANDOM}};
  image_1_371 = _RAND_947[3:0];
  _RAND_948 = {1{`RANDOM}};
  image_1_372 = _RAND_948[3:0];
  _RAND_949 = {1{`RANDOM}};
  image_1_373 = _RAND_949[3:0];
  _RAND_950 = {1{`RANDOM}};
  image_1_374 = _RAND_950[3:0];
  _RAND_951 = {1{`RANDOM}};
  image_1_375 = _RAND_951[3:0];
  _RAND_952 = {1{`RANDOM}};
  image_1_376 = _RAND_952[3:0];
  _RAND_953 = {1{`RANDOM}};
  image_1_377 = _RAND_953[3:0];
  _RAND_954 = {1{`RANDOM}};
  image_1_378 = _RAND_954[3:0];
  _RAND_955 = {1{`RANDOM}};
  image_1_379 = _RAND_955[3:0];
  _RAND_956 = {1{`RANDOM}};
  image_1_380 = _RAND_956[3:0];
  _RAND_957 = {1{`RANDOM}};
  image_1_381 = _RAND_957[3:0];
  _RAND_958 = {1{`RANDOM}};
  image_1_382 = _RAND_958[3:0];
  _RAND_959 = {1{`RANDOM}};
  image_1_383 = _RAND_959[3:0];
  _RAND_960 = {1{`RANDOM}};
  image_1_384 = _RAND_960[3:0];
  _RAND_961 = {1{`RANDOM}};
  image_1_385 = _RAND_961[3:0];
  _RAND_962 = {1{`RANDOM}};
  image_1_386 = _RAND_962[3:0];
  _RAND_963 = {1{`RANDOM}};
  image_1_387 = _RAND_963[3:0];
  _RAND_964 = {1{`RANDOM}};
  image_1_388 = _RAND_964[3:0];
  _RAND_965 = {1{`RANDOM}};
  image_1_389 = _RAND_965[3:0];
  _RAND_966 = {1{`RANDOM}};
  image_1_390 = _RAND_966[3:0];
  _RAND_967 = {1{`RANDOM}};
  image_1_391 = _RAND_967[3:0];
  _RAND_968 = {1{`RANDOM}};
  image_1_392 = _RAND_968[3:0];
  _RAND_969 = {1{`RANDOM}};
  image_1_393 = _RAND_969[3:0];
  _RAND_970 = {1{`RANDOM}};
  image_1_394 = _RAND_970[3:0];
  _RAND_971 = {1{`RANDOM}};
  image_1_395 = _RAND_971[3:0];
  _RAND_972 = {1{`RANDOM}};
  image_1_396 = _RAND_972[3:0];
  _RAND_973 = {1{`RANDOM}};
  image_1_397 = _RAND_973[3:0];
  _RAND_974 = {1{`RANDOM}};
  image_1_398 = _RAND_974[3:0];
  _RAND_975 = {1{`RANDOM}};
  image_1_399 = _RAND_975[3:0];
  _RAND_976 = {1{`RANDOM}};
  image_1_400 = _RAND_976[3:0];
  _RAND_977 = {1{`RANDOM}};
  image_1_401 = _RAND_977[3:0];
  _RAND_978 = {1{`RANDOM}};
  image_1_402 = _RAND_978[3:0];
  _RAND_979 = {1{`RANDOM}};
  image_1_403 = _RAND_979[3:0];
  _RAND_980 = {1{`RANDOM}};
  image_1_404 = _RAND_980[3:0];
  _RAND_981 = {1{`RANDOM}};
  image_1_405 = _RAND_981[3:0];
  _RAND_982 = {1{`RANDOM}};
  image_1_406 = _RAND_982[3:0];
  _RAND_983 = {1{`RANDOM}};
  image_1_407 = _RAND_983[3:0];
  _RAND_984 = {1{`RANDOM}};
  image_1_408 = _RAND_984[3:0];
  _RAND_985 = {1{`RANDOM}};
  image_1_409 = _RAND_985[3:0];
  _RAND_986 = {1{`RANDOM}};
  image_1_410 = _RAND_986[3:0];
  _RAND_987 = {1{`RANDOM}};
  image_1_411 = _RAND_987[3:0];
  _RAND_988 = {1{`RANDOM}};
  image_1_412 = _RAND_988[3:0];
  _RAND_989 = {1{`RANDOM}};
  image_1_413 = _RAND_989[3:0];
  _RAND_990 = {1{`RANDOM}};
  image_1_414 = _RAND_990[3:0];
  _RAND_991 = {1{`RANDOM}};
  image_1_415 = _RAND_991[3:0];
  _RAND_992 = {1{`RANDOM}};
  image_1_416 = _RAND_992[3:0];
  _RAND_993 = {1{`RANDOM}};
  image_1_417 = _RAND_993[3:0];
  _RAND_994 = {1{`RANDOM}};
  image_1_418 = _RAND_994[3:0];
  _RAND_995 = {1{`RANDOM}};
  image_1_419 = _RAND_995[3:0];
  _RAND_996 = {1{`RANDOM}};
  image_1_420 = _RAND_996[3:0];
  _RAND_997 = {1{`RANDOM}};
  image_1_421 = _RAND_997[3:0];
  _RAND_998 = {1{`RANDOM}};
  image_1_422 = _RAND_998[3:0];
  _RAND_999 = {1{`RANDOM}};
  image_1_423 = _RAND_999[3:0];
  _RAND_1000 = {1{`RANDOM}};
  image_1_424 = _RAND_1000[3:0];
  _RAND_1001 = {1{`RANDOM}};
  image_1_425 = _RAND_1001[3:0];
  _RAND_1002 = {1{`RANDOM}};
  image_1_426 = _RAND_1002[3:0];
  _RAND_1003 = {1{`RANDOM}};
  image_1_427 = _RAND_1003[3:0];
  _RAND_1004 = {1{`RANDOM}};
  image_1_428 = _RAND_1004[3:0];
  _RAND_1005 = {1{`RANDOM}};
  image_1_429 = _RAND_1005[3:0];
  _RAND_1006 = {1{`RANDOM}};
  image_1_430 = _RAND_1006[3:0];
  _RAND_1007 = {1{`RANDOM}};
  image_1_431 = _RAND_1007[3:0];
  _RAND_1008 = {1{`RANDOM}};
  image_1_432 = _RAND_1008[3:0];
  _RAND_1009 = {1{`RANDOM}};
  image_1_433 = _RAND_1009[3:0];
  _RAND_1010 = {1{`RANDOM}};
  image_1_434 = _RAND_1010[3:0];
  _RAND_1011 = {1{`RANDOM}};
  image_1_435 = _RAND_1011[3:0];
  _RAND_1012 = {1{`RANDOM}};
  image_1_436 = _RAND_1012[3:0];
  _RAND_1013 = {1{`RANDOM}};
  image_1_437 = _RAND_1013[3:0];
  _RAND_1014 = {1{`RANDOM}};
  image_1_438 = _RAND_1014[3:0];
  _RAND_1015 = {1{`RANDOM}};
  image_1_439 = _RAND_1015[3:0];
  _RAND_1016 = {1{`RANDOM}};
  image_1_440 = _RAND_1016[3:0];
  _RAND_1017 = {1{`RANDOM}};
  image_1_441 = _RAND_1017[3:0];
  _RAND_1018 = {1{`RANDOM}};
  image_1_442 = _RAND_1018[3:0];
  _RAND_1019 = {1{`RANDOM}};
  image_1_443 = _RAND_1019[3:0];
  _RAND_1020 = {1{`RANDOM}};
  image_1_444 = _RAND_1020[3:0];
  _RAND_1021 = {1{`RANDOM}};
  image_1_445 = _RAND_1021[3:0];
  _RAND_1022 = {1{`RANDOM}};
  image_1_446 = _RAND_1022[3:0];
  _RAND_1023 = {1{`RANDOM}};
  image_1_447 = _RAND_1023[3:0];
  _RAND_1024 = {1{`RANDOM}};
  image_1_448 = _RAND_1024[3:0];
  _RAND_1025 = {1{`RANDOM}};
  image_1_449 = _RAND_1025[3:0];
  _RAND_1026 = {1{`RANDOM}};
  image_1_450 = _RAND_1026[3:0];
  _RAND_1027 = {1{`RANDOM}};
  image_1_451 = _RAND_1027[3:0];
  _RAND_1028 = {1{`RANDOM}};
  image_1_452 = _RAND_1028[3:0];
  _RAND_1029 = {1{`RANDOM}};
  image_1_453 = _RAND_1029[3:0];
  _RAND_1030 = {1{`RANDOM}};
  image_1_454 = _RAND_1030[3:0];
  _RAND_1031 = {1{`RANDOM}};
  image_1_455 = _RAND_1031[3:0];
  _RAND_1032 = {1{`RANDOM}};
  image_1_456 = _RAND_1032[3:0];
  _RAND_1033 = {1{`RANDOM}};
  image_1_457 = _RAND_1033[3:0];
  _RAND_1034 = {1{`RANDOM}};
  image_1_458 = _RAND_1034[3:0];
  _RAND_1035 = {1{`RANDOM}};
  image_1_459 = _RAND_1035[3:0];
  _RAND_1036 = {1{`RANDOM}};
  image_1_460 = _RAND_1036[3:0];
  _RAND_1037 = {1{`RANDOM}};
  image_1_461 = _RAND_1037[3:0];
  _RAND_1038 = {1{`RANDOM}};
  image_1_462 = _RAND_1038[3:0];
  _RAND_1039 = {1{`RANDOM}};
  image_1_463 = _RAND_1039[3:0];
  _RAND_1040 = {1{`RANDOM}};
  image_1_464 = _RAND_1040[3:0];
  _RAND_1041 = {1{`RANDOM}};
  image_1_465 = _RAND_1041[3:0];
  _RAND_1042 = {1{`RANDOM}};
  image_1_466 = _RAND_1042[3:0];
  _RAND_1043 = {1{`RANDOM}};
  image_1_467 = _RAND_1043[3:0];
  _RAND_1044 = {1{`RANDOM}};
  image_1_468 = _RAND_1044[3:0];
  _RAND_1045 = {1{`RANDOM}};
  image_1_469 = _RAND_1045[3:0];
  _RAND_1046 = {1{`RANDOM}};
  image_1_470 = _RAND_1046[3:0];
  _RAND_1047 = {1{`RANDOM}};
  image_1_471 = _RAND_1047[3:0];
  _RAND_1048 = {1{`RANDOM}};
  image_1_472 = _RAND_1048[3:0];
  _RAND_1049 = {1{`RANDOM}};
  image_1_473 = _RAND_1049[3:0];
  _RAND_1050 = {1{`RANDOM}};
  image_1_474 = _RAND_1050[3:0];
  _RAND_1051 = {1{`RANDOM}};
  image_1_475 = _RAND_1051[3:0];
  _RAND_1052 = {1{`RANDOM}};
  image_1_476 = _RAND_1052[3:0];
  _RAND_1053 = {1{`RANDOM}};
  image_1_477 = _RAND_1053[3:0];
  _RAND_1054 = {1{`RANDOM}};
  image_1_478 = _RAND_1054[3:0];
  _RAND_1055 = {1{`RANDOM}};
  image_1_479 = _RAND_1055[3:0];
  _RAND_1056 = {1{`RANDOM}};
  image_1_480 = _RAND_1056[3:0];
  _RAND_1057 = {1{`RANDOM}};
  image_1_481 = _RAND_1057[3:0];
  _RAND_1058 = {1{`RANDOM}};
  image_1_482 = _RAND_1058[3:0];
  _RAND_1059 = {1{`RANDOM}};
  image_1_483 = _RAND_1059[3:0];
  _RAND_1060 = {1{`RANDOM}};
  image_1_484 = _RAND_1060[3:0];
  _RAND_1061 = {1{`RANDOM}};
  image_1_485 = _RAND_1061[3:0];
  _RAND_1062 = {1{`RANDOM}};
  image_1_486 = _RAND_1062[3:0];
  _RAND_1063 = {1{`RANDOM}};
  image_1_487 = _RAND_1063[3:0];
  _RAND_1064 = {1{`RANDOM}};
  image_1_488 = _RAND_1064[3:0];
  _RAND_1065 = {1{`RANDOM}};
  image_1_489 = _RAND_1065[3:0];
  _RAND_1066 = {1{`RANDOM}};
  image_1_490 = _RAND_1066[3:0];
  _RAND_1067 = {1{`RANDOM}};
  image_1_491 = _RAND_1067[3:0];
  _RAND_1068 = {1{`RANDOM}};
  image_1_492 = _RAND_1068[3:0];
  _RAND_1069 = {1{`RANDOM}};
  image_1_493 = _RAND_1069[3:0];
  _RAND_1070 = {1{`RANDOM}};
  image_1_494 = _RAND_1070[3:0];
  _RAND_1071 = {1{`RANDOM}};
  image_1_495 = _RAND_1071[3:0];
  _RAND_1072 = {1{`RANDOM}};
  image_1_496 = _RAND_1072[3:0];
  _RAND_1073 = {1{`RANDOM}};
  image_1_497 = _RAND_1073[3:0];
  _RAND_1074 = {1{`RANDOM}};
  image_1_498 = _RAND_1074[3:0];
  _RAND_1075 = {1{`RANDOM}};
  image_1_499 = _RAND_1075[3:0];
  _RAND_1076 = {1{`RANDOM}};
  image_1_500 = _RAND_1076[3:0];
  _RAND_1077 = {1{`RANDOM}};
  image_1_501 = _RAND_1077[3:0];
  _RAND_1078 = {1{`RANDOM}};
  image_1_502 = _RAND_1078[3:0];
  _RAND_1079 = {1{`RANDOM}};
  image_1_503 = _RAND_1079[3:0];
  _RAND_1080 = {1{`RANDOM}};
  image_1_504 = _RAND_1080[3:0];
  _RAND_1081 = {1{`RANDOM}};
  image_1_505 = _RAND_1081[3:0];
  _RAND_1082 = {1{`RANDOM}};
  image_1_506 = _RAND_1082[3:0];
  _RAND_1083 = {1{`RANDOM}};
  image_1_507 = _RAND_1083[3:0];
  _RAND_1084 = {1{`RANDOM}};
  image_1_508 = _RAND_1084[3:0];
  _RAND_1085 = {1{`RANDOM}};
  image_1_509 = _RAND_1085[3:0];
  _RAND_1086 = {1{`RANDOM}};
  image_1_510 = _RAND_1086[3:0];
  _RAND_1087 = {1{`RANDOM}};
  image_1_511 = _RAND_1087[3:0];
  _RAND_1088 = {1{`RANDOM}};
  image_1_512 = _RAND_1088[3:0];
  _RAND_1089 = {1{`RANDOM}};
  image_1_513 = _RAND_1089[3:0];
  _RAND_1090 = {1{`RANDOM}};
  image_1_514 = _RAND_1090[3:0];
  _RAND_1091 = {1{`RANDOM}};
  image_1_515 = _RAND_1091[3:0];
  _RAND_1092 = {1{`RANDOM}};
  image_1_516 = _RAND_1092[3:0];
  _RAND_1093 = {1{`RANDOM}};
  image_1_517 = _RAND_1093[3:0];
  _RAND_1094 = {1{`RANDOM}};
  image_1_518 = _RAND_1094[3:0];
  _RAND_1095 = {1{`RANDOM}};
  image_1_519 = _RAND_1095[3:0];
  _RAND_1096 = {1{`RANDOM}};
  image_1_520 = _RAND_1096[3:0];
  _RAND_1097 = {1{`RANDOM}};
  image_1_521 = _RAND_1097[3:0];
  _RAND_1098 = {1{`RANDOM}};
  image_1_522 = _RAND_1098[3:0];
  _RAND_1099 = {1{`RANDOM}};
  image_1_523 = _RAND_1099[3:0];
  _RAND_1100 = {1{`RANDOM}};
  image_1_524 = _RAND_1100[3:0];
  _RAND_1101 = {1{`RANDOM}};
  image_1_525 = _RAND_1101[3:0];
  _RAND_1102 = {1{`RANDOM}};
  image_1_526 = _RAND_1102[3:0];
  _RAND_1103 = {1{`RANDOM}};
  image_1_527 = _RAND_1103[3:0];
  _RAND_1104 = {1{`RANDOM}};
  image_1_528 = _RAND_1104[3:0];
  _RAND_1105 = {1{`RANDOM}};
  image_1_529 = _RAND_1105[3:0];
  _RAND_1106 = {1{`RANDOM}};
  image_1_530 = _RAND_1106[3:0];
  _RAND_1107 = {1{`RANDOM}};
  image_1_531 = _RAND_1107[3:0];
  _RAND_1108 = {1{`RANDOM}};
  image_1_532 = _RAND_1108[3:0];
  _RAND_1109 = {1{`RANDOM}};
  image_1_533 = _RAND_1109[3:0];
  _RAND_1110 = {1{`RANDOM}};
  image_1_534 = _RAND_1110[3:0];
  _RAND_1111 = {1{`RANDOM}};
  image_1_535 = _RAND_1111[3:0];
  _RAND_1112 = {1{`RANDOM}};
  image_1_536 = _RAND_1112[3:0];
  _RAND_1113 = {1{`RANDOM}};
  image_1_537 = _RAND_1113[3:0];
  _RAND_1114 = {1{`RANDOM}};
  image_1_538 = _RAND_1114[3:0];
  _RAND_1115 = {1{`RANDOM}};
  image_1_539 = _RAND_1115[3:0];
  _RAND_1116 = {1{`RANDOM}};
  image_1_540 = _RAND_1116[3:0];
  _RAND_1117 = {1{`RANDOM}};
  image_1_541 = _RAND_1117[3:0];
  _RAND_1118 = {1{`RANDOM}};
  image_1_542 = _RAND_1118[3:0];
  _RAND_1119 = {1{`RANDOM}};
  image_1_543 = _RAND_1119[3:0];
  _RAND_1120 = {1{`RANDOM}};
  image_1_544 = _RAND_1120[3:0];
  _RAND_1121 = {1{`RANDOM}};
  image_1_545 = _RAND_1121[3:0];
  _RAND_1122 = {1{`RANDOM}};
  image_1_546 = _RAND_1122[3:0];
  _RAND_1123 = {1{`RANDOM}};
  image_1_547 = _RAND_1123[3:0];
  _RAND_1124 = {1{`RANDOM}};
  image_1_548 = _RAND_1124[3:0];
  _RAND_1125 = {1{`RANDOM}};
  image_1_549 = _RAND_1125[3:0];
  _RAND_1126 = {1{`RANDOM}};
  image_1_550 = _RAND_1126[3:0];
  _RAND_1127 = {1{`RANDOM}};
  image_1_551 = _RAND_1127[3:0];
  _RAND_1128 = {1{`RANDOM}};
  image_1_552 = _RAND_1128[3:0];
  _RAND_1129 = {1{`RANDOM}};
  image_1_553 = _RAND_1129[3:0];
  _RAND_1130 = {1{`RANDOM}};
  image_1_554 = _RAND_1130[3:0];
  _RAND_1131 = {1{`RANDOM}};
  image_1_555 = _RAND_1131[3:0];
  _RAND_1132 = {1{`RANDOM}};
  image_1_556 = _RAND_1132[3:0];
  _RAND_1133 = {1{`RANDOM}};
  image_1_557 = _RAND_1133[3:0];
  _RAND_1134 = {1{`RANDOM}};
  image_1_558 = _RAND_1134[3:0];
  _RAND_1135 = {1{`RANDOM}};
  image_1_559 = _RAND_1135[3:0];
  _RAND_1136 = {1{`RANDOM}};
  image_1_560 = _RAND_1136[3:0];
  _RAND_1137 = {1{`RANDOM}};
  image_1_561 = _RAND_1137[3:0];
  _RAND_1138 = {1{`RANDOM}};
  image_1_562 = _RAND_1138[3:0];
  _RAND_1139 = {1{`RANDOM}};
  image_1_563 = _RAND_1139[3:0];
  _RAND_1140 = {1{`RANDOM}};
  image_1_564 = _RAND_1140[3:0];
  _RAND_1141 = {1{`RANDOM}};
  image_1_565 = _RAND_1141[3:0];
  _RAND_1142 = {1{`RANDOM}};
  image_1_566 = _RAND_1142[3:0];
  _RAND_1143 = {1{`RANDOM}};
  image_1_567 = _RAND_1143[3:0];
  _RAND_1144 = {1{`RANDOM}};
  image_1_568 = _RAND_1144[3:0];
  _RAND_1145 = {1{`RANDOM}};
  image_1_569 = _RAND_1145[3:0];
  _RAND_1146 = {1{`RANDOM}};
  image_1_570 = _RAND_1146[3:0];
  _RAND_1147 = {1{`RANDOM}};
  image_1_571 = _RAND_1147[3:0];
  _RAND_1148 = {1{`RANDOM}};
  image_1_572 = _RAND_1148[3:0];
  _RAND_1149 = {1{`RANDOM}};
  image_1_573 = _RAND_1149[3:0];
  _RAND_1150 = {1{`RANDOM}};
  image_1_574 = _RAND_1150[3:0];
  _RAND_1151 = {1{`RANDOM}};
  image_1_575 = _RAND_1151[3:0];
  _RAND_1152 = {1{`RANDOM}};
  image_2_0 = _RAND_1152[3:0];
  _RAND_1153 = {1{`RANDOM}};
  image_2_1 = _RAND_1153[3:0];
  _RAND_1154 = {1{`RANDOM}};
  image_2_2 = _RAND_1154[3:0];
  _RAND_1155 = {1{`RANDOM}};
  image_2_3 = _RAND_1155[3:0];
  _RAND_1156 = {1{`RANDOM}};
  image_2_4 = _RAND_1156[3:0];
  _RAND_1157 = {1{`RANDOM}};
  image_2_5 = _RAND_1157[3:0];
  _RAND_1158 = {1{`RANDOM}};
  image_2_6 = _RAND_1158[3:0];
  _RAND_1159 = {1{`RANDOM}};
  image_2_7 = _RAND_1159[3:0];
  _RAND_1160 = {1{`RANDOM}};
  image_2_8 = _RAND_1160[3:0];
  _RAND_1161 = {1{`RANDOM}};
  image_2_9 = _RAND_1161[3:0];
  _RAND_1162 = {1{`RANDOM}};
  image_2_10 = _RAND_1162[3:0];
  _RAND_1163 = {1{`RANDOM}};
  image_2_11 = _RAND_1163[3:0];
  _RAND_1164 = {1{`RANDOM}};
  image_2_12 = _RAND_1164[3:0];
  _RAND_1165 = {1{`RANDOM}};
  image_2_13 = _RAND_1165[3:0];
  _RAND_1166 = {1{`RANDOM}};
  image_2_14 = _RAND_1166[3:0];
  _RAND_1167 = {1{`RANDOM}};
  image_2_15 = _RAND_1167[3:0];
  _RAND_1168 = {1{`RANDOM}};
  image_2_16 = _RAND_1168[3:0];
  _RAND_1169 = {1{`RANDOM}};
  image_2_17 = _RAND_1169[3:0];
  _RAND_1170 = {1{`RANDOM}};
  image_2_18 = _RAND_1170[3:0];
  _RAND_1171 = {1{`RANDOM}};
  image_2_19 = _RAND_1171[3:0];
  _RAND_1172 = {1{`RANDOM}};
  image_2_20 = _RAND_1172[3:0];
  _RAND_1173 = {1{`RANDOM}};
  image_2_21 = _RAND_1173[3:0];
  _RAND_1174 = {1{`RANDOM}};
  image_2_22 = _RAND_1174[3:0];
  _RAND_1175 = {1{`RANDOM}};
  image_2_23 = _RAND_1175[3:0];
  _RAND_1176 = {1{`RANDOM}};
  image_2_24 = _RAND_1176[3:0];
  _RAND_1177 = {1{`RANDOM}};
  image_2_25 = _RAND_1177[3:0];
  _RAND_1178 = {1{`RANDOM}};
  image_2_26 = _RAND_1178[3:0];
  _RAND_1179 = {1{`RANDOM}};
  image_2_27 = _RAND_1179[3:0];
  _RAND_1180 = {1{`RANDOM}};
  image_2_28 = _RAND_1180[3:0];
  _RAND_1181 = {1{`RANDOM}};
  image_2_29 = _RAND_1181[3:0];
  _RAND_1182 = {1{`RANDOM}};
  image_2_30 = _RAND_1182[3:0];
  _RAND_1183 = {1{`RANDOM}};
  image_2_31 = _RAND_1183[3:0];
  _RAND_1184 = {1{`RANDOM}};
  image_2_32 = _RAND_1184[3:0];
  _RAND_1185 = {1{`RANDOM}};
  image_2_33 = _RAND_1185[3:0];
  _RAND_1186 = {1{`RANDOM}};
  image_2_34 = _RAND_1186[3:0];
  _RAND_1187 = {1{`RANDOM}};
  image_2_35 = _RAND_1187[3:0];
  _RAND_1188 = {1{`RANDOM}};
  image_2_36 = _RAND_1188[3:0];
  _RAND_1189 = {1{`RANDOM}};
  image_2_37 = _RAND_1189[3:0];
  _RAND_1190 = {1{`RANDOM}};
  image_2_38 = _RAND_1190[3:0];
  _RAND_1191 = {1{`RANDOM}};
  image_2_39 = _RAND_1191[3:0];
  _RAND_1192 = {1{`RANDOM}};
  image_2_40 = _RAND_1192[3:0];
  _RAND_1193 = {1{`RANDOM}};
  image_2_41 = _RAND_1193[3:0];
  _RAND_1194 = {1{`RANDOM}};
  image_2_42 = _RAND_1194[3:0];
  _RAND_1195 = {1{`RANDOM}};
  image_2_43 = _RAND_1195[3:0];
  _RAND_1196 = {1{`RANDOM}};
  image_2_44 = _RAND_1196[3:0];
  _RAND_1197 = {1{`RANDOM}};
  image_2_45 = _RAND_1197[3:0];
  _RAND_1198 = {1{`RANDOM}};
  image_2_46 = _RAND_1198[3:0];
  _RAND_1199 = {1{`RANDOM}};
  image_2_47 = _RAND_1199[3:0];
  _RAND_1200 = {1{`RANDOM}};
  image_2_48 = _RAND_1200[3:0];
  _RAND_1201 = {1{`RANDOM}};
  image_2_49 = _RAND_1201[3:0];
  _RAND_1202 = {1{`RANDOM}};
  image_2_50 = _RAND_1202[3:0];
  _RAND_1203 = {1{`RANDOM}};
  image_2_51 = _RAND_1203[3:0];
  _RAND_1204 = {1{`RANDOM}};
  image_2_52 = _RAND_1204[3:0];
  _RAND_1205 = {1{`RANDOM}};
  image_2_53 = _RAND_1205[3:0];
  _RAND_1206 = {1{`RANDOM}};
  image_2_54 = _RAND_1206[3:0];
  _RAND_1207 = {1{`RANDOM}};
  image_2_55 = _RAND_1207[3:0];
  _RAND_1208 = {1{`RANDOM}};
  image_2_56 = _RAND_1208[3:0];
  _RAND_1209 = {1{`RANDOM}};
  image_2_57 = _RAND_1209[3:0];
  _RAND_1210 = {1{`RANDOM}};
  image_2_58 = _RAND_1210[3:0];
  _RAND_1211 = {1{`RANDOM}};
  image_2_59 = _RAND_1211[3:0];
  _RAND_1212 = {1{`RANDOM}};
  image_2_60 = _RAND_1212[3:0];
  _RAND_1213 = {1{`RANDOM}};
  image_2_61 = _RAND_1213[3:0];
  _RAND_1214 = {1{`RANDOM}};
  image_2_62 = _RAND_1214[3:0];
  _RAND_1215 = {1{`RANDOM}};
  image_2_63 = _RAND_1215[3:0];
  _RAND_1216 = {1{`RANDOM}};
  image_2_64 = _RAND_1216[3:0];
  _RAND_1217 = {1{`RANDOM}};
  image_2_65 = _RAND_1217[3:0];
  _RAND_1218 = {1{`RANDOM}};
  image_2_66 = _RAND_1218[3:0];
  _RAND_1219 = {1{`RANDOM}};
  image_2_67 = _RAND_1219[3:0];
  _RAND_1220 = {1{`RANDOM}};
  image_2_68 = _RAND_1220[3:0];
  _RAND_1221 = {1{`RANDOM}};
  image_2_69 = _RAND_1221[3:0];
  _RAND_1222 = {1{`RANDOM}};
  image_2_70 = _RAND_1222[3:0];
  _RAND_1223 = {1{`RANDOM}};
  image_2_71 = _RAND_1223[3:0];
  _RAND_1224 = {1{`RANDOM}};
  image_2_72 = _RAND_1224[3:0];
  _RAND_1225 = {1{`RANDOM}};
  image_2_73 = _RAND_1225[3:0];
  _RAND_1226 = {1{`RANDOM}};
  image_2_74 = _RAND_1226[3:0];
  _RAND_1227 = {1{`RANDOM}};
  image_2_75 = _RAND_1227[3:0];
  _RAND_1228 = {1{`RANDOM}};
  image_2_76 = _RAND_1228[3:0];
  _RAND_1229 = {1{`RANDOM}};
  image_2_77 = _RAND_1229[3:0];
  _RAND_1230 = {1{`RANDOM}};
  image_2_78 = _RAND_1230[3:0];
  _RAND_1231 = {1{`RANDOM}};
  image_2_79 = _RAND_1231[3:0];
  _RAND_1232 = {1{`RANDOM}};
  image_2_80 = _RAND_1232[3:0];
  _RAND_1233 = {1{`RANDOM}};
  image_2_81 = _RAND_1233[3:0];
  _RAND_1234 = {1{`RANDOM}};
  image_2_82 = _RAND_1234[3:0];
  _RAND_1235 = {1{`RANDOM}};
  image_2_83 = _RAND_1235[3:0];
  _RAND_1236 = {1{`RANDOM}};
  image_2_84 = _RAND_1236[3:0];
  _RAND_1237 = {1{`RANDOM}};
  image_2_85 = _RAND_1237[3:0];
  _RAND_1238 = {1{`RANDOM}};
  image_2_86 = _RAND_1238[3:0];
  _RAND_1239 = {1{`RANDOM}};
  image_2_87 = _RAND_1239[3:0];
  _RAND_1240 = {1{`RANDOM}};
  image_2_88 = _RAND_1240[3:0];
  _RAND_1241 = {1{`RANDOM}};
  image_2_89 = _RAND_1241[3:0];
  _RAND_1242 = {1{`RANDOM}};
  image_2_90 = _RAND_1242[3:0];
  _RAND_1243 = {1{`RANDOM}};
  image_2_91 = _RAND_1243[3:0];
  _RAND_1244 = {1{`RANDOM}};
  image_2_92 = _RAND_1244[3:0];
  _RAND_1245 = {1{`RANDOM}};
  image_2_93 = _RAND_1245[3:0];
  _RAND_1246 = {1{`RANDOM}};
  image_2_94 = _RAND_1246[3:0];
  _RAND_1247 = {1{`RANDOM}};
  image_2_95 = _RAND_1247[3:0];
  _RAND_1248 = {1{`RANDOM}};
  image_2_96 = _RAND_1248[3:0];
  _RAND_1249 = {1{`RANDOM}};
  image_2_97 = _RAND_1249[3:0];
  _RAND_1250 = {1{`RANDOM}};
  image_2_98 = _RAND_1250[3:0];
  _RAND_1251 = {1{`RANDOM}};
  image_2_99 = _RAND_1251[3:0];
  _RAND_1252 = {1{`RANDOM}};
  image_2_100 = _RAND_1252[3:0];
  _RAND_1253 = {1{`RANDOM}};
  image_2_101 = _RAND_1253[3:0];
  _RAND_1254 = {1{`RANDOM}};
  image_2_102 = _RAND_1254[3:0];
  _RAND_1255 = {1{`RANDOM}};
  image_2_103 = _RAND_1255[3:0];
  _RAND_1256 = {1{`RANDOM}};
  image_2_104 = _RAND_1256[3:0];
  _RAND_1257 = {1{`RANDOM}};
  image_2_105 = _RAND_1257[3:0];
  _RAND_1258 = {1{`RANDOM}};
  image_2_106 = _RAND_1258[3:0];
  _RAND_1259 = {1{`RANDOM}};
  image_2_107 = _RAND_1259[3:0];
  _RAND_1260 = {1{`RANDOM}};
  image_2_108 = _RAND_1260[3:0];
  _RAND_1261 = {1{`RANDOM}};
  image_2_109 = _RAND_1261[3:0];
  _RAND_1262 = {1{`RANDOM}};
  image_2_110 = _RAND_1262[3:0];
  _RAND_1263 = {1{`RANDOM}};
  image_2_111 = _RAND_1263[3:0];
  _RAND_1264 = {1{`RANDOM}};
  image_2_112 = _RAND_1264[3:0];
  _RAND_1265 = {1{`RANDOM}};
  image_2_113 = _RAND_1265[3:0];
  _RAND_1266 = {1{`RANDOM}};
  image_2_114 = _RAND_1266[3:0];
  _RAND_1267 = {1{`RANDOM}};
  image_2_115 = _RAND_1267[3:0];
  _RAND_1268 = {1{`RANDOM}};
  image_2_116 = _RAND_1268[3:0];
  _RAND_1269 = {1{`RANDOM}};
  image_2_117 = _RAND_1269[3:0];
  _RAND_1270 = {1{`RANDOM}};
  image_2_118 = _RAND_1270[3:0];
  _RAND_1271 = {1{`RANDOM}};
  image_2_119 = _RAND_1271[3:0];
  _RAND_1272 = {1{`RANDOM}};
  image_2_120 = _RAND_1272[3:0];
  _RAND_1273 = {1{`RANDOM}};
  image_2_121 = _RAND_1273[3:0];
  _RAND_1274 = {1{`RANDOM}};
  image_2_122 = _RAND_1274[3:0];
  _RAND_1275 = {1{`RANDOM}};
  image_2_123 = _RAND_1275[3:0];
  _RAND_1276 = {1{`RANDOM}};
  image_2_124 = _RAND_1276[3:0];
  _RAND_1277 = {1{`RANDOM}};
  image_2_125 = _RAND_1277[3:0];
  _RAND_1278 = {1{`RANDOM}};
  image_2_126 = _RAND_1278[3:0];
  _RAND_1279 = {1{`RANDOM}};
  image_2_127 = _RAND_1279[3:0];
  _RAND_1280 = {1{`RANDOM}};
  image_2_128 = _RAND_1280[3:0];
  _RAND_1281 = {1{`RANDOM}};
  image_2_129 = _RAND_1281[3:0];
  _RAND_1282 = {1{`RANDOM}};
  image_2_130 = _RAND_1282[3:0];
  _RAND_1283 = {1{`RANDOM}};
  image_2_131 = _RAND_1283[3:0];
  _RAND_1284 = {1{`RANDOM}};
  image_2_132 = _RAND_1284[3:0];
  _RAND_1285 = {1{`RANDOM}};
  image_2_133 = _RAND_1285[3:0];
  _RAND_1286 = {1{`RANDOM}};
  image_2_134 = _RAND_1286[3:0];
  _RAND_1287 = {1{`RANDOM}};
  image_2_135 = _RAND_1287[3:0];
  _RAND_1288 = {1{`RANDOM}};
  image_2_136 = _RAND_1288[3:0];
  _RAND_1289 = {1{`RANDOM}};
  image_2_137 = _RAND_1289[3:0];
  _RAND_1290 = {1{`RANDOM}};
  image_2_138 = _RAND_1290[3:0];
  _RAND_1291 = {1{`RANDOM}};
  image_2_139 = _RAND_1291[3:0];
  _RAND_1292 = {1{`RANDOM}};
  image_2_140 = _RAND_1292[3:0];
  _RAND_1293 = {1{`RANDOM}};
  image_2_141 = _RAND_1293[3:0];
  _RAND_1294 = {1{`RANDOM}};
  image_2_142 = _RAND_1294[3:0];
  _RAND_1295 = {1{`RANDOM}};
  image_2_143 = _RAND_1295[3:0];
  _RAND_1296 = {1{`RANDOM}};
  image_2_144 = _RAND_1296[3:0];
  _RAND_1297 = {1{`RANDOM}};
  image_2_145 = _RAND_1297[3:0];
  _RAND_1298 = {1{`RANDOM}};
  image_2_146 = _RAND_1298[3:0];
  _RAND_1299 = {1{`RANDOM}};
  image_2_147 = _RAND_1299[3:0];
  _RAND_1300 = {1{`RANDOM}};
  image_2_148 = _RAND_1300[3:0];
  _RAND_1301 = {1{`RANDOM}};
  image_2_149 = _RAND_1301[3:0];
  _RAND_1302 = {1{`RANDOM}};
  image_2_150 = _RAND_1302[3:0];
  _RAND_1303 = {1{`RANDOM}};
  image_2_151 = _RAND_1303[3:0];
  _RAND_1304 = {1{`RANDOM}};
  image_2_152 = _RAND_1304[3:0];
  _RAND_1305 = {1{`RANDOM}};
  image_2_153 = _RAND_1305[3:0];
  _RAND_1306 = {1{`RANDOM}};
  image_2_154 = _RAND_1306[3:0];
  _RAND_1307 = {1{`RANDOM}};
  image_2_155 = _RAND_1307[3:0];
  _RAND_1308 = {1{`RANDOM}};
  image_2_156 = _RAND_1308[3:0];
  _RAND_1309 = {1{`RANDOM}};
  image_2_157 = _RAND_1309[3:0];
  _RAND_1310 = {1{`RANDOM}};
  image_2_158 = _RAND_1310[3:0];
  _RAND_1311 = {1{`RANDOM}};
  image_2_159 = _RAND_1311[3:0];
  _RAND_1312 = {1{`RANDOM}};
  image_2_160 = _RAND_1312[3:0];
  _RAND_1313 = {1{`RANDOM}};
  image_2_161 = _RAND_1313[3:0];
  _RAND_1314 = {1{`RANDOM}};
  image_2_162 = _RAND_1314[3:0];
  _RAND_1315 = {1{`RANDOM}};
  image_2_163 = _RAND_1315[3:0];
  _RAND_1316 = {1{`RANDOM}};
  image_2_164 = _RAND_1316[3:0];
  _RAND_1317 = {1{`RANDOM}};
  image_2_165 = _RAND_1317[3:0];
  _RAND_1318 = {1{`RANDOM}};
  image_2_166 = _RAND_1318[3:0];
  _RAND_1319 = {1{`RANDOM}};
  image_2_167 = _RAND_1319[3:0];
  _RAND_1320 = {1{`RANDOM}};
  image_2_168 = _RAND_1320[3:0];
  _RAND_1321 = {1{`RANDOM}};
  image_2_169 = _RAND_1321[3:0];
  _RAND_1322 = {1{`RANDOM}};
  image_2_170 = _RAND_1322[3:0];
  _RAND_1323 = {1{`RANDOM}};
  image_2_171 = _RAND_1323[3:0];
  _RAND_1324 = {1{`RANDOM}};
  image_2_172 = _RAND_1324[3:0];
  _RAND_1325 = {1{`RANDOM}};
  image_2_173 = _RAND_1325[3:0];
  _RAND_1326 = {1{`RANDOM}};
  image_2_174 = _RAND_1326[3:0];
  _RAND_1327 = {1{`RANDOM}};
  image_2_175 = _RAND_1327[3:0];
  _RAND_1328 = {1{`RANDOM}};
  image_2_176 = _RAND_1328[3:0];
  _RAND_1329 = {1{`RANDOM}};
  image_2_177 = _RAND_1329[3:0];
  _RAND_1330 = {1{`RANDOM}};
  image_2_178 = _RAND_1330[3:0];
  _RAND_1331 = {1{`RANDOM}};
  image_2_179 = _RAND_1331[3:0];
  _RAND_1332 = {1{`RANDOM}};
  image_2_180 = _RAND_1332[3:0];
  _RAND_1333 = {1{`RANDOM}};
  image_2_181 = _RAND_1333[3:0];
  _RAND_1334 = {1{`RANDOM}};
  image_2_182 = _RAND_1334[3:0];
  _RAND_1335 = {1{`RANDOM}};
  image_2_183 = _RAND_1335[3:0];
  _RAND_1336 = {1{`RANDOM}};
  image_2_184 = _RAND_1336[3:0];
  _RAND_1337 = {1{`RANDOM}};
  image_2_185 = _RAND_1337[3:0];
  _RAND_1338 = {1{`RANDOM}};
  image_2_186 = _RAND_1338[3:0];
  _RAND_1339 = {1{`RANDOM}};
  image_2_187 = _RAND_1339[3:0];
  _RAND_1340 = {1{`RANDOM}};
  image_2_188 = _RAND_1340[3:0];
  _RAND_1341 = {1{`RANDOM}};
  image_2_189 = _RAND_1341[3:0];
  _RAND_1342 = {1{`RANDOM}};
  image_2_190 = _RAND_1342[3:0];
  _RAND_1343 = {1{`RANDOM}};
  image_2_191 = _RAND_1343[3:0];
  _RAND_1344 = {1{`RANDOM}};
  image_2_192 = _RAND_1344[3:0];
  _RAND_1345 = {1{`RANDOM}};
  image_2_193 = _RAND_1345[3:0];
  _RAND_1346 = {1{`RANDOM}};
  image_2_194 = _RAND_1346[3:0];
  _RAND_1347 = {1{`RANDOM}};
  image_2_195 = _RAND_1347[3:0];
  _RAND_1348 = {1{`RANDOM}};
  image_2_196 = _RAND_1348[3:0];
  _RAND_1349 = {1{`RANDOM}};
  image_2_197 = _RAND_1349[3:0];
  _RAND_1350 = {1{`RANDOM}};
  image_2_198 = _RAND_1350[3:0];
  _RAND_1351 = {1{`RANDOM}};
  image_2_199 = _RAND_1351[3:0];
  _RAND_1352 = {1{`RANDOM}};
  image_2_200 = _RAND_1352[3:0];
  _RAND_1353 = {1{`RANDOM}};
  image_2_201 = _RAND_1353[3:0];
  _RAND_1354 = {1{`RANDOM}};
  image_2_202 = _RAND_1354[3:0];
  _RAND_1355 = {1{`RANDOM}};
  image_2_203 = _RAND_1355[3:0];
  _RAND_1356 = {1{`RANDOM}};
  image_2_204 = _RAND_1356[3:0];
  _RAND_1357 = {1{`RANDOM}};
  image_2_205 = _RAND_1357[3:0];
  _RAND_1358 = {1{`RANDOM}};
  image_2_206 = _RAND_1358[3:0];
  _RAND_1359 = {1{`RANDOM}};
  image_2_207 = _RAND_1359[3:0];
  _RAND_1360 = {1{`RANDOM}};
  image_2_208 = _RAND_1360[3:0];
  _RAND_1361 = {1{`RANDOM}};
  image_2_209 = _RAND_1361[3:0];
  _RAND_1362 = {1{`RANDOM}};
  image_2_210 = _RAND_1362[3:0];
  _RAND_1363 = {1{`RANDOM}};
  image_2_211 = _RAND_1363[3:0];
  _RAND_1364 = {1{`RANDOM}};
  image_2_212 = _RAND_1364[3:0];
  _RAND_1365 = {1{`RANDOM}};
  image_2_213 = _RAND_1365[3:0];
  _RAND_1366 = {1{`RANDOM}};
  image_2_214 = _RAND_1366[3:0];
  _RAND_1367 = {1{`RANDOM}};
  image_2_215 = _RAND_1367[3:0];
  _RAND_1368 = {1{`RANDOM}};
  image_2_216 = _RAND_1368[3:0];
  _RAND_1369 = {1{`RANDOM}};
  image_2_217 = _RAND_1369[3:0];
  _RAND_1370 = {1{`RANDOM}};
  image_2_218 = _RAND_1370[3:0];
  _RAND_1371 = {1{`RANDOM}};
  image_2_219 = _RAND_1371[3:0];
  _RAND_1372 = {1{`RANDOM}};
  image_2_220 = _RAND_1372[3:0];
  _RAND_1373 = {1{`RANDOM}};
  image_2_221 = _RAND_1373[3:0];
  _RAND_1374 = {1{`RANDOM}};
  image_2_222 = _RAND_1374[3:0];
  _RAND_1375 = {1{`RANDOM}};
  image_2_223 = _RAND_1375[3:0];
  _RAND_1376 = {1{`RANDOM}};
  image_2_224 = _RAND_1376[3:0];
  _RAND_1377 = {1{`RANDOM}};
  image_2_225 = _RAND_1377[3:0];
  _RAND_1378 = {1{`RANDOM}};
  image_2_226 = _RAND_1378[3:0];
  _RAND_1379 = {1{`RANDOM}};
  image_2_227 = _RAND_1379[3:0];
  _RAND_1380 = {1{`RANDOM}};
  image_2_228 = _RAND_1380[3:0];
  _RAND_1381 = {1{`RANDOM}};
  image_2_229 = _RAND_1381[3:0];
  _RAND_1382 = {1{`RANDOM}};
  image_2_230 = _RAND_1382[3:0];
  _RAND_1383 = {1{`RANDOM}};
  image_2_231 = _RAND_1383[3:0];
  _RAND_1384 = {1{`RANDOM}};
  image_2_232 = _RAND_1384[3:0];
  _RAND_1385 = {1{`RANDOM}};
  image_2_233 = _RAND_1385[3:0];
  _RAND_1386 = {1{`RANDOM}};
  image_2_234 = _RAND_1386[3:0];
  _RAND_1387 = {1{`RANDOM}};
  image_2_235 = _RAND_1387[3:0];
  _RAND_1388 = {1{`RANDOM}};
  image_2_236 = _RAND_1388[3:0];
  _RAND_1389 = {1{`RANDOM}};
  image_2_237 = _RAND_1389[3:0];
  _RAND_1390 = {1{`RANDOM}};
  image_2_238 = _RAND_1390[3:0];
  _RAND_1391 = {1{`RANDOM}};
  image_2_239 = _RAND_1391[3:0];
  _RAND_1392 = {1{`RANDOM}};
  image_2_240 = _RAND_1392[3:0];
  _RAND_1393 = {1{`RANDOM}};
  image_2_241 = _RAND_1393[3:0];
  _RAND_1394 = {1{`RANDOM}};
  image_2_242 = _RAND_1394[3:0];
  _RAND_1395 = {1{`RANDOM}};
  image_2_243 = _RAND_1395[3:0];
  _RAND_1396 = {1{`RANDOM}};
  image_2_244 = _RAND_1396[3:0];
  _RAND_1397 = {1{`RANDOM}};
  image_2_245 = _RAND_1397[3:0];
  _RAND_1398 = {1{`RANDOM}};
  image_2_246 = _RAND_1398[3:0];
  _RAND_1399 = {1{`RANDOM}};
  image_2_247 = _RAND_1399[3:0];
  _RAND_1400 = {1{`RANDOM}};
  image_2_248 = _RAND_1400[3:0];
  _RAND_1401 = {1{`RANDOM}};
  image_2_249 = _RAND_1401[3:0];
  _RAND_1402 = {1{`RANDOM}};
  image_2_250 = _RAND_1402[3:0];
  _RAND_1403 = {1{`RANDOM}};
  image_2_251 = _RAND_1403[3:0];
  _RAND_1404 = {1{`RANDOM}};
  image_2_252 = _RAND_1404[3:0];
  _RAND_1405 = {1{`RANDOM}};
  image_2_253 = _RAND_1405[3:0];
  _RAND_1406 = {1{`RANDOM}};
  image_2_254 = _RAND_1406[3:0];
  _RAND_1407 = {1{`RANDOM}};
  image_2_255 = _RAND_1407[3:0];
  _RAND_1408 = {1{`RANDOM}};
  image_2_256 = _RAND_1408[3:0];
  _RAND_1409 = {1{`RANDOM}};
  image_2_257 = _RAND_1409[3:0];
  _RAND_1410 = {1{`RANDOM}};
  image_2_258 = _RAND_1410[3:0];
  _RAND_1411 = {1{`RANDOM}};
  image_2_259 = _RAND_1411[3:0];
  _RAND_1412 = {1{`RANDOM}};
  image_2_260 = _RAND_1412[3:0];
  _RAND_1413 = {1{`RANDOM}};
  image_2_261 = _RAND_1413[3:0];
  _RAND_1414 = {1{`RANDOM}};
  image_2_262 = _RAND_1414[3:0];
  _RAND_1415 = {1{`RANDOM}};
  image_2_263 = _RAND_1415[3:0];
  _RAND_1416 = {1{`RANDOM}};
  image_2_264 = _RAND_1416[3:0];
  _RAND_1417 = {1{`RANDOM}};
  image_2_265 = _RAND_1417[3:0];
  _RAND_1418 = {1{`RANDOM}};
  image_2_266 = _RAND_1418[3:0];
  _RAND_1419 = {1{`RANDOM}};
  image_2_267 = _RAND_1419[3:0];
  _RAND_1420 = {1{`RANDOM}};
  image_2_268 = _RAND_1420[3:0];
  _RAND_1421 = {1{`RANDOM}};
  image_2_269 = _RAND_1421[3:0];
  _RAND_1422 = {1{`RANDOM}};
  image_2_270 = _RAND_1422[3:0];
  _RAND_1423 = {1{`RANDOM}};
  image_2_271 = _RAND_1423[3:0];
  _RAND_1424 = {1{`RANDOM}};
  image_2_272 = _RAND_1424[3:0];
  _RAND_1425 = {1{`RANDOM}};
  image_2_273 = _RAND_1425[3:0];
  _RAND_1426 = {1{`RANDOM}};
  image_2_274 = _RAND_1426[3:0];
  _RAND_1427 = {1{`RANDOM}};
  image_2_275 = _RAND_1427[3:0];
  _RAND_1428 = {1{`RANDOM}};
  image_2_276 = _RAND_1428[3:0];
  _RAND_1429 = {1{`RANDOM}};
  image_2_277 = _RAND_1429[3:0];
  _RAND_1430 = {1{`RANDOM}};
  image_2_278 = _RAND_1430[3:0];
  _RAND_1431 = {1{`RANDOM}};
  image_2_279 = _RAND_1431[3:0];
  _RAND_1432 = {1{`RANDOM}};
  image_2_280 = _RAND_1432[3:0];
  _RAND_1433 = {1{`RANDOM}};
  image_2_281 = _RAND_1433[3:0];
  _RAND_1434 = {1{`RANDOM}};
  image_2_282 = _RAND_1434[3:0];
  _RAND_1435 = {1{`RANDOM}};
  image_2_283 = _RAND_1435[3:0];
  _RAND_1436 = {1{`RANDOM}};
  image_2_284 = _RAND_1436[3:0];
  _RAND_1437 = {1{`RANDOM}};
  image_2_285 = _RAND_1437[3:0];
  _RAND_1438 = {1{`RANDOM}};
  image_2_286 = _RAND_1438[3:0];
  _RAND_1439 = {1{`RANDOM}};
  image_2_287 = _RAND_1439[3:0];
  _RAND_1440 = {1{`RANDOM}};
  image_2_288 = _RAND_1440[3:0];
  _RAND_1441 = {1{`RANDOM}};
  image_2_289 = _RAND_1441[3:0];
  _RAND_1442 = {1{`RANDOM}};
  image_2_290 = _RAND_1442[3:0];
  _RAND_1443 = {1{`RANDOM}};
  image_2_291 = _RAND_1443[3:0];
  _RAND_1444 = {1{`RANDOM}};
  image_2_292 = _RAND_1444[3:0];
  _RAND_1445 = {1{`RANDOM}};
  image_2_293 = _RAND_1445[3:0];
  _RAND_1446 = {1{`RANDOM}};
  image_2_294 = _RAND_1446[3:0];
  _RAND_1447 = {1{`RANDOM}};
  image_2_295 = _RAND_1447[3:0];
  _RAND_1448 = {1{`RANDOM}};
  image_2_296 = _RAND_1448[3:0];
  _RAND_1449 = {1{`RANDOM}};
  image_2_297 = _RAND_1449[3:0];
  _RAND_1450 = {1{`RANDOM}};
  image_2_298 = _RAND_1450[3:0];
  _RAND_1451 = {1{`RANDOM}};
  image_2_299 = _RAND_1451[3:0];
  _RAND_1452 = {1{`RANDOM}};
  image_2_300 = _RAND_1452[3:0];
  _RAND_1453 = {1{`RANDOM}};
  image_2_301 = _RAND_1453[3:0];
  _RAND_1454 = {1{`RANDOM}};
  image_2_302 = _RAND_1454[3:0];
  _RAND_1455 = {1{`RANDOM}};
  image_2_303 = _RAND_1455[3:0];
  _RAND_1456 = {1{`RANDOM}};
  image_2_304 = _RAND_1456[3:0];
  _RAND_1457 = {1{`RANDOM}};
  image_2_305 = _RAND_1457[3:0];
  _RAND_1458 = {1{`RANDOM}};
  image_2_306 = _RAND_1458[3:0];
  _RAND_1459 = {1{`RANDOM}};
  image_2_307 = _RAND_1459[3:0];
  _RAND_1460 = {1{`RANDOM}};
  image_2_308 = _RAND_1460[3:0];
  _RAND_1461 = {1{`RANDOM}};
  image_2_309 = _RAND_1461[3:0];
  _RAND_1462 = {1{`RANDOM}};
  image_2_310 = _RAND_1462[3:0];
  _RAND_1463 = {1{`RANDOM}};
  image_2_311 = _RAND_1463[3:0];
  _RAND_1464 = {1{`RANDOM}};
  image_2_312 = _RAND_1464[3:0];
  _RAND_1465 = {1{`RANDOM}};
  image_2_313 = _RAND_1465[3:0];
  _RAND_1466 = {1{`RANDOM}};
  image_2_314 = _RAND_1466[3:0];
  _RAND_1467 = {1{`RANDOM}};
  image_2_315 = _RAND_1467[3:0];
  _RAND_1468 = {1{`RANDOM}};
  image_2_316 = _RAND_1468[3:0];
  _RAND_1469 = {1{`RANDOM}};
  image_2_317 = _RAND_1469[3:0];
  _RAND_1470 = {1{`RANDOM}};
  image_2_318 = _RAND_1470[3:0];
  _RAND_1471 = {1{`RANDOM}};
  image_2_319 = _RAND_1471[3:0];
  _RAND_1472 = {1{`RANDOM}};
  image_2_320 = _RAND_1472[3:0];
  _RAND_1473 = {1{`RANDOM}};
  image_2_321 = _RAND_1473[3:0];
  _RAND_1474 = {1{`RANDOM}};
  image_2_322 = _RAND_1474[3:0];
  _RAND_1475 = {1{`RANDOM}};
  image_2_323 = _RAND_1475[3:0];
  _RAND_1476 = {1{`RANDOM}};
  image_2_324 = _RAND_1476[3:0];
  _RAND_1477 = {1{`RANDOM}};
  image_2_325 = _RAND_1477[3:0];
  _RAND_1478 = {1{`RANDOM}};
  image_2_326 = _RAND_1478[3:0];
  _RAND_1479 = {1{`RANDOM}};
  image_2_327 = _RAND_1479[3:0];
  _RAND_1480 = {1{`RANDOM}};
  image_2_328 = _RAND_1480[3:0];
  _RAND_1481 = {1{`RANDOM}};
  image_2_329 = _RAND_1481[3:0];
  _RAND_1482 = {1{`RANDOM}};
  image_2_330 = _RAND_1482[3:0];
  _RAND_1483 = {1{`RANDOM}};
  image_2_331 = _RAND_1483[3:0];
  _RAND_1484 = {1{`RANDOM}};
  image_2_332 = _RAND_1484[3:0];
  _RAND_1485 = {1{`RANDOM}};
  image_2_333 = _RAND_1485[3:0];
  _RAND_1486 = {1{`RANDOM}};
  image_2_334 = _RAND_1486[3:0];
  _RAND_1487 = {1{`RANDOM}};
  image_2_335 = _RAND_1487[3:0];
  _RAND_1488 = {1{`RANDOM}};
  image_2_336 = _RAND_1488[3:0];
  _RAND_1489 = {1{`RANDOM}};
  image_2_337 = _RAND_1489[3:0];
  _RAND_1490 = {1{`RANDOM}};
  image_2_338 = _RAND_1490[3:0];
  _RAND_1491 = {1{`RANDOM}};
  image_2_339 = _RAND_1491[3:0];
  _RAND_1492 = {1{`RANDOM}};
  image_2_340 = _RAND_1492[3:0];
  _RAND_1493 = {1{`RANDOM}};
  image_2_341 = _RAND_1493[3:0];
  _RAND_1494 = {1{`RANDOM}};
  image_2_342 = _RAND_1494[3:0];
  _RAND_1495 = {1{`RANDOM}};
  image_2_343 = _RAND_1495[3:0];
  _RAND_1496 = {1{`RANDOM}};
  image_2_344 = _RAND_1496[3:0];
  _RAND_1497 = {1{`RANDOM}};
  image_2_345 = _RAND_1497[3:0];
  _RAND_1498 = {1{`RANDOM}};
  image_2_346 = _RAND_1498[3:0];
  _RAND_1499 = {1{`RANDOM}};
  image_2_347 = _RAND_1499[3:0];
  _RAND_1500 = {1{`RANDOM}};
  image_2_348 = _RAND_1500[3:0];
  _RAND_1501 = {1{`RANDOM}};
  image_2_349 = _RAND_1501[3:0];
  _RAND_1502 = {1{`RANDOM}};
  image_2_350 = _RAND_1502[3:0];
  _RAND_1503 = {1{`RANDOM}};
  image_2_351 = _RAND_1503[3:0];
  _RAND_1504 = {1{`RANDOM}};
  image_2_352 = _RAND_1504[3:0];
  _RAND_1505 = {1{`RANDOM}};
  image_2_353 = _RAND_1505[3:0];
  _RAND_1506 = {1{`RANDOM}};
  image_2_354 = _RAND_1506[3:0];
  _RAND_1507 = {1{`RANDOM}};
  image_2_355 = _RAND_1507[3:0];
  _RAND_1508 = {1{`RANDOM}};
  image_2_356 = _RAND_1508[3:0];
  _RAND_1509 = {1{`RANDOM}};
  image_2_357 = _RAND_1509[3:0];
  _RAND_1510 = {1{`RANDOM}};
  image_2_358 = _RAND_1510[3:0];
  _RAND_1511 = {1{`RANDOM}};
  image_2_359 = _RAND_1511[3:0];
  _RAND_1512 = {1{`RANDOM}};
  image_2_360 = _RAND_1512[3:0];
  _RAND_1513 = {1{`RANDOM}};
  image_2_361 = _RAND_1513[3:0];
  _RAND_1514 = {1{`RANDOM}};
  image_2_362 = _RAND_1514[3:0];
  _RAND_1515 = {1{`RANDOM}};
  image_2_363 = _RAND_1515[3:0];
  _RAND_1516 = {1{`RANDOM}};
  image_2_364 = _RAND_1516[3:0];
  _RAND_1517 = {1{`RANDOM}};
  image_2_365 = _RAND_1517[3:0];
  _RAND_1518 = {1{`RANDOM}};
  image_2_366 = _RAND_1518[3:0];
  _RAND_1519 = {1{`RANDOM}};
  image_2_367 = _RAND_1519[3:0];
  _RAND_1520 = {1{`RANDOM}};
  image_2_368 = _RAND_1520[3:0];
  _RAND_1521 = {1{`RANDOM}};
  image_2_369 = _RAND_1521[3:0];
  _RAND_1522 = {1{`RANDOM}};
  image_2_370 = _RAND_1522[3:0];
  _RAND_1523 = {1{`RANDOM}};
  image_2_371 = _RAND_1523[3:0];
  _RAND_1524 = {1{`RANDOM}};
  image_2_372 = _RAND_1524[3:0];
  _RAND_1525 = {1{`RANDOM}};
  image_2_373 = _RAND_1525[3:0];
  _RAND_1526 = {1{`RANDOM}};
  image_2_374 = _RAND_1526[3:0];
  _RAND_1527 = {1{`RANDOM}};
  image_2_375 = _RAND_1527[3:0];
  _RAND_1528 = {1{`RANDOM}};
  image_2_376 = _RAND_1528[3:0];
  _RAND_1529 = {1{`RANDOM}};
  image_2_377 = _RAND_1529[3:0];
  _RAND_1530 = {1{`RANDOM}};
  image_2_378 = _RAND_1530[3:0];
  _RAND_1531 = {1{`RANDOM}};
  image_2_379 = _RAND_1531[3:0];
  _RAND_1532 = {1{`RANDOM}};
  image_2_380 = _RAND_1532[3:0];
  _RAND_1533 = {1{`RANDOM}};
  image_2_381 = _RAND_1533[3:0];
  _RAND_1534 = {1{`RANDOM}};
  image_2_382 = _RAND_1534[3:0];
  _RAND_1535 = {1{`RANDOM}};
  image_2_383 = _RAND_1535[3:0];
  _RAND_1536 = {1{`RANDOM}};
  image_2_384 = _RAND_1536[3:0];
  _RAND_1537 = {1{`RANDOM}};
  image_2_385 = _RAND_1537[3:0];
  _RAND_1538 = {1{`RANDOM}};
  image_2_386 = _RAND_1538[3:0];
  _RAND_1539 = {1{`RANDOM}};
  image_2_387 = _RAND_1539[3:0];
  _RAND_1540 = {1{`RANDOM}};
  image_2_388 = _RAND_1540[3:0];
  _RAND_1541 = {1{`RANDOM}};
  image_2_389 = _RAND_1541[3:0];
  _RAND_1542 = {1{`RANDOM}};
  image_2_390 = _RAND_1542[3:0];
  _RAND_1543 = {1{`RANDOM}};
  image_2_391 = _RAND_1543[3:0];
  _RAND_1544 = {1{`RANDOM}};
  image_2_392 = _RAND_1544[3:0];
  _RAND_1545 = {1{`RANDOM}};
  image_2_393 = _RAND_1545[3:0];
  _RAND_1546 = {1{`RANDOM}};
  image_2_394 = _RAND_1546[3:0];
  _RAND_1547 = {1{`RANDOM}};
  image_2_395 = _RAND_1547[3:0];
  _RAND_1548 = {1{`RANDOM}};
  image_2_396 = _RAND_1548[3:0];
  _RAND_1549 = {1{`RANDOM}};
  image_2_397 = _RAND_1549[3:0];
  _RAND_1550 = {1{`RANDOM}};
  image_2_398 = _RAND_1550[3:0];
  _RAND_1551 = {1{`RANDOM}};
  image_2_399 = _RAND_1551[3:0];
  _RAND_1552 = {1{`RANDOM}};
  image_2_400 = _RAND_1552[3:0];
  _RAND_1553 = {1{`RANDOM}};
  image_2_401 = _RAND_1553[3:0];
  _RAND_1554 = {1{`RANDOM}};
  image_2_402 = _RAND_1554[3:0];
  _RAND_1555 = {1{`RANDOM}};
  image_2_403 = _RAND_1555[3:0];
  _RAND_1556 = {1{`RANDOM}};
  image_2_404 = _RAND_1556[3:0];
  _RAND_1557 = {1{`RANDOM}};
  image_2_405 = _RAND_1557[3:0];
  _RAND_1558 = {1{`RANDOM}};
  image_2_406 = _RAND_1558[3:0];
  _RAND_1559 = {1{`RANDOM}};
  image_2_407 = _RAND_1559[3:0];
  _RAND_1560 = {1{`RANDOM}};
  image_2_408 = _RAND_1560[3:0];
  _RAND_1561 = {1{`RANDOM}};
  image_2_409 = _RAND_1561[3:0];
  _RAND_1562 = {1{`RANDOM}};
  image_2_410 = _RAND_1562[3:0];
  _RAND_1563 = {1{`RANDOM}};
  image_2_411 = _RAND_1563[3:0];
  _RAND_1564 = {1{`RANDOM}};
  image_2_412 = _RAND_1564[3:0];
  _RAND_1565 = {1{`RANDOM}};
  image_2_413 = _RAND_1565[3:0];
  _RAND_1566 = {1{`RANDOM}};
  image_2_414 = _RAND_1566[3:0];
  _RAND_1567 = {1{`RANDOM}};
  image_2_415 = _RAND_1567[3:0];
  _RAND_1568 = {1{`RANDOM}};
  image_2_416 = _RAND_1568[3:0];
  _RAND_1569 = {1{`RANDOM}};
  image_2_417 = _RAND_1569[3:0];
  _RAND_1570 = {1{`RANDOM}};
  image_2_418 = _RAND_1570[3:0];
  _RAND_1571 = {1{`RANDOM}};
  image_2_419 = _RAND_1571[3:0];
  _RAND_1572 = {1{`RANDOM}};
  image_2_420 = _RAND_1572[3:0];
  _RAND_1573 = {1{`RANDOM}};
  image_2_421 = _RAND_1573[3:0];
  _RAND_1574 = {1{`RANDOM}};
  image_2_422 = _RAND_1574[3:0];
  _RAND_1575 = {1{`RANDOM}};
  image_2_423 = _RAND_1575[3:0];
  _RAND_1576 = {1{`RANDOM}};
  image_2_424 = _RAND_1576[3:0];
  _RAND_1577 = {1{`RANDOM}};
  image_2_425 = _RAND_1577[3:0];
  _RAND_1578 = {1{`RANDOM}};
  image_2_426 = _RAND_1578[3:0];
  _RAND_1579 = {1{`RANDOM}};
  image_2_427 = _RAND_1579[3:0];
  _RAND_1580 = {1{`RANDOM}};
  image_2_428 = _RAND_1580[3:0];
  _RAND_1581 = {1{`RANDOM}};
  image_2_429 = _RAND_1581[3:0];
  _RAND_1582 = {1{`RANDOM}};
  image_2_430 = _RAND_1582[3:0];
  _RAND_1583 = {1{`RANDOM}};
  image_2_431 = _RAND_1583[3:0];
  _RAND_1584 = {1{`RANDOM}};
  image_2_432 = _RAND_1584[3:0];
  _RAND_1585 = {1{`RANDOM}};
  image_2_433 = _RAND_1585[3:0];
  _RAND_1586 = {1{`RANDOM}};
  image_2_434 = _RAND_1586[3:0];
  _RAND_1587 = {1{`RANDOM}};
  image_2_435 = _RAND_1587[3:0];
  _RAND_1588 = {1{`RANDOM}};
  image_2_436 = _RAND_1588[3:0];
  _RAND_1589 = {1{`RANDOM}};
  image_2_437 = _RAND_1589[3:0];
  _RAND_1590 = {1{`RANDOM}};
  image_2_438 = _RAND_1590[3:0];
  _RAND_1591 = {1{`RANDOM}};
  image_2_439 = _RAND_1591[3:0];
  _RAND_1592 = {1{`RANDOM}};
  image_2_440 = _RAND_1592[3:0];
  _RAND_1593 = {1{`RANDOM}};
  image_2_441 = _RAND_1593[3:0];
  _RAND_1594 = {1{`RANDOM}};
  image_2_442 = _RAND_1594[3:0];
  _RAND_1595 = {1{`RANDOM}};
  image_2_443 = _RAND_1595[3:0];
  _RAND_1596 = {1{`RANDOM}};
  image_2_444 = _RAND_1596[3:0];
  _RAND_1597 = {1{`RANDOM}};
  image_2_445 = _RAND_1597[3:0];
  _RAND_1598 = {1{`RANDOM}};
  image_2_446 = _RAND_1598[3:0];
  _RAND_1599 = {1{`RANDOM}};
  image_2_447 = _RAND_1599[3:0];
  _RAND_1600 = {1{`RANDOM}};
  image_2_448 = _RAND_1600[3:0];
  _RAND_1601 = {1{`RANDOM}};
  image_2_449 = _RAND_1601[3:0];
  _RAND_1602 = {1{`RANDOM}};
  image_2_450 = _RAND_1602[3:0];
  _RAND_1603 = {1{`RANDOM}};
  image_2_451 = _RAND_1603[3:0];
  _RAND_1604 = {1{`RANDOM}};
  image_2_452 = _RAND_1604[3:0];
  _RAND_1605 = {1{`RANDOM}};
  image_2_453 = _RAND_1605[3:0];
  _RAND_1606 = {1{`RANDOM}};
  image_2_454 = _RAND_1606[3:0];
  _RAND_1607 = {1{`RANDOM}};
  image_2_455 = _RAND_1607[3:0];
  _RAND_1608 = {1{`RANDOM}};
  image_2_456 = _RAND_1608[3:0];
  _RAND_1609 = {1{`RANDOM}};
  image_2_457 = _RAND_1609[3:0];
  _RAND_1610 = {1{`RANDOM}};
  image_2_458 = _RAND_1610[3:0];
  _RAND_1611 = {1{`RANDOM}};
  image_2_459 = _RAND_1611[3:0];
  _RAND_1612 = {1{`RANDOM}};
  image_2_460 = _RAND_1612[3:0];
  _RAND_1613 = {1{`RANDOM}};
  image_2_461 = _RAND_1613[3:0];
  _RAND_1614 = {1{`RANDOM}};
  image_2_462 = _RAND_1614[3:0];
  _RAND_1615 = {1{`RANDOM}};
  image_2_463 = _RAND_1615[3:0];
  _RAND_1616 = {1{`RANDOM}};
  image_2_464 = _RAND_1616[3:0];
  _RAND_1617 = {1{`RANDOM}};
  image_2_465 = _RAND_1617[3:0];
  _RAND_1618 = {1{`RANDOM}};
  image_2_466 = _RAND_1618[3:0];
  _RAND_1619 = {1{`RANDOM}};
  image_2_467 = _RAND_1619[3:0];
  _RAND_1620 = {1{`RANDOM}};
  image_2_468 = _RAND_1620[3:0];
  _RAND_1621 = {1{`RANDOM}};
  image_2_469 = _RAND_1621[3:0];
  _RAND_1622 = {1{`RANDOM}};
  image_2_470 = _RAND_1622[3:0];
  _RAND_1623 = {1{`RANDOM}};
  image_2_471 = _RAND_1623[3:0];
  _RAND_1624 = {1{`RANDOM}};
  image_2_472 = _RAND_1624[3:0];
  _RAND_1625 = {1{`RANDOM}};
  image_2_473 = _RAND_1625[3:0];
  _RAND_1626 = {1{`RANDOM}};
  image_2_474 = _RAND_1626[3:0];
  _RAND_1627 = {1{`RANDOM}};
  image_2_475 = _RAND_1627[3:0];
  _RAND_1628 = {1{`RANDOM}};
  image_2_476 = _RAND_1628[3:0];
  _RAND_1629 = {1{`RANDOM}};
  image_2_477 = _RAND_1629[3:0];
  _RAND_1630 = {1{`RANDOM}};
  image_2_478 = _RAND_1630[3:0];
  _RAND_1631 = {1{`RANDOM}};
  image_2_479 = _RAND_1631[3:0];
  _RAND_1632 = {1{`RANDOM}};
  image_2_480 = _RAND_1632[3:0];
  _RAND_1633 = {1{`RANDOM}};
  image_2_481 = _RAND_1633[3:0];
  _RAND_1634 = {1{`RANDOM}};
  image_2_482 = _RAND_1634[3:0];
  _RAND_1635 = {1{`RANDOM}};
  image_2_483 = _RAND_1635[3:0];
  _RAND_1636 = {1{`RANDOM}};
  image_2_484 = _RAND_1636[3:0];
  _RAND_1637 = {1{`RANDOM}};
  image_2_485 = _RAND_1637[3:0];
  _RAND_1638 = {1{`RANDOM}};
  image_2_486 = _RAND_1638[3:0];
  _RAND_1639 = {1{`RANDOM}};
  image_2_487 = _RAND_1639[3:0];
  _RAND_1640 = {1{`RANDOM}};
  image_2_488 = _RAND_1640[3:0];
  _RAND_1641 = {1{`RANDOM}};
  image_2_489 = _RAND_1641[3:0];
  _RAND_1642 = {1{`RANDOM}};
  image_2_490 = _RAND_1642[3:0];
  _RAND_1643 = {1{`RANDOM}};
  image_2_491 = _RAND_1643[3:0];
  _RAND_1644 = {1{`RANDOM}};
  image_2_492 = _RAND_1644[3:0];
  _RAND_1645 = {1{`RANDOM}};
  image_2_493 = _RAND_1645[3:0];
  _RAND_1646 = {1{`RANDOM}};
  image_2_494 = _RAND_1646[3:0];
  _RAND_1647 = {1{`RANDOM}};
  image_2_495 = _RAND_1647[3:0];
  _RAND_1648 = {1{`RANDOM}};
  image_2_496 = _RAND_1648[3:0];
  _RAND_1649 = {1{`RANDOM}};
  image_2_497 = _RAND_1649[3:0];
  _RAND_1650 = {1{`RANDOM}};
  image_2_498 = _RAND_1650[3:0];
  _RAND_1651 = {1{`RANDOM}};
  image_2_499 = _RAND_1651[3:0];
  _RAND_1652 = {1{`RANDOM}};
  image_2_500 = _RAND_1652[3:0];
  _RAND_1653 = {1{`RANDOM}};
  image_2_501 = _RAND_1653[3:0];
  _RAND_1654 = {1{`RANDOM}};
  image_2_502 = _RAND_1654[3:0];
  _RAND_1655 = {1{`RANDOM}};
  image_2_503 = _RAND_1655[3:0];
  _RAND_1656 = {1{`RANDOM}};
  image_2_504 = _RAND_1656[3:0];
  _RAND_1657 = {1{`RANDOM}};
  image_2_505 = _RAND_1657[3:0];
  _RAND_1658 = {1{`RANDOM}};
  image_2_506 = _RAND_1658[3:0];
  _RAND_1659 = {1{`RANDOM}};
  image_2_507 = _RAND_1659[3:0];
  _RAND_1660 = {1{`RANDOM}};
  image_2_508 = _RAND_1660[3:0];
  _RAND_1661 = {1{`RANDOM}};
  image_2_509 = _RAND_1661[3:0];
  _RAND_1662 = {1{`RANDOM}};
  image_2_510 = _RAND_1662[3:0];
  _RAND_1663 = {1{`RANDOM}};
  image_2_511 = _RAND_1663[3:0];
  _RAND_1664 = {1{`RANDOM}};
  image_2_512 = _RAND_1664[3:0];
  _RAND_1665 = {1{`RANDOM}};
  image_2_513 = _RAND_1665[3:0];
  _RAND_1666 = {1{`RANDOM}};
  image_2_514 = _RAND_1666[3:0];
  _RAND_1667 = {1{`RANDOM}};
  image_2_515 = _RAND_1667[3:0];
  _RAND_1668 = {1{`RANDOM}};
  image_2_516 = _RAND_1668[3:0];
  _RAND_1669 = {1{`RANDOM}};
  image_2_517 = _RAND_1669[3:0];
  _RAND_1670 = {1{`RANDOM}};
  image_2_518 = _RAND_1670[3:0];
  _RAND_1671 = {1{`RANDOM}};
  image_2_519 = _RAND_1671[3:0];
  _RAND_1672 = {1{`RANDOM}};
  image_2_520 = _RAND_1672[3:0];
  _RAND_1673 = {1{`RANDOM}};
  image_2_521 = _RAND_1673[3:0];
  _RAND_1674 = {1{`RANDOM}};
  image_2_522 = _RAND_1674[3:0];
  _RAND_1675 = {1{`RANDOM}};
  image_2_523 = _RAND_1675[3:0];
  _RAND_1676 = {1{`RANDOM}};
  image_2_524 = _RAND_1676[3:0];
  _RAND_1677 = {1{`RANDOM}};
  image_2_525 = _RAND_1677[3:0];
  _RAND_1678 = {1{`RANDOM}};
  image_2_526 = _RAND_1678[3:0];
  _RAND_1679 = {1{`RANDOM}};
  image_2_527 = _RAND_1679[3:0];
  _RAND_1680 = {1{`RANDOM}};
  image_2_528 = _RAND_1680[3:0];
  _RAND_1681 = {1{`RANDOM}};
  image_2_529 = _RAND_1681[3:0];
  _RAND_1682 = {1{`RANDOM}};
  image_2_530 = _RAND_1682[3:0];
  _RAND_1683 = {1{`RANDOM}};
  image_2_531 = _RAND_1683[3:0];
  _RAND_1684 = {1{`RANDOM}};
  image_2_532 = _RAND_1684[3:0];
  _RAND_1685 = {1{`RANDOM}};
  image_2_533 = _RAND_1685[3:0];
  _RAND_1686 = {1{`RANDOM}};
  image_2_534 = _RAND_1686[3:0];
  _RAND_1687 = {1{`RANDOM}};
  image_2_535 = _RAND_1687[3:0];
  _RAND_1688 = {1{`RANDOM}};
  image_2_536 = _RAND_1688[3:0];
  _RAND_1689 = {1{`RANDOM}};
  image_2_537 = _RAND_1689[3:0];
  _RAND_1690 = {1{`RANDOM}};
  image_2_538 = _RAND_1690[3:0];
  _RAND_1691 = {1{`RANDOM}};
  image_2_539 = _RAND_1691[3:0];
  _RAND_1692 = {1{`RANDOM}};
  image_2_540 = _RAND_1692[3:0];
  _RAND_1693 = {1{`RANDOM}};
  image_2_541 = _RAND_1693[3:0];
  _RAND_1694 = {1{`RANDOM}};
  image_2_542 = _RAND_1694[3:0];
  _RAND_1695 = {1{`RANDOM}};
  image_2_543 = _RAND_1695[3:0];
  _RAND_1696 = {1{`RANDOM}};
  image_2_544 = _RAND_1696[3:0];
  _RAND_1697 = {1{`RANDOM}};
  image_2_545 = _RAND_1697[3:0];
  _RAND_1698 = {1{`RANDOM}};
  image_2_546 = _RAND_1698[3:0];
  _RAND_1699 = {1{`RANDOM}};
  image_2_547 = _RAND_1699[3:0];
  _RAND_1700 = {1{`RANDOM}};
  image_2_548 = _RAND_1700[3:0];
  _RAND_1701 = {1{`RANDOM}};
  image_2_549 = _RAND_1701[3:0];
  _RAND_1702 = {1{`RANDOM}};
  image_2_550 = _RAND_1702[3:0];
  _RAND_1703 = {1{`RANDOM}};
  image_2_551 = _RAND_1703[3:0];
  _RAND_1704 = {1{`RANDOM}};
  image_2_552 = _RAND_1704[3:0];
  _RAND_1705 = {1{`RANDOM}};
  image_2_553 = _RAND_1705[3:0];
  _RAND_1706 = {1{`RANDOM}};
  image_2_554 = _RAND_1706[3:0];
  _RAND_1707 = {1{`RANDOM}};
  image_2_555 = _RAND_1707[3:0];
  _RAND_1708 = {1{`RANDOM}};
  image_2_556 = _RAND_1708[3:0];
  _RAND_1709 = {1{`RANDOM}};
  image_2_557 = _RAND_1709[3:0];
  _RAND_1710 = {1{`RANDOM}};
  image_2_558 = _RAND_1710[3:0];
  _RAND_1711 = {1{`RANDOM}};
  image_2_559 = _RAND_1711[3:0];
  _RAND_1712 = {1{`RANDOM}};
  image_2_560 = _RAND_1712[3:0];
  _RAND_1713 = {1{`RANDOM}};
  image_2_561 = _RAND_1713[3:0];
  _RAND_1714 = {1{`RANDOM}};
  image_2_562 = _RAND_1714[3:0];
  _RAND_1715 = {1{`RANDOM}};
  image_2_563 = _RAND_1715[3:0];
  _RAND_1716 = {1{`RANDOM}};
  image_2_564 = _RAND_1716[3:0];
  _RAND_1717 = {1{`RANDOM}};
  image_2_565 = _RAND_1717[3:0];
  _RAND_1718 = {1{`RANDOM}};
  image_2_566 = _RAND_1718[3:0];
  _RAND_1719 = {1{`RANDOM}};
  image_2_567 = _RAND_1719[3:0];
  _RAND_1720 = {1{`RANDOM}};
  image_2_568 = _RAND_1720[3:0];
  _RAND_1721 = {1{`RANDOM}};
  image_2_569 = _RAND_1721[3:0];
  _RAND_1722 = {1{`RANDOM}};
  image_2_570 = _RAND_1722[3:0];
  _RAND_1723 = {1{`RANDOM}};
  image_2_571 = _RAND_1723[3:0];
  _RAND_1724 = {1{`RANDOM}};
  image_2_572 = _RAND_1724[3:0];
  _RAND_1725 = {1{`RANDOM}};
  image_2_573 = _RAND_1725[3:0];
  _RAND_1726 = {1{`RANDOM}};
  image_2_574 = _RAND_1726[3:0];
  _RAND_1727 = {1{`RANDOM}};
  image_2_575 = _RAND_1727[3:0];
  _RAND_1728 = {1{`RANDOM}};
  pixelIndex = _RAND_1728[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      image_0_0 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h0 == _T_37[9:0]) begin
        image_0_0 <= io_pixelVal_in_0_7;
      end else if (10'h0 == _T_34[9:0]) begin
        image_0_0 <= io_pixelVal_in_0_6;
      end else if (10'h0 == _T_31[9:0]) begin
        image_0_0 <= io_pixelVal_in_0_5;
      end else if (10'h0 == _T_28[9:0]) begin
        image_0_0 <= io_pixelVal_in_0_4;
      end else if (10'h0 == _T_25[9:0]) begin
        image_0_0 <= io_pixelVal_in_0_3;
      end else if (10'h0 == _T_22[9:0]) begin
        image_0_0 <= io_pixelVal_in_0_2;
      end else if (10'h0 == _T_19[9:0]) begin
        image_0_0 <= io_pixelVal_in_0_1;
      end else if (10'h0 == _T_15[9:0]) begin
        image_0_0 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_1 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1 == _T_37[9:0]) begin
        image_0_1 <= io_pixelVal_in_0_7;
      end else if (10'h1 == _T_34[9:0]) begin
        image_0_1 <= io_pixelVal_in_0_6;
      end else if (10'h1 == _T_31[9:0]) begin
        image_0_1 <= io_pixelVal_in_0_5;
      end else if (10'h1 == _T_28[9:0]) begin
        image_0_1 <= io_pixelVal_in_0_4;
      end else if (10'h1 == _T_25[9:0]) begin
        image_0_1 <= io_pixelVal_in_0_3;
      end else if (10'h1 == _T_22[9:0]) begin
        image_0_1 <= io_pixelVal_in_0_2;
      end else if (10'h1 == _T_19[9:0]) begin
        image_0_1 <= io_pixelVal_in_0_1;
      end else if (10'h1 == _T_15[9:0]) begin
        image_0_1 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_2 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h2 == _T_37[9:0]) begin
        image_0_2 <= io_pixelVal_in_0_7;
      end else if (10'h2 == _T_34[9:0]) begin
        image_0_2 <= io_pixelVal_in_0_6;
      end else if (10'h2 == _T_31[9:0]) begin
        image_0_2 <= io_pixelVal_in_0_5;
      end else if (10'h2 == _T_28[9:0]) begin
        image_0_2 <= io_pixelVal_in_0_4;
      end else if (10'h2 == _T_25[9:0]) begin
        image_0_2 <= io_pixelVal_in_0_3;
      end else if (10'h2 == _T_22[9:0]) begin
        image_0_2 <= io_pixelVal_in_0_2;
      end else if (10'h2 == _T_19[9:0]) begin
        image_0_2 <= io_pixelVal_in_0_1;
      end else if (10'h2 == _T_15[9:0]) begin
        image_0_2 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_3 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h3 == _T_37[9:0]) begin
        image_0_3 <= io_pixelVal_in_0_7;
      end else if (10'h3 == _T_34[9:0]) begin
        image_0_3 <= io_pixelVal_in_0_6;
      end else if (10'h3 == _T_31[9:0]) begin
        image_0_3 <= io_pixelVal_in_0_5;
      end else if (10'h3 == _T_28[9:0]) begin
        image_0_3 <= io_pixelVal_in_0_4;
      end else if (10'h3 == _T_25[9:0]) begin
        image_0_3 <= io_pixelVal_in_0_3;
      end else if (10'h3 == _T_22[9:0]) begin
        image_0_3 <= io_pixelVal_in_0_2;
      end else if (10'h3 == _T_19[9:0]) begin
        image_0_3 <= io_pixelVal_in_0_1;
      end else if (10'h3 == _T_15[9:0]) begin
        image_0_3 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_4 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h4 == _T_37[9:0]) begin
        image_0_4 <= io_pixelVal_in_0_7;
      end else if (10'h4 == _T_34[9:0]) begin
        image_0_4 <= io_pixelVal_in_0_6;
      end else if (10'h4 == _T_31[9:0]) begin
        image_0_4 <= io_pixelVal_in_0_5;
      end else if (10'h4 == _T_28[9:0]) begin
        image_0_4 <= io_pixelVal_in_0_4;
      end else if (10'h4 == _T_25[9:0]) begin
        image_0_4 <= io_pixelVal_in_0_3;
      end else if (10'h4 == _T_22[9:0]) begin
        image_0_4 <= io_pixelVal_in_0_2;
      end else if (10'h4 == _T_19[9:0]) begin
        image_0_4 <= io_pixelVal_in_0_1;
      end else if (10'h4 == _T_15[9:0]) begin
        image_0_4 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_5 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h5 == _T_37[9:0]) begin
        image_0_5 <= io_pixelVal_in_0_7;
      end else if (10'h5 == _T_34[9:0]) begin
        image_0_5 <= io_pixelVal_in_0_6;
      end else if (10'h5 == _T_31[9:0]) begin
        image_0_5 <= io_pixelVal_in_0_5;
      end else if (10'h5 == _T_28[9:0]) begin
        image_0_5 <= io_pixelVal_in_0_4;
      end else if (10'h5 == _T_25[9:0]) begin
        image_0_5 <= io_pixelVal_in_0_3;
      end else if (10'h5 == _T_22[9:0]) begin
        image_0_5 <= io_pixelVal_in_0_2;
      end else if (10'h5 == _T_19[9:0]) begin
        image_0_5 <= io_pixelVal_in_0_1;
      end else if (10'h5 == _T_15[9:0]) begin
        image_0_5 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_6 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h6 == _T_37[9:0]) begin
        image_0_6 <= io_pixelVal_in_0_7;
      end else if (10'h6 == _T_34[9:0]) begin
        image_0_6 <= io_pixelVal_in_0_6;
      end else if (10'h6 == _T_31[9:0]) begin
        image_0_6 <= io_pixelVal_in_0_5;
      end else if (10'h6 == _T_28[9:0]) begin
        image_0_6 <= io_pixelVal_in_0_4;
      end else if (10'h6 == _T_25[9:0]) begin
        image_0_6 <= io_pixelVal_in_0_3;
      end else if (10'h6 == _T_22[9:0]) begin
        image_0_6 <= io_pixelVal_in_0_2;
      end else if (10'h6 == _T_19[9:0]) begin
        image_0_6 <= io_pixelVal_in_0_1;
      end else if (10'h6 == _T_15[9:0]) begin
        image_0_6 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_7 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h7 == _T_37[9:0]) begin
        image_0_7 <= io_pixelVal_in_0_7;
      end else if (10'h7 == _T_34[9:0]) begin
        image_0_7 <= io_pixelVal_in_0_6;
      end else if (10'h7 == _T_31[9:0]) begin
        image_0_7 <= io_pixelVal_in_0_5;
      end else if (10'h7 == _T_28[9:0]) begin
        image_0_7 <= io_pixelVal_in_0_4;
      end else if (10'h7 == _T_25[9:0]) begin
        image_0_7 <= io_pixelVal_in_0_3;
      end else if (10'h7 == _T_22[9:0]) begin
        image_0_7 <= io_pixelVal_in_0_2;
      end else if (10'h7 == _T_19[9:0]) begin
        image_0_7 <= io_pixelVal_in_0_1;
      end else if (10'h7 == _T_15[9:0]) begin
        image_0_7 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_8 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h8 == _T_37[9:0]) begin
        image_0_8 <= io_pixelVal_in_0_7;
      end else if (10'h8 == _T_34[9:0]) begin
        image_0_8 <= io_pixelVal_in_0_6;
      end else if (10'h8 == _T_31[9:0]) begin
        image_0_8 <= io_pixelVal_in_0_5;
      end else if (10'h8 == _T_28[9:0]) begin
        image_0_8 <= io_pixelVal_in_0_4;
      end else if (10'h8 == _T_25[9:0]) begin
        image_0_8 <= io_pixelVal_in_0_3;
      end else if (10'h8 == _T_22[9:0]) begin
        image_0_8 <= io_pixelVal_in_0_2;
      end else if (10'h8 == _T_19[9:0]) begin
        image_0_8 <= io_pixelVal_in_0_1;
      end else if (10'h8 == _T_15[9:0]) begin
        image_0_8 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_9 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h9 == _T_37[9:0]) begin
        image_0_9 <= io_pixelVal_in_0_7;
      end else if (10'h9 == _T_34[9:0]) begin
        image_0_9 <= io_pixelVal_in_0_6;
      end else if (10'h9 == _T_31[9:0]) begin
        image_0_9 <= io_pixelVal_in_0_5;
      end else if (10'h9 == _T_28[9:0]) begin
        image_0_9 <= io_pixelVal_in_0_4;
      end else if (10'h9 == _T_25[9:0]) begin
        image_0_9 <= io_pixelVal_in_0_3;
      end else if (10'h9 == _T_22[9:0]) begin
        image_0_9 <= io_pixelVal_in_0_2;
      end else if (10'h9 == _T_19[9:0]) begin
        image_0_9 <= io_pixelVal_in_0_1;
      end else if (10'h9 == _T_15[9:0]) begin
        image_0_9 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_10 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'ha == _T_37[9:0]) begin
        image_0_10 <= io_pixelVal_in_0_7;
      end else if (10'ha == _T_34[9:0]) begin
        image_0_10 <= io_pixelVal_in_0_6;
      end else if (10'ha == _T_31[9:0]) begin
        image_0_10 <= io_pixelVal_in_0_5;
      end else if (10'ha == _T_28[9:0]) begin
        image_0_10 <= io_pixelVal_in_0_4;
      end else if (10'ha == _T_25[9:0]) begin
        image_0_10 <= io_pixelVal_in_0_3;
      end else if (10'ha == _T_22[9:0]) begin
        image_0_10 <= io_pixelVal_in_0_2;
      end else if (10'ha == _T_19[9:0]) begin
        image_0_10 <= io_pixelVal_in_0_1;
      end else if (10'ha == _T_15[9:0]) begin
        image_0_10 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_11 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hb == _T_37[9:0]) begin
        image_0_11 <= io_pixelVal_in_0_7;
      end else if (10'hb == _T_34[9:0]) begin
        image_0_11 <= io_pixelVal_in_0_6;
      end else if (10'hb == _T_31[9:0]) begin
        image_0_11 <= io_pixelVal_in_0_5;
      end else if (10'hb == _T_28[9:0]) begin
        image_0_11 <= io_pixelVal_in_0_4;
      end else if (10'hb == _T_25[9:0]) begin
        image_0_11 <= io_pixelVal_in_0_3;
      end else if (10'hb == _T_22[9:0]) begin
        image_0_11 <= io_pixelVal_in_0_2;
      end else if (10'hb == _T_19[9:0]) begin
        image_0_11 <= io_pixelVal_in_0_1;
      end else if (10'hb == _T_15[9:0]) begin
        image_0_11 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_12 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hc == _T_37[9:0]) begin
        image_0_12 <= io_pixelVal_in_0_7;
      end else if (10'hc == _T_34[9:0]) begin
        image_0_12 <= io_pixelVal_in_0_6;
      end else if (10'hc == _T_31[9:0]) begin
        image_0_12 <= io_pixelVal_in_0_5;
      end else if (10'hc == _T_28[9:0]) begin
        image_0_12 <= io_pixelVal_in_0_4;
      end else if (10'hc == _T_25[9:0]) begin
        image_0_12 <= io_pixelVal_in_0_3;
      end else if (10'hc == _T_22[9:0]) begin
        image_0_12 <= io_pixelVal_in_0_2;
      end else if (10'hc == _T_19[9:0]) begin
        image_0_12 <= io_pixelVal_in_0_1;
      end else if (10'hc == _T_15[9:0]) begin
        image_0_12 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_13 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hd == _T_37[9:0]) begin
        image_0_13 <= io_pixelVal_in_0_7;
      end else if (10'hd == _T_34[9:0]) begin
        image_0_13 <= io_pixelVal_in_0_6;
      end else if (10'hd == _T_31[9:0]) begin
        image_0_13 <= io_pixelVal_in_0_5;
      end else if (10'hd == _T_28[9:0]) begin
        image_0_13 <= io_pixelVal_in_0_4;
      end else if (10'hd == _T_25[9:0]) begin
        image_0_13 <= io_pixelVal_in_0_3;
      end else if (10'hd == _T_22[9:0]) begin
        image_0_13 <= io_pixelVal_in_0_2;
      end else if (10'hd == _T_19[9:0]) begin
        image_0_13 <= io_pixelVal_in_0_1;
      end else if (10'hd == _T_15[9:0]) begin
        image_0_13 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_14 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'he == _T_37[9:0]) begin
        image_0_14 <= io_pixelVal_in_0_7;
      end else if (10'he == _T_34[9:0]) begin
        image_0_14 <= io_pixelVal_in_0_6;
      end else if (10'he == _T_31[9:0]) begin
        image_0_14 <= io_pixelVal_in_0_5;
      end else if (10'he == _T_28[9:0]) begin
        image_0_14 <= io_pixelVal_in_0_4;
      end else if (10'he == _T_25[9:0]) begin
        image_0_14 <= io_pixelVal_in_0_3;
      end else if (10'he == _T_22[9:0]) begin
        image_0_14 <= io_pixelVal_in_0_2;
      end else if (10'he == _T_19[9:0]) begin
        image_0_14 <= io_pixelVal_in_0_1;
      end else if (10'he == _T_15[9:0]) begin
        image_0_14 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_15 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hf == _T_37[9:0]) begin
        image_0_15 <= io_pixelVal_in_0_7;
      end else if (10'hf == _T_34[9:0]) begin
        image_0_15 <= io_pixelVal_in_0_6;
      end else if (10'hf == _T_31[9:0]) begin
        image_0_15 <= io_pixelVal_in_0_5;
      end else if (10'hf == _T_28[9:0]) begin
        image_0_15 <= io_pixelVal_in_0_4;
      end else if (10'hf == _T_25[9:0]) begin
        image_0_15 <= io_pixelVal_in_0_3;
      end else if (10'hf == _T_22[9:0]) begin
        image_0_15 <= io_pixelVal_in_0_2;
      end else if (10'hf == _T_19[9:0]) begin
        image_0_15 <= io_pixelVal_in_0_1;
      end else if (10'hf == _T_15[9:0]) begin
        image_0_15 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_16 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h10 == _T_37[9:0]) begin
        image_0_16 <= io_pixelVal_in_0_7;
      end else if (10'h10 == _T_34[9:0]) begin
        image_0_16 <= io_pixelVal_in_0_6;
      end else if (10'h10 == _T_31[9:0]) begin
        image_0_16 <= io_pixelVal_in_0_5;
      end else if (10'h10 == _T_28[9:0]) begin
        image_0_16 <= io_pixelVal_in_0_4;
      end else if (10'h10 == _T_25[9:0]) begin
        image_0_16 <= io_pixelVal_in_0_3;
      end else if (10'h10 == _T_22[9:0]) begin
        image_0_16 <= io_pixelVal_in_0_2;
      end else if (10'h10 == _T_19[9:0]) begin
        image_0_16 <= io_pixelVal_in_0_1;
      end else if (10'h10 == _T_15[9:0]) begin
        image_0_16 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_17 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h11 == _T_37[9:0]) begin
        image_0_17 <= io_pixelVal_in_0_7;
      end else if (10'h11 == _T_34[9:0]) begin
        image_0_17 <= io_pixelVal_in_0_6;
      end else if (10'h11 == _T_31[9:0]) begin
        image_0_17 <= io_pixelVal_in_0_5;
      end else if (10'h11 == _T_28[9:0]) begin
        image_0_17 <= io_pixelVal_in_0_4;
      end else if (10'h11 == _T_25[9:0]) begin
        image_0_17 <= io_pixelVal_in_0_3;
      end else if (10'h11 == _T_22[9:0]) begin
        image_0_17 <= io_pixelVal_in_0_2;
      end else if (10'h11 == _T_19[9:0]) begin
        image_0_17 <= io_pixelVal_in_0_1;
      end else if (10'h11 == _T_15[9:0]) begin
        image_0_17 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_18 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h12 == _T_37[9:0]) begin
        image_0_18 <= io_pixelVal_in_0_7;
      end else if (10'h12 == _T_34[9:0]) begin
        image_0_18 <= io_pixelVal_in_0_6;
      end else if (10'h12 == _T_31[9:0]) begin
        image_0_18 <= io_pixelVal_in_0_5;
      end else if (10'h12 == _T_28[9:0]) begin
        image_0_18 <= io_pixelVal_in_0_4;
      end else if (10'h12 == _T_25[9:0]) begin
        image_0_18 <= io_pixelVal_in_0_3;
      end else if (10'h12 == _T_22[9:0]) begin
        image_0_18 <= io_pixelVal_in_0_2;
      end else if (10'h12 == _T_19[9:0]) begin
        image_0_18 <= io_pixelVal_in_0_1;
      end else if (10'h12 == _T_15[9:0]) begin
        image_0_18 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_19 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h13 == _T_37[9:0]) begin
        image_0_19 <= io_pixelVal_in_0_7;
      end else if (10'h13 == _T_34[9:0]) begin
        image_0_19 <= io_pixelVal_in_0_6;
      end else if (10'h13 == _T_31[9:0]) begin
        image_0_19 <= io_pixelVal_in_0_5;
      end else if (10'h13 == _T_28[9:0]) begin
        image_0_19 <= io_pixelVal_in_0_4;
      end else if (10'h13 == _T_25[9:0]) begin
        image_0_19 <= io_pixelVal_in_0_3;
      end else if (10'h13 == _T_22[9:0]) begin
        image_0_19 <= io_pixelVal_in_0_2;
      end else if (10'h13 == _T_19[9:0]) begin
        image_0_19 <= io_pixelVal_in_0_1;
      end else if (10'h13 == _T_15[9:0]) begin
        image_0_19 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_20 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h14 == _T_37[9:0]) begin
        image_0_20 <= io_pixelVal_in_0_7;
      end else if (10'h14 == _T_34[9:0]) begin
        image_0_20 <= io_pixelVal_in_0_6;
      end else if (10'h14 == _T_31[9:0]) begin
        image_0_20 <= io_pixelVal_in_0_5;
      end else if (10'h14 == _T_28[9:0]) begin
        image_0_20 <= io_pixelVal_in_0_4;
      end else if (10'h14 == _T_25[9:0]) begin
        image_0_20 <= io_pixelVal_in_0_3;
      end else if (10'h14 == _T_22[9:0]) begin
        image_0_20 <= io_pixelVal_in_0_2;
      end else if (10'h14 == _T_19[9:0]) begin
        image_0_20 <= io_pixelVal_in_0_1;
      end else if (10'h14 == _T_15[9:0]) begin
        image_0_20 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_21 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h15 == _T_37[9:0]) begin
        image_0_21 <= io_pixelVal_in_0_7;
      end else if (10'h15 == _T_34[9:0]) begin
        image_0_21 <= io_pixelVal_in_0_6;
      end else if (10'h15 == _T_31[9:0]) begin
        image_0_21 <= io_pixelVal_in_0_5;
      end else if (10'h15 == _T_28[9:0]) begin
        image_0_21 <= io_pixelVal_in_0_4;
      end else if (10'h15 == _T_25[9:0]) begin
        image_0_21 <= io_pixelVal_in_0_3;
      end else if (10'h15 == _T_22[9:0]) begin
        image_0_21 <= io_pixelVal_in_0_2;
      end else if (10'h15 == _T_19[9:0]) begin
        image_0_21 <= io_pixelVal_in_0_1;
      end else if (10'h15 == _T_15[9:0]) begin
        image_0_21 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_22 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h16 == _T_37[9:0]) begin
        image_0_22 <= io_pixelVal_in_0_7;
      end else if (10'h16 == _T_34[9:0]) begin
        image_0_22 <= io_pixelVal_in_0_6;
      end else if (10'h16 == _T_31[9:0]) begin
        image_0_22 <= io_pixelVal_in_0_5;
      end else if (10'h16 == _T_28[9:0]) begin
        image_0_22 <= io_pixelVal_in_0_4;
      end else if (10'h16 == _T_25[9:0]) begin
        image_0_22 <= io_pixelVal_in_0_3;
      end else if (10'h16 == _T_22[9:0]) begin
        image_0_22 <= io_pixelVal_in_0_2;
      end else if (10'h16 == _T_19[9:0]) begin
        image_0_22 <= io_pixelVal_in_0_1;
      end else if (10'h16 == _T_15[9:0]) begin
        image_0_22 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_23 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h17 == _T_37[9:0]) begin
        image_0_23 <= io_pixelVal_in_0_7;
      end else if (10'h17 == _T_34[9:0]) begin
        image_0_23 <= io_pixelVal_in_0_6;
      end else if (10'h17 == _T_31[9:0]) begin
        image_0_23 <= io_pixelVal_in_0_5;
      end else if (10'h17 == _T_28[9:0]) begin
        image_0_23 <= io_pixelVal_in_0_4;
      end else if (10'h17 == _T_25[9:0]) begin
        image_0_23 <= io_pixelVal_in_0_3;
      end else if (10'h17 == _T_22[9:0]) begin
        image_0_23 <= io_pixelVal_in_0_2;
      end else if (10'h17 == _T_19[9:0]) begin
        image_0_23 <= io_pixelVal_in_0_1;
      end else if (10'h17 == _T_15[9:0]) begin
        image_0_23 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_24 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h18 == _T_37[9:0]) begin
        image_0_24 <= io_pixelVal_in_0_7;
      end else if (10'h18 == _T_34[9:0]) begin
        image_0_24 <= io_pixelVal_in_0_6;
      end else if (10'h18 == _T_31[9:0]) begin
        image_0_24 <= io_pixelVal_in_0_5;
      end else if (10'h18 == _T_28[9:0]) begin
        image_0_24 <= io_pixelVal_in_0_4;
      end else if (10'h18 == _T_25[9:0]) begin
        image_0_24 <= io_pixelVal_in_0_3;
      end else if (10'h18 == _T_22[9:0]) begin
        image_0_24 <= io_pixelVal_in_0_2;
      end else if (10'h18 == _T_19[9:0]) begin
        image_0_24 <= io_pixelVal_in_0_1;
      end else if (10'h18 == _T_15[9:0]) begin
        image_0_24 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_25 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h19 == _T_37[9:0]) begin
        image_0_25 <= io_pixelVal_in_0_7;
      end else if (10'h19 == _T_34[9:0]) begin
        image_0_25 <= io_pixelVal_in_0_6;
      end else if (10'h19 == _T_31[9:0]) begin
        image_0_25 <= io_pixelVal_in_0_5;
      end else if (10'h19 == _T_28[9:0]) begin
        image_0_25 <= io_pixelVal_in_0_4;
      end else if (10'h19 == _T_25[9:0]) begin
        image_0_25 <= io_pixelVal_in_0_3;
      end else if (10'h19 == _T_22[9:0]) begin
        image_0_25 <= io_pixelVal_in_0_2;
      end else if (10'h19 == _T_19[9:0]) begin
        image_0_25 <= io_pixelVal_in_0_1;
      end else if (10'h19 == _T_15[9:0]) begin
        image_0_25 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_26 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1a == _T_37[9:0]) begin
        image_0_26 <= io_pixelVal_in_0_7;
      end else if (10'h1a == _T_34[9:0]) begin
        image_0_26 <= io_pixelVal_in_0_6;
      end else if (10'h1a == _T_31[9:0]) begin
        image_0_26 <= io_pixelVal_in_0_5;
      end else if (10'h1a == _T_28[9:0]) begin
        image_0_26 <= io_pixelVal_in_0_4;
      end else if (10'h1a == _T_25[9:0]) begin
        image_0_26 <= io_pixelVal_in_0_3;
      end else if (10'h1a == _T_22[9:0]) begin
        image_0_26 <= io_pixelVal_in_0_2;
      end else if (10'h1a == _T_19[9:0]) begin
        image_0_26 <= io_pixelVal_in_0_1;
      end else if (10'h1a == _T_15[9:0]) begin
        image_0_26 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_27 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1b == _T_37[9:0]) begin
        image_0_27 <= io_pixelVal_in_0_7;
      end else if (10'h1b == _T_34[9:0]) begin
        image_0_27 <= io_pixelVal_in_0_6;
      end else if (10'h1b == _T_31[9:0]) begin
        image_0_27 <= io_pixelVal_in_0_5;
      end else if (10'h1b == _T_28[9:0]) begin
        image_0_27 <= io_pixelVal_in_0_4;
      end else if (10'h1b == _T_25[9:0]) begin
        image_0_27 <= io_pixelVal_in_0_3;
      end else if (10'h1b == _T_22[9:0]) begin
        image_0_27 <= io_pixelVal_in_0_2;
      end else if (10'h1b == _T_19[9:0]) begin
        image_0_27 <= io_pixelVal_in_0_1;
      end else if (10'h1b == _T_15[9:0]) begin
        image_0_27 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_28 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1c == _T_37[9:0]) begin
        image_0_28 <= io_pixelVal_in_0_7;
      end else if (10'h1c == _T_34[9:0]) begin
        image_0_28 <= io_pixelVal_in_0_6;
      end else if (10'h1c == _T_31[9:0]) begin
        image_0_28 <= io_pixelVal_in_0_5;
      end else if (10'h1c == _T_28[9:0]) begin
        image_0_28 <= io_pixelVal_in_0_4;
      end else if (10'h1c == _T_25[9:0]) begin
        image_0_28 <= io_pixelVal_in_0_3;
      end else if (10'h1c == _T_22[9:0]) begin
        image_0_28 <= io_pixelVal_in_0_2;
      end else if (10'h1c == _T_19[9:0]) begin
        image_0_28 <= io_pixelVal_in_0_1;
      end else if (10'h1c == _T_15[9:0]) begin
        image_0_28 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_29 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1d == _T_37[9:0]) begin
        image_0_29 <= io_pixelVal_in_0_7;
      end else if (10'h1d == _T_34[9:0]) begin
        image_0_29 <= io_pixelVal_in_0_6;
      end else if (10'h1d == _T_31[9:0]) begin
        image_0_29 <= io_pixelVal_in_0_5;
      end else if (10'h1d == _T_28[9:0]) begin
        image_0_29 <= io_pixelVal_in_0_4;
      end else if (10'h1d == _T_25[9:0]) begin
        image_0_29 <= io_pixelVal_in_0_3;
      end else if (10'h1d == _T_22[9:0]) begin
        image_0_29 <= io_pixelVal_in_0_2;
      end else if (10'h1d == _T_19[9:0]) begin
        image_0_29 <= io_pixelVal_in_0_1;
      end else if (10'h1d == _T_15[9:0]) begin
        image_0_29 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_30 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1e == _T_37[9:0]) begin
        image_0_30 <= io_pixelVal_in_0_7;
      end else if (10'h1e == _T_34[9:0]) begin
        image_0_30 <= io_pixelVal_in_0_6;
      end else if (10'h1e == _T_31[9:0]) begin
        image_0_30 <= io_pixelVal_in_0_5;
      end else if (10'h1e == _T_28[9:0]) begin
        image_0_30 <= io_pixelVal_in_0_4;
      end else if (10'h1e == _T_25[9:0]) begin
        image_0_30 <= io_pixelVal_in_0_3;
      end else if (10'h1e == _T_22[9:0]) begin
        image_0_30 <= io_pixelVal_in_0_2;
      end else if (10'h1e == _T_19[9:0]) begin
        image_0_30 <= io_pixelVal_in_0_1;
      end else if (10'h1e == _T_15[9:0]) begin
        image_0_30 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_31 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1f == _T_37[9:0]) begin
        image_0_31 <= io_pixelVal_in_0_7;
      end else if (10'h1f == _T_34[9:0]) begin
        image_0_31 <= io_pixelVal_in_0_6;
      end else if (10'h1f == _T_31[9:0]) begin
        image_0_31 <= io_pixelVal_in_0_5;
      end else if (10'h1f == _T_28[9:0]) begin
        image_0_31 <= io_pixelVal_in_0_4;
      end else if (10'h1f == _T_25[9:0]) begin
        image_0_31 <= io_pixelVal_in_0_3;
      end else if (10'h1f == _T_22[9:0]) begin
        image_0_31 <= io_pixelVal_in_0_2;
      end else if (10'h1f == _T_19[9:0]) begin
        image_0_31 <= io_pixelVal_in_0_1;
      end else if (10'h1f == _T_15[9:0]) begin
        image_0_31 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_32 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h20 == _T_37[9:0]) begin
        image_0_32 <= io_pixelVal_in_0_7;
      end else if (10'h20 == _T_34[9:0]) begin
        image_0_32 <= io_pixelVal_in_0_6;
      end else if (10'h20 == _T_31[9:0]) begin
        image_0_32 <= io_pixelVal_in_0_5;
      end else if (10'h20 == _T_28[9:0]) begin
        image_0_32 <= io_pixelVal_in_0_4;
      end else if (10'h20 == _T_25[9:0]) begin
        image_0_32 <= io_pixelVal_in_0_3;
      end else if (10'h20 == _T_22[9:0]) begin
        image_0_32 <= io_pixelVal_in_0_2;
      end else if (10'h20 == _T_19[9:0]) begin
        image_0_32 <= io_pixelVal_in_0_1;
      end else if (10'h20 == _T_15[9:0]) begin
        image_0_32 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_33 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h21 == _T_37[9:0]) begin
        image_0_33 <= io_pixelVal_in_0_7;
      end else if (10'h21 == _T_34[9:0]) begin
        image_0_33 <= io_pixelVal_in_0_6;
      end else if (10'h21 == _T_31[9:0]) begin
        image_0_33 <= io_pixelVal_in_0_5;
      end else if (10'h21 == _T_28[9:0]) begin
        image_0_33 <= io_pixelVal_in_0_4;
      end else if (10'h21 == _T_25[9:0]) begin
        image_0_33 <= io_pixelVal_in_0_3;
      end else if (10'h21 == _T_22[9:0]) begin
        image_0_33 <= io_pixelVal_in_0_2;
      end else if (10'h21 == _T_19[9:0]) begin
        image_0_33 <= io_pixelVal_in_0_1;
      end else if (10'h21 == _T_15[9:0]) begin
        image_0_33 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_34 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h22 == _T_37[9:0]) begin
        image_0_34 <= io_pixelVal_in_0_7;
      end else if (10'h22 == _T_34[9:0]) begin
        image_0_34 <= io_pixelVal_in_0_6;
      end else if (10'h22 == _T_31[9:0]) begin
        image_0_34 <= io_pixelVal_in_0_5;
      end else if (10'h22 == _T_28[9:0]) begin
        image_0_34 <= io_pixelVal_in_0_4;
      end else if (10'h22 == _T_25[9:0]) begin
        image_0_34 <= io_pixelVal_in_0_3;
      end else if (10'h22 == _T_22[9:0]) begin
        image_0_34 <= io_pixelVal_in_0_2;
      end else if (10'h22 == _T_19[9:0]) begin
        image_0_34 <= io_pixelVal_in_0_1;
      end else if (10'h22 == _T_15[9:0]) begin
        image_0_34 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_35 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h23 == _T_37[9:0]) begin
        image_0_35 <= io_pixelVal_in_0_7;
      end else if (10'h23 == _T_34[9:0]) begin
        image_0_35 <= io_pixelVal_in_0_6;
      end else if (10'h23 == _T_31[9:0]) begin
        image_0_35 <= io_pixelVal_in_0_5;
      end else if (10'h23 == _T_28[9:0]) begin
        image_0_35 <= io_pixelVal_in_0_4;
      end else if (10'h23 == _T_25[9:0]) begin
        image_0_35 <= io_pixelVal_in_0_3;
      end else if (10'h23 == _T_22[9:0]) begin
        image_0_35 <= io_pixelVal_in_0_2;
      end else if (10'h23 == _T_19[9:0]) begin
        image_0_35 <= io_pixelVal_in_0_1;
      end else if (10'h23 == _T_15[9:0]) begin
        image_0_35 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_36 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h24 == _T_37[9:0]) begin
        image_0_36 <= io_pixelVal_in_0_7;
      end else if (10'h24 == _T_34[9:0]) begin
        image_0_36 <= io_pixelVal_in_0_6;
      end else if (10'h24 == _T_31[9:0]) begin
        image_0_36 <= io_pixelVal_in_0_5;
      end else if (10'h24 == _T_28[9:0]) begin
        image_0_36 <= io_pixelVal_in_0_4;
      end else if (10'h24 == _T_25[9:0]) begin
        image_0_36 <= io_pixelVal_in_0_3;
      end else if (10'h24 == _T_22[9:0]) begin
        image_0_36 <= io_pixelVal_in_0_2;
      end else if (10'h24 == _T_19[9:0]) begin
        image_0_36 <= io_pixelVal_in_0_1;
      end else if (10'h24 == _T_15[9:0]) begin
        image_0_36 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_37 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h25 == _T_37[9:0]) begin
        image_0_37 <= io_pixelVal_in_0_7;
      end else if (10'h25 == _T_34[9:0]) begin
        image_0_37 <= io_pixelVal_in_0_6;
      end else if (10'h25 == _T_31[9:0]) begin
        image_0_37 <= io_pixelVal_in_0_5;
      end else if (10'h25 == _T_28[9:0]) begin
        image_0_37 <= io_pixelVal_in_0_4;
      end else if (10'h25 == _T_25[9:0]) begin
        image_0_37 <= io_pixelVal_in_0_3;
      end else if (10'h25 == _T_22[9:0]) begin
        image_0_37 <= io_pixelVal_in_0_2;
      end else if (10'h25 == _T_19[9:0]) begin
        image_0_37 <= io_pixelVal_in_0_1;
      end else if (10'h25 == _T_15[9:0]) begin
        image_0_37 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_38 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h26 == _T_37[9:0]) begin
        image_0_38 <= io_pixelVal_in_0_7;
      end else if (10'h26 == _T_34[9:0]) begin
        image_0_38 <= io_pixelVal_in_0_6;
      end else if (10'h26 == _T_31[9:0]) begin
        image_0_38 <= io_pixelVal_in_0_5;
      end else if (10'h26 == _T_28[9:0]) begin
        image_0_38 <= io_pixelVal_in_0_4;
      end else if (10'h26 == _T_25[9:0]) begin
        image_0_38 <= io_pixelVal_in_0_3;
      end else if (10'h26 == _T_22[9:0]) begin
        image_0_38 <= io_pixelVal_in_0_2;
      end else if (10'h26 == _T_19[9:0]) begin
        image_0_38 <= io_pixelVal_in_0_1;
      end else if (10'h26 == _T_15[9:0]) begin
        image_0_38 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_39 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h27 == _T_37[9:0]) begin
        image_0_39 <= io_pixelVal_in_0_7;
      end else if (10'h27 == _T_34[9:0]) begin
        image_0_39 <= io_pixelVal_in_0_6;
      end else if (10'h27 == _T_31[9:0]) begin
        image_0_39 <= io_pixelVal_in_0_5;
      end else if (10'h27 == _T_28[9:0]) begin
        image_0_39 <= io_pixelVal_in_0_4;
      end else if (10'h27 == _T_25[9:0]) begin
        image_0_39 <= io_pixelVal_in_0_3;
      end else if (10'h27 == _T_22[9:0]) begin
        image_0_39 <= io_pixelVal_in_0_2;
      end else if (10'h27 == _T_19[9:0]) begin
        image_0_39 <= io_pixelVal_in_0_1;
      end else if (10'h27 == _T_15[9:0]) begin
        image_0_39 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_40 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h28 == _T_37[9:0]) begin
        image_0_40 <= io_pixelVal_in_0_7;
      end else if (10'h28 == _T_34[9:0]) begin
        image_0_40 <= io_pixelVal_in_0_6;
      end else if (10'h28 == _T_31[9:0]) begin
        image_0_40 <= io_pixelVal_in_0_5;
      end else if (10'h28 == _T_28[9:0]) begin
        image_0_40 <= io_pixelVal_in_0_4;
      end else if (10'h28 == _T_25[9:0]) begin
        image_0_40 <= io_pixelVal_in_0_3;
      end else if (10'h28 == _T_22[9:0]) begin
        image_0_40 <= io_pixelVal_in_0_2;
      end else if (10'h28 == _T_19[9:0]) begin
        image_0_40 <= io_pixelVal_in_0_1;
      end else if (10'h28 == _T_15[9:0]) begin
        image_0_40 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_41 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h29 == _T_37[9:0]) begin
        image_0_41 <= io_pixelVal_in_0_7;
      end else if (10'h29 == _T_34[9:0]) begin
        image_0_41 <= io_pixelVal_in_0_6;
      end else if (10'h29 == _T_31[9:0]) begin
        image_0_41 <= io_pixelVal_in_0_5;
      end else if (10'h29 == _T_28[9:0]) begin
        image_0_41 <= io_pixelVal_in_0_4;
      end else if (10'h29 == _T_25[9:0]) begin
        image_0_41 <= io_pixelVal_in_0_3;
      end else if (10'h29 == _T_22[9:0]) begin
        image_0_41 <= io_pixelVal_in_0_2;
      end else if (10'h29 == _T_19[9:0]) begin
        image_0_41 <= io_pixelVal_in_0_1;
      end else if (10'h29 == _T_15[9:0]) begin
        image_0_41 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_42 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h2a == _T_37[9:0]) begin
        image_0_42 <= io_pixelVal_in_0_7;
      end else if (10'h2a == _T_34[9:0]) begin
        image_0_42 <= io_pixelVal_in_0_6;
      end else if (10'h2a == _T_31[9:0]) begin
        image_0_42 <= io_pixelVal_in_0_5;
      end else if (10'h2a == _T_28[9:0]) begin
        image_0_42 <= io_pixelVal_in_0_4;
      end else if (10'h2a == _T_25[9:0]) begin
        image_0_42 <= io_pixelVal_in_0_3;
      end else if (10'h2a == _T_22[9:0]) begin
        image_0_42 <= io_pixelVal_in_0_2;
      end else if (10'h2a == _T_19[9:0]) begin
        image_0_42 <= io_pixelVal_in_0_1;
      end else if (10'h2a == _T_15[9:0]) begin
        image_0_42 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_43 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h2b == _T_37[9:0]) begin
        image_0_43 <= io_pixelVal_in_0_7;
      end else if (10'h2b == _T_34[9:0]) begin
        image_0_43 <= io_pixelVal_in_0_6;
      end else if (10'h2b == _T_31[9:0]) begin
        image_0_43 <= io_pixelVal_in_0_5;
      end else if (10'h2b == _T_28[9:0]) begin
        image_0_43 <= io_pixelVal_in_0_4;
      end else if (10'h2b == _T_25[9:0]) begin
        image_0_43 <= io_pixelVal_in_0_3;
      end else if (10'h2b == _T_22[9:0]) begin
        image_0_43 <= io_pixelVal_in_0_2;
      end else if (10'h2b == _T_19[9:0]) begin
        image_0_43 <= io_pixelVal_in_0_1;
      end else if (10'h2b == _T_15[9:0]) begin
        image_0_43 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_44 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h2c == _T_37[9:0]) begin
        image_0_44 <= io_pixelVal_in_0_7;
      end else if (10'h2c == _T_34[9:0]) begin
        image_0_44 <= io_pixelVal_in_0_6;
      end else if (10'h2c == _T_31[9:0]) begin
        image_0_44 <= io_pixelVal_in_0_5;
      end else if (10'h2c == _T_28[9:0]) begin
        image_0_44 <= io_pixelVal_in_0_4;
      end else if (10'h2c == _T_25[9:0]) begin
        image_0_44 <= io_pixelVal_in_0_3;
      end else if (10'h2c == _T_22[9:0]) begin
        image_0_44 <= io_pixelVal_in_0_2;
      end else if (10'h2c == _T_19[9:0]) begin
        image_0_44 <= io_pixelVal_in_0_1;
      end else if (10'h2c == _T_15[9:0]) begin
        image_0_44 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_45 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h2d == _T_37[9:0]) begin
        image_0_45 <= io_pixelVal_in_0_7;
      end else if (10'h2d == _T_34[9:0]) begin
        image_0_45 <= io_pixelVal_in_0_6;
      end else if (10'h2d == _T_31[9:0]) begin
        image_0_45 <= io_pixelVal_in_0_5;
      end else if (10'h2d == _T_28[9:0]) begin
        image_0_45 <= io_pixelVal_in_0_4;
      end else if (10'h2d == _T_25[9:0]) begin
        image_0_45 <= io_pixelVal_in_0_3;
      end else if (10'h2d == _T_22[9:0]) begin
        image_0_45 <= io_pixelVal_in_0_2;
      end else if (10'h2d == _T_19[9:0]) begin
        image_0_45 <= io_pixelVal_in_0_1;
      end else if (10'h2d == _T_15[9:0]) begin
        image_0_45 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_46 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h2e == _T_37[9:0]) begin
        image_0_46 <= io_pixelVal_in_0_7;
      end else if (10'h2e == _T_34[9:0]) begin
        image_0_46 <= io_pixelVal_in_0_6;
      end else if (10'h2e == _T_31[9:0]) begin
        image_0_46 <= io_pixelVal_in_0_5;
      end else if (10'h2e == _T_28[9:0]) begin
        image_0_46 <= io_pixelVal_in_0_4;
      end else if (10'h2e == _T_25[9:0]) begin
        image_0_46 <= io_pixelVal_in_0_3;
      end else if (10'h2e == _T_22[9:0]) begin
        image_0_46 <= io_pixelVal_in_0_2;
      end else if (10'h2e == _T_19[9:0]) begin
        image_0_46 <= io_pixelVal_in_0_1;
      end else if (10'h2e == _T_15[9:0]) begin
        image_0_46 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_47 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h2f == _T_37[9:0]) begin
        image_0_47 <= io_pixelVal_in_0_7;
      end else if (10'h2f == _T_34[9:0]) begin
        image_0_47 <= io_pixelVal_in_0_6;
      end else if (10'h2f == _T_31[9:0]) begin
        image_0_47 <= io_pixelVal_in_0_5;
      end else if (10'h2f == _T_28[9:0]) begin
        image_0_47 <= io_pixelVal_in_0_4;
      end else if (10'h2f == _T_25[9:0]) begin
        image_0_47 <= io_pixelVal_in_0_3;
      end else if (10'h2f == _T_22[9:0]) begin
        image_0_47 <= io_pixelVal_in_0_2;
      end else if (10'h2f == _T_19[9:0]) begin
        image_0_47 <= io_pixelVal_in_0_1;
      end else if (10'h2f == _T_15[9:0]) begin
        image_0_47 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_48 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h30 == _T_37[9:0]) begin
        image_0_48 <= io_pixelVal_in_0_7;
      end else if (10'h30 == _T_34[9:0]) begin
        image_0_48 <= io_pixelVal_in_0_6;
      end else if (10'h30 == _T_31[9:0]) begin
        image_0_48 <= io_pixelVal_in_0_5;
      end else if (10'h30 == _T_28[9:0]) begin
        image_0_48 <= io_pixelVal_in_0_4;
      end else if (10'h30 == _T_25[9:0]) begin
        image_0_48 <= io_pixelVal_in_0_3;
      end else if (10'h30 == _T_22[9:0]) begin
        image_0_48 <= io_pixelVal_in_0_2;
      end else if (10'h30 == _T_19[9:0]) begin
        image_0_48 <= io_pixelVal_in_0_1;
      end else if (10'h30 == _T_15[9:0]) begin
        image_0_48 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_49 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h31 == _T_37[9:0]) begin
        image_0_49 <= io_pixelVal_in_0_7;
      end else if (10'h31 == _T_34[9:0]) begin
        image_0_49 <= io_pixelVal_in_0_6;
      end else if (10'h31 == _T_31[9:0]) begin
        image_0_49 <= io_pixelVal_in_0_5;
      end else if (10'h31 == _T_28[9:0]) begin
        image_0_49 <= io_pixelVal_in_0_4;
      end else if (10'h31 == _T_25[9:0]) begin
        image_0_49 <= io_pixelVal_in_0_3;
      end else if (10'h31 == _T_22[9:0]) begin
        image_0_49 <= io_pixelVal_in_0_2;
      end else if (10'h31 == _T_19[9:0]) begin
        image_0_49 <= io_pixelVal_in_0_1;
      end else if (10'h31 == _T_15[9:0]) begin
        image_0_49 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_50 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h32 == _T_37[9:0]) begin
        image_0_50 <= io_pixelVal_in_0_7;
      end else if (10'h32 == _T_34[9:0]) begin
        image_0_50 <= io_pixelVal_in_0_6;
      end else if (10'h32 == _T_31[9:0]) begin
        image_0_50 <= io_pixelVal_in_0_5;
      end else if (10'h32 == _T_28[9:0]) begin
        image_0_50 <= io_pixelVal_in_0_4;
      end else if (10'h32 == _T_25[9:0]) begin
        image_0_50 <= io_pixelVal_in_0_3;
      end else if (10'h32 == _T_22[9:0]) begin
        image_0_50 <= io_pixelVal_in_0_2;
      end else if (10'h32 == _T_19[9:0]) begin
        image_0_50 <= io_pixelVal_in_0_1;
      end else if (10'h32 == _T_15[9:0]) begin
        image_0_50 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_51 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h33 == _T_37[9:0]) begin
        image_0_51 <= io_pixelVal_in_0_7;
      end else if (10'h33 == _T_34[9:0]) begin
        image_0_51 <= io_pixelVal_in_0_6;
      end else if (10'h33 == _T_31[9:0]) begin
        image_0_51 <= io_pixelVal_in_0_5;
      end else if (10'h33 == _T_28[9:0]) begin
        image_0_51 <= io_pixelVal_in_0_4;
      end else if (10'h33 == _T_25[9:0]) begin
        image_0_51 <= io_pixelVal_in_0_3;
      end else if (10'h33 == _T_22[9:0]) begin
        image_0_51 <= io_pixelVal_in_0_2;
      end else if (10'h33 == _T_19[9:0]) begin
        image_0_51 <= io_pixelVal_in_0_1;
      end else if (10'h33 == _T_15[9:0]) begin
        image_0_51 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_52 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h34 == _T_37[9:0]) begin
        image_0_52 <= io_pixelVal_in_0_7;
      end else if (10'h34 == _T_34[9:0]) begin
        image_0_52 <= io_pixelVal_in_0_6;
      end else if (10'h34 == _T_31[9:0]) begin
        image_0_52 <= io_pixelVal_in_0_5;
      end else if (10'h34 == _T_28[9:0]) begin
        image_0_52 <= io_pixelVal_in_0_4;
      end else if (10'h34 == _T_25[9:0]) begin
        image_0_52 <= io_pixelVal_in_0_3;
      end else if (10'h34 == _T_22[9:0]) begin
        image_0_52 <= io_pixelVal_in_0_2;
      end else if (10'h34 == _T_19[9:0]) begin
        image_0_52 <= io_pixelVal_in_0_1;
      end else if (10'h34 == _T_15[9:0]) begin
        image_0_52 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_53 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h35 == _T_37[9:0]) begin
        image_0_53 <= io_pixelVal_in_0_7;
      end else if (10'h35 == _T_34[9:0]) begin
        image_0_53 <= io_pixelVal_in_0_6;
      end else if (10'h35 == _T_31[9:0]) begin
        image_0_53 <= io_pixelVal_in_0_5;
      end else if (10'h35 == _T_28[9:0]) begin
        image_0_53 <= io_pixelVal_in_0_4;
      end else if (10'h35 == _T_25[9:0]) begin
        image_0_53 <= io_pixelVal_in_0_3;
      end else if (10'h35 == _T_22[9:0]) begin
        image_0_53 <= io_pixelVal_in_0_2;
      end else if (10'h35 == _T_19[9:0]) begin
        image_0_53 <= io_pixelVal_in_0_1;
      end else if (10'h35 == _T_15[9:0]) begin
        image_0_53 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_54 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h36 == _T_37[9:0]) begin
        image_0_54 <= io_pixelVal_in_0_7;
      end else if (10'h36 == _T_34[9:0]) begin
        image_0_54 <= io_pixelVal_in_0_6;
      end else if (10'h36 == _T_31[9:0]) begin
        image_0_54 <= io_pixelVal_in_0_5;
      end else if (10'h36 == _T_28[9:0]) begin
        image_0_54 <= io_pixelVal_in_0_4;
      end else if (10'h36 == _T_25[9:0]) begin
        image_0_54 <= io_pixelVal_in_0_3;
      end else if (10'h36 == _T_22[9:0]) begin
        image_0_54 <= io_pixelVal_in_0_2;
      end else if (10'h36 == _T_19[9:0]) begin
        image_0_54 <= io_pixelVal_in_0_1;
      end else if (10'h36 == _T_15[9:0]) begin
        image_0_54 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_55 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h37 == _T_37[9:0]) begin
        image_0_55 <= io_pixelVal_in_0_7;
      end else if (10'h37 == _T_34[9:0]) begin
        image_0_55 <= io_pixelVal_in_0_6;
      end else if (10'h37 == _T_31[9:0]) begin
        image_0_55 <= io_pixelVal_in_0_5;
      end else if (10'h37 == _T_28[9:0]) begin
        image_0_55 <= io_pixelVal_in_0_4;
      end else if (10'h37 == _T_25[9:0]) begin
        image_0_55 <= io_pixelVal_in_0_3;
      end else if (10'h37 == _T_22[9:0]) begin
        image_0_55 <= io_pixelVal_in_0_2;
      end else if (10'h37 == _T_19[9:0]) begin
        image_0_55 <= io_pixelVal_in_0_1;
      end else if (10'h37 == _T_15[9:0]) begin
        image_0_55 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_56 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h38 == _T_37[9:0]) begin
        image_0_56 <= io_pixelVal_in_0_7;
      end else if (10'h38 == _T_34[9:0]) begin
        image_0_56 <= io_pixelVal_in_0_6;
      end else if (10'h38 == _T_31[9:0]) begin
        image_0_56 <= io_pixelVal_in_0_5;
      end else if (10'h38 == _T_28[9:0]) begin
        image_0_56 <= io_pixelVal_in_0_4;
      end else if (10'h38 == _T_25[9:0]) begin
        image_0_56 <= io_pixelVal_in_0_3;
      end else if (10'h38 == _T_22[9:0]) begin
        image_0_56 <= io_pixelVal_in_0_2;
      end else if (10'h38 == _T_19[9:0]) begin
        image_0_56 <= io_pixelVal_in_0_1;
      end else if (10'h38 == _T_15[9:0]) begin
        image_0_56 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_57 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h39 == _T_37[9:0]) begin
        image_0_57 <= io_pixelVal_in_0_7;
      end else if (10'h39 == _T_34[9:0]) begin
        image_0_57 <= io_pixelVal_in_0_6;
      end else if (10'h39 == _T_31[9:0]) begin
        image_0_57 <= io_pixelVal_in_0_5;
      end else if (10'h39 == _T_28[9:0]) begin
        image_0_57 <= io_pixelVal_in_0_4;
      end else if (10'h39 == _T_25[9:0]) begin
        image_0_57 <= io_pixelVal_in_0_3;
      end else if (10'h39 == _T_22[9:0]) begin
        image_0_57 <= io_pixelVal_in_0_2;
      end else if (10'h39 == _T_19[9:0]) begin
        image_0_57 <= io_pixelVal_in_0_1;
      end else if (10'h39 == _T_15[9:0]) begin
        image_0_57 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_58 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h3a == _T_37[9:0]) begin
        image_0_58 <= io_pixelVal_in_0_7;
      end else if (10'h3a == _T_34[9:0]) begin
        image_0_58 <= io_pixelVal_in_0_6;
      end else if (10'h3a == _T_31[9:0]) begin
        image_0_58 <= io_pixelVal_in_0_5;
      end else if (10'h3a == _T_28[9:0]) begin
        image_0_58 <= io_pixelVal_in_0_4;
      end else if (10'h3a == _T_25[9:0]) begin
        image_0_58 <= io_pixelVal_in_0_3;
      end else if (10'h3a == _T_22[9:0]) begin
        image_0_58 <= io_pixelVal_in_0_2;
      end else if (10'h3a == _T_19[9:0]) begin
        image_0_58 <= io_pixelVal_in_0_1;
      end else if (10'h3a == _T_15[9:0]) begin
        image_0_58 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_59 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h3b == _T_37[9:0]) begin
        image_0_59 <= io_pixelVal_in_0_7;
      end else if (10'h3b == _T_34[9:0]) begin
        image_0_59 <= io_pixelVal_in_0_6;
      end else if (10'h3b == _T_31[9:0]) begin
        image_0_59 <= io_pixelVal_in_0_5;
      end else if (10'h3b == _T_28[9:0]) begin
        image_0_59 <= io_pixelVal_in_0_4;
      end else if (10'h3b == _T_25[9:0]) begin
        image_0_59 <= io_pixelVal_in_0_3;
      end else if (10'h3b == _T_22[9:0]) begin
        image_0_59 <= io_pixelVal_in_0_2;
      end else if (10'h3b == _T_19[9:0]) begin
        image_0_59 <= io_pixelVal_in_0_1;
      end else if (10'h3b == _T_15[9:0]) begin
        image_0_59 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_60 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h3c == _T_37[9:0]) begin
        image_0_60 <= io_pixelVal_in_0_7;
      end else if (10'h3c == _T_34[9:0]) begin
        image_0_60 <= io_pixelVal_in_0_6;
      end else if (10'h3c == _T_31[9:0]) begin
        image_0_60 <= io_pixelVal_in_0_5;
      end else if (10'h3c == _T_28[9:0]) begin
        image_0_60 <= io_pixelVal_in_0_4;
      end else if (10'h3c == _T_25[9:0]) begin
        image_0_60 <= io_pixelVal_in_0_3;
      end else if (10'h3c == _T_22[9:0]) begin
        image_0_60 <= io_pixelVal_in_0_2;
      end else if (10'h3c == _T_19[9:0]) begin
        image_0_60 <= io_pixelVal_in_0_1;
      end else if (10'h3c == _T_15[9:0]) begin
        image_0_60 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_61 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h3d == _T_37[9:0]) begin
        image_0_61 <= io_pixelVal_in_0_7;
      end else if (10'h3d == _T_34[9:0]) begin
        image_0_61 <= io_pixelVal_in_0_6;
      end else if (10'h3d == _T_31[9:0]) begin
        image_0_61 <= io_pixelVal_in_0_5;
      end else if (10'h3d == _T_28[9:0]) begin
        image_0_61 <= io_pixelVal_in_0_4;
      end else if (10'h3d == _T_25[9:0]) begin
        image_0_61 <= io_pixelVal_in_0_3;
      end else if (10'h3d == _T_22[9:0]) begin
        image_0_61 <= io_pixelVal_in_0_2;
      end else if (10'h3d == _T_19[9:0]) begin
        image_0_61 <= io_pixelVal_in_0_1;
      end else if (10'h3d == _T_15[9:0]) begin
        image_0_61 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_62 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h3e == _T_37[9:0]) begin
        image_0_62 <= io_pixelVal_in_0_7;
      end else if (10'h3e == _T_34[9:0]) begin
        image_0_62 <= io_pixelVal_in_0_6;
      end else if (10'h3e == _T_31[9:0]) begin
        image_0_62 <= io_pixelVal_in_0_5;
      end else if (10'h3e == _T_28[9:0]) begin
        image_0_62 <= io_pixelVal_in_0_4;
      end else if (10'h3e == _T_25[9:0]) begin
        image_0_62 <= io_pixelVal_in_0_3;
      end else if (10'h3e == _T_22[9:0]) begin
        image_0_62 <= io_pixelVal_in_0_2;
      end else if (10'h3e == _T_19[9:0]) begin
        image_0_62 <= io_pixelVal_in_0_1;
      end else if (10'h3e == _T_15[9:0]) begin
        image_0_62 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_63 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h3f == _T_37[9:0]) begin
        image_0_63 <= io_pixelVal_in_0_7;
      end else if (10'h3f == _T_34[9:0]) begin
        image_0_63 <= io_pixelVal_in_0_6;
      end else if (10'h3f == _T_31[9:0]) begin
        image_0_63 <= io_pixelVal_in_0_5;
      end else if (10'h3f == _T_28[9:0]) begin
        image_0_63 <= io_pixelVal_in_0_4;
      end else if (10'h3f == _T_25[9:0]) begin
        image_0_63 <= io_pixelVal_in_0_3;
      end else if (10'h3f == _T_22[9:0]) begin
        image_0_63 <= io_pixelVal_in_0_2;
      end else if (10'h3f == _T_19[9:0]) begin
        image_0_63 <= io_pixelVal_in_0_1;
      end else if (10'h3f == _T_15[9:0]) begin
        image_0_63 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_64 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h40 == _T_37[9:0]) begin
        image_0_64 <= io_pixelVal_in_0_7;
      end else if (10'h40 == _T_34[9:0]) begin
        image_0_64 <= io_pixelVal_in_0_6;
      end else if (10'h40 == _T_31[9:0]) begin
        image_0_64 <= io_pixelVal_in_0_5;
      end else if (10'h40 == _T_28[9:0]) begin
        image_0_64 <= io_pixelVal_in_0_4;
      end else if (10'h40 == _T_25[9:0]) begin
        image_0_64 <= io_pixelVal_in_0_3;
      end else if (10'h40 == _T_22[9:0]) begin
        image_0_64 <= io_pixelVal_in_0_2;
      end else if (10'h40 == _T_19[9:0]) begin
        image_0_64 <= io_pixelVal_in_0_1;
      end else if (10'h40 == _T_15[9:0]) begin
        image_0_64 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_65 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h41 == _T_37[9:0]) begin
        image_0_65 <= io_pixelVal_in_0_7;
      end else if (10'h41 == _T_34[9:0]) begin
        image_0_65 <= io_pixelVal_in_0_6;
      end else if (10'h41 == _T_31[9:0]) begin
        image_0_65 <= io_pixelVal_in_0_5;
      end else if (10'h41 == _T_28[9:0]) begin
        image_0_65 <= io_pixelVal_in_0_4;
      end else if (10'h41 == _T_25[9:0]) begin
        image_0_65 <= io_pixelVal_in_0_3;
      end else if (10'h41 == _T_22[9:0]) begin
        image_0_65 <= io_pixelVal_in_0_2;
      end else if (10'h41 == _T_19[9:0]) begin
        image_0_65 <= io_pixelVal_in_0_1;
      end else if (10'h41 == _T_15[9:0]) begin
        image_0_65 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_66 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h42 == _T_37[9:0]) begin
        image_0_66 <= io_pixelVal_in_0_7;
      end else if (10'h42 == _T_34[9:0]) begin
        image_0_66 <= io_pixelVal_in_0_6;
      end else if (10'h42 == _T_31[9:0]) begin
        image_0_66 <= io_pixelVal_in_0_5;
      end else if (10'h42 == _T_28[9:0]) begin
        image_0_66 <= io_pixelVal_in_0_4;
      end else if (10'h42 == _T_25[9:0]) begin
        image_0_66 <= io_pixelVal_in_0_3;
      end else if (10'h42 == _T_22[9:0]) begin
        image_0_66 <= io_pixelVal_in_0_2;
      end else if (10'h42 == _T_19[9:0]) begin
        image_0_66 <= io_pixelVal_in_0_1;
      end else if (10'h42 == _T_15[9:0]) begin
        image_0_66 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_67 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h43 == _T_37[9:0]) begin
        image_0_67 <= io_pixelVal_in_0_7;
      end else if (10'h43 == _T_34[9:0]) begin
        image_0_67 <= io_pixelVal_in_0_6;
      end else if (10'h43 == _T_31[9:0]) begin
        image_0_67 <= io_pixelVal_in_0_5;
      end else if (10'h43 == _T_28[9:0]) begin
        image_0_67 <= io_pixelVal_in_0_4;
      end else if (10'h43 == _T_25[9:0]) begin
        image_0_67 <= io_pixelVal_in_0_3;
      end else if (10'h43 == _T_22[9:0]) begin
        image_0_67 <= io_pixelVal_in_0_2;
      end else if (10'h43 == _T_19[9:0]) begin
        image_0_67 <= io_pixelVal_in_0_1;
      end else if (10'h43 == _T_15[9:0]) begin
        image_0_67 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_68 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h44 == _T_37[9:0]) begin
        image_0_68 <= io_pixelVal_in_0_7;
      end else if (10'h44 == _T_34[9:0]) begin
        image_0_68 <= io_pixelVal_in_0_6;
      end else if (10'h44 == _T_31[9:0]) begin
        image_0_68 <= io_pixelVal_in_0_5;
      end else if (10'h44 == _T_28[9:0]) begin
        image_0_68 <= io_pixelVal_in_0_4;
      end else if (10'h44 == _T_25[9:0]) begin
        image_0_68 <= io_pixelVal_in_0_3;
      end else if (10'h44 == _T_22[9:0]) begin
        image_0_68 <= io_pixelVal_in_0_2;
      end else if (10'h44 == _T_19[9:0]) begin
        image_0_68 <= io_pixelVal_in_0_1;
      end else if (10'h44 == _T_15[9:0]) begin
        image_0_68 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_69 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h45 == _T_37[9:0]) begin
        image_0_69 <= io_pixelVal_in_0_7;
      end else if (10'h45 == _T_34[9:0]) begin
        image_0_69 <= io_pixelVal_in_0_6;
      end else if (10'h45 == _T_31[9:0]) begin
        image_0_69 <= io_pixelVal_in_0_5;
      end else if (10'h45 == _T_28[9:0]) begin
        image_0_69 <= io_pixelVal_in_0_4;
      end else if (10'h45 == _T_25[9:0]) begin
        image_0_69 <= io_pixelVal_in_0_3;
      end else if (10'h45 == _T_22[9:0]) begin
        image_0_69 <= io_pixelVal_in_0_2;
      end else if (10'h45 == _T_19[9:0]) begin
        image_0_69 <= io_pixelVal_in_0_1;
      end else if (10'h45 == _T_15[9:0]) begin
        image_0_69 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_70 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h46 == _T_37[9:0]) begin
        image_0_70 <= io_pixelVal_in_0_7;
      end else if (10'h46 == _T_34[9:0]) begin
        image_0_70 <= io_pixelVal_in_0_6;
      end else if (10'h46 == _T_31[9:0]) begin
        image_0_70 <= io_pixelVal_in_0_5;
      end else if (10'h46 == _T_28[9:0]) begin
        image_0_70 <= io_pixelVal_in_0_4;
      end else if (10'h46 == _T_25[9:0]) begin
        image_0_70 <= io_pixelVal_in_0_3;
      end else if (10'h46 == _T_22[9:0]) begin
        image_0_70 <= io_pixelVal_in_0_2;
      end else if (10'h46 == _T_19[9:0]) begin
        image_0_70 <= io_pixelVal_in_0_1;
      end else if (10'h46 == _T_15[9:0]) begin
        image_0_70 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_71 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h47 == _T_37[9:0]) begin
        image_0_71 <= io_pixelVal_in_0_7;
      end else if (10'h47 == _T_34[9:0]) begin
        image_0_71 <= io_pixelVal_in_0_6;
      end else if (10'h47 == _T_31[9:0]) begin
        image_0_71 <= io_pixelVal_in_0_5;
      end else if (10'h47 == _T_28[9:0]) begin
        image_0_71 <= io_pixelVal_in_0_4;
      end else if (10'h47 == _T_25[9:0]) begin
        image_0_71 <= io_pixelVal_in_0_3;
      end else if (10'h47 == _T_22[9:0]) begin
        image_0_71 <= io_pixelVal_in_0_2;
      end else if (10'h47 == _T_19[9:0]) begin
        image_0_71 <= io_pixelVal_in_0_1;
      end else if (10'h47 == _T_15[9:0]) begin
        image_0_71 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_72 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h48 == _T_37[9:0]) begin
        image_0_72 <= io_pixelVal_in_0_7;
      end else if (10'h48 == _T_34[9:0]) begin
        image_0_72 <= io_pixelVal_in_0_6;
      end else if (10'h48 == _T_31[9:0]) begin
        image_0_72 <= io_pixelVal_in_0_5;
      end else if (10'h48 == _T_28[9:0]) begin
        image_0_72 <= io_pixelVal_in_0_4;
      end else if (10'h48 == _T_25[9:0]) begin
        image_0_72 <= io_pixelVal_in_0_3;
      end else if (10'h48 == _T_22[9:0]) begin
        image_0_72 <= io_pixelVal_in_0_2;
      end else if (10'h48 == _T_19[9:0]) begin
        image_0_72 <= io_pixelVal_in_0_1;
      end else if (10'h48 == _T_15[9:0]) begin
        image_0_72 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_73 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h49 == _T_37[9:0]) begin
        image_0_73 <= io_pixelVal_in_0_7;
      end else if (10'h49 == _T_34[9:0]) begin
        image_0_73 <= io_pixelVal_in_0_6;
      end else if (10'h49 == _T_31[9:0]) begin
        image_0_73 <= io_pixelVal_in_0_5;
      end else if (10'h49 == _T_28[9:0]) begin
        image_0_73 <= io_pixelVal_in_0_4;
      end else if (10'h49 == _T_25[9:0]) begin
        image_0_73 <= io_pixelVal_in_0_3;
      end else if (10'h49 == _T_22[9:0]) begin
        image_0_73 <= io_pixelVal_in_0_2;
      end else if (10'h49 == _T_19[9:0]) begin
        image_0_73 <= io_pixelVal_in_0_1;
      end else if (10'h49 == _T_15[9:0]) begin
        image_0_73 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_74 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h4a == _T_37[9:0]) begin
        image_0_74 <= io_pixelVal_in_0_7;
      end else if (10'h4a == _T_34[9:0]) begin
        image_0_74 <= io_pixelVal_in_0_6;
      end else if (10'h4a == _T_31[9:0]) begin
        image_0_74 <= io_pixelVal_in_0_5;
      end else if (10'h4a == _T_28[9:0]) begin
        image_0_74 <= io_pixelVal_in_0_4;
      end else if (10'h4a == _T_25[9:0]) begin
        image_0_74 <= io_pixelVal_in_0_3;
      end else if (10'h4a == _T_22[9:0]) begin
        image_0_74 <= io_pixelVal_in_0_2;
      end else if (10'h4a == _T_19[9:0]) begin
        image_0_74 <= io_pixelVal_in_0_1;
      end else if (10'h4a == _T_15[9:0]) begin
        image_0_74 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_75 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h4b == _T_37[9:0]) begin
        image_0_75 <= io_pixelVal_in_0_7;
      end else if (10'h4b == _T_34[9:0]) begin
        image_0_75 <= io_pixelVal_in_0_6;
      end else if (10'h4b == _T_31[9:0]) begin
        image_0_75 <= io_pixelVal_in_0_5;
      end else if (10'h4b == _T_28[9:0]) begin
        image_0_75 <= io_pixelVal_in_0_4;
      end else if (10'h4b == _T_25[9:0]) begin
        image_0_75 <= io_pixelVal_in_0_3;
      end else if (10'h4b == _T_22[9:0]) begin
        image_0_75 <= io_pixelVal_in_0_2;
      end else if (10'h4b == _T_19[9:0]) begin
        image_0_75 <= io_pixelVal_in_0_1;
      end else if (10'h4b == _T_15[9:0]) begin
        image_0_75 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_76 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h4c == _T_37[9:0]) begin
        image_0_76 <= io_pixelVal_in_0_7;
      end else if (10'h4c == _T_34[9:0]) begin
        image_0_76 <= io_pixelVal_in_0_6;
      end else if (10'h4c == _T_31[9:0]) begin
        image_0_76 <= io_pixelVal_in_0_5;
      end else if (10'h4c == _T_28[9:0]) begin
        image_0_76 <= io_pixelVal_in_0_4;
      end else if (10'h4c == _T_25[9:0]) begin
        image_0_76 <= io_pixelVal_in_0_3;
      end else if (10'h4c == _T_22[9:0]) begin
        image_0_76 <= io_pixelVal_in_0_2;
      end else if (10'h4c == _T_19[9:0]) begin
        image_0_76 <= io_pixelVal_in_0_1;
      end else if (10'h4c == _T_15[9:0]) begin
        image_0_76 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_77 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h4d == _T_37[9:0]) begin
        image_0_77 <= io_pixelVal_in_0_7;
      end else if (10'h4d == _T_34[9:0]) begin
        image_0_77 <= io_pixelVal_in_0_6;
      end else if (10'h4d == _T_31[9:0]) begin
        image_0_77 <= io_pixelVal_in_0_5;
      end else if (10'h4d == _T_28[9:0]) begin
        image_0_77 <= io_pixelVal_in_0_4;
      end else if (10'h4d == _T_25[9:0]) begin
        image_0_77 <= io_pixelVal_in_0_3;
      end else if (10'h4d == _T_22[9:0]) begin
        image_0_77 <= io_pixelVal_in_0_2;
      end else if (10'h4d == _T_19[9:0]) begin
        image_0_77 <= io_pixelVal_in_0_1;
      end else if (10'h4d == _T_15[9:0]) begin
        image_0_77 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_78 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h4e == _T_37[9:0]) begin
        image_0_78 <= io_pixelVal_in_0_7;
      end else if (10'h4e == _T_34[9:0]) begin
        image_0_78 <= io_pixelVal_in_0_6;
      end else if (10'h4e == _T_31[9:0]) begin
        image_0_78 <= io_pixelVal_in_0_5;
      end else if (10'h4e == _T_28[9:0]) begin
        image_0_78 <= io_pixelVal_in_0_4;
      end else if (10'h4e == _T_25[9:0]) begin
        image_0_78 <= io_pixelVal_in_0_3;
      end else if (10'h4e == _T_22[9:0]) begin
        image_0_78 <= io_pixelVal_in_0_2;
      end else if (10'h4e == _T_19[9:0]) begin
        image_0_78 <= io_pixelVal_in_0_1;
      end else if (10'h4e == _T_15[9:0]) begin
        image_0_78 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_79 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h4f == _T_37[9:0]) begin
        image_0_79 <= io_pixelVal_in_0_7;
      end else if (10'h4f == _T_34[9:0]) begin
        image_0_79 <= io_pixelVal_in_0_6;
      end else if (10'h4f == _T_31[9:0]) begin
        image_0_79 <= io_pixelVal_in_0_5;
      end else if (10'h4f == _T_28[9:0]) begin
        image_0_79 <= io_pixelVal_in_0_4;
      end else if (10'h4f == _T_25[9:0]) begin
        image_0_79 <= io_pixelVal_in_0_3;
      end else if (10'h4f == _T_22[9:0]) begin
        image_0_79 <= io_pixelVal_in_0_2;
      end else if (10'h4f == _T_19[9:0]) begin
        image_0_79 <= io_pixelVal_in_0_1;
      end else if (10'h4f == _T_15[9:0]) begin
        image_0_79 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_80 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h50 == _T_37[9:0]) begin
        image_0_80 <= io_pixelVal_in_0_7;
      end else if (10'h50 == _T_34[9:0]) begin
        image_0_80 <= io_pixelVal_in_0_6;
      end else if (10'h50 == _T_31[9:0]) begin
        image_0_80 <= io_pixelVal_in_0_5;
      end else if (10'h50 == _T_28[9:0]) begin
        image_0_80 <= io_pixelVal_in_0_4;
      end else if (10'h50 == _T_25[9:0]) begin
        image_0_80 <= io_pixelVal_in_0_3;
      end else if (10'h50 == _T_22[9:0]) begin
        image_0_80 <= io_pixelVal_in_0_2;
      end else if (10'h50 == _T_19[9:0]) begin
        image_0_80 <= io_pixelVal_in_0_1;
      end else if (10'h50 == _T_15[9:0]) begin
        image_0_80 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_81 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h51 == _T_37[9:0]) begin
        image_0_81 <= io_pixelVal_in_0_7;
      end else if (10'h51 == _T_34[9:0]) begin
        image_0_81 <= io_pixelVal_in_0_6;
      end else if (10'h51 == _T_31[9:0]) begin
        image_0_81 <= io_pixelVal_in_0_5;
      end else if (10'h51 == _T_28[9:0]) begin
        image_0_81 <= io_pixelVal_in_0_4;
      end else if (10'h51 == _T_25[9:0]) begin
        image_0_81 <= io_pixelVal_in_0_3;
      end else if (10'h51 == _T_22[9:0]) begin
        image_0_81 <= io_pixelVal_in_0_2;
      end else if (10'h51 == _T_19[9:0]) begin
        image_0_81 <= io_pixelVal_in_0_1;
      end else if (10'h51 == _T_15[9:0]) begin
        image_0_81 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_82 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h52 == _T_37[9:0]) begin
        image_0_82 <= io_pixelVal_in_0_7;
      end else if (10'h52 == _T_34[9:0]) begin
        image_0_82 <= io_pixelVal_in_0_6;
      end else if (10'h52 == _T_31[9:0]) begin
        image_0_82 <= io_pixelVal_in_0_5;
      end else if (10'h52 == _T_28[9:0]) begin
        image_0_82 <= io_pixelVal_in_0_4;
      end else if (10'h52 == _T_25[9:0]) begin
        image_0_82 <= io_pixelVal_in_0_3;
      end else if (10'h52 == _T_22[9:0]) begin
        image_0_82 <= io_pixelVal_in_0_2;
      end else if (10'h52 == _T_19[9:0]) begin
        image_0_82 <= io_pixelVal_in_0_1;
      end else if (10'h52 == _T_15[9:0]) begin
        image_0_82 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_83 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h53 == _T_37[9:0]) begin
        image_0_83 <= io_pixelVal_in_0_7;
      end else if (10'h53 == _T_34[9:0]) begin
        image_0_83 <= io_pixelVal_in_0_6;
      end else if (10'h53 == _T_31[9:0]) begin
        image_0_83 <= io_pixelVal_in_0_5;
      end else if (10'h53 == _T_28[9:0]) begin
        image_0_83 <= io_pixelVal_in_0_4;
      end else if (10'h53 == _T_25[9:0]) begin
        image_0_83 <= io_pixelVal_in_0_3;
      end else if (10'h53 == _T_22[9:0]) begin
        image_0_83 <= io_pixelVal_in_0_2;
      end else if (10'h53 == _T_19[9:0]) begin
        image_0_83 <= io_pixelVal_in_0_1;
      end else if (10'h53 == _T_15[9:0]) begin
        image_0_83 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_84 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h54 == _T_37[9:0]) begin
        image_0_84 <= io_pixelVal_in_0_7;
      end else if (10'h54 == _T_34[9:0]) begin
        image_0_84 <= io_pixelVal_in_0_6;
      end else if (10'h54 == _T_31[9:0]) begin
        image_0_84 <= io_pixelVal_in_0_5;
      end else if (10'h54 == _T_28[9:0]) begin
        image_0_84 <= io_pixelVal_in_0_4;
      end else if (10'h54 == _T_25[9:0]) begin
        image_0_84 <= io_pixelVal_in_0_3;
      end else if (10'h54 == _T_22[9:0]) begin
        image_0_84 <= io_pixelVal_in_0_2;
      end else if (10'h54 == _T_19[9:0]) begin
        image_0_84 <= io_pixelVal_in_0_1;
      end else if (10'h54 == _T_15[9:0]) begin
        image_0_84 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_85 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h55 == _T_37[9:0]) begin
        image_0_85 <= io_pixelVal_in_0_7;
      end else if (10'h55 == _T_34[9:0]) begin
        image_0_85 <= io_pixelVal_in_0_6;
      end else if (10'h55 == _T_31[9:0]) begin
        image_0_85 <= io_pixelVal_in_0_5;
      end else if (10'h55 == _T_28[9:0]) begin
        image_0_85 <= io_pixelVal_in_0_4;
      end else if (10'h55 == _T_25[9:0]) begin
        image_0_85 <= io_pixelVal_in_0_3;
      end else if (10'h55 == _T_22[9:0]) begin
        image_0_85 <= io_pixelVal_in_0_2;
      end else if (10'h55 == _T_19[9:0]) begin
        image_0_85 <= io_pixelVal_in_0_1;
      end else if (10'h55 == _T_15[9:0]) begin
        image_0_85 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_86 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h56 == _T_37[9:0]) begin
        image_0_86 <= io_pixelVal_in_0_7;
      end else if (10'h56 == _T_34[9:0]) begin
        image_0_86 <= io_pixelVal_in_0_6;
      end else if (10'h56 == _T_31[9:0]) begin
        image_0_86 <= io_pixelVal_in_0_5;
      end else if (10'h56 == _T_28[9:0]) begin
        image_0_86 <= io_pixelVal_in_0_4;
      end else if (10'h56 == _T_25[9:0]) begin
        image_0_86 <= io_pixelVal_in_0_3;
      end else if (10'h56 == _T_22[9:0]) begin
        image_0_86 <= io_pixelVal_in_0_2;
      end else if (10'h56 == _T_19[9:0]) begin
        image_0_86 <= io_pixelVal_in_0_1;
      end else if (10'h56 == _T_15[9:0]) begin
        image_0_86 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_87 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h57 == _T_37[9:0]) begin
        image_0_87 <= io_pixelVal_in_0_7;
      end else if (10'h57 == _T_34[9:0]) begin
        image_0_87 <= io_pixelVal_in_0_6;
      end else if (10'h57 == _T_31[9:0]) begin
        image_0_87 <= io_pixelVal_in_0_5;
      end else if (10'h57 == _T_28[9:0]) begin
        image_0_87 <= io_pixelVal_in_0_4;
      end else if (10'h57 == _T_25[9:0]) begin
        image_0_87 <= io_pixelVal_in_0_3;
      end else if (10'h57 == _T_22[9:0]) begin
        image_0_87 <= io_pixelVal_in_0_2;
      end else if (10'h57 == _T_19[9:0]) begin
        image_0_87 <= io_pixelVal_in_0_1;
      end else if (10'h57 == _T_15[9:0]) begin
        image_0_87 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_88 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h58 == _T_37[9:0]) begin
        image_0_88 <= io_pixelVal_in_0_7;
      end else if (10'h58 == _T_34[9:0]) begin
        image_0_88 <= io_pixelVal_in_0_6;
      end else if (10'h58 == _T_31[9:0]) begin
        image_0_88 <= io_pixelVal_in_0_5;
      end else if (10'h58 == _T_28[9:0]) begin
        image_0_88 <= io_pixelVal_in_0_4;
      end else if (10'h58 == _T_25[9:0]) begin
        image_0_88 <= io_pixelVal_in_0_3;
      end else if (10'h58 == _T_22[9:0]) begin
        image_0_88 <= io_pixelVal_in_0_2;
      end else if (10'h58 == _T_19[9:0]) begin
        image_0_88 <= io_pixelVal_in_0_1;
      end else if (10'h58 == _T_15[9:0]) begin
        image_0_88 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_89 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h59 == _T_37[9:0]) begin
        image_0_89 <= io_pixelVal_in_0_7;
      end else if (10'h59 == _T_34[9:0]) begin
        image_0_89 <= io_pixelVal_in_0_6;
      end else if (10'h59 == _T_31[9:0]) begin
        image_0_89 <= io_pixelVal_in_0_5;
      end else if (10'h59 == _T_28[9:0]) begin
        image_0_89 <= io_pixelVal_in_0_4;
      end else if (10'h59 == _T_25[9:0]) begin
        image_0_89 <= io_pixelVal_in_0_3;
      end else if (10'h59 == _T_22[9:0]) begin
        image_0_89 <= io_pixelVal_in_0_2;
      end else if (10'h59 == _T_19[9:0]) begin
        image_0_89 <= io_pixelVal_in_0_1;
      end else if (10'h59 == _T_15[9:0]) begin
        image_0_89 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_90 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h5a == _T_37[9:0]) begin
        image_0_90 <= io_pixelVal_in_0_7;
      end else if (10'h5a == _T_34[9:0]) begin
        image_0_90 <= io_pixelVal_in_0_6;
      end else if (10'h5a == _T_31[9:0]) begin
        image_0_90 <= io_pixelVal_in_0_5;
      end else if (10'h5a == _T_28[9:0]) begin
        image_0_90 <= io_pixelVal_in_0_4;
      end else if (10'h5a == _T_25[9:0]) begin
        image_0_90 <= io_pixelVal_in_0_3;
      end else if (10'h5a == _T_22[9:0]) begin
        image_0_90 <= io_pixelVal_in_0_2;
      end else if (10'h5a == _T_19[9:0]) begin
        image_0_90 <= io_pixelVal_in_0_1;
      end else if (10'h5a == _T_15[9:0]) begin
        image_0_90 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_91 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h5b == _T_37[9:0]) begin
        image_0_91 <= io_pixelVal_in_0_7;
      end else if (10'h5b == _T_34[9:0]) begin
        image_0_91 <= io_pixelVal_in_0_6;
      end else if (10'h5b == _T_31[9:0]) begin
        image_0_91 <= io_pixelVal_in_0_5;
      end else if (10'h5b == _T_28[9:0]) begin
        image_0_91 <= io_pixelVal_in_0_4;
      end else if (10'h5b == _T_25[9:0]) begin
        image_0_91 <= io_pixelVal_in_0_3;
      end else if (10'h5b == _T_22[9:0]) begin
        image_0_91 <= io_pixelVal_in_0_2;
      end else if (10'h5b == _T_19[9:0]) begin
        image_0_91 <= io_pixelVal_in_0_1;
      end else if (10'h5b == _T_15[9:0]) begin
        image_0_91 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_92 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h5c == _T_37[9:0]) begin
        image_0_92 <= io_pixelVal_in_0_7;
      end else if (10'h5c == _T_34[9:0]) begin
        image_0_92 <= io_pixelVal_in_0_6;
      end else if (10'h5c == _T_31[9:0]) begin
        image_0_92 <= io_pixelVal_in_0_5;
      end else if (10'h5c == _T_28[9:0]) begin
        image_0_92 <= io_pixelVal_in_0_4;
      end else if (10'h5c == _T_25[9:0]) begin
        image_0_92 <= io_pixelVal_in_0_3;
      end else if (10'h5c == _T_22[9:0]) begin
        image_0_92 <= io_pixelVal_in_0_2;
      end else if (10'h5c == _T_19[9:0]) begin
        image_0_92 <= io_pixelVal_in_0_1;
      end else if (10'h5c == _T_15[9:0]) begin
        image_0_92 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_93 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h5d == _T_37[9:0]) begin
        image_0_93 <= io_pixelVal_in_0_7;
      end else if (10'h5d == _T_34[9:0]) begin
        image_0_93 <= io_pixelVal_in_0_6;
      end else if (10'h5d == _T_31[9:0]) begin
        image_0_93 <= io_pixelVal_in_0_5;
      end else if (10'h5d == _T_28[9:0]) begin
        image_0_93 <= io_pixelVal_in_0_4;
      end else if (10'h5d == _T_25[9:0]) begin
        image_0_93 <= io_pixelVal_in_0_3;
      end else if (10'h5d == _T_22[9:0]) begin
        image_0_93 <= io_pixelVal_in_0_2;
      end else if (10'h5d == _T_19[9:0]) begin
        image_0_93 <= io_pixelVal_in_0_1;
      end else if (10'h5d == _T_15[9:0]) begin
        image_0_93 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_94 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h5e == _T_37[9:0]) begin
        image_0_94 <= io_pixelVal_in_0_7;
      end else if (10'h5e == _T_34[9:0]) begin
        image_0_94 <= io_pixelVal_in_0_6;
      end else if (10'h5e == _T_31[9:0]) begin
        image_0_94 <= io_pixelVal_in_0_5;
      end else if (10'h5e == _T_28[9:0]) begin
        image_0_94 <= io_pixelVal_in_0_4;
      end else if (10'h5e == _T_25[9:0]) begin
        image_0_94 <= io_pixelVal_in_0_3;
      end else if (10'h5e == _T_22[9:0]) begin
        image_0_94 <= io_pixelVal_in_0_2;
      end else if (10'h5e == _T_19[9:0]) begin
        image_0_94 <= io_pixelVal_in_0_1;
      end else if (10'h5e == _T_15[9:0]) begin
        image_0_94 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_95 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h5f == _T_37[9:0]) begin
        image_0_95 <= io_pixelVal_in_0_7;
      end else if (10'h5f == _T_34[9:0]) begin
        image_0_95 <= io_pixelVal_in_0_6;
      end else if (10'h5f == _T_31[9:0]) begin
        image_0_95 <= io_pixelVal_in_0_5;
      end else if (10'h5f == _T_28[9:0]) begin
        image_0_95 <= io_pixelVal_in_0_4;
      end else if (10'h5f == _T_25[9:0]) begin
        image_0_95 <= io_pixelVal_in_0_3;
      end else if (10'h5f == _T_22[9:0]) begin
        image_0_95 <= io_pixelVal_in_0_2;
      end else if (10'h5f == _T_19[9:0]) begin
        image_0_95 <= io_pixelVal_in_0_1;
      end else if (10'h5f == _T_15[9:0]) begin
        image_0_95 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_96 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h60 == _T_37[9:0]) begin
        image_0_96 <= io_pixelVal_in_0_7;
      end else if (10'h60 == _T_34[9:0]) begin
        image_0_96 <= io_pixelVal_in_0_6;
      end else if (10'h60 == _T_31[9:0]) begin
        image_0_96 <= io_pixelVal_in_0_5;
      end else if (10'h60 == _T_28[9:0]) begin
        image_0_96 <= io_pixelVal_in_0_4;
      end else if (10'h60 == _T_25[9:0]) begin
        image_0_96 <= io_pixelVal_in_0_3;
      end else if (10'h60 == _T_22[9:0]) begin
        image_0_96 <= io_pixelVal_in_0_2;
      end else if (10'h60 == _T_19[9:0]) begin
        image_0_96 <= io_pixelVal_in_0_1;
      end else if (10'h60 == _T_15[9:0]) begin
        image_0_96 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_97 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h61 == _T_37[9:0]) begin
        image_0_97 <= io_pixelVal_in_0_7;
      end else if (10'h61 == _T_34[9:0]) begin
        image_0_97 <= io_pixelVal_in_0_6;
      end else if (10'h61 == _T_31[9:0]) begin
        image_0_97 <= io_pixelVal_in_0_5;
      end else if (10'h61 == _T_28[9:0]) begin
        image_0_97 <= io_pixelVal_in_0_4;
      end else if (10'h61 == _T_25[9:0]) begin
        image_0_97 <= io_pixelVal_in_0_3;
      end else if (10'h61 == _T_22[9:0]) begin
        image_0_97 <= io_pixelVal_in_0_2;
      end else if (10'h61 == _T_19[9:0]) begin
        image_0_97 <= io_pixelVal_in_0_1;
      end else if (10'h61 == _T_15[9:0]) begin
        image_0_97 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_98 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h62 == _T_37[9:0]) begin
        image_0_98 <= io_pixelVal_in_0_7;
      end else if (10'h62 == _T_34[9:0]) begin
        image_0_98 <= io_pixelVal_in_0_6;
      end else if (10'h62 == _T_31[9:0]) begin
        image_0_98 <= io_pixelVal_in_0_5;
      end else if (10'h62 == _T_28[9:0]) begin
        image_0_98 <= io_pixelVal_in_0_4;
      end else if (10'h62 == _T_25[9:0]) begin
        image_0_98 <= io_pixelVal_in_0_3;
      end else if (10'h62 == _T_22[9:0]) begin
        image_0_98 <= io_pixelVal_in_0_2;
      end else if (10'h62 == _T_19[9:0]) begin
        image_0_98 <= io_pixelVal_in_0_1;
      end else if (10'h62 == _T_15[9:0]) begin
        image_0_98 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_99 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h63 == _T_37[9:0]) begin
        image_0_99 <= io_pixelVal_in_0_7;
      end else if (10'h63 == _T_34[9:0]) begin
        image_0_99 <= io_pixelVal_in_0_6;
      end else if (10'h63 == _T_31[9:0]) begin
        image_0_99 <= io_pixelVal_in_0_5;
      end else if (10'h63 == _T_28[9:0]) begin
        image_0_99 <= io_pixelVal_in_0_4;
      end else if (10'h63 == _T_25[9:0]) begin
        image_0_99 <= io_pixelVal_in_0_3;
      end else if (10'h63 == _T_22[9:0]) begin
        image_0_99 <= io_pixelVal_in_0_2;
      end else if (10'h63 == _T_19[9:0]) begin
        image_0_99 <= io_pixelVal_in_0_1;
      end else if (10'h63 == _T_15[9:0]) begin
        image_0_99 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_100 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h64 == _T_37[9:0]) begin
        image_0_100 <= io_pixelVal_in_0_7;
      end else if (10'h64 == _T_34[9:0]) begin
        image_0_100 <= io_pixelVal_in_0_6;
      end else if (10'h64 == _T_31[9:0]) begin
        image_0_100 <= io_pixelVal_in_0_5;
      end else if (10'h64 == _T_28[9:0]) begin
        image_0_100 <= io_pixelVal_in_0_4;
      end else if (10'h64 == _T_25[9:0]) begin
        image_0_100 <= io_pixelVal_in_0_3;
      end else if (10'h64 == _T_22[9:0]) begin
        image_0_100 <= io_pixelVal_in_0_2;
      end else if (10'h64 == _T_19[9:0]) begin
        image_0_100 <= io_pixelVal_in_0_1;
      end else if (10'h64 == _T_15[9:0]) begin
        image_0_100 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_101 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h65 == _T_37[9:0]) begin
        image_0_101 <= io_pixelVal_in_0_7;
      end else if (10'h65 == _T_34[9:0]) begin
        image_0_101 <= io_pixelVal_in_0_6;
      end else if (10'h65 == _T_31[9:0]) begin
        image_0_101 <= io_pixelVal_in_0_5;
      end else if (10'h65 == _T_28[9:0]) begin
        image_0_101 <= io_pixelVal_in_0_4;
      end else if (10'h65 == _T_25[9:0]) begin
        image_0_101 <= io_pixelVal_in_0_3;
      end else if (10'h65 == _T_22[9:0]) begin
        image_0_101 <= io_pixelVal_in_0_2;
      end else if (10'h65 == _T_19[9:0]) begin
        image_0_101 <= io_pixelVal_in_0_1;
      end else if (10'h65 == _T_15[9:0]) begin
        image_0_101 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_102 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h66 == _T_37[9:0]) begin
        image_0_102 <= io_pixelVal_in_0_7;
      end else if (10'h66 == _T_34[9:0]) begin
        image_0_102 <= io_pixelVal_in_0_6;
      end else if (10'h66 == _T_31[9:0]) begin
        image_0_102 <= io_pixelVal_in_0_5;
      end else if (10'h66 == _T_28[9:0]) begin
        image_0_102 <= io_pixelVal_in_0_4;
      end else if (10'h66 == _T_25[9:0]) begin
        image_0_102 <= io_pixelVal_in_0_3;
      end else if (10'h66 == _T_22[9:0]) begin
        image_0_102 <= io_pixelVal_in_0_2;
      end else if (10'h66 == _T_19[9:0]) begin
        image_0_102 <= io_pixelVal_in_0_1;
      end else if (10'h66 == _T_15[9:0]) begin
        image_0_102 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_103 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h67 == _T_37[9:0]) begin
        image_0_103 <= io_pixelVal_in_0_7;
      end else if (10'h67 == _T_34[9:0]) begin
        image_0_103 <= io_pixelVal_in_0_6;
      end else if (10'h67 == _T_31[9:0]) begin
        image_0_103 <= io_pixelVal_in_0_5;
      end else if (10'h67 == _T_28[9:0]) begin
        image_0_103 <= io_pixelVal_in_0_4;
      end else if (10'h67 == _T_25[9:0]) begin
        image_0_103 <= io_pixelVal_in_0_3;
      end else if (10'h67 == _T_22[9:0]) begin
        image_0_103 <= io_pixelVal_in_0_2;
      end else if (10'h67 == _T_19[9:0]) begin
        image_0_103 <= io_pixelVal_in_0_1;
      end else if (10'h67 == _T_15[9:0]) begin
        image_0_103 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_104 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h68 == _T_37[9:0]) begin
        image_0_104 <= io_pixelVal_in_0_7;
      end else if (10'h68 == _T_34[9:0]) begin
        image_0_104 <= io_pixelVal_in_0_6;
      end else if (10'h68 == _T_31[9:0]) begin
        image_0_104 <= io_pixelVal_in_0_5;
      end else if (10'h68 == _T_28[9:0]) begin
        image_0_104 <= io_pixelVal_in_0_4;
      end else if (10'h68 == _T_25[9:0]) begin
        image_0_104 <= io_pixelVal_in_0_3;
      end else if (10'h68 == _T_22[9:0]) begin
        image_0_104 <= io_pixelVal_in_0_2;
      end else if (10'h68 == _T_19[9:0]) begin
        image_0_104 <= io_pixelVal_in_0_1;
      end else if (10'h68 == _T_15[9:0]) begin
        image_0_104 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_105 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h69 == _T_37[9:0]) begin
        image_0_105 <= io_pixelVal_in_0_7;
      end else if (10'h69 == _T_34[9:0]) begin
        image_0_105 <= io_pixelVal_in_0_6;
      end else if (10'h69 == _T_31[9:0]) begin
        image_0_105 <= io_pixelVal_in_0_5;
      end else if (10'h69 == _T_28[9:0]) begin
        image_0_105 <= io_pixelVal_in_0_4;
      end else if (10'h69 == _T_25[9:0]) begin
        image_0_105 <= io_pixelVal_in_0_3;
      end else if (10'h69 == _T_22[9:0]) begin
        image_0_105 <= io_pixelVal_in_0_2;
      end else if (10'h69 == _T_19[9:0]) begin
        image_0_105 <= io_pixelVal_in_0_1;
      end else if (10'h69 == _T_15[9:0]) begin
        image_0_105 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_106 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h6a == _T_37[9:0]) begin
        image_0_106 <= io_pixelVal_in_0_7;
      end else if (10'h6a == _T_34[9:0]) begin
        image_0_106 <= io_pixelVal_in_0_6;
      end else if (10'h6a == _T_31[9:0]) begin
        image_0_106 <= io_pixelVal_in_0_5;
      end else if (10'h6a == _T_28[9:0]) begin
        image_0_106 <= io_pixelVal_in_0_4;
      end else if (10'h6a == _T_25[9:0]) begin
        image_0_106 <= io_pixelVal_in_0_3;
      end else if (10'h6a == _T_22[9:0]) begin
        image_0_106 <= io_pixelVal_in_0_2;
      end else if (10'h6a == _T_19[9:0]) begin
        image_0_106 <= io_pixelVal_in_0_1;
      end else if (10'h6a == _T_15[9:0]) begin
        image_0_106 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_107 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h6b == _T_37[9:0]) begin
        image_0_107 <= io_pixelVal_in_0_7;
      end else if (10'h6b == _T_34[9:0]) begin
        image_0_107 <= io_pixelVal_in_0_6;
      end else if (10'h6b == _T_31[9:0]) begin
        image_0_107 <= io_pixelVal_in_0_5;
      end else if (10'h6b == _T_28[9:0]) begin
        image_0_107 <= io_pixelVal_in_0_4;
      end else if (10'h6b == _T_25[9:0]) begin
        image_0_107 <= io_pixelVal_in_0_3;
      end else if (10'h6b == _T_22[9:0]) begin
        image_0_107 <= io_pixelVal_in_0_2;
      end else if (10'h6b == _T_19[9:0]) begin
        image_0_107 <= io_pixelVal_in_0_1;
      end else if (10'h6b == _T_15[9:0]) begin
        image_0_107 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_108 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h6c == _T_37[9:0]) begin
        image_0_108 <= io_pixelVal_in_0_7;
      end else if (10'h6c == _T_34[9:0]) begin
        image_0_108 <= io_pixelVal_in_0_6;
      end else if (10'h6c == _T_31[9:0]) begin
        image_0_108 <= io_pixelVal_in_0_5;
      end else if (10'h6c == _T_28[9:0]) begin
        image_0_108 <= io_pixelVal_in_0_4;
      end else if (10'h6c == _T_25[9:0]) begin
        image_0_108 <= io_pixelVal_in_0_3;
      end else if (10'h6c == _T_22[9:0]) begin
        image_0_108 <= io_pixelVal_in_0_2;
      end else if (10'h6c == _T_19[9:0]) begin
        image_0_108 <= io_pixelVal_in_0_1;
      end else if (10'h6c == _T_15[9:0]) begin
        image_0_108 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_109 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h6d == _T_37[9:0]) begin
        image_0_109 <= io_pixelVal_in_0_7;
      end else if (10'h6d == _T_34[9:0]) begin
        image_0_109 <= io_pixelVal_in_0_6;
      end else if (10'h6d == _T_31[9:0]) begin
        image_0_109 <= io_pixelVal_in_0_5;
      end else if (10'h6d == _T_28[9:0]) begin
        image_0_109 <= io_pixelVal_in_0_4;
      end else if (10'h6d == _T_25[9:0]) begin
        image_0_109 <= io_pixelVal_in_0_3;
      end else if (10'h6d == _T_22[9:0]) begin
        image_0_109 <= io_pixelVal_in_0_2;
      end else if (10'h6d == _T_19[9:0]) begin
        image_0_109 <= io_pixelVal_in_0_1;
      end else if (10'h6d == _T_15[9:0]) begin
        image_0_109 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_110 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h6e == _T_37[9:0]) begin
        image_0_110 <= io_pixelVal_in_0_7;
      end else if (10'h6e == _T_34[9:0]) begin
        image_0_110 <= io_pixelVal_in_0_6;
      end else if (10'h6e == _T_31[9:0]) begin
        image_0_110 <= io_pixelVal_in_0_5;
      end else if (10'h6e == _T_28[9:0]) begin
        image_0_110 <= io_pixelVal_in_0_4;
      end else if (10'h6e == _T_25[9:0]) begin
        image_0_110 <= io_pixelVal_in_0_3;
      end else if (10'h6e == _T_22[9:0]) begin
        image_0_110 <= io_pixelVal_in_0_2;
      end else if (10'h6e == _T_19[9:0]) begin
        image_0_110 <= io_pixelVal_in_0_1;
      end else if (10'h6e == _T_15[9:0]) begin
        image_0_110 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_111 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h6f == _T_37[9:0]) begin
        image_0_111 <= io_pixelVal_in_0_7;
      end else if (10'h6f == _T_34[9:0]) begin
        image_0_111 <= io_pixelVal_in_0_6;
      end else if (10'h6f == _T_31[9:0]) begin
        image_0_111 <= io_pixelVal_in_0_5;
      end else if (10'h6f == _T_28[9:0]) begin
        image_0_111 <= io_pixelVal_in_0_4;
      end else if (10'h6f == _T_25[9:0]) begin
        image_0_111 <= io_pixelVal_in_0_3;
      end else if (10'h6f == _T_22[9:0]) begin
        image_0_111 <= io_pixelVal_in_0_2;
      end else if (10'h6f == _T_19[9:0]) begin
        image_0_111 <= io_pixelVal_in_0_1;
      end else if (10'h6f == _T_15[9:0]) begin
        image_0_111 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_112 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h70 == _T_37[9:0]) begin
        image_0_112 <= io_pixelVal_in_0_7;
      end else if (10'h70 == _T_34[9:0]) begin
        image_0_112 <= io_pixelVal_in_0_6;
      end else if (10'h70 == _T_31[9:0]) begin
        image_0_112 <= io_pixelVal_in_0_5;
      end else if (10'h70 == _T_28[9:0]) begin
        image_0_112 <= io_pixelVal_in_0_4;
      end else if (10'h70 == _T_25[9:0]) begin
        image_0_112 <= io_pixelVal_in_0_3;
      end else if (10'h70 == _T_22[9:0]) begin
        image_0_112 <= io_pixelVal_in_0_2;
      end else if (10'h70 == _T_19[9:0]) begin
        image_0_112 <= io_pixelVal_in_0_1;
      end else if (10'h70 == _T_15[9:0]) begin
        image_0_112 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_113 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h71 == _T_37[9:0]) begin
        image_0_113 <= io_pixelVal_in_0_7;
      end else if (10'h71 == _T_34[9:0]) begin
        image_0_113 <= io_pixelVal_in_0_6;
      end else if (10'h71 == _T_31[9:0]) begin
        image_0_113 <= io_pixelVal_in_0_5;
      end else if (10'h71 == _T_28[9:0]) begin
        image_0_113 <= io_pixelVal_in_0_4;
      end else if (10'h71 == _T_25[9:0]) begin
        image_0_113 <= io_pixelVal_in_0_3;
      end else if (10'h71 == _T_22[9:0]) begin
        image_0_113 <= io_pixelVal_in_0_2;
      end else if (10'h71 == _T_19[9:0]) begin
        image_0_113 <= io_pixelVal_in_0_1;
      end else if (10'h71 == _T_15[9:0]) begin
        image_0_113 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_114 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h72 == _T_37[9:0]) begin
        image_0_114 <= io_pixelVal_in_0_7;
      end else if (10'h72 == _T_34[9:0]) begin
        image_0_114 <= io_pixelVal_in_0_6;
      end else if (10'h72 == _T_31[9:0]) begin
        image_0_114 <= io_pixelVal_in_0_5;
      end else if (10'h72 == _T_28[9:0]) begin
        image_0_114 <= io_pixelVal_in_0_4;
      end else if (10'h72 == _T_25[9:0]) begin
        image_0_114 <= io_pixelVal_in_0_3;
      end else if (10'h72 == _T_22[9:0]) begin
        image_0_114 <= io_pixelVal_in_0_2;
      end else if (10'h72 == _T_19[9:0]) begin
        image_0_114 <= io_pixelVal_in_0_1;
      end else if (10'h72 == _T_15[9:0]) begin
        image_0_114 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_115 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h73 == _T_37[9:0]) begin
        image_0_115 <= io_pixelVal_in_0_7;
      end else if (10'h73 == _T_34[9:0]) begin
        image_0_115 <= io_pixelVal_in_0_6;
      end else if (10'h73 == _T_31[9:0]) begin
        image_0_115 <= io_pixelVal_in_0_5;
      end else if (10'h73 == _T_28[9:0]) begin
        image_0_115 <= io_pixelVal_in_0_4;
      end else if (10'h73 == _T_25[9:0]) begin
        image_0_115 <= io_pixelVal_in_0_3;
      end else if (10'h73 == _T_22[9:0]) begin
        image_0_115 <= io_pixelVal_in_0_2;
      end else if (10'h73 == _T_19[9:0]) begin
        image_0_115 <= io_pixelVal_in_0_1;
      end else if (10'h73 == _T_15[9:0]) begin
        image_0_115 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_116 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h74 == _T_37[9:0]) begin
        image_0_116 <= io_pixelVal_in_0_7;
      end else if (10'h74 == _T_34[9:0]) begin
        image_0_116 <= io_pixelVal_in_0_6;
      end else if (10'h74 == _T_31[9:0]) begin
        image_0_116 <= io_pixelVal_in_0_5;
      end else if (10'h74 == _T_28[9:0]) begin
        image_0_116 <= io_pixelVal_in_0_4;
      end else if (10'h74 == _T_25[9:0]) begin
        image_0_116 <= io_pixelVal_in_0_3;
      end else if (10'h74 == _T_22[9:0]) begin
        image_0_116 <= io_pixelVal_in_0_2;
      end else if (10'h74 == _T_19[9:0]) begin
        image_0_116 <= io_pixelVal_in_0_1;
      end else if (10'h74 == _T_15[9:0]) begin
        image_0_116 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_117 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h75 == _T_37[9:0]) begin
        image_0_117 <= io_pixelVal_in_0_7;
      end else if (10'h75 == _T_34[9:0]) begin
        image_0_117 <= io_pixelVal_in_0_6;
      end else if (10'h75 == _T_31[9:0]) begin
        image_0_117 <= io_pixelVal_in_0_5;
      end else if (10'h75 == _T_28[9:0]) begin
        image_0_117 <= io_pixelVal_in_0_4;
      end else if (10'h75 == _T_25[9:0]) begin
        image_0_117 <= io_pixelVal_in_0_3;
      end else if (10'h75 == _T_22[9:0]) begin
        image_0_117 <= io_pixelVal_in_0_2;
      end else if (10'h75 == _T_19[9:0]) begin
        image_0_117 <= io_pixelVal_in_0_1;
      end else if (10'h75 == _T_15[9:0]) begin
        image_0_117 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_118 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h76 == _T_37[9:0]) begin
        image_0_118 <= io_pixelVal_in_0_7;
      end else if (10'h76 == _T_34[9:0]) begin
        image_0_118 <= io_pixelVal_in_0_6;
      end else if (10'h76 == _T_31[9:0]) begin
        image_0_118 <= io_pixelVal_in_0_5;
      end else if (10'h76 == _T_28[9:0]) begin
        image_0_118 <= io_pixelVal_in_0_4;
      end else if (10'h76 == _T_25[9:0]) begin
        image_0_118 <= io_pixelVal_in_0_3;
      end else if (10'h76 == _T_22[9:0]) begin
        image_0_118 <= io_pixelVal_in_0_2;
      end else if (10'h76 == _T_19[9:0]) begin
        image_0_118 <= io_pixelVal_in_0_1;
      end else if (10'h76 == _T_15[9:0]) begin
        image_0_118 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_119 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h77 == _T_37[9:0]) begin
        image_0_119 <= io_pixelVal_in_0_7;
      end else if (10'h77 == _T_34[9:0]) begin
        image_0_119 <= io_pixelVal_in_0_6;
      end else if (10'h77 == _T_31[9:0]) begin
        image_0_119 <= io_pixelVal_in_0_5;
      end else if (10'h77 == _T_28[9:0]) begin
        image_0_119 <= io_pixelVal_in_0_4;
      end else if (10'h77 == _T_25[9:0]) begin
        image_0_119 <= io_pixelVal_in_0_3;
      end else if (10'h77 == _T_22[9:0]) begin
        image_0_119 <= io_pixelVal_in_0_2;
      end else if (10'h77 == _T_19[9:0]) begin
        image_0_119 <= io_pixelVal_in_0_1;
      end else if (10'h77 == _T_15[9:0]) begin
        image_0_119 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_120 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h78 == _T_37[9:0]) begin
        image_0_120 <= io_pixelVal_in_0_7;
      end else if (10'h78 == _T_34[9:0]) begin
        image_0_120 <= io_pixelVal_in_0_6;
      end else if (10'h78 == _T_31[9:0]) begin
        image_0_120 <= io_pixelVal_in_0_5;
      end else if (10'h78 == _T_28[9:0]) begin
        image_0_120 <= io_pixelVal_in_0_4;
      end else if (10'h78 == _T_25[9:0]) begin
        image_0_120 <= io_pixelVal_in_0_3;
      end else if (10'h78 == _T_22[9:0]) begin
        image_0_120 <= io_pixelVal_in_0_2;
      end else if (10'h78 == _T_19[9:0]) begin
        image_0_120 <= io_pixelVal_in_0_1;
      end else if (10'h78 == _T_15[9:0]) begin
        image_0_120 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_121 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h79 == _T_37[9:0]) begin
        image_0_121 <= io_pixelVal_in_0_7;
      end else if (10'h79 == _T_34[9:0]) begin
        image_0_121 <= io_pixelVal_in_0_6;
      end else if (10'h79 == _T_31[9:0]) begin
        image_0_121 <= io_pixelVal_in_0_5;
      end else if (10'h79 == _T_28[9:0]) begin
        image_0_121 <= io_pixelVal_in_0_4;
      end else if (10'h79 == _T_25[9:0]) begin
        image_0_121 <= io_pixelVal_in_0_3;
      end else if (10'h79 == _T_22[9:0]) begin
        image_0_121 <= io_pixelVal_in_0_2;
      end else if (10'h79 == _T_19[9:0]) begin
        image_0_121 <= io_pixelVal_in_0_1;
      end else if (10'h79 == _T_15[9:0]) begin
        image_0_121 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_122 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h7a == _T_37[9:0]) begin
        image_0_122 <= io_pixelVal_in_0_7;
      end else if (10'h7a == _T_34[9:0]) begin
        image_0_122 <= io_pixelVal_in_0_6;
      end else if (10'h7a == _T_31[9:0]) begin
        image_0_122 <= io_pixelVal_in_0_5;
      end else if (10'h7a == _T_28[9:0]) begin
        image_0_122 <= io_pixelVal_in_0_4;
      end else if (10'h7a == _T_25[9:0]) begin
        image_0_122 <= io_pixelVal_in_0_3;
      end else if (10'h7a == _T_22[9:0]) begin
        image_0_122 <= io_pixelVal_in_0_2;
      end else if (10'h7a == _T_19[9:0]) begin
        image_0_122 <= io_pixelVal_in_0_1;
      end else if (10'h7a == _T_15[9:0]) begin
        image_0_122 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_123 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h7b == _T_37[9:0]) begin
        image_0_123 <= io_pixelVal_in_0_7;
      end else if (10'h7b == _T_34[9:0]) begin
        image_0_123 <= io_pixelVal_in_0_6;
      end else if (10'h7b == _T_31[9:0]) begin
        image_0_123 <= io_pixelVal_in_0_5;
      end else if (10'h7b == _T_28[9:0]) begin
        image_0_123 <= io_pixelVal_in_0_4;
      end else if (10'h7b == _T_25[9:0]) begin
        image_0_123 <= io_pixelVal_in_0_3;
      end else if (10'h7b == _T_22[9:0]) begin
        image_0_123 <= io_pixelVal_in_0_2;
      end else if (10'h7b == _T_19[9:0]) begin
        image_0_123 <= io_pixelVal_in_0_1;
      end else if (10'h7b == _T_15[9:0]) begin
        image_0_123 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_124 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h7c == _T_37[9:0]) begin
        image_0_124 <= io_pixelVal_in_0_7;
      end else if (10'h7c == _T_34[9:0]) begin
        image_0_124 <= io_pixelVal_in_0_6;
      end else if (10'h7c == _T_31[9:0]) begin
        image_0_124 <= io_pixelVal_in_0_5;
      end else if (10'h7c == _T_28[9:0]) begin
        image_0_124 <= io_pixelVal_in_0_4;
      end else if (10'h7c == _T_25[9:0]) begin
        image_0_124 <= io_pixelVal_in_0_3;
      end else if (10'h7c == _T_22[9:0]) begin
        image_0_124 <= io_pixelVal_in_0_2;
      end else if (10'h7c == _T_19[9:0]) begin
        image_0_124 <= io_pixelVal_in_0_1;
      end else if (10'h7c == _T_15[9:0]) begin
        image_0_124 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_125 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h7d == _T_37[9:0]) begin
        image_0_125 <= io_pixelVal_in_0_7;
      end else if (10'h7d == _T_34[9:0]) begin
        image_0_125 <= io_pixelVal_in_0_6;
      end else if (10'h7d == _T_31[9:0]) begin
        image_0_125 <= io_pixelVal_in_0_5;
      end else if (10'h7d == _T_28[9:0]) begin
        image_0_125 <= io_pixelVal_in_0_4;
      end else if (10'h7d == _T_25[9:0]) begin
        image_0_125 <= io_pixelVal_in_0_3;
      end else if (10'h7d == _T_22[9:0]) begin
        image_0_125 <= io_pixelVal_in_0_2;
      end else if (10'h7d == _T_19[9:0]) begin
        image_0_125 <= io_pixelVal_in_0_1;
      end else if (10'h7d == _T_15[9:0]) begin
        image_0_125 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_126 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h7e == _T_37[9:0]) begin
        image_0_126 <= io_pixelVal_in_0_7;
      end else if (10'h7e == _T_34[9:0]) begin
        image_0_126 <= io_pixelVal_in_0_6;
      end else if (10'h7e == _T_31[9:0]) begin
        image_0_126 <= io_pixelVal_in_0_5;
      end else if (10'h7e == _T_28[9:0]) begin
        image_0_126 <= io_pixelVal_in_0_4;
      end else if (10'h7e == _T_25[9:0]) begin
        image_0_126 <= io_pixelVal_in_0_3;
      end else if (10'h7e == _T_22[9:0]) begin
        image_0_126 <= io_pixelVal_in_0_2;
      end else if (10'h7e == _T_19[9:0]) begin
        image_0_126 <= io_pixelVal_in_0_1;
      end else if (10'h7e == _T_15[9:0]) begin
        image_0_126 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_127 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h7f == _T_37[9:0]) begin
        image_0_127 <= io_pixelVal_in_0_7;
      end else if (10'h7f == _T_34[9:0]) begin
        image_0_127 <= io_pixelVal_in_0_6;
      end else if (10'h7f == _T_31[9:0]) begin
        image_0_127 <= io_pixelVal_in_0_5;
      end else if (10'h7f == _T_28[9:0]) begin
        image_0_127 <= io_pixelVal_in_0_4;
      end else if (10'h7f == _T_25[9:0]) begin
        image_0_127 <= io_pixelVal_in_0_3;
      end else if (10'h7f == _T_22[9:0]) begin
        image_0_127 <= io_pixelVal_in_0_2;
      end else if (10'h7f == _T_19[9:0]) begin
        image_0_127 <= io_pixelVal_in_0_1;
      end else if (10'h7f == _T_15[9:0]) begin
        image_0_127 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_128 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h80 == _T_37[9:0]) begin
        image_0_128 <= io_pixelVal_in_0_7;
      end else if (10'h80 == _T_34[9:0]) begin
        image_0_128 <= io_pixelVal_in_0_6;
      end else if (10'h80 == _T_31[9:0]) begin
        image_0_128 <= io_pixelVal_in_0_5;
      end else if (10'h80 == _T_28[9:0]) begin
        image_0_128 <= io_pixelVal_in_0_4;
      end else if (10'h80 == _T_25[9:0]) begin
        image_0_128 <= io_pixelVal_in_0_3;
      end else if (10'h80 == _T_22[9:0]) begin
        image_0_128 <= io_pixelVal_in_0_2;
      end else if (10'h80 == _T_19[9:0]) begin
        image_0_128 <= io_pixelVal_in_0_1;
      end else if (10'h80 == _T_15[9:0]) begin
        image_0_128 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_129 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h81 == _T_37[9:0]) begin
        image_0_129 <= io_pixelVal_in_0_7;
      end else if (10'h81 == _T_34[9:0]) begin
        image_0_129 <= io_pixelVal_in_0_6;
      end else if (10'h81 == _T_31[9:0]) begin
        image_0_129 <= io_pixelVal_in_0_5;
      end else if (10'h81 == _T_28[9:0]) begin
        image_0_129 <= io_pixelVal_in_0_4;
      end else if (10'h81 == _T_25[9:0]) begin
        image_0_129 <= io_pixelVal_in_0_3;
      end else if (10'h81 == _T_22[9:0]) begin
        image_0_129 <= io_pixelVal_in_0_2;
      end else if (10'h81 == _T_19[9:0]) begin
        image_0_129 <= io_pixelVal_in_0_1;
      end else if (10'h81 == _T_15[9:0]) begin
        image_0_129 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_130 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h82 == _T_37[9:0]) begin
        image_0_130 <= io_pixelVal_in_0_7;
      end else if (10'h82 == _T_34[9:0]) begin
        image_0_130 <= io_pixelVal_in_0_6;
      end else if (10'h82 == _T_31[9:0]) begin
        image_0_130 <= io_pixelVal_in_0_5;
      end else if (10'h82 == _T_28[9:0]) begin
        image_0_130 <= io_pixelVal_in_0_4;
      end else if (10'h82 == _T_25[9:0]) begin
        image_0_130 <= io_pixelVal_in_0_3;
      end else if (10'h82 == _T_22[9:0]) begin
        image_0_130 <= io_pixelVal_in_0_2;
      end else if (10'h82 == _T_19[9:0]) begin
        image_0_130 <= io_pixelVal_in_0_1;
      end else if (10'h82 == _T_15[9:0]) begin
        image_0_130 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_131 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h83 == _T_37[9:0]) begin
        image_0_131 <= io_pixelVal_in_0_7;
      end else if (10'h83 == _T_34[9:0]) begin
        image_0_131 <= io_pixelVal_in_0_6;
      end else if (10'h83 == _T_31[9:0]) begin
        image_0_131 <= io_pixelVal_in_0_5;
      end else if (10'h83 == _T_28[9:0]) begin
        image_0_131 <= io_pixelVal_in_0_4;
      end else if (10'h83 == _T_25[9:0]) begin
        image_0_131 <= io_pixelVal_in_0_3;
      end else if (10'h83 == _T_22[9:0]) begin
        image_0_131 <= io_pixelVal_in_0_2;
      end else if (10'h83 == _T_19[9:0]) begin
        image_0_131 <= io_pixelVal_in_0_1;
      end else if (10'h83 == _T_15[9:0]) begin
        image_0_131 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_132 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h84 == _T_37[9:0]) begin
        image_0_132 <= io_pixelVal_in_0_7;
      end else if (10'h84 == _T_34[9:0]) begin
        image_0_132 <= io_pixelVal_in_0_6;
      end else if (10'h84 == _T_31[9:0]) begin
        image_0_132 <= io_pixelVal_in_0_5;
      end else if (10'h84 == _T_28[9:0]) begin
        image_0_132 <= io_pixelVal_in_0_4;
      end else if (10'h84 == _T_25[9:0]) begin
        image_0_132 <= io_pixelVal_in_0_3;
      end else if (10'h84 == _T_22[9:0]) begin
        image_0_132 <= io_pixelVal_in_0_2;
      end else if (10'h84 == _T_19[9:0]) begin
        image_0_132 <= io_pixelVal_in_0_1;
      end else if (10'h84 == _T_15[9:0]) begin
        image_0_132 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_133 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h85 == _T_37[9:0]) begin
        image_0_133 <= io_pixelVal_in_0_7;
      end else if (10'h85 == _T_34[9:0]) begin
        image_0_133 <= io_pixelVal_in_0_6;
      end else if (10'h85 == _T_31[9:0]) begin
        image_0_133 <= io_pixelVal_in_0_5;
      end else if (10'h85 == _T_28[9:0]) begin
        image_0_133 <= io_pixelVal_in_0_4;
      end else if (10'h85 == _T_25[9:0]) begin
        image_0_133 <= io_pixelVal_in_0_3;
      end else if (10'h85 == _T_22[9:0]) begin
        image_0_133 <= io_pixelVal_in_0_2;
      end else if (10'h85 == _T_19[9:0]) begin
        image_0_133 <= io_pixelVal_in_0_1;
      end else if (10'h85 == _T_15[9:0]) begin
        image_0_133 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_134 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h86 == _T_37[9:0]) begin
        image_0_134 <= io_pixelVal_in_0_7;
      end else if (10'h86 == _T_34[9:0]) begin
        image_0_134 <= io_pixelVal_in_0_6;
      end else if (10'h86 == _T_31[9:0]) begin
        image_0_134 <= io_pixelVal_in_0_5;
      end else if (10'h86 == _T_28[9:0]) begin
        image_0_134 <= io_pixelVal_in_0_4;
      end else if (10'h86 == _T_25[9:0]) begin
        image_0_134 <= io_pixelVal_in_0_3;
      end else if (10'h86 == _T_22[9:0]) begin
        image_0_134 <= io_pixelVal_in_0_2;
      end else if (10'h86 == _T_19[9:0]) begin
        image_0_134 <= io_pixelVal_in_0_1;
      end else if (10'h86 == _T_15[9:0]) begin
        image_0_134 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_135 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h87 == _T_37[9:0]) begin
        image_0_135 <= io_pixelVal_in_0_7;
      end else if (10'h87 == _T_34[9:0]) begin
        image_0_135 <= io_pixelVal_in_0_6;
      end else if (10'h87 == _T_31[9:0]) begin
        image_0_135 <= io_pixelVal_in_0_5;
      end else if (10'h87 == _T_28[9:0]) begin
        image_0_135 <= io_pixelVal_in_0_4;
      end else if (10'h87 == _T_25[9:0]) begin
        image_0_135 <= io_pixelVal_in_0_3;
      end else if (10'h87 == _T_22[9:0]) begin
        image_0_135 <= io_pixelVal_in_0_2;
      end else if (10'h87 == _T_19[9:0]) begin
        image_0_135 <= io_pixelVal_in_0_1;
      end else if (10'h87 == _T_15[9:0]) begin
        image_0_135 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_136 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h88 == _T_37[9:0]) begin
        image_0_136 <= io_pixelVal_in_0_7;
      end else if (10'h88 == _T_34[9:0]) begin
        image_0_136 <= io_pixelVal_in_0_6;
      end else if (10'h88 == _T_31[9:0]) begin
        image_0_136 <= io_pixelVal_in_0_5;
      end else if (10'h88 == _T_28[9:0]) begin
        image_0_136 <= io_pixelVal_in_0_4;
      end else if (10'h88 == _T_25[9:0]) begin
        image_0_136 <= io_pixelVal_in_0_3;
      end else if (10'h88 == _T_22[9:0]) begin
        image_0_136 <= io_pixelVal_in_0_2;
      end else if (10'h88 == _T_19[9:0]) begin
        image_0_136 <= io_pixelVal_in_0_1;
      end else if (10'h88 == _T_15[9:0]) begin
        image_0_136 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_137 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h89 == _T_37[9:0]) begin
        image_0_137 <= io_pixelVal_in_0_7;
      end else if (10'h89 == _T_34[9:0]) begin
        image_0_137 <= io_pixelVal_in_0_6;
      end else if (10'h89 == _T_31[9:0]) begin
        image_0_137 <= io_pixelVal_in_0_5;
      end else if (10'h89 == _T_28[9:0]) begin
        image_0_137 <= io_pixelVal_in_0_4;
      end else if (10'h89 == _T_25[9:0]) begin
        image_0_137 <= io_pixelVal_in_0_3;
      end else if (10'h89 == _T_22[9:0]) begin
        image_0_137 <= io_pixelVal_in_0_2;
      end else if (10'h89 == _T_19[9:0]) begin
        image_0_137 <= io_pixelVal_in_0_1;
      end else if (10'h89 == _T_15[9:0]) begin
        image_0_137 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_138 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h8a == _T_37[9:0]) begin
        image_0_138 <= io_pixelVal_in_0_7;
      end else if (10'h8a == _T_34[9:0]) begin
        image_0_138 <= io_pixelVal_in_0_6;
      end else if (10'h8a == _T_31[9:0]) begin
        image_0_138 <= io_pixelVal_in_0_5;
      end else if (10'h8a == _T_28[9:0]) begin
        image_0_138 <= io_pixelVal_in_0_4;
      end else if (10'h8a == _T_25[9:0]) begin
        image_0_138 <= io_pixelVal_in_0_3;
      end else if (10'h8a == _T_22[9:0]) begin
        image_0_138 <= io_pixelVal_in_0_2;
      end else if (10'h8a == _T_19[9:0]) begin
        image_0_138 <= io_pixelVal_in_0_1;
      end else if (10'h8a == _T_15[9:0]) begin
        image_0_138 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_139 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h8b == _T_37[9:0]) begin
        image_0_139 <= io_pixelVal_in_0_7;
      end else if (10'h8b == _T_34[9:0]) begin
        image_0_139 <= io_pixelVal_in_0_6;
      end else if (10'h8b == _T_31[9:0]) begin
        image_0_139 <= io_pixelVal_in_0_5;
      end else if (10'h8b == _T_28[9:0]) begin
        image_0_139 <= io_pixelVal_in_0_4;
      end else if (10'h8b == _T_25[9:0]) begin
        image_0_139 <= io_pixelVal_in_0_3;
      end else if (10'h8b == _T_22[9:0]) begin
        image_0_139 <= io_pixelVal_in_0_2;
      end else if (10'h8b == _T_19[9:0]) begin
        image_0_139 <= io_pixelVal_in_0_1;
      end else if (10'h8b == _T_15[9:0]) begin
        image_0_139 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_140 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h8c == _T_37[9:0]) begin
        image_0_140 <= io_pixelVal_in_0_7;
      end else if (10'h8c == _T_34[9:0]) begin
        image_0_140 <= io_pixelVal_in_0_6;
      end else if (10'h8c == _T_31[9:0]) begin
        image_0_140 <= io_pixelVal_in_0_5;
      end else if (10'h8c == _T_28[9:0]) begin
        image_0_140 <= io_pixelVal_in_0_4;
      end else if (10'h8c == _T_25[9:0]) begin
        image_0_140 <= io_pixelVal_in_0_3;
      end else if (10'h8c == _T_22[9:0]) begin
        image_0_140 <= io_pixelVal_in_0_2;
      end else if (10'h8c == _T_19[9:0]) begin
        image_0_140 <= io_pixelVal_in_0_1;
      end else if (10'h8c == _T_15[9:0]) begin
        image_0_140 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_141 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h8d == _T_37[9:0]) begin
        image_0_141 <= io_pixelVal_in_0_7;
      end else if (10'h8d == _T_34[9:0]) begin
        image_0_141 <= io_pixelVal_in_0_6;
      end else if (10'h8d == _T_31[9:0]) begin
        image_0_141 <= io_pixelVal_in_0_5;
      end else if (10'h8d == _T_28[9:0]) begin
        image_0_141 <= io_pixelVal_in_0_4;
      end else if (10'h8d == _T_25[9:0]) begin
        image_0_141 <= io_pixelVal_in_0_3;
      end else if (10'h8d == _T_22[9:0]) begin
        image_0_141 <= io_pixelVal_in_0_2;
      end else if (10'h8d == _T_19[9:0]) begin
        image_0_141 <= io_pixelVal_in_0_1;
      end else if (10'h8d == _T_15[9:0]) begin
        image_0_141 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_142 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h8e == _T_37[9:0]) begin
        image_0_142 <= io_pixelVal_in_0_7;
      end else if (10'h8e == _T_34[9:0]) begin
        image_0_142 <= io_pixelVal_in_0_6;
      end else if (10'h8e == _T_31[9:0]) begin
        image_0_142 <= io_pixelVal_in_0_5;
      end else if (10'h8e == _T_28[9:0]) begin
        image_0_142 <= io_pixelVal_in_0_4;
      end else if (10'h8e == _T_25[9:0]) begin
        image_0_142 <= io_pixelVal_in_0_3;
      end else if (10'h8e == _T_22[9:0]) begin
        image_0_142 <= io_pixelVal_in_0_2;
      end else if (10'h8e == _T_19[9:0]) begin
        image_0_142 <= io_pixelVal_in_0_1;
      end else if (10'h8e == _T_15[9:0]) begin
        image_0_142 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_143 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h8f == _T_37[9:0]) begin
        image_0_143 <= io_pixelVal_in_0_7;
      end else if (10'h8f == _T_34[9:0]) begin
        image_0_143 <= io_pixelVal_in_0_6;
      end else if (10'h8f == _T_31[9:0]) begin
        image_0_143 <= io_pixelVal_in_0_5;
      end else if (10'h8f == _T_28[9:0]) begin
        image_0_143 <= io_pixelVal_in_0_4;
      end else if (10'h8f == _T_25[9:0]) begin
        image_0_143 <= io_pixelVal_in_0_3;
      end else if (10'h8f == _T_22[9:0]) begin
        image_0_143 <= io_pixelVal_in_0_2;
      end else if (10'h8f == _T_19[9:0]) begin
        image_0_143 <= io_pixelVal_in_0_1;
      end else if (10'h8f == _T_15[9:0]) begin
        image_0_143 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_144 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h90 == _T_37[9:0]) begin
        image_0_144 <= io_pixelVal_in_0_7;
      end else if (10'h90 == _T_34[9:0]) begin
        image_0_144 <= io_pixelVal_in_0_6;
      end else if (10'h90 == _T_31[9:0]) begin
        image_0_144 <= io_pixelVal_in_0_5;
      end else if (10'h90 == _T_28[9:0]) begin
        image_0_144 <= io_pixelVal_in_0_4;
      end else if (10'h90 == _T_25[9:0]) begin
        image_0_144 <= io_pixelVal_in_0_3;
      end else if (10'h90 == _T_22[9:0]) begin
        image_0_144 <= io_pixelVal_in_0_2;
      end else if (10'h90 == _T_19[9:0]) begin
        image_0_144 <= io_pixelVal_in_0_1;
      end else if (10'h90 == _T_15[9:0]) begin
        image_0_144 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_145 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h91 == _T_37[9:0]) begin
        image_0_145 <= io_pixelVal_in_0_7;
      end else if (10'h91 == _T_34[9:0]) begin
        image_0_145 <= io_pixelVal_in_0_6;
      end else if (10'h91 == _T_31[9:0]) begin
        image_0_145 <= io_pixelVal_in_0_5;
      end else if (10'h91 == _T_28[9:0]) begin
        image_0_145 <= io_pixelVal_in_0_4;
      end else if (10'h91 == _T_25[9:0]) begin
        image_0_145 <= io_pixelVal_in_0_3;
      end else if (10'h91 == _T_22[9:0]) begin
        image_0_145 <= io_pixelVal_in_0_2;
      end else if (10'h91 == _T_19[9:0]) begin
        image_0_145 <= io_pixelVal_in_0_1;
      end else if (10'h91 == _T_15[9:0]) begin
        image_0_145 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_146 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h92 == _T_37[9:0]) begin
        image_0_146 <= io_pixelVal_in_0_7;
      end else if (10'h92 == _T_34[9:0]) begin
        image_0_146 <= io_pixelVal_in_0_6;
      end else if (10'h92 == _T_31[9:0]) begin
        image_0_146 <= io_pixelVal_in_0_5;
      end else if (10'h92 == _T_28[9:0]) begin
        image_0_146 <= io_pixelVal_in_0_4;
      end else if (10'h92 == _T_25[9:0]) begin
        image_0_146 <= io_pixelVal_in_0_3;
      end else if (10'h92 == _T_22[9:0]) begin
        image_0_146 <= io_pixelVal_in_0_2;
      end else if (10'h92 == _T_19[9:0]) begin
        image_0_146 <= io_pixelVal_in_0_1;
      end else if (10'h92 == _T_15[9:0]) begin
        image_0_146 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_147 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h93 == _T_37[9:0]) begin
        image_0_147 <= io_pixelVal_in_0_7;
      end else if (10'h93 == _T_34[9:0]) begin
        image_0_147 <= io_pixelVal_in_0_6;
      end else if (10'h93 == _T_31[9:0]) begin
        image_0_147 <= io_pixelVal_in_0_5;
      end else if (10'h93 == _T_28[9:0]) begin
        image_0_147 <= io_pixelVal_in_0_4;
      end else if (10'h93 == _T_25[9:0]) begin
        image_0_147 <= io_pixelVal_in_0_3;
      end else if (10'h93 == _T_22[9:0]) begin
        image_0_147 <= io_pixelVal_in_0_2;
      end else if (10'h93 == _T_19[9:0]) begin
        image_0_147 <= io_pixelVal_in_0_1;
      end else if (10'h93 == _T_15[9:0]) begin
        image_0_147 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_148 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h94 == _T_37[9:0]) begin
        image_0_148 <= io_pixelVal_in_0_7;
      end else if (10'h94 == _T_34[9:0]) begin
        image_0_148 <= io_pixelVal_in_0_6;
      end else if (10'h94 == _T_31[9:0]) begin
        image_0_148 <= io_pixelVal_in_0_5;
      end else if (10'h94 == _T_28[9:0]) begin
        image_0_148 <= io_pixelVal_in_0_4;
      end else if (10'h94 == _T_25[9:0]) begin
        image_0_148 <= io_pixelVal_in_0_3;
      end else if (10'h94 == _T_22[9:0]) begin
        image_0_148 <= io_pixelVal_in_0_2;
      end else if (10'h94 == _T_19[9:0]) begin
        image_0_148 <= io_pixelVal_in_0_1;
      end else if (10'h94 == _T_15[9:0]) begin
        image_0_148 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_149 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h95 == _T_37[9:0]) begin
        image_0_149 <= io_pixelVal_in_0_7;
      end else if (10'h95 == _T_34[9:0]) begin
        image_0_149 <= io_pixelVal_in_0_6;
      end else if (10'h95 == _T_31[9:0]) begin
        image_0_149 <= io_pixelVal_in_0_5;
      end else if (10'h95 == _T_28[9:0]) begin
        image_0_149 <= io_pixelVal_in_0_4;
      end else if (10'h95 == _T_25[9:0]) begin
        image_0_149 <= io_pixelVal_in_0_3;
      end else if (10'h95 == _T_22[9:0]) begin
        image_0_149 <= io_pixelVal_in_0_2;
      end else if (10'h95 == _T_19[9:0]) begin
        image_0_149 <= io_pixelVal_in_0_1;
      end else if (10'h95 == _T_15[9:0]) begin
        image_0_149 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_150 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h96 == _T_37[9:0]) begin
        image_0_150 <= io_pixelVal_in_0_7;
      end else if (10'h96 == _T_34[9:0]) begin
        image_0_150 <= io_pixelVal_in_0_6;
      end else if (10'h96 == _T_31[9:0]) begin
        image_0_150 <= io_pixelVal_in_0_5;
      end else if (10'h96 == _T_28[9:0]) begin
        image_0_150 <= io_pixelVal_in_0_4;
      end else if (10'h96 == _T_25[9:0]) begin
        image_0_150 <= io_pixelVal_in_0_3;
      end else if (10'h96 == _T_22[9:0]) begin
        image_0_150 <= io_pixelVal_in_0_2;
      end else if (10'h96 == _T_19[9:0]) begin
        image_0_150 <= io_pixelVal_in_0_1;
      end else if (10'h96 == _T_15[9:0]) begin
        image_0_150 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_151 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h97 == _T_37[9:0]) begin
        image_0_151 <= io_pixelVal_in_0_7;
      end else if (10'h97 == _T_34[9:0]) begin
        image_0_151 <= io_pixelVal_in_0_6;
      end else if (10'h97 == _T_31[9:0]) begin
        image_0_151 <= io_pixelVal_in_0_5;
      end else if (10'h97 == _T_28[9:0]) begin
        image_0_151 <= io_pixelVal_in_0_4;
      end else if (10'h97 == _T_25[9:0]) begin
        image_0_151 <= io_pixelVal_in_0_3;
      end else if (10'h97 == _T_22[9:0]) begin
        image_0_151 <= io_pixelVal_in_0_2;
      end else if (10'h97 == _T_19[9:0]) begin
        image_0_151 <= io_pixelVal_in_0_1;
      end else if (10'h97 == _T_15[9:0]) begin
        image_0_151 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_152 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h98 == _T_37[9:0]) begin
        image_0_152 <= io_pixelVal_in_0_7;
      end else if (10'h98 == _T_34[9:0]) begin
        image_0_152 <= io_pixelVal_in_0_6;
      end else if (10'h98 == _T_31[9:0]) begin
        image_0_152 <= io_pixelVal_in_0_5;
      end else if (10'h98 == _T_28[9:0]) begin
        image_0_152 <= io_pixelVal_in_0_4;
      end else if (10'h98 == _T_25[9:0]) begin
        image_0_152 <= io_pixelVal_in_0_3;
      end else if (10'h98 == _T_22[9:0]) begin
        image_0_152 <= io_pixelVal_in_0_2;
      end else if (10'h98 == _T_19[9:0]) begin
        image_0_152 <= io_pixelVal_in_0_1;
      end else if (10'h98 == _T_15[9:0]) begin
        image_0_152 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_153 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h99 == _T_37[9:0]) begin
        image_0_153 <= io_pixelVal_in_0_7;
      end else if (10'h99 == _T_34[9:0]) begin
        image_0_153 <= io_pixelVal_in_0_6;
      end else if (10'h99 == _T_31[9:0]) begin
        image_0_153 <= io_pixelVal_in_0_5;
      end else if (10'h99 == _T_28[9:0]) begin
        image_0_153 <= io_pixelVal_in_0_4;
      end else if (10'h99 == _T_25[9:0]) begin
        image_0_153 <= io_pixelVal_in_0_3;
      end else if (10'h99 == _T_22[9:0]) begin
        image_0_153 <= io_pixelVal_in_0_2;
      end else if (10'h99 == _T_19[9:0]) begin
        image_0_153 <= io_pixelVal_in_0_1;
      end else if (10'h99 == _T_15[9:0]) begin
        image_0_153 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_154 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h9a == _T_37[9:0]) begin
        image_0_154 <= io_pixelVal_in_0_7;
      end else if (10'h9a == _T_34[9:0]) begin
        image_0_154 <= io_pixelVal_in_0_6;
      end else if (10'h9a == _T_31[9:0]) begin
        image_0_154 <= io_pixelVal_in_0_5;
      end else if (10'h9a == _T_28[9:0]) begin
        image_0_154 <= io_pixelVal_in_0_4;
      end else if (10'h9a == _T_25[9:0]) begin
        image_0_154 <= io_pixelVal_in_0_3;
      end else if (10'h9a == _T_22[9:0]) begin
        image_0_154 <= io_pixelVal_in_0_2;
      end else if (10'h9a == _T_19[9:0]) begin
        image_0_154 <= io_pixelVal_in_0_1;
      end else if (10'h9a == _T_15[9:0]) begin
        image_0_154 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_155 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h9b == _T_37[9:0]) begin
        image_0_155 <= io_pixelVal_in_0_7;
      end else if (10'h9b == _T_34[9:0]) begin
        image_0_155 <= io_pixelVal_in_0_6;
      end else if (10'h9b == _T_31[9:0]) begin
        image_0_155 <= io_pixelVal_in_0_5;
      end else if (10'h9b == _T_28[9:0]) begin
        image_0_155 <= io_pixelVal_in_0_4;
      end else if (10'h9b == _T_25[9:0]) begin
        image_0_155 <= io_pixelVal_in_0_3;
      end else if (10'h9b == _T_22[9:0]) begin
        image_0_155 <= io_pixelVal_in_0_2;
      end else if (10'h9b == _T_19[9:0]) begin
        image_0_155 <= io_pixelVal_in_0_1;
      end else if (10'h9b == _T_15[9:0]) begin
        image_0_155 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_156 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h9c == _T_37[9:0]) begin
        image_0_156 <= io_pixelVal_in_0_7;
      end else if (10'h9c == _T_34[9:0]) begin
        image_0_156 <= io_pixelVal_in_0_6;
      end else if (10'h9c == _T_31[9:0]) begin
        image_0_156 <= io_pixelVal_in_0_5;
      end else if (10'h9c == _T_28[9:0]) begin
        image_0_156 <= io_pixelVal_in_0_4;
      end else if (10'h9c == _T_25[9:0]) begin
        image_0_156 <= io_pixelVal_in_0_3;
      end else if (10'h9c == _T_22[9:0]) begin
        image_0_156 <= io_pixelVal_in_0_2;
      end else if (10'h9c == _T_19[9:0]) begin
        image_0_156 <= io_pixelVal_in_0_1;
      end else if (10'h9c == _T_15[9:0]) begin
        image_0_156 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_157 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h9d == _T_37[9:0]) begin
        image_0_157 <= io_pixelVal_in_0_7;
      end else if (10'h9d == _T_34[9:0]) begin
        image_0_157 <= io_pixelVal_in_0_6;
      end else if (10'h9d == _T_31[9:0]) begin
        image_0_157 <= io_pixelVal_in_0_5;
      end else if (10'h9d == _T_28[9:0]) begin
        image_0_157 <= io_pixelVal_in_0_4;
      end else if (10'h9d == _T_25[9:0]) begin
        image_0_157 <= io_pixelVal_in_0_3;
      end else if (10'h9d == _T_22[9:0]) begin
        image_0_157 <= io_pixelVal_in_0_2;
      end else if (10'h9d == _T_19[9:0]) begin
        image_0_157 <= io_pixelVal_in_0_1;
      end else if (10'h9d == _T_15[9:0]) begin
        image_0_157 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_158 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h9e == _T_37[9:0]) begin
        image_0_158 <= io_pixelVal_in_0_7;
      end else if (10'h9e == _T_34[9:0]) begin
        image_0_158 <= io_pixelVal_in_0_6;
      end else if (10'h9e == _T_31[9:0]) begin
        image_0_158 <= io_pixelVal_in_0_5;
      end else if (10'h9e == _T_28[9:0]) begin
        image_0_158 <= io_pixelVal_in_0_4;
      end else if (10'h9e == _T_25[9:0]) begin
        image_0_158 <= io_pixelVal_in_0_3;
      end else if (10'h9e == _T_22[9:0]) begin
        image_0_158 <= io_pixelVal_in_0_2;
      end else if (10'h9e == _T_19[9:0]) begin
        image_0_158 <= io_pixelVal_in_0_1;
      end else if (10'h9e == _T_15[9:0]) begin
        image_0_158 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_159 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h9f == _T_37[9:0]) begin
        image_0_159 <= io_pixelVal_in_0_7;
      end else if (10'h9f == _T_34[9:0]) begin
        image_0_159 <= io_pixelVal_in_0_6;
      end else if (10'h9f == _T_31[9:0]) begin
        image_0_159 <= io_pixelVal_in_0_5;
      end else if (10'h9f == _T_28[9:0]) begin
        image_0_159 <= io_pixelVal_in_0_4;
      end else if (10'h9f == _T_25[9:0]) begin
        image_0_159 <= io_pixelVal_in_0_3;
      end else if (10'h9f == _T_22[9:0]) begin
        image_0_159 <= io_pixelVal_in_0_2;
      end else if (10'h9f == _T_19[9:0]) begin
        image_0_159 <= io_pixelVal_in_0_1;
      end else if (10'h9f == _T_15[9:0]) begin
        image_0_159 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_160 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'ha0 == _T_37[9:0]) begin
        image_0_160 <= io_pixelVal_in_0_7;
      end else if (10'ha0 == _T_34[9:0]) begin
        image_0_160 <= io_pixelVal_in_0_6;
      end else if (10'ha0 == _T_31[9:0]) begin
        image_0_160 <= io_pixelVal_in_0_5;
      end else if (10'ha0 == _T_28[9:0]) begin
        image_0_160 <= io_pixelVal_in_0_4;
      end else if (10'ha0 == _T_25[9:0]) begin
        image_0_160 <= io_pixelVal_in_0_3;
      end else if (10'ha0 == _T_22[9:0]) begin
        image_0_160 <= io_pixelVal_in_0_2;
      end else if (10'ha0 == _T_19[9:0]) begin
        image_0_160 <= io_pixelVal_in_0_1;
      end else if (10'ha0 == _T_15[9:0]) begin
        image_0_160 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_161 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'ha1 == _T_37[9:0]) begin
        image_0_161 <= io_pixelVal_in_0_7;
      end else if (10'ha1 == _T_34[9:0]) begin
        image_0_161 <= io_pixelVal_in_0_6;
      end else if (10'ha1 == _T_31[9:0]) begin
        image_0_161 <= io_pixelVal_in_0_5;
      end else if (10'ha1 == _T_28[9:0]) begin
        image_0_161 <= io_pixelVal_in_0_4;
      end else if (10'ha1 == _T_25[9:0]) begin
        image_0_161 <= io_pixelVal_in_0_3;
      end else if (10'ha1 == _T_22[9:0]) begin
        image_0_161 <= io_pixelVal_in_0_2;
      end else if (10'ha1 == _T_19[9:0]) begin
        image_0_161 <= io_pixelVal_in_0_1;
      end else if (10'ha1 == _T_15[9:0]) begin
        image_0_161 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_162 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'ha2 == _T_37[9:0]) begin
        image_0_162 <= io_pixelVal_in_0_7;
      end else if (10'ha2 == _T_34[9:0]) begin
        image_0_162 <= io_pixelVal_in_0_6;
      end else if (10'ha2 == _T_31[9:0]) begin
        image_0_162 <= io_pixelVal_in_0_5;
      end else if (10'ha2 == _T_28[9:0]) begin
        image_0_162 <= io_pixelVal_in_0_4;
      end else if (10'ha2 == _T_25[9:0]) begin
        image_0_162 <= io_pixelVal_in_0_3;
      end else if (10'ha2 == _T_22[9:0]) begin
        image_0_162 <= io_pixelVal_in_0_2;
      end else if (10'ha2 == _T_19[9:0]) begin
        image_0_162 <= io_pixelVal_in_0_1;
      end else if (10'ha2 == _T_15[9:0]) begin
        image_0_162 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_163 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'ha3 == _T_37[9:0]) begin
        image_0_163 <= io_pixelVal_in_0_7;
      end else if (10'ha3 == _T_34[9:0]) begin
        image_0_163 <= io_pixelVal_in_0_6;
      end else if (10'ha3 == _T_31[9:0]) begin
        image_0_163 <= io_pixelVal_in_0_5;
      end else if (10'ha3 == _T_28[9:0]) begin
        image_0_163 <= io_pixelVal_in_0_4;
      end else if (10'ha3 == _T_25[9:0]) begin
        image_0_163 <= io_pixelVal_in_0_3;
      end else if (10'ha3 == _T_22[9:0]) begin
        image_0_163 <= io_pixelVal_in_0_2;
      end else if (10'ha3 == _T_19[9:0]) begin
        image_0_163 <= io_pixelVal_in_0_1;
      end else if (10'ha3 == _T_15[9:0]) begin
        image_0_163 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_164 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'ha4 == _T_37[9:0]) begin
        image_0_164 <= io_pixelVal_in_0_7;
      end else if (10'ha4 == _T_34[9:0]) begin
        image_0_164 <= io_pixelVal_in_0_6;
      end else if (10'ha4 == _T_31[9:0]) begin
        image_0_164 <= io_pixelVal_in_0_5;
      end else if (10'ha4 == _T_28[9:0]) begin
        image_0_164 <= io_pixelVal_in_0_4;
      end else if (10'ha4 == _T_25[9:0]) begin
        image_0_164 <= io_pixelVal_in_0_3;
      end else if (10'ha4 == _T_22[9:0]) begin
        image_0_164 <= io_pixelVal_in_0_2;
      end else if (10'ha4 == _T_19[9:0]) begin
        image_0_164 <= io_pixelVal_in_0_1;
      end else if (10'ha4 == _T_15[9:0]) begin
        image_0_164 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_165 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'ha5 == _T_37[9:0]) begin
        image_0_165 <= io_pixelVal_in_0_7;
      end else if (10'ha5 == _T_34[9:0]) begin
        image_0_165 <= io_pixelVal_in_0_6;
      end else if (10'ha5 == _T_31[9:0]) begin
        image_0_165 <= io_pixelVal_in_0_5;
      end else if (10'ha5 == _T_28[9:0]) begin
        image_0_165 <= io_pixelVal_in_0_4;
      end else if (10'ha5 == _T_25[9:0]) begin
        image_0_165 <= io_pixelVal_in_0_3;
      end else if (10'ha5 == _T_22[9:0]) begin
        image_0_165 <= io_pixelVal_in_0_2;
      end else if (10'ha5 == _T_19[9:0]) begin
        image_0_165 <= io_pixelVal_in_0_1;
      end else if (10'ha5 == _T_15[9:0]) begin
        image_0_165 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_166 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'ha6 == _T_37[9:0]) begin
        image_0_166 <= io_pixelVal_in_0_7;
      end else if (10'ha6 == _T_34[9:0]) begin
        image_0_166 <= io_pixelVal_in_0_6;
      end else if (10'ha6 == _T_31[9:0]) begin
        image_0_166 <= io_pixelVal_in_0_5;
      end else if (10'ha6 == _T_28[9:0]) begin
        image_0_166 <= io_pixelVal_in_0_4;
      end else if (10'ha6 == _T_25[9:0]) begin
        image_0_166 <= io_pixelVal_in_0_3;
      end else if (10'ha6 == _T_22[9:0]) begin
        image_0_166 <= io_pixelVal_in_0_2;
      end else if (10'ha6 == _T_19[9:0]) begin
        image_0_166 <= io_pixelVal_in_0_1;
      end else if (10'ha6 == _T_15[9:0]) begin
        image_0_166 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_167 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'ha7 == _T_37[9:0]) begin
        image_0_167 <= io_pixelVal_in_0_7;
      end else if (10'ha7 == _T_34[9:0]) begin
        image_0_167 <= io_pixelVal_in_0_6;
      end else if (10'ha7 == _T_31[9:0]) begin
        image_0_167 <= io_pixelVal_in_0_5;
      end else if (10'ha7 == _T_28[9:0]) begin
        image_0_167 <= io_pixelVal_in_0_4;
      end else if (10'ha7 == _T_25[9:0]) begin
        image_0_167 <= io_pixelVal_in_0_3;
      end else if (10'ha7 == _T_22[9:0]) begin
        image_0_167 <= io_pixelVal_in_0_2;
      end else if (10'ha7 == _T_19[9:0]) begin
        image_0_167 <= io_pixelVal_in_0_1;
      end else if (10'ha7 == _T_15[9:0]) begin
        image_0_167 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_168 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'ha8 == _T_37[9:0]) begin
        image_0_168 <= io_pixelVal_in_0_7;
      end else if (10'ha8 == _T_34[9:0]) begin
        image_0_168 <= io_pixelVal_in_0_6;
      end else if (10'ha8 == _T_31[9:0]) begin
        image_0_168 <= io_pixelVal_in_0_5;
      end else if (10'ha8 == _T_28[9:0]) begin
        image_0_168 <= io_pixelVal_in_0_4;
      end else if (10'ha8 == _T_25[9:0]) begin
        image_0_168 <= io_pixelVal_in_0_3;
      end else if (10'ha8 == _T_22[9:0]) begin
        image_0_168 <= io_pixelVal_in_0_2;
      end else if (10'ha8 == _T_19[9:0]) begin
        image_0_168 <= io_pixelVal_in_0_1;
      end else if (10'ha8 == _T_15[9:0]) begin
        image_0_168 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_169 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'ha9 == _T_37[9:0]) begin
        image_0_169 <= io_pixelVal_in_0_7;
      end else if (10'ha9 == _T_34[9:0]) begin
        image_0_169 <= io_pixelVal_in_0_6;
      end else if (10'ha9 == _T_31[9:0]) begin
        image_0_169 <= io_pixelVal_in_0_5;
      end else if (10'ha9 == _T_28[9:0]) begin
        image_0_169 <= io_pixelVal_in_0_4;
      end else if (10'ha9 == _T_25[9:0]) begin
        image_0_169 <= io_pixelVal_in_0_3;
      end else if (10'ha9 == _T_22[9:0]) begin
        image_0_169 <= io_pixelVal_in_0_2;
      end else if (10'ha9 == _T_19[9:0]) begin
        image_0_169 <= io_pixelVal_in_0_1;
      end else if (10'ha9 == _T_15[9:0]) begin
        image_0_169 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_170 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'haa == _T_37[9:0]) begin
        image_0_170 <= io_pixelVal_in_0_7;
      end else if (10'haa == _T_34[9:0]) begin
        image_0_170 <= io_pixelVal_in_0_6;
      end else if (10'haa == _T_31[9:0]) begin
        image_0_170 <= io_pixelVal_in_0_5;
      end else if (10'haa == _T_28[9:0]) begin
        image_0_170 <= io_pixelVal_in_0_4;
      end else if (10'haa == _T_25[9:0]) begin
        image_0_170 <= io_pixelVal_in_0_3;
      end else if (10'haa == _T_22[9:0]) begin
        image_0_170 <= io_pixelVal_in_0_2;
      end else if (10'haa == _T_19[9:0]) begin
        image_0_170 <= io_pixelVal_in_0_1;
      end else if (10'haa == _T_15[9:0]) begin
        image_0_170 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_171 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hab == _T_37[9:0]) begin
        image_0_171 <= io_pixelVal_in_0_7;
      end else if (10'hab == _T_34[9:0]) begin
        image_0_171 <= io_pixelVal_in_0_6;
      end else if (10'hab == _T_31[9:0]) begin
        image_0_171 <= io_pixelVal_in_0_5;
      end else if (10'hab == _T_28[9:0]) begin
        image_0_171 <= io_pixelVal_in_0_4;
      end else if (10'hab == _T_25[9:0]) begin
        image_0_171 <= io_pixelVal_in_0_3;
      end else if (10'hab == _T_22[9:0]) begin
        image_0_171 <= io_pixelVal_in_0_2;
      end else if (10'hab == _T_19[9:0]) begin
        image_0_171 <= io_pixelVal_in_0_1;
      end else if (10'hab == _T_15[9:0]) begin
        image_0_171 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_172 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hac == _T_37[9:0]) begin
        image_0_172 <= io_pixelVal_in_0_7;
      end else if (10'hac == _T_34[9:0]) begin
        image_0_172 <= io_pixelVal_in_0_6;
      end else if (10'hac == _T_31[9:0]) begin
        image_0_172 <= io_pixelVal_in_0_5;
      end else if (10'hac == _T_28[9:0]) begin
        image_0_172 <= io_pixelVal_in_0_4;
      end else if (10'hac == _T_25[9:0]) begin
        image_0_172 <= io_pixelVal_in_0_3;
      end else if (10'hac == _T_22[9:0]) begin
        image_0_172 <= io_pixelVal_in_0_2;
      end else if (10'hac == _T_19[9:0]) begin
        image_0_172 <= io_pixelVal_in_0_1;
      end else if (10'hac == _T_15[9:0]) begin
        image_0_172 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_173 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'had == _T_37[9:0]) begin
        image_0_173 <= io_pixelVal_in_0_7;
      end else if (10'had == _T_34[9:0]) begin
        image_0_173 <= io_pixelVal_in_0_6;
      end else if (10'had == _T_31[9:0]) begin
        image_0_173 <= io_pixelVal_in_0_5;
      end else if (10'had == _T_28[9:0]) begin
        image_0_173 <= io_pixelVal_in_0_4;
      end else if (10'had == _T_25[9:0]) begin
        image_0_173 <= io_pixelVal_in_0_3;
      end else if (10'had == _T_22[9:0]) begin
        image_0_173 <= io_pixelVal_in_0_2;
      end else if (10'had == _T_19[9:0]) begin
        image_0_173 <= io_pixelVal_in_0_1;
      end else if (10'had == _T_15[9:0]) begin
        image_0_173 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_174 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hae == _T_37[9:0]) begin
        image_0_174 <= io_pixelVal_in_0_7;
      end else if (10'hae == _T_34[9:0]) begin
        image_0_174 <= io_pixelVal_in_0_6;
      end else if (10'hae == _T_31[9:0]) begin
        image_0_174 <= io_pixelVal_in_0_5;
      end else if (10'hae == _T_28[9:0]) begin
        image_0_174 <= io_pixelVal_in_0_4;
      end else if (10'hae == _T_25[9:0]) begin
        image_0_174 <= io_pixelVal_in_0_3;
      end else if (10'hae == _T_22[9:0]) begin
        image_0_174 <= io_pixelVal_in_0_2;
      end else if (10'hae == _T_19[9:0]) begin
        image_0_174 <= io_pixelVal_in_0_1;
      end else if (10'hae == _T_15[9:0]) begin
        image_0_174 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_175 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'haf == _T_37[9:0]) begin
        image_0_175 <= io_pixelVal_in_0_7;
      end else if (10'haf == _T_34[9:0]) begin
        image_0_175 <= io_pixelVal_in_0_6;
      end else if (10'haf == _T_31[9:0]) begin
        image_0_175 <= io_pixelVal_in_0_5;
      end else if (10'haf == _T_28[9:0]) begin
        image_0_175 <= io_pixelVal_in_0_4;
      end else if (10'haf == _T_25[9:0]) begin
        image_0_175 <= io_pixelVal_in_0_3;
      end else if (10'haf == _T_22[9:0]) begin
        image_0_175 <= io_pixelVal_in_0_2;
      end else if (10'haf == _T_19[9:0]) begin
        image_0_175 <= io_pixelVal_in_0_1;
      end else if (10'haf == _T_15[9:0]) begin
        image_0_175 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_176 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hb0 == _T_37[9:0]) begin
        image_0_176 <= io_pixelVal_in_0_7;
      end else if (10'hb0 == _T_34[9:0]) begin
        image_0_176 <= io_pixelVal_in_0_6;
      end else if (10'hb0 == _T_31[9:0]) begin
        image_0_176 <= io_pixelVal_in_0_5;
      end else if (10'hb0 == _T_28[9:0]) begin
        image_0_176 <= io_pixelVal_in_0_4;
      end else if (10'hb0 == _T_25[9:0]) begin
        image_0_176 <= io_pixelVal_in_0_3;
      end else if (10'hb0 == _T_22[9:0]) begin
        image_0_176 <= io_pixelVal_in_0_2;
      end else if (10'hb0 == _T_19[9:0]) begin
        image_0_176 <= io_pixelVal_in_0_1;
      end else if (10'hb0 == _T_15[9:0]) begin
        image_0_176 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_177 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hb1 == _T_37[9:0]) begin
        image_0_177 <= io_pixelVal_in_0_7;
      end else if (10'hb1 == _T_34[9:0]) begin
        image_0_177 <= io_pixelVal_in_0_6;
      end else if (10'hb1 == _T_31[9:0]) begin
        image_0_177 <= io_pixelVal_in_0_5;
      end else if (10'hb1 == _T_28[9:0]) begin
        image_0_177 <= io_pixelVal_in_0_4;
      end else if (10'hb1 == _T_25[9:0]) begin
        image_0_177 <= io_pixelVal_in_0_3;
      end else if (10'hb1 == _T_22[9:0]) begin
        image_0_177 <= io_pixelVal_in_0_2;
      end else if (10'hb1 == _T_19[9:0]) begin
        image_0_177 <= io_pixelVal_in_0_1;
      end else if (10'hb1 == _T_15[9:0]) begin
        image_0_177 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_178 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hb2 == _T_37[9:0]) begin
        image_0_178 <= io_pixelVal_in_0_7;
      end else if (10'hb2 == _T_34[9:0]) begin
        image_0_178 <= io_pixelVal_in_0_6;
      end else if (10'hb2 == _T_31[9:0]) begin
        image_0_178 <= io_pixelVal_in_0_5;
      end else if (10'hb2 == _T_28[9:0]) begin
        image_0_178 <= io_pixelVal_in_0_4;
      end else if (10'hb2 == _T_25[9:0]) begin
        image_0_178 <= io_pixelVal_in_0_3;
      end else if (10'hb2 == _T_22[9:0]) begin
        image_0_178 <= io_pixelVal_in_0_2;
      end else if (10'hb2 == _T_19[9:0]) begin
        image_0_178 <= io_pixelVal_in_0_1;
      end else if (10'hb2 == _T_15[9:0]) begin
        image_0_178 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_179 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hb3 == _T_37[9:0]) begin
        image_0_179 <= io_pixelVal_in_0_7;
      end else if (10'hb3 == _T_34[9:0]) begin
        image_0_179 <= io_pixelVal_in_0_6;
      end else if (10'hb3 == _T_31[9:0]) begin
        image_0_179 <= io_pixelVal_in_0_5;
      end else if (10'hb3 == _T_28[9:0]) begin
        image_0_179 <= io_pixelVal_in_0_4;
      end else if (10'hb3 == _T_25[9:0]) begin
        image_0_179 <= io_pixelVal_in_0_3;
      end else if (10'hb3 == _T_22[9:0]) begin
        image_0_179 <= io_pixelVal_in_0_2;
      end else if (10'hb3 == _T_19[9:0]) begin
        image_0_179 <= io_pixelVal_in_0_1;
      end else if (10'hb3 == _T_15[9:0]) begin
        image_0_179 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_180 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hb4 == _T_37[9:0]) begin
        image_0_180 <= io_pixelVal_in_0_7;
      end else if (10'hb4 == _T_34[9:0]) begin
        image_0_180 <= io_pixelVal_in_0_6;
      end else if (10'hb4 == _T_31[9:0]) begin
        image_0_180 <= io_pixelVal_in_0_5;
      end else if (10'hb4 == _T_28[9:0]) begin
        image_0_180 <= io_pixelVal_in_0_4;
      end else if (10'hb4 == _T_25[9:0]) begin
        image_0_180 <= io_pixelVal_in_0_3;
      end else if (10'hb4 == _T_22[9:0]) begin
        image_0_180 <= io_pixelVal_in_0_2;
      end else if (10'hb4 == _T_19[9:0]) begin
        image_0_180 <= io_pixelVal_in_0_1;
      end else if (10'hb4 == _T_15[9:0]) begin
        image_0_180 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_181 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hb5 == _T_37[9:0]) begin
        image_0_181 <= io_pixelVal_in_0_7;
      end else if (10'hb5 == _T_34[9:0]) begin
        image_0_181 <= io_pixelVal_in_0_6;
      end else if (10'hb5 == _T_31[9:0]) begin
        image_0_181 <= io_pixelVal_in_0_5;
      end else if (10'hb5 == _T_28[9:0]) begin
        image_0_181 <= io_pixelVal_in_0_4;
      end else if (10'hb5 == _T_25[9:0]) begin
        image_0_181 <= io_pixelVal_in_0_3;
      end else if (10'hb5 == _T_22[9:0]) begin
        image_0_181 <= io_pixelVal_in_0_2;
      end else if (10'hb5 == _T_19[9:0]) begin
        image_0_181 <= io_pixelVal_in_0_1;
      end else if (10'hb5 == _T_15[9:0]) begin
        image_0_181 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_182 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hb6 == _T_37[9:0]) begin
        image_0_182 <= io_pixelVal_in_0_7;
      end else if (10'hb6 == _T_34[9:0]) begin
        image_0_182 <= io_pixelVal_in_0_6;
      end else if (10'hb6 == _T_31[9:0]) begin
        image_0_182 <= io_pixelVal_in_0_5;
      end else if (10'hb6 == _T_28[9:0]) begin
        image_0_182 <= io_pixelVal_in_0_4;
      end else if (10'hb6 == _T_25[9:0]) begin
        image_0_182 <= io_pixelVal_in_0_3;
      end else if (10'hb6 == _T_22[9:0]) begin
        image_0_182 <= io_pixelVal_in_0_2;
      end else if (10'hb6 == _T_19[9:0]) begin
        image_0_182 <= io_pixelVal_in_0_1;
      end else if (10'hb6 == _T_15[9:0]) begin
        image_0_182 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_183 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hb7 == _T_37[9:0]) begin
        image_0_183 <= io_pixelVal_in_0_7;
      end else if (10'hb7 == _T_34[9:0]) begin
        image_0_183 <= io_pixelVal_in_0_6;
      end else if (10'hb7 == _T_31[9:0]) begin
        image_0_183 <= io_pixelVal_in_0_5;
      end else if (10'hb7 == _T_28[9:0]) begin
        image_0_183 <= io_pixelVal_in_0_4;
      end else if (10'hb7 == _T_25[9:0]) begin
        image_0_183 <= io_pixelVal_in_0_3;
      end else if (10'hb7 == _T_22[9:0]) begin
        image_0_183 <= io_pixelVal_in_0_2;
      end else if (10'hb7 == _T_19[9:0]) begin
        image_0_183 <= io_pixelVal_in_0_1;
      end else if (10'hb7 == _T_15[9:0]) begin
        image_0_183 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_184 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hb8 == _T_37[9:0]) begin
        image_0_184 <= io_pixelVal_in_0_7;
      end else if (10'hb8 == _T_34[9:0]) begin
        image_0_184 <= io_pixelVal_in_0_6;
      end else if (10'hb8 == _T_31[9:0]) begin
        image_0_184 <= io_pixelVal_in_0_5;
      end else if (10'hb8 == _T_28[9:0]) begin
        image_0_184 <= io_pixelVal_in_0_4;
      end else if (10'hb8 == _T_25[9:0]) begin
        image_0_184 <= io_pixelVal_in_0_3;
      end else if (10'hb8 == _T_22[9:0]) begin
        image_0_184 <= io_pixelVal_in_0_2;
      end else if (10'hb8 == _T_19[9:0]) begin
        image_0_184 <= io_pixelVal_in_0_1;
      end else if (10'hb8 == _T_15[9:0]) begin
        image_0_184 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_185 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hb9 == _T_37[9:0]) begin
        image_0_185 <= io_pixelVal_in_0_7;
      end else if (10'hb9 == _T_34[9:0]) begin
        image_0_185 <= io_pixelVal_in_0_6;
      end else if (10'hb9 == _T_31[9:0]) begin
        image_0_185 <= io_pixelVal_in_0_5;
      end else if (10'hb9 == _T_28[9:0]) begin
        image_0_185 <= io_pixelVal_in_0_4;
      end else if (10'hb9 == _T_25[9:0]) begin
        image_0_185 <= io_pixelVal_in_0_3;
      end else if (10'hb9 == _T_22[9:0]) begin
        image_0_185 <= io_pixelVal_in_0_2;
      end else if (10'hb9 == _T_19[9:0]) begin
        image_0_185 <= io_pixelVal_in_0_1;
      end else if (10'hb9 == _T_15[9:0]) begin
        image_0_185 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_186 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hba == _T_37[9:0]) begin
        image_0_186 <= io_pixelVal_in_0_7;
      end else if (10'hba == _T_34[9:0]) begin
        image_0_186 <= io_pixelVal_in_0_6;
      end else if (10'hba == _T_31[9:0]) begin
        image_0_186 <= io_pixelVal_in_0_5;
      end else if (10'hba == _T_28[9:0]) begin
        image_0_186 <= io_pixelVal_in_0_4;
      end else if (10'hba == _T_25[9:0]) begin
        image_0_186 <= io_pixelVal_in_0_3;
      end else if (10'hba == _T_22[9:0]) begin
        image_0_186 <= io_pixelVal_in_0_2;
      end else if (10'hba == _T_19[9:0]) begin
        image_0_186 <= io_pixelVal_in_0_1;
      end else if (10'hba == _T_15[9:0]) begin
        image_0_186 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_187 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hbb == _T_37[9:0]) begin
        image_0_187 <= io_pixelVal_in_0_7;
      end else if (10'hbb == _T_34[9:0]) begin
        image_0_187 <= io_pixelVal_in_0_6;
      end else if (10'hbb == _T_31[9:0]) begin
        image_0_187 <= io_pixelVal_in_0_5;
      end else if (10'hbb == _T_28[9:0]) begin
        image_0_187 <= io_pixelVal_in_0_4;
      end else if (10'hbb == _T_25[9:0]) begin
        image_0_187 <= io_pixelVal_in_0_3;
      end else if (10'hbb == _T_22[9:0]) begin
        image_0_187 <= io_pixelVal_in_0_2;
      end else if (10'hbb == _T_19[9:0]) begin
        image_0_187 <= io_pixelVal_in_0_1;
      end else if (10'hbb == _T_15[9:0]) begin
        image_0_187 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_188 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hbc == _T_37[9:0]) begin
        image_0_188 <= io_pixelVal_in_0_7;
      end else if (10'hbc == _T_34[9:0]) begin
        image_0_188 <= io_pixelVal_in_0_6;
      end else if (10'hbc == _T_31[9:0]) begin
        image_0_188 <= io_pixelVal_in_0_5;
      end else if (10'hbc == _T_28[9:0]) begin
        image_0_188 <= io_pixelVal_in_0_4;
      end else if (10'hbc == _T_25[9:0]) begin
        image_0_188 <= io_pixelVal_in_0_3;
      end else if (10'hbc == _T_22[9:0]) begin
        image_0_188 <= io_pixelVal_in_0_2;
      end else if (10'hbc == _T_19[9:0]) begin
        image_0_188 <= io_pixelVal_in_0_1;
      end else if (10'hbc == _T_15[9:0]) begin
        image_0_188 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_189 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hbd == _T_37[9:0]) begin
        image_0_189 <= io_pixelVal_in_0_7;
      end else if (10'hbd == _T_34[9:0]) begin
        image_0_189 <= io_pixelVal_in_0_6;
      end else if (10'hbd == _T_31[9:0]) begin
        image_0_189 <= io_pixelVal_in_0_5;
      end else if (10'hbd == _T_28[9:0]) begin
        image_0_189 <= io_pixelVal_in_0_4;
      end else if (10'hbd == _T_25[9:0]) begin
        image_0_189 <= io_pixelVal_in_0_3;
      end else if (10'hbd == _T_22[9:0]) begin
        image_0_189 <= io_pixelVal_in_0_2;
      end else if (10'hbd == _T_19[9:0]) begin
        image_0_189 <= io_pixelVal_in_0_1;
      end else if (10'hbd == _T_15[9:0]) begin
        image_0_189 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_190 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hbe == _T_37[9:0]) begin
        image_0_190 <= io_pixelVal_in_0_7;
      end else if (10'hbe == _T_34[9:0]) begin
        image_0_190 <= io_pixelVal_in_0_6;
      end else if (10'hbe == _T_31[9:0]) begin
        image_0_190 <= io_pixelVal_in_0_5;
      end else if (10'hbe == _T_28[9:0]) begin
        image_0_190 <= io_pixelVal_in_0_4;
      end else if (10'hbe == _T_25[9:0]) begin
        image_0_190 <= io_pixelVal_in_0_3;
      end else if (10'hbe == _T_22[9:0]) begin
        image_0_190 <= io_pixelVal_in_0_2;
      end else if (10'hbe == _T_19[9:0]) begin
        image_0_190 <= io_pixelVal_in_0_1;
      end else if (10'hbe == _T_15[9:0]) begin
        image_0_190 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_191 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hbf == _T_37[9:0]) begin
        image_0_191 <= io_pixelVal_in_0_7;
      end else if (10'hbf == _T_34[9:0]) begin
        image_0_191 <= io_pixelVal_in_0_6;
      end else if (10'hbf == _T_31[9:0]) begin
        image_0_191 <= io_pixelVal_in_0_5;
      end else if (10'hbf == _T_28[9:0]) begin
        image_0_191 <= io_pixelVal_in_0_4;
      end else if (10'hbf == _T_25[9:0]) begin
        image_0_191 <= io_pixelVal_in_0_3;
      end else if (10'hbf == _T_22[9:0]) begin
        image_0_191 <= io_pixelVal_in_0_2;
      end else if (10'hbf == _T_19[9:0]) begin
        image_0_191 <= io_pixelVal_in_0_1;
      end else if (10'hbf == _T_15[9:0]) begin
        image_0_191 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_192 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hc0 == _T_37[9:0]) begin
        image_0_192 <= io_pixelVal_in_0_7;
      end else if (10'hc0 == _T_34[9:0]) begin
        image_0_192 <= io_pixelVal_in_0_6;
      end else if (10'hc0 == _T_31[9:0]) begin
        image_0_192 <= io_pixelVal_in_0_5;
      end else if (10'hc0 == _T_28[9:0]) begin
        image_0_192 <= io_pixelVal_in_0_4;
      end else if (10'hc0 == _T_25[9:0]) begin
        image_0_192 <= io_pixelVal_in_0_3;
      end else if (10'hc0 == _T_22[9:0]) begin
        image_0_192 <= io_pixelVal_in_0_2;
      end else if (10'hc0 == _T_19[9:0]) begin
        image_0_192 <= io_pixelVal_in_0_1;
      end else if (10'hc0 == _T_15[9:0]) begin
        image_0_192 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_193 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hc1 == _T_37[9:0]) begin
        image_0_193 <= io_pixelVal_in_0_7;
      end else if (10'hc1 == _T_34[9:0]) begin
        image_0_193 <= io_pixelVal_in_0_6;
      end else if (10'hc1 == _T_31[9:0]) begin
        image_0_193 <= io_pixelVal_in_0_5;
      end else if (10'hc1 == _T_28[9:0]) begin
        image_0_193 <= io_pixelVal_in_0_4;
      end else if (10'hc1 == _T_25[9:0]) begin
        image_0_193 <= io_pixelVal_in_0_3;
      end else if (10'hc1 == _T_22[9:0]) begin
        image_0_193 <= io_pixelVal_in_0_2;
      end else if (10'hc1 == _T_19[9:0]) begin
        image_0_193 <= io_pixelVal_in_0_1;
      end else if (10'hc1 == _T_15[9:0]) begin
        image_0_193 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_194 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hc2 == _T_37[9:0]) begin
        image_0_194 <= io_pixelVal_in_0_7;
      end else if (10'hc2 == _T_34[9:0]) begin
        image_0_194 <= io_pixelVal_in_0_6;
      end else if (10'hc2 == _T_31[9:0]) begin
        image_0_194 <= io_pixelVal_in_0_5;
      end else if (10'hc2 == _T_28[9:0]) begin
        image_0_194 <= io_pixelVal_in_0_4;
      end else if (10'hc2 == _T_25[9:0]) begin
        image_0_194 <= io_pixelVal_in_0_3;
      end else if (10'hc2 == _T_22[9:0]) begin
        image_0_194 <= io_pixelVal_in_0_2;
      end else if (10'hc2 == _T_19[9:0]) begin
        image_0_194 <= io_pixelVal_in_0_1;
      end else if (10'hc2 == _T_15[9:0]) begin
        image_0_194 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_195 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hc3 == _T_37[9:0]) begin
        image_0_195 <= io_pixelVal_in_0_7;
      end else if (10'hc3 == _T_34[9:0]) begin
        image_0_195 <= io_pixelVal_in_0_6;
      end else if (10'hc3 == _T_31[9:0]) begin
        image_0_195 <= io_pixelVal_in_0_5;
      end else if (10'hc3 == _T_28[9:0]) begin
        image_0_195 <= io_pixelVal_in_0_4;
      end else if (10'hc3 == _T_25[9:0]) begin
        image_0_195 <= io_pixelVal_in_0_3;
      end else if (10'hc3 == _T_22[9:0]) begin
        image_0_195 <= io_pixelVal_in_0_2;
      end else if (10'hc3 == _T_19[9:0]) begin
        image_0_195 <= io_pixelVal_in_0_1;
      end else if (10'hc3 == _T_15[9:0]) begin
        image_0_195 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_196 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hc4 == _T_37[9:0]) begin
        image_0_196 <= io_pixelVal_in_0_7;
      end else if (10'hc4 == _T_34[9:0]) begin
        image_0_196 <= io_pixelVal_in_0_6;
      end else if (10'hc4 == _T_31[9:0]) begin
        image_0_196 <= io_pixelVal_in_0_5;
      end else if (10'hc4 == _T_28[9:0]) begin
        image_0_196 <= io_pixelVal_in_0_4;
      end else if (10'hc4 == _T_25[9:0]) begin
        image_0_196 <= io_pixelVal_in_0_3;
      end else if (10'hc4 == _T_22[9:0]) begin
        image_0_196 <= io_pixelVal_in_0_2;
      end else if (10'hc4 == _T_19[9:0]) begin
        image_0_196 <= io_pixelVal_in_0_1;
      end else if (10'hc4 == _T_15[9:0]) begin
        image_0_196 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_197 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hc5 == _T_37[9:0]) begin
        image_0_197 <= io_pixelVal_in_0_7;
      end else if (10'hc5 == _T_34[9:0]) begin
        image_0_197 <= io_pixelVal_in_0_6;
      end else if (10'hc5 == _T_31[9:0]) begin
        image_0_197 <= io_pixelVal_in_0_5;
      end else if (10'hc5 == _T_28[9:0]) begin
        image_0_197 <= io_pixelVal_in_0_4;
      end else if (10'hc5 == _T_25[9:0]) begin
        image_0_197 <= io_pixelVal_in_0_3;
      end else if (10'hc5 == _T_22[9:0]) begin
        image_0_197 <= io_pixelVal_in_0_2;
      end else if (10'hc5 == _T_19[9:0]) begin
        image_0_197 <= io_pixelVal_in_0_1;
      end else if (10'hc5 == _T_15[9:0]) begin
        image_0_197 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_198 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hc6 == _T_37[9:0]) begin
        image_0_198 <= io_pixelVal_in_0_7;
      end else if (10'hc6 == _T_34[9:0]) begin
        image_0_198 <= io_pixelVal_in_0_6;
      end else if (10'hc6 == _T_31[9:0]) begin
        image_0_198 <= io_pixelVal_in_0_5;
      end else if (10'hc6 == _T_28[9:0]) begin
        image_0_198 <= io_pixelVal_in_0_4;
      end else if (10'hc6 == _T_25[9:0]) begin
        image_0_198 <= io_pixelVal_in_0_3;
      end else if (10'hc6 == _T_22[9:0]) begin
        image_0_198 <= io_pixelVal_in_0_2;
      end else if (10'hc6 == _T_19[9:0]) begin
        image_0_198 <= io_pixelVal_in_0_1;
      end else if (10'hc6 == _T_15[9:0]) begin
        image_0_198 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_199 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hc7 == _T_37[9:0]) begin
        image_0_199 <= io_pixelVal_in_0_7;
      end else if (10'hc7 == _T_34[9:0]) begin
        image_0_199 <= io_pixelVal_in_0_6;
      end else if (10'hc7 == _T_31[9:0]) begin
        image_0_199 <= io_pixelVal_in_0_5;
      end else if (10'hc7 == _T_28[9:0]) begin
        image_0_199 <= io_pixelVal_in_0_4;
      end else if (10'hc7 == _T_25[9:0]) begin
        image_0_199 <= io_pixelVal_in_0_3;
      end else if (10'hc7 == _T_22[9:0]) begin
        image_0_199 <= io_pixelVal_in_0_2;
      end else if (10'hc7 == _T_19[9:0]) begin
        image_0_199 <= io_pixelVal_in_0_1;
      end else if (10'hc7 == _T_15[9:0]) begin
        image_0_199 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_200 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hc8 == _T_37[9:0]) begin
        image_0_200 <= io_pixelVal_in_0_7;
      end else if (10'hc8 == _T_34[9:0]) begin
        image_0_200 <= io_pixelVal_in_0_6;
      end else if (10'hc8 == _T_31[9:0]) begin
        image_0_200 <= io_pixelVal_in_0_5;
      end else if (10'hc8 == _T_28[9:0]) begin
        image_0_200 <= io_pixelVal_in_0_4;
      end else if (10'hc8 == _T_25[9:0]) begin
        image_0_200 <= io_pixelVal_in_0_3;
      end else if (10'hc8 == _T_22[9:0]) begin
        image_0_200 <= io_pixelVal_in_0_2;
      end else if (10'hc8 == _T_19[9:0]) begin
        image_0_200 <= io_pixelVal_in_0_1;
      end else if (10'hc8 == _T_15[9:0]) begin
        image_0_200 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_201 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hc9 == _T_37[9:0]) begin
        image_0_201 <= io_pixelVal_in_0_7;
      end else if (10'hc9 == _T_34[9:0]) begin
        image_0_201 <= io_pixelVal_in_0_6;
      end else if (10'hc9 == _T_31[9:0]) begin
        image_0_201 <= io_pixelVal_in_0_5;
      end else if (10'hc9 == _T_28[9:0]) begin
        image_0_201 <= io_pixelVal_in_0_4;
      end else if (10'hc9 == _T_25[9:0]) begin
        image_0_201 <= io_pixelVal_in_0_3;
      end else if (10'hc9 == _T_22[9:0]) begin
        image_0_201 <= io_pixelVal_in_0_2;
      end else if (10'hc9 == _T_19[9:0]) begin
        image_0_201 <= io_pixelVal_in_0_1;
      end else if (10'hc9 == _T_15[9:0]) begin
        image_0_201 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_202 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hca == _T_37[9:0]) begin
        image_0_202 <= io_pixelVal_in_0_7;
      end else if (10'hca == _T_34[9:0]) begin
        image_0_202 <= io_pixelVal_in_0_6;
      end else if (10'hca == _T_31[9:0]) begin
        image_0_202 <= io_pixelVal_in_0_5;
      end else if (10'hca == _T_28[9:0]) begin
        image_0_202 <= io_pixelVal_in_0_4;
      end else if (10'hca == _T_25[9:0]) begin
        image_0_202 <= io_pixelVal_in_0_3;
      end else if (10'hca == _T_22[9:0]) begin
        image_0_202 <= io_pixelVal_in_0_2;
      end else if (10'hca == _T_19[9:0]) begin
        image_0_202 <= io_pixelVal_in_0_1;
      end else if (10'hca == _T_15[9:0]) begin
        image_0_202 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_203 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hcb == _T_37[9:0]) begin
        image_0_203 <= io_pixelVal_in_0_7;
      end else if (10'hcb == _T_34[9:0]) begin
        image_0_203 <= io_pixelVal_in_0_6;
      end else if (10'hcb == _T_31[9:0]) begin
        image_0_203 <= io_pixelVal_in_0_5;
      end else if (10'hcb == _T_28[9:0]) begin
        image_0_203 <= io_pixelVal_in_0_4;
      end else if (10'hcb == _T_25[9:0]) begin
        image_0_203 <= io_pixelVal_in_0_3;
      end else if (10'hcb == _T_22[9:0]) begin
        image_0_203 <= io_pixelVal_in_0_2;
      end else if (10'hcb == _T_19[9:0]) begin
        image_0_203 <= io_pixelVal_in_0_1;
      end else if (10'hcb == _T_15[9:0]) begin
        image_0_203 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_204 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hcc == _T_37[9:0]) begin
        image_0_204 <= io_pixelVal_in_0_7;
      end else if (10'hcc == _T_34[9:0]) begin
        image_0_204 <= io_pixelVal_in_0_6;
      end else if (10'hcc == _T_31[9:0]) begin
        image_0_204 <= io_pixelVal_in_0_5;
      end else if (10'hcc == _T_28[9:0]) begin
        image_0_204 <= io_pixelVal_in_0_4;
      end else if (10'hcc == _T_25[9:0]) begin
        image_0_204 <= io_pixelVal_in_0_3;
      end else if (10'hcc == _T_22[9:0]) begin
        image_0_204 <= io_pixelVal_in_0_2;
      end else if (10'hcc == _T_19[9:0]) begin
        image_0_204 <= io_pixelVal_in_0_1;
      end else if (10'hcc == _T_15[9:0]) begin
        image_0_204 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_205 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hcd == _T_37[9:0]) begin
        image_0_205 <= io_pixelVal_in_0_7;
      end else if (10'hcd == _T_34[9:0]) begin
        image_0_205 <= io_pixelVal_in_0_6;
      end else if (10'hcd == _T_31[9:0]) begin
        image_0_205 <= io_pixelVal_in_0_5;
      end else if (10'hcd == _T_28[9:0]) begin
        image_0_205 <= io_pixelVal_in_0_4;
      end else if (10'hcd == _T_25[9:0]) begin
        image_0_205 <= io_pixelVal_in_0_3;
      end else if (10'hcd == _T_22[9:0]) begin
        image_0_205 <= io_pixelVal_in_0_2;
      end else if (10'hcd == _T_19[9:0]) begin
        image_0_205 <= io_pixelVal_in_0_1;
      end else if (10'hcd == _T_15[9:0]) begin
        image_0_205 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_206 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hce == _T_37[9:0]) begin
        image_0_206 <= io_pixelVal_in_0_7;
      end else if (10'hce == _T_34[9:0]) begin
        image_0_206 <= io_pixelVal_in_0_6;
      end else if (10'hce == _T_31[9:0]) begin
        image_0_206 <= io_pixelVal_in_0_5;
      end else if (10'hce == _T_28[9:0]) begin
        image_0_206 <= io_pixelVal_in_0_4;
      end else if (10'hce == _T_25[9:0]) begin
        image_0_206 <= io_pixelVal_in_0_3;
      end else if (10'hce == _T_22[9:0]) begin
        image_0_206 <= io_pixelVal_in_0_2;
      end else if (10'hce == _T_19[9:0]) begin
        image_0_206 <= io_pixelVal_in_0_1;
      end else if (10'hce == _T_15[9:0]) begin
        image_0_206 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_207 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hcf == _T_37[9:0]) begin
        image_0_207 <= io_pixelVal_in_0_7;
      end else if (10'hcf == _T_34[9:0]) begin
        image_0_207 <= io_pixelVal_in_0_6;
      end else if (10'hcf == _T_31[9:0]) begin
        image_0_207 <= io_pixelVal_in_0_5;
      end else if (10'hcf == _T_28[9:0]) begin
        image_0_207 <= io_pixelVal_in_0_4;
      end else if (10'hcf == _T_25[9:0]) begin
        image_0_207 <= io_pixelVal_in_0_3;
      end else if (10'hcf == _T_22[9:0]) begin
        image_0_207 <= io_pixelVal_in_0_2;
      end else if (10'hcf == _T_19[9:0]) begin
        image_0_207 <= io_pixelVal_in_0_1;
      end else if (10'hcf == _T_15[9:0]) begin
        image_0_207 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_208 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hd0 == _T_37[9:0]) begin
        image_0_208 <= io_pixelVal_in_0_7;
      end else if (10'hd0 == _T_34[9:0]) begin
        image_0_208 <= io_pixelVal_in_0_6;
      end else if (10'hd0 == _T_31[9:0]) begin
        image_0_208 <= io_pixelVal_in_0_5;
      end else if (10'hd0 == _T_28[9:0]) begin
        image_0_208 <= io_pixelVal_in_0_4;
      end else if (10'hd0 == _T_25[9:0]) begin
        image_0_208 <= io_pixelVal_in_0_3;
      end else if (10'hd0 == _T_22[9:0]) begin
        image_0_208 <= io_pixelVal_in_0_2;
      end else if (10'hd0 == _T_19[9:0]) begin
        image_0_208 <= io_pixelVal_in_0_1;
      end else if (10'hd0 == _T_15[9:0]) begin
        image_0_208 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_209 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hd1 == _T_37[9:0]) begin
        image_0_209 <= io_pixelVal_in_0_7;
      end else if (10'hd1 == _T_34[9:0]) begin
        image_0_209 <= io_pixelVal_in_0_6;
      end else if (10'hd1 == _T_31[9:0]) begin
        image_0_209 <= io_pixelVal_in_0_5;
      end else if (10'hd1 == _T_28[9:0]) begin
        image_0_209 <= io_pixelVal_in_0_4;
      end else if (10'hd1 == _T_25[9:0]) begin
        image_0_209 <= io_pixelVal_in_0_3;
      end else if (10'hd1 == _T_22[9:0]) begin
        image_0_209 <= io_pixelVal_in_0_2;
      end else if (10'hd1 == _T_19[9:0]) begin
        image_0_209 <= io_pixelVal_in_0_1;
      end else if (10'hd1 == _T_15[9:0]) begin
        image_0_209 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_210 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hd2 == _T_37[9:0]) begin
        image_0_210 <= io_pixelVal_in_0_7;
      end else if (10'hd2 == _T_34[9:0]) begin
        image_0_210 <= io_pixelVal_in_0_6;
      end else if (10'hd2 == _T_31[9:0]) begin
        image_0_210 <= io_pixelVal_in_0_5;
      end else if (10'hd2 == _T_28[9:0]) begin
        image_0_210 <= io_pixelVal_in_0_4;
      end else if (10'hd2 == _T_25[9:0]) begin
        image_0_210 <= io_pixelVal_in_0_3;
      end else if (10'hd2 == _T_22[9:0]) begin
        image_0_210 <= io_pixelVal_in_0_2;
      end else if (10'hd2 == _T_19[9:0]) begin
        image_0_210 <= io_pixelVal_in_0_1;
      end else if (10'hd2 == _T_15[9:0]) begin
        image_0_210 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_211 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hd3 == _T_37[9:0]) begin
        image_0_211 <= io_pixelVal_in_0_7;
      end else if (10'hd3 == _T_34[9:0]) begin
        image_0_211 <= io_pixelVal_in_0_6;
      end else if (10'hd3 == _T_31[9:0]) begin
        image_0_211 <= io_pixelVal_in_0_5;
      end else if (10'hd3 == _T_28[9:0]) begin
        image_0_211 <= io_pixelVal_in_0_4;
      end else if (10'hd3 == _T_25[9:0]) begin
        image_0_211 <= io_pixelVal_in_0_3;
      end else if (10'hd3 == _T_22[9:0]) begin
        image_0_211 <= io_pixelVal_in_0_2;
      end else if (10'hd3 == _T_19[9:0]) begin
        image_0_211 <= io_pixelVal_in_0_1;
      end else if (10'hd3 == _T_15[9:0]) begin
        image_0_211 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_212 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hd4 == _T_37[9:0]) begin
        image_0_212 <= io_pixelVal_in_0_7;
      end else if (10'hd4 == _T_34[9:0]) begin
        image_0_212 <= io_pixelVal_in_0_6;
      end else if (10'hd4 == _T_31[9:0]) begin
        image_0_212 <= io_pixelVal_in_0_5;
      end else if (10'hd4 == _T_28[9:0]) begin
        image_0_212 <= io_pixelVal_in_0_4;
      end else if (10'hd4 == _T_25[9:0]) begin
        image_0_212 <= io_pixelVal_in_0_3;
      end else if (10'hd4 == _T_22[9:0]) begin
        image_0_212 <= io_pixelVal_in_0_2;
      end else if (10'hd4 == _T_19[9:0]) begin
        image_0_212 <= io_pixelVal_in_0_1;
      end else if (10'hd4 == _T_15[9:0]) begin
        image_0_212 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_213 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hd5 == _T_37[9:0]) begin
        image_0_213 <= io_pixelVal_in_0_7;
      end else if (10'hd5 == _T_34[9:0]) begin
        image_0_213 <= io_pixelVal_in_0_6;
      end else if (10'hd5 == _T_31[9:0]) begin
        image_0_213 <= io_pixelVal_in_0_5;
      end else if (10'hd5 == _T_28[9:0]) begin
        image_0_213 <= io_pixelVal_in_0_4;
      end else if (10'hd5 == _T_25[9:0]) begin
        image_0_213 <= io_pixelVal_in_0_3;
      end else if (10'hd5 == _T_22[9:0]) begin
        image_0_213 <= io_pixelVal_in_0_2;
      end else if (10'hd5 == _T_19[9:0]) begin
        image_0_213 <= io_pixelVal_in_0_1;
      end else if (10'hd5 == _T_15[9:0]) begin
        image_0_213 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_214 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hd6 == _T_37[9:0]) begin
        image_0_214 <= io_pixelVal_in_0_7;
      end else if (10'hd6 == _T_34[9:0]) begin
        image_0_214 <= io_pixelVal_in_0_6;
      end else if (10'hd6 == _T_31[9:0]) begin
        image_0_214 <= io_pixelVal_in_0_5;
      end else if (10'hd6 == _T_28[9:0]) begin
        image_0_214 <= io_pixelVal_in_0_4;
      end else if (10'hd6 == _T_25[9:0]) begin
        image_0_214 <= io_pixelVal_in_0_3;
      end else if (10'hd6 == _T_22[9:0]) begin
        image_0_214 <= io_pixelVal_in_0_2;
      end else if (10'hd6 == _T_19[9:0]) begin
        image_0_214 <= io_pixelVal_in_0_1;
      end else if (10'hd6 == _T_15[9:0]) begin
        image_0_214 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_215 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hd7 == _T_37[9:0]) begin
        image_0_215 <= io_pixelVal_in_0_7;
      end else if (10'hd7 == _T_34[9:0]) begin
        image_0_215 <= io_pixelVal_in_0_6;
      end else if (10'hd7 == _T_31[9:0]) begin
        image_0_215 <= io_pixelVal_in_0_5;
      end else if (10'hd7 == _T_28[9:0]) begin
        image_0_215 <= io_pixelVal_in_0_4;
      end else if (10'hd7 == _T_25[9:0]) begin
        image_0_215 <= io_pixelVal_in_0_3;
      end else if (10'hd7 == _T_22[9:0]) begin
        image_0_215 <= io_pixelVal_in_0_2;
      end else if (10'hd7 == _T_19[9:0]) begin
        image_0_215 <= io_pixelVal_in_0_1;
      end else if (10'hd7 == _T_15[9:0]) begin
        image_0_215 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_216 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hd8 == _T_37[9:0]) begin
        image_0_216 <= io_pixelVal_in_0_7;
      end else if (10'hd8 == _T_34[9:0]) begin
        image_0_216 <= io_pixelVal_in_0_6;
      end else if (10'hd8 == _T_31[9:0]) begin
        image_0_216 <= io_pixelVal_in_0_5;
      end else if (10'hd8 == _T_28[9:0]) begin
        image_0_216 <= io_pixelVal_in_0_4;
      end else if (10'hd8 == _T_25[9:0]) begin
        image_0_216 <= io_pixelVal_in_0_3;
      end else if (10'hd8 == _T_22[9:0]) begin
        image_0_216 <= io_pixelVal_in_0_2;
      end else if (10'hd8 == _T_19[9:0]) begin
        image_0_216 <= io_pixelVal_in_0_1;
      end else if (10'hd8 == _T_15[9:0]) begin
        image_0_216 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_217 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hd9 == _T_37[9:0]) begin
        image_0_217 <= io_pixelVal_in_0_7;
      end else if (10'hd9 == _T_34[9:0]) begin
        image_0_217 <= io_pixelVal_in_0_6;
      end else if (10'hd9 == _T_31[9:0]) begin
        image_0_217 <= io_pixelVal_in_0_5;
      end else if (10'hd9 == _T_28[9:0]) begin
        image_0_217 <= io_pixelVal_in_0_4;
      end else if (10'hd9 == _T_25[9:0]) begin
        image_0_217 <= io_pixelVal_in_0_3;
      end else if (10'hd9 == _T_22[9:0]) begin
        image_0_217 <= io_pixelVal_in_0_2;
      end else if (10'hd9 == _T_19[9:0]) begin
        image_0_217 <= io_pixelVal_in_0_1;
      end else if (10'hd9 == _T_15[9:0]) begin
        image_0_217 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_218 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hda == _T_37[9:0]) begin
        image_0_218 <= io_pixelVal_in_0_7;
      end else if (10'hda == _T_34[9:0]) begin
        image_0_218 <= io_pixelVal_in_0_6;
      end else if (10'hda == _T_31[9:0]) begin
        image_0_218 <= io_pixelVal_in_0_5;
      end else if (10'hda == _T_28[9:0]) begin
        image_0_218 <= io_pixelVal_in_0_4;
      end else if (10'hda == _T_25[9:0]) begin
        image_0_218 <= io_pixelVal_in_0_3;
      end else if (10'hda == _T_22[9:0]) begin
        image_0_218 <= io_pixelVal_in_0_2;
      end else if (10'hda == _T_19[9:0]) begin
        image_0_218 <= io_pixelVal_in_0_1;
      end else if (10'hda == _T_15[9:0]) begin
        image_0_218 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_219 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hdb == _T_37[9:0]) begin
        image_0_219 <= io_pixelVal_in_0_7;
      end else if (10'hdb == _T_34[9:0]) begin
        image_0_219 <= io_pixelVal_in_0_6;
      end else if (10'hdb == _T_31[9:0]) begin
        image_0_219 <= io_pixelVal_in_0_5;
      end else if (10'hdb == _T_28[9:0]) begin
        image_0_219 <= io_pixelVal_in_0_4;
      end else if (10'hdb == _T_25[9:0]) begin
        image_0_219 <= io_pixelVal_in_0_3;
      end else if (10'hdb == _T_22[9:0]) begin
        image_0_219 <= io_pixelVal_in_0_2;
      end else if (10'hdb == _T_19[9:0]) begin
        image_0_219 <= io_pixelVal_in_0_1;
      end else if (10'hdb == _T_15[9:0]) begin
        image_0_219 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_220 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hdc == _T_37[9:0]) begin
        image_0_220 <= io_pixelVal_in_0_7;
      end else if (10'hdc == _T_34[9:0]) begin
        image_0_220 <= io_pixelVal_in_0_6;
      end else if (10'hdc == _T_31[9:0]) begin
        image_0_220 <= io_pixelVal_in_0_5;
      end else if (10'hdc == _T_28[9:0]) begin
        image_0_220 <= io_pixelVal_in_0_4;
      end else if (10'hdc == _T_25[9:0]) begin
        image_0_220 <= io_pixelVal_in_0_3;
      end else if (10'hdc == _T_22[9:0]) begin
        image_0_220 <= io_pixelVal_in_0_2;
      end else if (10'hdc == _T_19[9:0]) begin
        image_0_220 <= io_pixelVal_in_0_1;
      end else if (10'hdc == _T_15[9:0]) begin
        image_0_220 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_221 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hdd == _T_37[9:0]) begin
        image_0_221 <= io_pixelVal_in_0_7;
      end else if (10'hdd == _T_34[9:0]) begin
        image_0_221 <= io_pixelVal_in_0_6;
      end else if (10'hdd == _T_31[9:0]) begin
        image_0_221 <= io_pixelVal_in_0_5;
      end else if (10'hdd == _T_28[9:0]) begin
        image_0_221 <= io_pixelVal_in_0_4;
      end else if (10'hdd == _T_25[9:0]) begin
        image_0_221 <= io_pixelVal_in_0_3;
      end else if (10'hdd == _T_22[9:0]) begin
        image_0_221 <= io_pixelVal_in_0_2;
      end else if (10'hdd == _T_19[9:0]) begin
        image_0_221 <= io_pixelVal_in_0_1;
      end else if (10'hdd == _T_15[9:0]) begin
        image_0_221 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_222 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hde == _T_37[9:0]) begin
        image_0_222 <= io_pixelVal_in_0_7;
      end else if (10'hde == _T_34[9:0]) begin
        image_0_222 <= io_pixelVal_in_0_6;
      end else if (10'hde == _T_31[9:0]) begin
        image_0_222 <= io_pixelVal_in_0_5;
      end else if (10'hde == _T_28[9:0]) begin
        image_0_222 <= io_pixelVal_in_0_4;
      end else if (10'hde == _T_25[9:0]) begin
        image_0_222 <= io_pixelVal_in_0_3;
      end else if (10'hde == _T_22[9:0]) begin
        image_0_222 <= io_pixelVal_in_0_2;
      end else if (10'hde == _T_19[9:0]) begin
        image_0_222 <= io_pixelVal_in_0_1;
      end else if (10'hde == _T_15[9:0]) begin
        image_0_222 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_223 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hdf == _T_37[9:0]) begin
        image_0_223 <= io_pixelVal_in_0_7;
      end else if (10'hdf == _T_34[9:0]) begin
        image_0_223 <= io_pixelVal_in_0_6;
      end else if (10'hdf == _T_31[9:0]) begin
        image_0_223 <= io_pixelVal_in_0_5;
      end else if (10'hdf == _T_28[9:0]) begin
        image_0_223 <= io_pixelVal_in_0_4;
      end else if (10'hdf == _T_25[9:0]) begin
        image_0_223 <= io_pixelVal_in_0_3;
      end else if (10'hdf == _T_22[9:0]) begin
        image_0_223 <= io_pixelVal_in_0_2;
      end else if (10'hdf == _T_19[9:0]) begin
        image_0_223 <= io_pixelVal_in_0_1;
      end else if (10'hdf == _T_15[9:0]) begin
        image_0_223 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_224 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'he0 == _T_37[9:0]) begin
        image_0_224 <= io_pixelVal_in_0_7;
      end else if (10'he0 == _T_34[9:0]) begin
        image_0_224 <= io_pixelVal_in_0_6;
      end else if (10'he0 == _T_31[9:0]) begin
        image_0_224 <= io_pixelVal_in_0_5;
      end else if (10'he0 == _T_28[9:0]) begin
        image_0_224 <= io_pixelVal_in_0_4;
      end else if (10'he0 == _T_25[9:0]) begin
        image_0_224 <= io_pixelVal_in_0_3;
      end else if (10'he0 == _T_22[9:0]) begin
        image_0_224 <= io_pixelVal_in_0_2;
      end else if (10'he0 == _T_19[9:0]) begin
        image_0_224 <= io_pixelVal_in_0_1;
      end else if (10'he0 == _T_15[9:0]) begin
        image_0_224 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_225 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'he1 == _T_37[9:0]) begin
        image_0_225 <= io_pixelVal_in_0_7;
      end else if (10'he1 == _T_34[9:0]) begin
        image_0_225 <= io_pixelVal_in_0_6;
      end else if (10'he1 == _T_31[9:0]) begin
        image_0_225 <= io_pixelVal_in_0_5;
      end else if (10'he1 == _T_28[9:0]) begin
        image_0_225 <= io_pixelVal_in_0_4;
      end else if (10'he1 == _T_25[9:0]) begin
        image_0_225 <= io_pixelVal_in_0_3;
      end else if (10'he1 == _T_22[9:0]) begin
        image_0_225 <= io_pixelVal_in_0_2;
      end else if (10'he1 == _T_19[9:0]) begin
        image_0_225 <= io_pixelVal_in_0_1;
      end else if (10'he1 == _T_15[9:0]) begin
        image_0_225 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_226 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'he2 == _T_37[9:0]) begin
        image_0_226 <= io_pixelVal_in_0_7;
      end else if (10'he2 == _T_34[9:0]) begin
        image_0_226 <= io_pixelVal_in_0_6;
      end else if (10'he2 == _T_31[9:0]) begin
        image_0_226 <= io_pixelVal_in_0_5;
      end else if (10'he2 == _T_28[9:0]) begin
        image_0_226 <= io_pixelVal_in_0_4;
      end else if (10'he2 == _T_25[9:0]) begin
        image_0_226 <= io_pixelVal_in_0_3;
      end else if (10'he2 == _T_22[9:0]) begin
        image_0_226 <= io_pixelVal_in_0_2;
      end else if (10'he2 == _T_19[9:0]) begin
        image_0_226 <= io_pixelVal_in_0_1;
      end else if (10'he2 == _T_15[9:0]) begin
        image_0_226 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_227 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'he3 == _T_37[9:0]) begin
        image_0_227 <= io_pixelVal_in_0_7;
      end else if (10'he3 == _T_34[9:0]) begin
        image_0_227 <= io_pixelVal_in_0_6;
      end else if (10'he3 == _T_31[9:0]) begin
        image_0_227 <= io_pixelVal_in_0_5;
      end else if (10'he3 == _T_28[9:0]) begin
        image_0_227 <= io_pixelVal_in_0_4;
      end else if (10'he3 == _T_25[9:0]) begin
        image_0_227 <= io_pixelVal_in_0_3;
      end else if (10'he3 == _T_22[9:0]) begin
        image_0_227 <= io_pixelVal_in_0_2;
      end else if (10'he3 == _T_19[9:0]) begin
        image_0_227 <= io_pixelVal_in_0_1;
      end else if (10'he3 == _T_15[9:0]) begin
        image_0_227 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_228 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'he4 == _T_37[9:0]) begin
        image_0_228 <= io_pixelVal_in_0_7;
      end else if (10'he4 == _T_34[9:0]) begin
        image_0_228 <= io_pixelVal_in_0_6;
      end else if (10'he4 == _T_31[9:0]) begin
        image_0_228 <= io_pixelVal_in_0_5;
      end else if (10'he4 == _T_28[9:0]) begin
        image_0_228 <= io_pixelVal_in_0_4;
      end else if (10'he4 == _T_25[9:0]) begin
        image_0_228 <= io_pixelVal_in_0_3;
      end else if (10'he4 == _T_22[9:0]) begin
        image_0_228 <= io_pixelVal_in_0_2;
      end else if (10'he4 == _T_19[9:0]) begin
        image_0_228 <= io_pixelVal_in_0_1;
      end else if (10'he4 == _T_15[9:0]) begin
        image_0_228 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_229 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'he5 == _T_37[9:0]) begin
        image_0_229 <= io_pixelVal_in_0_7;
      end else if (10'he5 == _T_34[9:0]) begin
        image_0_229 <= io_pixelVal_in_0_6;
      end else if (10'he5 == _T_31[9:0]) begin
        image_0_229 <= io_pixelVal_in_0_5;
      end else if (10'he5 == _T_28[9:0]) begin
        image_0_229 <= io_pixelVal_in_0_4;
      end else if (10'he5 == _T_25[9:0]) begin
        image_0_229 <= io_pixelVal_in_0_3;
      end else if (10'he5 == _T_22[9:0]) begin
        image_0_229 <= io_pixelVal_in_0_2;
      end else if (10'he5 == _T_19[9:0]) begin
        image_0_229 <= io_pixelVal_in_0_1;
      end else if (10'he5 == _T_15[9:0]) begin
        image_0_229 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_230 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'he6 == _T_37[9:0]) begin
        image_0_230 <= io_pixelVal_in_0_7;
      end else if (10'he6 == _T_34[9:0]) begin
        image_0_230 <= io_pixelVal_in_0_6;
      end else if (10'he6 == _T_31[9:0]) begin
        image_0_230 <= io_pixelVal_in_0_5;
      end else if (10'he6 == _T_28[9:0]) begin
        image_0_230 <= io_pixelVal_in_0_4;
      end else if (10'he6 == _T_25[9:0]) begin
        image_0_230 <= io_pixelVal_in_0_3;
      end else if (10'he6 == _T_22[9:0]) begin
        image_0_230 <= io_pixelVal_in_0_2;
      end else if (10'he6 == _T_19[9:0]) begin
        image_0_230 <= io_pixelVal_in_0_1;
      end else if (10'he6 == _T_15[9:0]) begin
        image_0_230 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_231 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'he7 == _T_37[9:0]) begin
        image_0_231 <= io_pixelVal_in_0_7;
      end else if (10'he7 == _T_34[9:0]) begin
        image_0_231 <= io_pixelVal_in_0_6;
      end else if (10'he7 == _T_31[9:0]) begin
        image_0_231 <= io_pixelVal_in_0_5;
      end else if (10'he7 == _T_28[9:0]) begin
        image_0_231 <= io_pixelVal_in_0_4;
      end else if (10'he7 == _T_25[9:0]) begin
        image_0_231 <= io_pixelVal_in_0_3;
      end else if (10'he7 == _T_22[9:0]) begin
        image_0_231 <= io_pixelVal_in_0_2;
      end else if (10'he7 == _T_19[9:0]) begin
        image_0_231 <= io_pixelVal_in_0_1;
      end else if (10'he7 == _T_15[9:0]) begin
        image_0_231 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_232 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'he8 == _T_37[9:0]) begin
        image_0_232 <= io_pixelVal_in_0_7;
      end else if (10'he8 == _T_34[9:0]) begin
        image_0_232 <= io_pixelVal_in_0_6;
      end else if (10'he8 == _T_31[9:0]) begin
        image_0_232 <= io_pixelVal_in_0_5;
      end else if (10'he8 == _T_28[9:0]) begin
        image_0_232 <= io_pixelVal_in_0_4;
      end else if (10'he8 == _T_25[9:0]) begin
        image_0_232 <= io_pixelVal_in_0_3;
      end else if (10'he8 == _T_22[9:0]) begin
        image_0_232 <= io_pixelVal_in_0_2;
      end else if (10'he8 == _T_19[9:0]) begin
        image_0_232 <= io_pixelVal_in_0_1;
      end else if (10'he8 == _T_15[9:0]) begin
        image_0_232 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_233 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'he9 == _T_37[9:0]) begin
        image_0_233 <= io_pixelVal_in_0_7;
      end else if (10'he9 == _T_34[9:0]) begin
        image_0_233 <= io_pixelVal_in_0_6;
      end else if (10'he9 == _T_31[9:0]) begin
        image_0_233 <= io_pixelVal_in_0_5;
      end else if (10'he9 == _T_28[9:0]) begin
        image_0_233 <= io_pixelVal_in_0_4;
      end else if (10'he9 == _T_25[9:0]) begin
        image_0_233 <= io_pixelVal_in_0_3;
      end else if (10'he9 == _T_22[9:0]) begin
        image_0_233 <= io_pixelVal_in_0_2;
      end else if (10'he9 == _T_19[9:0]) begin
        image_0_233 <= io_pixelVal_in_0_1;
      end else if (10'he9 == _T_15[9:0]) begin
        image_0_233 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_234 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hea == _T_37[9:0]) begin
        image_0_234 <= io_pixelVal_in_0_7;
      end else if (10'hea == _T_34[9:0]) begin
        image_0_234 <= io_pixelVal_in_0_6;
      end else if (10'hea == _T_31[9:0]) begin
        image_0_234 <= io_pixelVal_in_0_5;
      end else if (10'hea == _T_28[9:0]) begin
        image_0_234 <= io_pixelVal_in_0_4;
      end else if (10'hea == _T_25[9:0]) begin
        image_0_234 <= io_pixelVal_in_0_3;
      end else if (10'hea == _T_22[9:0]) begin
        image_0_234 <= io_pixelVal_in_0_2;
      end else if (10'hea == _T_19[9:0]) begin
        image_0_234 <= io_pixelVal_in_0_1;
      end else if (10'hea == _T_15[9:0]) begin
        image_0_234 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_235 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'heb == _T_37[9:0]) begin
        image_0_235 <= io_pixelVal_in_0_7;
      end else if (10'heb == _T_34[9:0]) begin
        image_0_235 <= io_pixelVal_in_0_6;
      end else if (10'heb == _T_31[9:0]) begin
        image_0_235 <= io_pixelVal_in_0_5;
      end else if (10'heb == _T_28[9:0]) begin
        image_0_235 <= io_pixelVal_in_0_4;
      end else if (10'heb == _T_25[9:0]) begin
        image_0_235 <= io_pixelVal_in_0_3;
      end else if (10'heb == _T_22[9:0]) begin
        image_0_235 <= io_pixelVal_in_0_2;
      end else if (10'heb == _T_19[9:0]) begin
        image_0_235 <= io_pixelVal_in_0_1;
      end else if (10'heb == _T_15[9:0]) begin
        image_0_235 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_236 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hec == _T_37[9:0]) begin
        image_0_236 <= io_pixelVal_in_0_7;
      end else if (10'hec == _T_34[9:0]) begin
        image_0_236 <= io_pixelVal_in_0_6;
      end else if (10'hec == _T_31[9:0]) begin
        image_0_236 <= io_pixelVal_in_0_5;
      end else if (10'hec == _T_28[9:0]) begin
        image_0_236 <= io_pixelVal_in_0_4;
      end else if (10'hec == _T_25[9:0]) begin
        image_0_236 <= io_pixelVal_in_0_3;
      end else if (10'hec == _T_22[9:0]) begin
        image_0_236 <= io_pixelVal_in_0_2;
      end else if (10'hec == _T_19[9:0]) begin
        image_0_236 <= io_pixelVal_in_0_1;
      end else if (10'hec == _T_15[9:0]) begin
        image_0_236 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_237 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hed == _T_37[9:0]) begin
        image_0_237 <= io_pixelVal_in_0_7;
      end else if (10'hed == _T_34[9:0]) begin
        image_0_237 <= io_pixelVal_in_0_6;
      end else if (10'hed == _T_31[9:0]) begin
        image_0_237 <= io_pixelVal_in_0_5;
      end else if (10'hed == _T_28[9:0]) begin
        image_0_237 <= io_pixelVal_in_0_4;
      end else if (10'hed == _T_25[9:0]) begin
        image_0_237 <= io_pixelVal_in_0_3;
      end else if (10'hed == _T_22[9:0]) begin
        image_0_237 <= io_pixelVal_in_0_2;
      end else if (10'hed == _T_19[9:0]) begin
        image_0_237 <= io_pixelVal_in_0_1;
      end else if (10'hed == _T_15[9:0]) begin
        image_0_237 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_238 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hee == _T_37[9:0]) begin
        image_0_238 <= io_pixelVal_in_0_7;
      end else if (10'hee == _T_34[9:0]) begin
        image_0_238 <= io_pixelVal_in_0_6;
      end else if (10'hee == _T_31[9:0]) begin
        image_0_238 <= io_pixelVal_in_0_5;
      end else if (10'hee == _T_28[9:0]) begin
        image_0_238 <= io_pixelVal_in_0_4;
      end else if (10'hee == _T_25[9:0]) begin
        image_0_238 <= io_pixelVal_in_0_3;
      end else if (10'hee == _T_22[9:0]) begin
        image_0_238 <= io_pixelVal_in_0_2;
      end else if (10'hee == _T_19[9:0]) begin
        image_0_238 <= io_pixelVal_in_0_1;
      end else if (10'hee == _T_15[9:0]) begin
        image_0_238 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_239 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hef == _T_37[9:0]) begin
        image_0_239 <= io_pixelVal_in_0_7;
      end else if (10'hef == _T_34[9:0]) begin
        image_0_239 <= io_pixelVal_in_0_6;
      end else if (10'hef == _T_31[9:0]) begin
        image_0_239 <= io_pixelVal_in_0_5;
      end else if (10'hef == _T_28[9:0]) begin
        image_0_239 <= io_pixelVal_in_0_4;
      end else if (10'hef == _T_25[9:0]) begin
        image_0_239 <= io_pixelVal_in_0_3;
      end else if (10'hef == _T_22[9:0]) begin
        image_0_239 <= io_pixelVal_in_0_2;
      end else if (10'hef == _T_19[9:0]) begin
        image_0_239 <= io_pixelVal_in_0_1;
      end else if (10'hef == _T_15[9:0]) begin
        image_0_239 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_240 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hf0 == _T_37[9:0]) begin
        image_0_240 <= io_pixelVal_in_0_7;
      end else if (10'hf0 == _T_34[9:0]) begin
        image_0_240 <= io_pixelVal_in_0_6;
      end else if (10'hf0 == _T_31[9:0]) begin
        image_0_240 <= io_pixelVal_in_0_5;
      end else if (10'hf0 == _T_28[9:0]) begin
        image_0_240 <= io_pixelVal_in_0_4;
      end else if (10'hf0 == _T_25[9:0]) begin
        image_0_240 <= io_pixelVal_in_0_3;
      end else if (10'hf0 == _T_22[9:0]) begin
        image_0_240 <= io_pixelVal_in_0_2;
      end else if (10'hf0 == _T_19[9:0]) begin
        image_0_240 <= io_pixelVal_in_0_1;
      end else if (10'hf0 == _T_15[9:0]) begin
        image_0_240 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_241 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hf1 == _T_37[9:0]) begin
        image_0_241 <= io_pixelVal_in_0_7;
      end else if (10'hf1 == _T_34[9:0]) begin
        image_0_241 <= io_pixelVal_in_0_6;
      end else if (10'hf1 == _T_31[9:0]) begin
        image_0_241 <= io_pixelVal_in_0_5;
      end else if (10'hf1 == _T_28[9:0]) begin
        image_0_241 <= io_pixelVal_in_0_4;
      end else if (10'hf1 == _T_25[9:0]) begin
        image_0_241 <= io_pixelVal_in_0_3;
      end else if (10'hf1 == _T_22[9:0]) begin
        image_0_241 <= io_pixelVal_in_0_2;
      end else if (10'hf1 == _T_19[9:0]) begin
        image_0_241 <= io_pixelVal_in_0_1;
      end else if (10'hf1 == _T_15[9:0]) begin
        image_0_241 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_242 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hf2 == _T_37[9:0]) begin
        image_0_242 <= io_pixelVal_in_0_7;
      end else if (10'hf2 == _T_34[9:0]) begin
        image_0_242 <= io_pixelVal_in_0_6;
      end else if (10'hf2 == _T_31[9:0]) begin
        image_0_242 <= io_pixelVal_in_0_5;
      end else if (10'hf2 == _T_28[9:0]) begin
        image_0_242 <= io_pixelVal_in_0_4;
      end else if (10'hf2 == _T_25[9:0]) begin
        image_0_242 <= io_pixelVal_in_0_3;
      end else if (10'hf2 == _T_22[9:0]) begin
        image_0_242 <= io_pixelVal_in_0_2;
      end else if (10'hf2 == _T_19[9:0]) begin
        image_0_242 <= io_pixelVal_in_0_1;
      end else if (10'hf2 == _T_15[9:0]) begin
        image_0_242 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_243 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hf3 == _T_37[9:0]) begin
        image_0_243 <= io_pixelVal_in_0_7;
      end else if (10'hf3 == _T_34[9:0]) begin
        image_0_243 <= io_pixelVal_in_0_6;
      end else if (10'hf3 == _T_31[9:0]) begin
        image_0_243 <= io_pixelVal_in_0_5;
      end else if (10'hf3 == _T_28[9:0]) begin
        image_0_243 <= io_pixelVal_in_0_4;
      end else if (10'hf3 == _T_25[9:0]) begin
        image_0_243 <= io_pixelVal_in_0_3;
      end else if (10'hf3 == _T_22[9:0]) begin
        image_0_243 <= io_pixelVal_in_0_2;
      end else if (10'hf3 == _T_19[9:0]) begin
        image_0_243 <= io_pixelVal_in_0_1;
      end else if (10'hf3 == _T_15[9:0]) begin
        image_0_243 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_244 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hf4 == _T_37[9:0]) begin
        image_0_244 <= io_pixelVal_in_0_7;
      end else if (10'hf4 == _T_34[9:0]) begin
        image_0_244 <= io_pixelVal_in_0_6;
      end else if (10'hf4 == _T_31[9:0]) begin
        image_0_244 <= io_pixelVal_in_0_5;
      end else if (10'hf4 == _T_28[9:0]) begin
        image_0_244 <= io_pixelVal_in_0_4;
      end else if (10'hf4 == _T_25[9:0]) begin
        image_0_244 <= io_pixelVal_in_0_3;
      end else if (10'hf4 == _T_22[9:0]) begin
        image_0_244 <= io_pixelVal_in_0_2;
      end else if (10'hf4 == _T_19[9:0]) begin
        image_0_244 <= io_pixelVal_in_0_1;
      end else if (10'hf4 == _T_15[9:0]) begin
        image_0_244 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_245 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hf5 == _T_37[9:0]) begin
        image_0_245 <= io_pixelVal_in_0_7;
      end else if (10'hf5 == _T_34[9:0]) begin
        image_0_245 <= io_pixelVal_in_0_6;
      end else if (10'hf5 == _T_31[9:0]) begin
        image_0_245 <= io_pixelVal_in_0_5;
      end else if (10'hf5 == _T_28[9:0]) begin
        image_0_245 <= io_pixelVal_in_0_4;
      end else if (10'hf5 == _T_25[9:0]) begin
        image_0_245 <= io_pixelVal_in_0_3;
      end else if (10'hf5 == _T_22[9:0]) begin
        image_0_245 <= io_pixelVal_in_0_2;
      end else if (10'hf5 == _T_19[9:0]) begin
        image_0_245 <= io_pixelVal_in_0_1;
      end else if (10'hf5 == _T_15[9:0]) begin
        image_0_245 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_246 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hf6 == _T_37[9:0]) begin
        image_0_246 <= io_pixelVal_in_0_7;
      end else if (10'hf6 == _T_34[9:0]) begin
        image_0_246 <= io_pixelVal_in_0_6;
      end else if (10'hf6 == _T_31[9:0]) begin
        image_0_246 <= io_pixelVal_in_0_5;
      end else if (10'hf6 == _T_28[9:0]) begin
        image_0_246 <= io_pixelVal_in_0_4;
      end else if (10'hf6 == _T_25[9:0]) begin
        image_0_246 <= io_pixelVal_in_0_3;
      end else if (10'hf6 == _T_22[9:0]) begin
        image_0_246 <= io_pixelVal_in_0_2;
      end else if (10'hf6 == _T_19[9:0]) begin
        image_0_246 <= io_pixelVal_in_0_1;
      end else if (10'hf6 == _T_15[9:0]) begin
        image_0_246 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_247 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hf7 == _T_37[9:0]) begin
        image_0_247 <= io_pixelVal_in_0_7;
      end else if (10'hf7 == _T_34[9:0]) begin
        image_0_247 <= io_pixelVal_in_0_6;
      end else if (10'hf7 == _T_31[9:0]) begin
        image_0_247 <= io_pixelVal_in_0_5;
      end else if (10'hf7 == _T_28[9:0]) begin
        image_0_247 <= io_pixelVal_in_0_4;
      end else if (10'hf7 == _T_25[9:0]) begin
        image_0_247 <= io_pixelVal_in_0_3;
      end else if (10'hf7 == _T_22[9:0]) begin
        image_0_247 <= io_pixelVal_in_0_2;
      end else if (10'hf7 == _T_19[9:0]) begin
        image_0_247 <= io_pixelVal_in_0_1;
      end else if (10'hf7 == _T_15[9:0]) begin
        image_0_247 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_248 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hf8 == _T_37[9:0]) begin
        image_0_248 <= io_pixelVal_in_0_7;
      end else if (10'hf8 == _T_34[9:0]) begin
        image_0_248 <= io_pixelVal_in_0_6;
      end else if (10'hf8 == _T_31[9:0]) begin
        image_0_248 <= io_pixelVal_in_0_5;
      end else if (10'hf8 == _T_28[9:0]) begin
        image_0_248 <= io_pixelVal_in_0_4;
      end else if (10'hf8 == _T_25[9:0]) begin
        image_0_248 <= io_pixelVal_in_0_3;
      end else if (10'hf8 == _T_22[9:0]) begin
        image_0_248 <= io_pixelVal_in_0_2;
      end else if (10'hf8 == _T_19[9:0]) begin
        image_0_248 <= io_pixelVal_in_0_1;
      end else if (10'hf8 == _T_15[9:0]) begin
        image_0_248 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_249 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hf9 == _T_37[9:0]) begin
        image_0_249 <= io_pixelVal_in_0_7;
      end else if (10'hf9 == _T_34[9:0]) begin
        image_0_249 <= io_pixelVal_in_0_6;
      end else if (10'hf9 == _T_31[9:0]) begin
        image_0_249 <= io_pixelVal_in_0_5;
      end else if (10'hf9 == _T_28[9:0]) begin
        image_0_249 <= io_pixelVal_in_0_4;
      end else if (10'hf9 == _T_25[9:0]) begin
        image_0_249 <= io_pixelVal_in_0_3;
      end else if (10'hf9 == _T_22[9:0]) begin
        image_0_249 <= io_pixelVal_in_0_2;
      end else if (10'hf9 == _T_19[9:0]) begin
        image_0_249 <= io_pixelVal_in_0_1;
      end else if (10'hf9 == _T_15[9:0]) begin
        image_0_249 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_250 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hfa == _T_37[9:0]) begin
        image_0_250 <= io_pixelVal_in_0_7;
      end else if (10'hfa == _T_34[9:0]) begin
        image_0_250 <= io_pixelVal_in_0_6;
      end else if (10'hfa == _T_31[9:0]) begin
        image_0_250 <= io_pixelVal_in_0_5;
      end else if (10'hfa == _T_28[9:0]) begin
        image_0_250 <= io_pixelVal_in_0_4;
      end else if (10'hfa == _T_25[9:0]) begin
        image_0_250 <= io_pixelVal_in_0_3;
      end else if (10'hfa == _T_22[9:0]) begin
        image_0_250 <= io_pixelVal_in_0_2;
      end else if (10'hfa == _T_19[9:0]) begin
        image_0_250 <= io_pixelVal_in_0_1;
      end else if (10'hfa == _T_15[9:0]) begin
        image_0_250 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_251 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hfb == _T_37[9:0]) begin
        image_0_251 <= io_pixelVal_in_0_7;
      end else if (10'hfb == _T_34[9:0]) begin
        image_0_251 <= io_pixelVal_in_0_6;
      end else if (10'hfb == _T_31[9:0]) begin
        image_0_251 <= io_pixelVal_in_0_5;
      end else if (10'hfb == _T_28[9:0]) begin
        image_0_251 <= io_pixelVal_in_0_4;
      end else if (10'hfb == _T_25[9:0]) begin
        image_0_251 <= io_pixelVal_in_0_3;
      end else if (10'hfb == _T_22[9:0]) begin
        image_0_251 <= io_pixelVal_in_0_2;
      end else if (10'hfb == _T_19[9:0]) begin
        image_0_251 <= io_pixelVal_in_0_1;
      end else if (10'hfb == _T_15[9:0]) begin
        image_0_251 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_252 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hfc == _T_37[9:0]) begin
        image_0_252 <= io_pixelVal_in_0_7;
      end else if (10'hfc == _T_34[9:0]) begin
        image_0_252 <= io_pixelVal_in_0_6;
      end else if (10'hfc == _T_31[9:0]) begin
        image_0_252 <= io_pixelVal_in_0_5;
      end else if (10'hfc == _T_28[9:0]) begin
        image_0_252 <= io_pixelVal_in_0_4;
      end else if (10'hfc == _T_25[9:0]) begin
        image_0_252 <= io_pixelVal_in_0_3;
      end else if (10'hfc == _T_22[9:0]) begin
        image_0_252 <= io_pixelVal_in_0_2;
      end else if (10'hfc == _T_19[9:0]) begin
        image_0_252 <= io_pixelVal_in_0_1;
      end else if (10'hfc == _T_15[9:0]) begin
        image_0_252 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_253 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hfd == _T_37[9:0]) begin
        image_0_253 <= io_pixelVal_in_0_7;
      end else if (10'hfd == _T_34[9:0]) begin
        image_0_253 <= io_pixelVal_in_0_6;
      end else if (10'hfd == _T_31[9:0]) begin
        image_0_253 <= io_pixelVal_in_0_5;
      end else if (10'hfd == _T_28[9:0]) begin
        image_0_253 <= io_pixelVal_in_0_4;
      end else if (10'hfd == _T_25[9:0]) begin
        image_0_253 <= io_pixelVal_in_0_3;
      end else if (10'hfd == _T_22[9:0]) begin
        image_0_253 <= io_pixelVal_in_0_2;
      end else if (10'hfd == _T_19[9:0]) begin
        image_0_253 <= io_pixelVal_in_0_1;
      end else if (10'hfd == _T_15[9:0]) begin
        image_0_253 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_254 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hfe == _T_37[9:0]) begin
        image_0_254 <= io_pixelVal_in_0_7;
      end else if (10'hfe == _T_34[9:0]) begin
        image_0_254 <= io_pixelVal_in_0_6;
      end else if (10'hfe == _T_31[9:0]) begin
        image_0_254 <= io_pixelVal_in_0_5;
      end else if (10'hfe == _T_28[9:0]) begin
        image_0_254 <= io_pixelVal_in_0_4;
      end else if (10'hfe == _T_25[9:0]) begin
        image_0_254 <= io_pixelVal_in_0_3;
      end else if (10'hfe == _T_22[9:0]) begin
        image_0_254 <= io_pixelVal_in_0_2;
      end else if (10'hfe == _T_19[9:0]) begin
        image_0_254 <= io_pixelVal_in_0_1;
      end else if (10'hfe == _T_15[9:0]) begin
        image_0_254 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_255 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'hff == _T_37[9:0]) begin
        image_0_255 <= io_pixelVal_in_0_7;
      end else if (10'hff == _T_34[9:0]) begin
        image_0_255 <= io_pixelVal_in_0_6;
      end else if (10'hff == _T_31[9:0]) begin
        image_0_255 <= io_pixelVal_in_0_5;
      end else if (10'hff == _T_28[9:0]) begin
        image_0_255 <= io_pixelVal_in_0_4;
      end else if (10'hff == _T_25[9:0]) begin
        image_0_255 <= io_pixelVal_in_0_3;
      end else if (10'hff == _T_22[9:0]) begin
        image_0_255 <= io_pixelVal_in_0_2;
      end else if (10'hff == _T_19[9:0]) begin
        image_0_255 <= io_pixelVal_in_0_1;
      end else if (10'hff == _T_15[9:0]) begin
        image_0_255 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_256 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h100 == _T_37[9:0]) begin
        image_0_256 <= io_pixelVal_in_0_7;
      end else if (10'h100 == _T_34[9:0]) begin
        image_0_256 <= io_pixelVal_in_0_6;
      end else if (10'h100 == _T_31[9:0]) begin
        image_0_256 <= io_pixelVal_in_0_5;
      end else if (10'h100 == _T_28[9:0]) begin
        image_0_256 <= io_pixelVal_in_0_4;
      end else if (10'h100 == _T_25[9:0]) begin
        image_0_256 <= io_pixelVal_in_0_3;
      end else if (10'h100 == _T_22[9:0]) begin
        image_0_256 <= io_pixelVal_in_0_2;
      end else if (10'h100 == _T_19[9:0]) begin
        image_0_256 <= io_pixelVal_in_0_1;
      end else if (10'h100 == _T_15[9:0]) begin
        image_0_256 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_257 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h101 == _T_37[9:0]) begin
        image_0_257 <= io_pixelVal_in_0_7;
      end else if (10'h101 == _T_34[9:0]) begin
        image_0_257 <= io_pixelVal_in_0_6;
      end else if (10'h101 == _T_31[9:0]) begin
        image_0_257 <= io_pixelVal_in_0_5;
      end else if (10'h101 == _T_28[9:0]) begin
        image_0_257 <= io_pixelVal_in_0_4;
      end else if (10'h101 == _T_25[9:0]) begin
        image_0_257 <= io_pixelVal_in_0_3;
      end else if (10'h101 == _T_22[9:0]) begin
        image_0_257 <= io_pixelVal_in_0_2;
      end else if (10'h101 == _T_19[9:0]) begin
        image_0_257 <= io_pixelVal_in_0_1;
      end else if (10'h101 == _T_15[9:0]) begin
        image_0_257 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_258 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h102 == _T_37[9:0]) begin
        image_0_258 <= io_pixelVal_in_0_7;
      end else if (10'h102 == _T_34[9:0]) begin
        image_0_258 <= io_pixelVal_in_0_6;
      end else if (10'h102 == _T_31[9:0]) begin
        image_0_258 <= io_pixelVal_in_0_5;
      end else if (10'h102 == _T_28[9:0]) begin
        image_0_258 <= io_pixelVal_in_0_4;
      end else if (10'h102 == _T_25[9:0]) begin
        image_0_258 <= io_pixelVal_in_0_3;
      end else if (10'h102 == _T_22[9:0]) begin
        image_0_258 <= io_pixelVal_in_0_2;
      end else if (10'h102 == _T_19[9:0]) begin
        image_0_258 <= io_pixelVal_in_0_1;
      end else if (10'h102 == _T_15[9:0]) begin
        image_0_258 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_259 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h103 == _T_37[9:0]) begin
        image_0_259 <= io_pixelVal_in_0_7;
      end else if (10'h103 == _T_34[9:0]) begin
        image_0_259 <= io_pixelVal_in_0_6;
      end else if (10'h103 == _T_31[9:0]) begin
        image_0_259 <= io_pixelVal_in_0_5;
      end else if (10'h103 == _T_28[9:0]) begin
        image_0_259 <= io_pixelVal_in_0_4;
      end else if (10'h103 == _T_25[9:0]) begin
        image_0_259 <= io_pixelVal_in_0_3;
      end else if (10'h103 == _T_22[9:0]) begin
        image_0_259 <= io_pixelVal_in_0_2;
      end else if (10'h103 == _T_19[9:0]) begin
        image_0_259 <= io_pixelVal_in_0_1;
      end else if (10'h103 == _T_15[9:0]) begin
        image_0_259 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_260 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h104 == _T_37[9:0]) begin
        image_0_260 <= io_pixelVal_in_0_7;
      end else if (10'h104 == _T_34[9:0]) begin
        image_0_260 <= io_pixelVal_in_0_6;
      end else if (10'h104 == _T_31[9:0]) begin
        image_0_260 <= io_pixelVal_in_0_5;
      end else if (10'h104 == _T_28[9:0]) begin
        image_0_260 <= io_pixelVal_in_0_4;
      end else if (10'h104 == _T_25[9:0]) begin
        image_0_260 <= io_pixelVal_in_0_3;
      end else if (10'h104 == _T_22[9:0]) begin
        image_0_260 <= io_pixelVal_in_0_2;
      end else if (10'h104 == _T_19[9:0]) begin
        image_0_260 <= io_pixelVal_in_0_1;
      end else if (10'h104 == _T_15[9:0]) begin
        image_0_260 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_261 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h105 == _T_37[9:0]) begin
        image_0_261 <= io_pixelVal_in_0_7;
      end else if (10'h105 == _T_34[9:0]) begin
        image_0_261 <= io_pixelVal_in_0_6;
      end else if (10'h105 == _T_31[9:0]) begin
        image_0_261 <= io_pixelVal_in_0_5;
      end else if (10'h105 == _T_28[9:0]) begin
        image_0_261 <= io_pixelVal_in_0_4;
      end else if (10'h105 == _T_25[9:0]) begin
        image_0_261 <= io_pixelVal_in_0_3;
      end else if (10'h105 == _T_22[9:0]) begin
        image_0_261 <= io_pixelVal_in_0_2;
      end else if (10'h105 == _T_19[9:0]) begin
        image_0_261 <= io_pixelVal_in_0_1;
      end else if (10'h105 == _T_15[9:0]) begin
        image_0_261 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_262 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h106 == _T_37[9:0]) begin
        image_0_262 <= io_pixelVal_in_0_7;
      end else if (10'h106 == _T_34[9:0]) begin
        image_0_262 <= io_pixelVal_in_0_6;
      end else if (10'h106 == _T_31[9:0]) begin
        image_0_262 <= io_pixelVal_in_0_5;
      end else if (10'h106 == _T_28[9:0]) begin
        image_0_262 <= io_pixelVal_in_0_4;
      end else if (10'h106 == _T_25[9:0]) begin
        image_0_262 <= io_pixelVal_in_0_3;
      end else if (10'h106 == _T_22[9:0]) begin
        image_0_262 <= io_pixelVal_in_0_2;
      end else if (10'h106 == _T_19[9:0]) begin
        image_0_262 <= io_pixelVal_in_0_1;
      end else if (10'h106 == _T_15[9:0]) begin
        image_0_262 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_263 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h107 == _T_37[9:0]) begin
        image_0_263 <= io_pixelVal_in_0_7;
      end else if (10'h107 == _T_34[9:0]) begin
        image_0_263 <= io_pixelVal_in_0_6;
      end else if (10'h107 == _T_31[9:0]) begin
        image_0_263 <= io_pixelVal_in_0_5;
      end else if (10'h107 == _T_28[9:0]) begin
        image_0_263 <= io_pixelVal_in_0_4;
      end else if (10'h107 == _T_25[9:0]) begin
        image_0_263 <= io_pixelVal_in_0_3;
      end else if (10'h107 == _T_22[9:0]) begin
        image_0_263 <= io_pixelVal_in_0_2;
      end else if (10'h107 == _T_19[9:0]) begin
        image_0_263 <= io_pixelVal_in_0_1;
      end else if (10'h107 == _T_15[9:0]) begin
        image_0_263 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_264 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h108 == _T_37[9:0]) begin
        image_0_264 <= io_pixelVal_in_0_7;
      end else if (10'h108 == _T_34[9:0]) begin
        image_0_264 <= io_pixelVal_in_0_6;
      end else if (10'h108 == _T_31[9:0]) begin
        image_0_264 <= io_pixelVal_in_0_5;
      end else if (10'h108 == _T_28[9:0]) begin
        image_0_264 <= io_pixelVal_in_0_4;
      end else if (10'h108 == _T_25[9:0]) begin
        image_0_264 <= io_pixelVal_in_0_3;
      end else if (10'h108 == _T_22[9:0]) begin
        image_0_264 <= io_pixelVal_in_0_2;
      end else if (10'h108 == _T_19[9:0]) begin
        image_0_264 <= io_pixelVal_in_0_1;
      end else if (10'h108 == _T_15[9:0]) begin
        image_0_264 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_265 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h109 == _T_37[9:0]) begin
        image_0_265 <= io_pixelVal_in_0_7;
      end else if (10'h109 == _T_34[9:0]) begin
        image_0_265 <= io_pixelVal_in_0_6;
      end else if (10'h109 == _T_31[9:0]) begin
        image_0_265 <= io_pixelVal_in_0_5;
      end else if (10'h109 == _T_28[9:0]) begin
        image_0_265 <= io_pixelVal_in_0_4;
      end else if (10'h109 == _T_25[9:0]) begin
        image_0_265 <= io_pixelVal_in_0_3;
      end else if (10'h109 == _T_22[9:0]) begin
        image_0_265 <= io_pixelVal_in_0_2;
      end else if (10'h109 == _T_19[9:0]) begin
        image_0_265 <= io_pixelVal_in_0_1;
      end else if (10'h109 == _T_15[9:0]) begin
        image_0_265 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_266 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h10a == _T_37[9:0]) begin
        image_0_266 <= io_pixelVal_in_0_7;
      end else if (10'h10a == _T_34[9:0]) begin
        image_0_266 <= io_pixelVal_in_0_6;
      end else if (10'h10a == _T_31[9:0]) begin
        image_0_266 <= io_pixelVal_in_0_5;
      end else if (10'h10a == _T_28[9:0]) begin
        image_0_266 <= io_pixelVal_in_0_4;
      end else if (10'h10a == _T_25[9:0]) begin
        image_0_266 <= io_pixelVal_in_0_3;
      end else if (10'h10a == _T_22[9:0]) begin
        image_0_266 <= io_pixelVal_in_0_2;
      end else if (10'h10a == _T_19[9:0]) begin
        image_0_266 <= io_pixelVal_in_0_1;
      end else if (10'h10a == _T_15[9:0]) begin
        image_0_266 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_267 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h10b == _T_37[9:0]) begin
        image_0_267 <= io_pixelVal_in_0_7;
      end else if (10'h10b == _T_34[9:0]) begin
        image_0_267 <= io_pixelVal_in_0_6;
      end else if (10'h10b == _T_31[9:0]) begin
        image_0_267 <= io_pixelVal_in_0_5;
      end else if (10'h10b == _T_28[9:0]) begin
        image_0_267 <= io_pixelVal_in_0_4;
      end else if (10'h10b == _T_25[9:0]) begin
        image_0_267 <= io_pixelVal_in_0_3;
      end else if (10'h10b == _T_22[9:0]) begin
        image_0_267 <= io_pixelVal_in_0_2;
      end else if (10'h10b == _T_19[9:0]) begin
        image_0_267 <= io_pixelVal_in_0_1;
      end else if (10'h10b == _T_15[9:0]) begin
        image_0_267 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_268 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h10c == _T_37[9:0]) begin
        image_0_268 <= io_pixelVal_in_0_7;
      end else if (10'h10c == _T_34[9:0]) begin
        image_0_268 <= io_pixelVal_in_0_6;
      end else if (10'h10c == _T_31[9:0]) begin
        image_0_268 <= io_pixelVal_in_0_5;
      end else if (10'h10c == _T_28[9:0]) begin
        image_0_268 <= io_pixelVal_in_0_4;
      end else if (10'h10c == _T_25[9:0]) begin
        image_0_268 <= io_pixelVal_in_0_3;
      end else if (10'h10c == _T_22[9:0]) begin
        image_0_268 <= io_pixelVal_in_0_2;
      end else if (10'h10c == _T_19[9:0]) begin
        image_0_268 <= io_pixelVal_in_0_1;
      end else if (10'h10c == _T_15[9:0]) begin
        image_0_268 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_269 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h10d == _T_37[9:0]) begin
        image_0_269 <= io_pixelVal_in_0_7;
      end else if (10'h10d == _T_34[9:0]) begin
        image_0_269 <= io_pixelVal_in_0_6;
      end else if (10'h10d == _T_31[9:0]) begin
        image_0_269 <= io_pixelVal_in_0_5;
      end else if (10'h10d == _T_28[9:0]) begin
        image_0_269 <= io_pixelVal_in_0_4;
      end else if (10'h10d == _T_25[9:0]) begin
        image_0_269 <= io_pixelVal_in_0_3;
      end else if (10'h10d == _T_22[9:0]) begin
        image_0_269 <= io_pixelVal_in_0_2;
      end else if (10'h10d == _T_19[9:0]) begin
        image_0_269 <= io_pixelVal_in_0_1;
      end else if (10'h10d == _T_15[9:0]) begin
        image_0_269 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_270 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h10e == _T_37[9:0]) begin
        image_0_270 <= io_pixelVal_in_0_7;
      end else if (10'h10e == _T_34[9:0]) begin
        image_0_270 <= io_pixelVal_in_0_6;
      end else if (10'h10e == _T_31[9:0]) begin
        image_0_270 <= io_pixelVal_in_0_5;
      end else if (10'h10e == _T_28[9:0]) begin
        image_0_270 <= io_pixelVal_in_0_4;
      end else if (10'h10e == _T_25[9:0]) begin
        image_0_270 <= io_pixelVal_in_0_3;
      end else if (10'h10e == _T_22[9:0]) begin
        image_0_270 <= io_pixelVal_in_0_2;
      end else if (10'h10e == _T_19[9:0]) begin
        image_0_270 <= io_pixelVal_in_0_1;
      end else if (10'h10e == _T_15[9:0]) begin
        image_0_270 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_271 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h10f == _T_37[9:0]) begin
        image_0_271 <= io_pixelVal_in_0_7;
      end else if (10'h10f == _T_34[9:0]) begin
        image_0_271 <= io_pixelVal_in_0_6;
      end else if (10'h10f == _T_31[9:0]) begin
        image_0_271 <= io_pixelVal_in_0_5;
      end else if (10'h10f == _T_28[9:0]) begin
        image_0_271 <= io_pixelVal_in_0_4;
      end else if (10'h10f == _T_25[9:0]) begin
        image_0_271 <= io_pixelVal_in_0_3;
      end else if (10'h10f == _T_22[9:0]) begin
        image_0_271 <= io_pixelVal_in_0_2;
      end else if (10'h10f == _T_19[9:0]) begin
        image_0_271 <= io_pixelVal_in_0_1;
      end else if (10'h10f == _T_15[9:0]) begin
        image_0_271 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_272 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h110 == _T_37[9:0]) begin
        image_0_272 <= io_pixelVal_in_0_7;
      end else if (10'h110 == _T_34[9:0]) begin
        image_0_272 <= io_pixelVal_in_0_6;
      end else if (10'h110 == _T_31[9:0]) begin
        image_0_272 <= io_pixelVal_in_0_5;
      end else if (10'h110 == _T_28[9:0]) begin
        image_0_272 <= io_pixelVal_in_0_4;
      end else if (10'h110 == _T_25[9:0]) begin
        image_0_272 <= io_pixelVal_in_0_3;
      end else if (10'h110 == _T_22[9:0]) begin
        image_0_272 <= io_pixelVal_in_0_2;
      end else if (10'h110 == _T_19[9:0]) begin
        image_0_272 <= io_pixelVal_in_0_1;
      end else if (10'h110 == _T_15[9:0]) begin
        image_0_272 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_273 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h111 == _T_37[9:0]) begin
        image_0_273 <= io_pixelVal_in_0_7;
      end else if (10'h111 == _T_34[9:0]) begin
        image_0_273 <= io_pixelVal_in_0_6;
      end else if (10'h111 == _T_31[9:0]) begin
        image_0_273 <= io_pixelVal_in_0_5;
      end else if (10'h111 == _T_28[9:0]) begin
        image_0_273 <= io_pixelVal_in_0_4;
      end else if (10'h111 == _T_25[9:0]) begin
        image_0_273 <= io_pixelVal_in_0_3;
      end else if (10'h111 == _T_22[9:0]) begin
        image_0_273 <= io_pixelVal_in_0_2;
      end else if (10'h111 == _T_19[9:0]) begin
        image_0_273 <= io_pixelVal_in_0_1;
      end else if (10'h111 == _T_15[9:0]) begin
        image_0_273 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_274 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h112 == _T_37[9:0]) begin
        image_0_274 <= io_pixelVal_in_0_7;
      end else if (10'h112 == _T_34[9:0]) begin
        image_0_274 <= io_pixelVal_in_0_6;
      end else if (10'h112 == _T_31[9:0]) begin
        image_0_274 <= io_pixelVal_in_0_5;
      end else if (10'h112 == _T_28[9:0]) begin
        image_0_274 <= io_pixelVal_in_0_4;
      end else if (10'h112 == _T_25[9:0]) begin
        image_0_274 <= io_pixelVal_in_0_3;
      end else if (10'h112 == _T_22[9:0]) begin
        image_0_274 <= io_pixelVal_in_0_2;
      end else if (10'h112 == _T_19[9:0]) begin
        image_0_274 <= io_pixelVal_in_0_1;
      end else if (10'h112 == _T_15[9:0]) begin
        image_0_274 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_275 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h113 == _T_37[9:0]) begin
        image_0_275 <= io_pixelVal_in_0_7;
      end else if (10'h113 == _T_34[9:0]) begin
        image_0_275 <= io_pixelVal_in_0_6;
      end else if (10'h113 == _T_31[9:0]) begin
        image_0_275 <= io_pixelVal_in_0_5;
      end else if (10'h113 == _T_28[9:0]) begin
        image_0_275 <= io_pixelVal_in_0_4;
      end else if (10'h113 == _T_25[9:0]) begin
        image_0_275 <= io_pixelVal_in_0_3;
      end else if (10'h113 == _T_22[9:0]) begin
        image_0_275 <= io_pixelVal_in_0_2;
      end else if (10'h113 == _T_19[9:0]) begin
        image_0_275 <= io_pixelVal_in_0_1;
      end else if (10'h113 == _T_15[9:0]) begin
        image_0_275 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_276 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h114 == _T_37[9:0]) begin
        image_0_276 <= io_pixelVal_in_0_7;
      end else if (10'h114 == _T_34[9:0]) begin
        image_0_276 <= io_pixelVal_in_0_6;
      end else if (10'h114 == _T_31[9:0]) begin
        image_0_276 <= io_pixelVal_in_0_5;
      end else if (10'h114 == _T_28[9:0]) begin
        image_0_276 <= io_pixelVal_in_0_4;
      end else if (10'h114 == _T_25[9:0]) begin
        image_0_276 <= io_pixelVal_in_0_3;
      end else if (10'h114 == _T_22[9:0]) begin
        image_0_276 <= io_pixelVal_in_0_2;
      end else if (10'h114 == _T_19[9:0]) begin
        image_0_276 <= io_pixelVal_in_0_1;
      end else if (10'h114 == _T_15[9:0]) begin
        image_0_276 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_277 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h115 == _T_37[9:0]) begin
        image_0_277 <= io_pixelVal_in_0_7;
      end else if (10'h115 == _T_34[9:0]) begin
        image_0_277 <= io_pixelVal_in_0_6;
      end else if (10'h115 == _T_31[9:0]) begin
        image_0_277 <= io_pixelVal_in_0_5;
      end else if (10'h115 == _T_28[9:0]) begin
        image_0_277 <= io_pixelVal_in_0_4;
      end else if (10'h115 == _T_25[9:0]) begin
        image_0_277 <= io_pixelVal_in_0_3;
      end else if (10'h115 == _T_22[9:0]) begin
        image_0_277 <= io_pixelVal_in_0_2;
      end else if (10'h115 == _T_19[9:0]) begin
        image_0_277 <= io_pixelVal_in_0_1;
      end else if (10'h115 == _T_15[9:0]) begin
        image_0_277 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_278 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h116 == _T_37[9:0]) begin
        image_0_278 <= io_pixelVal_in_0_7;
      end else if (10'h116 == _T_34[9:0]) begin
        image_0_278 <= io_pixelVal_in_0_6;
      end else if (10'h116 == _T_31[9:0]) begin
        image_0_278 <= io_pixelVal_in_0_5;
      end else if (10'h116 == _T_28[9:0]) begin
        image_0_278 <= io_pixelVal_in_0_4;
      end else if (10'h116 == _T_25[9:0]) begin
        image_0_278 <= io_pixelVal_in_0_3;
      end else if (10'h116 == _T_22[9:0]) begin
        image_0_278 <= io_pixelVal_in_0_2;
      end else if (10'h116 == _T_19[9:0]) begin
        image_0_278 <= io_pixelVal_in_0_1;
      end else if (10'h116 == _T_15[9:0]) begin
        image_0_278 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_279 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h117 == _T_37[9:0]) begin
        image_0_279 <= io_pixelVal_in_0_7;
      end else if (10'h117 == _T_34[9:0]) begin
        image_0_279 <= io_pixelVal_in_0_6;
      end else if (10'h117 == _T_31[9:0]) begin
        image_0_279 <= io_pixelVal_in_0_5;
      end else if (10'h117 == _T_28[9:0]) begin
        image_0_279 <= io_pixelVal_in_0_4;
      end else if (10'h117 == _T_25[9:0]) begin
        image_0_279 <= io_pixelVal_in_0_3;
      end else if (10'h117 == _T_22[9:0]) begin
        image_0_279 <= io_pixelVal_in_0_2;
      end else if (10'h117 == _T_19[9:0]) begin
        image_0_279 <= io_pixelVal_in_0_1;
      end else if (10'h117 == _T_15[9:0]) begin
        image_0_279 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_280 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h118 == _T_37[9:0]) begin
        image_0_280 <= io_pixelVal_in_0_7;
      end else if (10'h118 == _T_34[9:0]) begin
        image_0_280 <= io_pixelVal_in_0_6;
      end else if (10'h118 == _T_31[9:0]) begin
        image_0_280 <= io_pixelVal_in_0_5;
      end else if (10'h118 == _T_28[9:0]) begin
        image_0_280 <= io_pixelVal_in_0_4;
      end else if (10'h118 == _T_25[9:0]) begin
        image_0_280 <= io_pixelVal_in_0_3;
      end else if (10'h118 == _T_22[9:0]) begin
        image_0_280 <= io_pixelVal_in_0_2;
      end else if (10'h118 == _T_19[9:0]) begin
        image_0_280 <= io_pixelVal_in_0_1;
      end else if (10'h118 == _T_15[9:0]) begin
        image_0_280 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_281 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h119 == _T_37[9:0]) begin
        image_0_281 <= io_pixelVal_in_0_7;
      end else if (10'h119 == _T_34[9:0]) begin
        image_0_281 <= io_pixelVal_in_0_6;
      end else if (10'h119 == _T_31[9:0]) begin
        image_0_281 <= io_pixelVal_in_0_5;
      end else if (10'h119 == _T_28[9:0]) begin
        image_0_281 <= io_pixelVal_in_0_4;
      end else if (10'h119 == _T_25[9:0]) begin
        image_0_281 <= io_pixelVal_in_0_3;
      end else if (10'h119 == _T_22[9:0]) begin
        image_0_281 <= io_pixelVal_in_0_2;
      end else if (10'h119 == _T_19[9:0]) begin
        image_0_281 <= io_pixelVal_in_0_1;
      end else if (10'h119 == _T_15[9:0]) begin
        image_0_281 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_282 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h11a == _T_37[9:0]) begin
        image_0_282 <= io_pixelVal_in_0_7;
      end else if (10'h11a == _T_34[9:0]) begin
        image_0_282 <= io_pixelVal_in_0_6;
      end else if (10'h11a == _T_31[9:0]) begin
        image_0_282 <= io_pixelVal_in_0_5;
      end else if (10'h11a == _T_28[9:0]) begin
        image_0_282 <= io_pixelVal_in_0_4;
      end else if (10'h11a == _T_25[9:0]) begin
        image_0_282 <= io_pixelVal_in_0_3;
      end else if (10'h11a == _T_22[9:0]) begin
        image_0_282 <= io_pixelVal_in_0_2;
      end else if (10'h11a == _T_19[9:0]) begin
        image_0_282 <= io_pixelVal_in_0_1;
      end else if (10'h11a == _T_15[9:0]) begin
        image_0_282 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_283 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h11b == _T_37[9:0]) begin
        image_0_283 <= io_pixelVal_in_0_7;
      end else if (10'h11b == _T_34[9:0]) begin
        image_0_283 <= io_pixelVal_in_0_6;
      end else if (10'h11b == _T_31[9:0]) begin
        image_0_283 <= io_pixelVal_in_0_5;
      end else if (10'h11b == _T_28[9:0]) begin
        image_0_283 <= io_pixelVal_in_0_4;
      end else if (10'h11b == _T_25[9:0]) begin
        image_0_283 <= io_pixelVal_in_0_3;
      end else if (10'h11b == _T_22[9:0]) begin
        image_0_283 <= io_pixelVal_in_0_2;
      end else if (10'h11b == _T_19[9:0]) begin
        image_0_283 <= io_pixelVal_in_0_1;
      end else if (10'h11b == _T_15[9:0]) begin
        image_0_283 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_284 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h11c == _T_37[9:0]) begin
        image_0_284 <= io_pixelVal_in_0_7;
      end else if (10'h11c == _T_34[9:0]) begin
        image_0_284 <= io_pixelVal_in_0_6;
      end else if (10'h11c == _T_31[9:0]) begin
        image_0_284 <= io_pixelVal_in_0_5;
      end else if (10'h11c == _T_28[9:0]) begin
        image_0_284 <= io_pixelVal_in_0_4;
      end else if (10'h11c == _T_25[9:0]) begin
        image_0_284 <= io_pixelVal_in_0_3;
      end else if (10'h11c == _T_22[9:0]) begin
        image_0_284 <= io_pixelVal_in_0_2;
      end else if (10'h11c == _T_19[9:0]) begin
        image_0_284 <= io_pixelVal_in_0_1;
      end else if (10'h11c == _T_15[9:0]) begin
        image_0_284 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_285 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h11d == _T_37[9:0]) begin
        image_0_285 <= io_pixelVal_in_0_7;
      end else if (10'h11d == _T_34[9:0]) begin
        image_0_285 <= io_pixelVal_in_0_6;
      end else if (10'h11d == _T_31[9:0]) begin
        image_0_285 <= io_pixelVal_in_0_5;
      end else if (10'h11d == _T_28[9:0]) begin
        image_0_285 <= io_pixelVal_in_0_4;
      end else if (10'h11d == _T_25[9:0]) begin
        image_0_285 <= io_pixelVal_in_0_3;
      end else if (10'h11d == _T_22[9:0]) begin
        image_0_285 <= io_pixelVal_in_0_2;
      end else if (10'h11d == _T_19[9:0]) begin
        image_0_285 <= io_pixelVal_in_0_1;
      end else if (10'h11d == _T_15[9:0]) begin
        image_0_285 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_286 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h11e == _T_37[9:0]) begin
        image_0_286 <= io_pixelVal_in_0_7;
      end else if (10'h11e == _T_34[9:0]) begin
        image_0_286 <= io_pixelVal_in_0_6;
      end else if (10'h11e == _T_31[9:0]) begin
        image_0_286 <= io_pixelVal_in_0_5;
      end else if (10'h11e == _T_28[9:0]) begin
        image_0_286 <= io_pixelVal_in_0_4;
      end else if (10'h11e == _T_25[9:0]) begin
        image_0_286 <= io_pixelVal_in_0_3;
      end else if (10'h11e == _T_22[9:0]) begin
        image_0_286 <= io_pixelVal_in_0_2;
      end else if (10'h11e == _T_19[9:0]) begin
        image_0_286 <= io_pixelVal_in_0_1;
      end else if (10'h11e == _T_15[9:0]) begin
        image_0_286 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_287 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h11f == _T_37[9:0]) begin
        image_0_287 <= io_pixelVal_in_0_7;
      end else if (10'h11f == _T_34[9:0]) begin
        image_0_287 <= io_pixelVal_in_0_6;
      end else if (10'h11f == _T_31[9:0]) begin
        image_0_287 <= io_pixelVal_in_0_5;
      end else if (10'h11f == _T_28[9:0]) begin
        image_0_287 <= io_pixelVal_in_0_4;
      end else if (10'h11f == _T_25[9:0]) begin
        image_0_287 <= io_pixelVal_in_0_3;
      end else if (10'h11f == _T_22[9:0]) begin
        image_0_287 <= io_pixelVal_in_0_2;
      end else if (10'h11f == _T_19[9:0]) begin
        image_0_287 <= io_pixelVal_in_0_1;
      end else if (10'h11f == _T_15[9:0]) begin
        image_0_287 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_288 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h120 == _T_37[9:0]) begin
        image_0_288 <= io_pixelVal_in_0_7;
      end else if (10'h120 == _T_34[9:0]) begin
        image_0_288 <= io_pixelVal_in_0_6;
      end else if (10'h120 == _T_31[9:0]) begin
        image_0_288 <= io_pixelVal_in_0_5;
      end else if (10'h120 == _T_28[9:0]) begin
        image_0_288 <= io_pixelVal_in_0_4;
      end else if (10'h120 == _T_25[9:0]) begin
        image_0_288 <= io_pixelVal_in_0_3;
      end else if (10'h120 == _T_22[9:0]) begin
        image_0_288 <= io_pixelVal_in_0_2;
      end else if (10'h120 == _T_19[9:0]) begin
        image_0_288 <= io_pixelVal_in_0_1;
      end else if (10'h120 == _T_15[9:0]) begin
        image_0_288 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_289 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h121 == _T_37[9:0]) begin
        image_0_289 <= io_pixelVal_in_0_7;
      end else if (10'h121 == _T_34[9:0]) begin
        image_0_289 <= io_pixelVal_in_0_6;
      end else if (10'h121 == _T_31[9:0]) begin
        image_0_289 <= io_pixelVal_in_0_5;
      end else if (10'h121 == _T_28[9:0]) begin
        image_0_289 <= io_pixelVal_in_0_4;
      end else if (10'h121 == _T_25[9:0]) begin
        image_0_289 <= io_pixelVal_in_0_3;
      end else if (10'h121 == _T_22[9:0]) begin
        image_0_289 <= io_pixelVal_in_0_2;
      end else if (10'h121 == _T_19[9:0]) begin
        image_0_289 <= io_pixelVal_in_0_1;
      end else if (10'h121 == _T_15[9:0]) begin
        image_0_289 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_290 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h122 == _T_37[9:0]) begin
        image_0_290 <= io_pixelVal_in_0_7;
      end else if (10'h122 == _T_34[9:0]) begin
        image_0_290 <= io_pixelVal_in_0_6;
      end else if (10'h122 == _T_31[9:0]) begin
        image_0_290 <= io_pixelVal_in_0_5;
      end else if (10'h122 == _T_28[9:0]) begin
        image_0_290 <= io_pixelVal_in_0_4;
      end else if (10'h122 == _T_25[9:0]) begin
        image_0_290 <= io_pixelVal_in_0_3;
      end else if (10'h122 == _T_22[9:0]) begin
        image_0_290 <= io_pixelVal_in_0_2;
      end else if (10'h122 == _T_19[9:0]) begin
        image_0_290 <= io_pixelVal_in_0_1;
      end else if (10'h122 == _T_15[9:0]) begin
        image_0_290 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_291 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h123 == _T_37[9:0]) begin
        image_0_291 <= io_pixelVal_in_0_7;
      end else if (10'h123 == _T_34[9:0]) begin
        image_0_291 <= io_pixelVal_in_0_6;
      end else if (10'h123 == _T_31[9:0]) begin
        image_0_291 <= io_pixelVal_in_0_5;
      end else if (10'h123 == _T_28[9:0]) begin
        image_0_291 <= io_pixelVal_in_0_4;
      end else if (10'h123 == _T_25[9:0]) begin
        image_0_291 <= io_pixelVal_in_0_3;
      end else if (10'h123 == _T_22[9:0]) begin
        image_0_291 <= io_pixelVal_in_0_2;
      end else if (10'h123 == _T_19[9:0]) begin
        image_0_291 <= io_pixelVal_in_0_1;
      end else if (10'h123 == _T_15[9:0]) begin
        image_0_291 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_292 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h124 == _T_37[9:0]) begin
        image_0_292 <= io_pixelVal_in_0_7;
      end else if (10'h124 == _T_34[9:0]) begin
        image_0_292 <= io_pixelVal_in_0_6;
      end else if (10'h124 == _T_31[9:0]) begin
        image_0_292 <= io_pixelVal_in_0_5;
      end else if (10'h124 == _T_28[9:0]) begin
        image_0_292 <= io_pixelVal_in_0_4;
      end else if (10'h124 == _T_25[9:0]) begin
        image_0_292 <= io_pixelVal_in_0_3;
      end else if (10'h124 == _T_22[9:0]) begin
        image_0_292 <= io_pixelVal_in_0_2;
      end else if (10'h124 == _T_19[9:0]) begin
        image_0_292 <= io_pixelVal_in_0_1;
      end else if (10'h124 == _T_15[9:0]) begin
        image_0_292 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_293 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h125 == _T_37[9:0]) begin
        image_0_293 <= io_pixelVal_in_0_7;
      end else if (10'h125 == _T_34[9:0]) begin
        image_0_293 <= io_pixelVal_in_0_6;
      end else if (10'h125 == _T_31[9:0]) begin
        image_0_293 <= io_pixelVal_in_0_5;
      end else if (10'h125 == _T_28[9:0]) begin
        image_0_293 <= io_pixelVal_in_0_4;
      end else if (10'h125 == _T_25[9:0]) begin
        image_0_293 <= io_pixelVal_in_0_3;
      end else if (10'h125 == _T_22[9:0]) begin
        image_0_293 <= io_pixelVal_in_0_2;
      end else if (10'h125 == _T_19[9:0]) begin
        image_0_293 <= io_pixelVal_in_0_1;
      end else if (10'h125 == _T_15[9:0]) begin
        image_0_293 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_294 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h126 == _T_37[9:0]) begin
        image_0_294 <= io_pixelVal_in_0_7;
      end else if (10'h126 == _T_34[9:0]) begin
        image_0_294 <= io_pixelVal_in_0_6;
      end else if (10'h126 == _T_31[9:0]) begin
        image_0_294 <= io_pixelVal_in_0_5;
      end else if (10'h126 == _T_28[9:0]) begin
        image_0_294 <= io_pixelVal_in_0_4;
      end else if (10'h126 == _T_25[9:0]) begin
        image_0_294 <= io_pixelVal_in_0_3;
      end else if (10'h126 == _T_22[9:0]) begin
        image_0_294 <= io_pixelVal_in_0_2;
      end else if (10'h126 == _T_19[9:0]) begin
        image_0_294 <= io_pixelVal_in_0_1;
      end else if (10'h126 == _T_15[9:0]) begin
        image_0_294 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_295 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h127 == _T_37[9:0]) begin
        image_0_295 <= io_pixelVal_in_0_7;
      end else if (10'h127 == _T_34[9:0]) begin
        image_0_295 <= io_pixelVal_in_0_6;
      end else if (10'h127 == _T_31[9:0]) begin
        image_0_295 <= io_pixelVal_in_0_5;
      end else if (10'h127 == _T_28[9:0]) begin
        image_0_295 <= io_pixelVal_in_0_4;
      end else if (10'h127 == _T_25[9:0]) begin
        image_0_295 <= io_pixelVal_in_0_3;
      end else if (10'h127 == _T_22[9:0]) begin
        image_0_295 <= io_pixelVal_in_0_2;
      end else if (10'h127 == _T_19[9:0]) begin
        image_0_295 <= io_pixelVal_in_0_1;
      end else if (10'h127 == _T_15[9:0]) begin
        image_0_295 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_296 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h128 == _T_37[9:0]) begin
        image_0_296 <= io_pixelVal_in_0_7;
      end else if (10'h128 == _T_34[9:0]) begin
        image_0_296 <= io_pixelVal_in_0_6;
      end else if (10'h128 == _T_31[9:0]) begin
        image_0_296 <= io_pixelVal_in_0_5;
      end else if (10'h128 == _T_28[9:0]) begin
        image_0_296 <= io_pixelVal_in_0_4;
      end else if (10'h128 == _T_25[9:0]) begin
        image_0_296 <= io_pixelVal_in_0_3;
      end else if (10'h128 == _T_22[9:0]) begin
        image_0_296 <= io_pixelVal_in_0_2;
      end else if (10'h128 == _T_19[9:0]) begin
        image_0_296 <= io_pixelVal_in_0_1;
      end else if (10'h128 == _T_15[9:0]) begin
        image_0_296 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_297 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h129 == _T_37[9:0]) begin
        image_0_297 <= io_pixelVal_in_0_7;
      end else if (10'h129 == _T_34[9:0]) begin
        image_0_297 <= io_pixelVal_in_0_6;
      end else if (10'h129 == _T_31[9:0]) begin
        image_0_297 <= io_pixelVal_in_0_5;
      end else if (10'h129 == _T_28[9:0]) begin
        image_0_297 <= io_pixelVal_in_0_4;
      end else if (10'h129 == _T_25[9:0]) begin
        image_0_297 <= io_pixelVal_in_0_3;
      end else if (10'h129 == _T_22[9:0]) begin
        image_0_297 <= io_pixelVal_in_0_2;
      end else if (10'h129 == _T_19[9:0]) begin
        image_0_297 <= io_pixelVal_in_0_1;
      end else if (10'h129 == _T_15[9:0]) begin
        image_0_297 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_298 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h12a == _T_37[9:0]) begin
        image_0_298 <= io_pixelVal_in_0_7;
      end else if (10'h12a == _T_34[9:0]) begin
        image_0_298 <= io_pixelVal_in_0_6;
      end else if (10'h12a == _T_31[9:0]) begin
        image_0_298 <= io_pixelVal_in_0_5;
      end else if (10'h12a == _T_28[9:0]) begin
        image_0_298 <= io_pixelVal_in_0_4;
      end else if (10'h12a == _T_25[9:0]) begin
        image_0_298 <= io_pixelVal_in_0_3;
      end else if (10'h12a == _T_22[9:0]) begin
        image_0_298 <= io_pixelVal_in_0_2;
      end else if (10'h12a == _T_19[9:0]) begin
        image_0_298 <= io_pixelVal_in_0_1;
      end else if (10'h12a == _T_15[9:0]) begin
        image_0_298 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_299 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h12b == _T_37[9:0]) begin
        image_0_299 <= io_pixelVal_in_0_7;
      end else if (10'h12b == _T_34[9:0]) begin
        image_0_299 <= io_pixelVal_in_0_6;
      end else if (10'h12b == _T_31[9:0]) begin
        image_0_299 <= io_pixelVal_in_0_5;
      end else if (10'h12b == _T_28[9:0]) begin
        image_0_299 <= io_pixelVal_in_0_4;
      end else if (10'h12b == _T_25[9:0]) begin
        image_0_299 <= io_pixelVal_in_0_3;
      end else if (10'h12b == _T_22[9:0]) begin
        image_0_299 <= io_pixelVal_in_0_2;
      end else if (10'h12b == _T_19[9:0]) begin
        image_0_299 <= io_pixelVal_in_0_1;
      end else if (10'h12b == _T_15[9:0]) begin
        image_0_299 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_300 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h12c == _T_37[9:0]) begin
        image_0_300 <= io_pixelVal_in_0_7;
      end else if (10'h12c == _T_34[9:0]) begin
        image_0_300 <= io_pixelVal_in_0_6;
      end else if (10'h12c == _T_31[9:0]) begin
        image_0_300 <= io_pixelVal_in_0_5;
      end else if (10'h12c == _T_28[9:0]) begin
        image_0_300 <= io_pixelVal_in_0_4;
      end else if (10'h12c == _T_25[9:0]) begin
        image_0_300 <= io_pixelVal_in_0_3;
      end else if (10'h12c == _T_22[9:0]) begin
        image_0_300 <= io_pixelVal_in_0_2;
      end else if (10'h12c == _T_19[9:0]) begin
        image_0_300 <= io_pixelVal_in_0_1;
      end else if (10'h12c == _T_15[9:0]) begin
        image_0_300 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_301 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h12d == _T_37[9:0]) begin
        image_0_301 <= io_pixelVal_in_0_7;
      end else if (10'h12d == _T_34[9:0]) begin
        image_0_301 <= io_pixelVal_in_0_6;
      end else if (10'h12d == _T_31[9:0]) begin
        image_0_301 <= io_pixelVal_in_0_5;
      end else if (10'h12d == _T_28[9:0]) begin
        image_0_301 <= io_pixelVal_in_0_4;
      end else if (10'h12d == _T_25[9:0]) begin
        image_0_301 <= io_pixelVal_in_0_3;
      end else if (10'h12d == _T_22[9:0]) begin
        image_0_301 <= io_pixelVal_in_0_2;
      end else if (10'h12d == _T_19[9:0]) begin
        image_0_301 <= io_pixelVal_in_0_1;
      end else if (10'h12d == _T_15[9:0]) begin
        image_0_301 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_302 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h12e == _T_37[9:0]) begin
        image_0_302 <= io_pixelVal_in_0_7;
      end else if (10'h12e == _T_34[9:0]) begin
        image_0_302 <= io_pixelVal_in_0_6;
      end else if (10'h12e == _T_31[9:0]) begin
        image_0_302 <= io_pixelVal_in_0_5;
      end else if (10'h12e == _T_28[9:0]) begin
        image_0_302 <= io_pixelVal_in_0_4;
      end else if (10'h12e == _T_25[9:0]) begin
        image_0_302 <= io_pixelVal_in_0_3;
      end else if (10'h12e == _T_22[9:0]) begin
        image_0_302 <= io_pixelVal_in_0_2;
      end else if (10'h12e == _T_19[9:0]) begin
        image_0_302 <= io_pixelVal_in_0_1;
      end else if (10'h12e == _T_15[9:0]) begin
        image_0_302 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_303 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h12f == _T_37[9:0]) begin
        image_0_303 <= io_pixelVal_in_0_7;
      end else if (10'h12f == _T_34[9:0]) begin
        image_0_303 <= io_pixelVal_in_0_6;
      end else if (10'h12f == _T_31[9:0]) begin
        image_0_303 <= io_pixelVal_in_0_5;
      end else if (10'h12f == _T_28[9:0]) begin
        image_0_303 <= io_pixelVal_in_0_4;
      end else if (10'h12f == _T_25[9:0]) begin
        image_0_303 <= io_pixelVal_in_0_3;
      end else if (10'h12f == _T_22[9:0]) begin
        image_0_303 <= io_pixelVal_in_0_2;
      end else if (10'h12f == _T_19[9:0]) begin
        image_0_303 <= io_pixelVal_in_0_1;
      end else if (10'h12f == _T_15[9:0]) begin
        image_0_303 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_304 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h130 == _T_37[9:0]) begin
        image_0_304 <= io_pixelVal_in_0_7;
      end else if (10'h130 == _T_34[9:0]) begin
        image_0_304 <= io_pixelVal_in_0_6;
      end else if (10'h130 == _T_31[9:0]) begin
        image_0_304 <= io_pixelVal_in_0_5;
      end else if (10'h130 == _T_28[9:0]) begin
        image_0_304 <= io_pixelVal_in_0_4;
      end else if (10'h130 == _T_25[9:0]) begin
        image_0_304 <= io_pixelVal_in_0_3;
      end else if (10'h130 == _T_22[9:0]) begin
        image_0_304 <= io_pixelVal_in_0_2;
      end else if (10'h130 == _T_19[9:0]) begin
        image_0_304 <= io_pixelVal_in_0_1;
      end else if (10'h130 == _T_15[9:0]) begin
        image_0_304 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_305 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h131 == _T_37[9:0]) begin
        image_0_305 <= io_pixelVal_in_0_7;
      end else if (10'h131 == _T_34[9:0]) begin
        image_0_305 <= io_pixelVal_in_0_6;
      end else if (10'h131 == _T_31[9:0]) begin
        image_0_305 <= io_pixelVal_in_0_5;
      end else if (10'h131 == _T_28[9:0]) begin
        image_0_305 <= io_pixelVal_in_0_4;
      end else if (10'h131 == _T_25[9:0]) begin
        image_0_305 <= io_pixelVal_in_0_3;
      end else if (10'h131 == _T_22[9:0]) begin
        image_0_305 <= io_pixelVal_in_0_2;
      end else if (10'h131 == _T_19[9:0]) begin
        image_0_305 <= io_pixelVal_in_0_1;
      end else if (10'h131 == _T_15[9:0]) begin
        image_0_305 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_306 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h132 == _T_37[9:0]) begin
        image_0_306 <= io_pixelVal_in_0_7;
      end else if (10'h132 == _T_34[9:0]) begin
        image_0_306 <= io_pixelVal_in_0_6;
      end else if (10'h132 == _T_31[9:0]) begin
        image_0_306 <= io_pixelVal_in_0_5;
      end else if (10'h132 == _T_28[9:0]) begin
        image_0_306 <= io_pixelVal_in_0_4;
      end else if (10'h132 == _T_25[9:0]) begin
        image_0_306 <= io_pixelVal_in_0_3;
      end else if (10'h132 == _T_22[9:0]) begin
        image_0_306 <= io_pixelVal_in_0_2;
      end else if (10'h132 == _T_19[9:0]) begin
        image_0_306 <= io_pixelVal_in_0_1;
      end else if (10'h132 == _T_15[9:0]) begin
        image_0_306 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_307 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h133 == _T_37[9:0]) begin
        image_0_307 <= io_pixelVal_in_0_7;
      end else if (10'h133 == _T_34[9:0]) begin
        image_0_307 <= io_pixelVal_in_0_6;
      end else if (10'h133 == _T_31[9:0]) begin
        image_0_307 <= io_pixelVal_in_0_5;
      end else if (10'h133 == _T_28[9:0]) begin
        image_0_307 <= io_pixelVal_in_0_4;
      end else if (10'h133 == _T_25[9:0]) begin
        image_0_307 <= io_pixelVal_in_0_3;
      end else if (10'h133 == _T_22[9:0]) begin
        image_0_307 <= io_pixelVal_in_0_2;
      end else if (10'h133 == _T_19[9:0]) begin
        image_0_307 <= io_pixelVal_in_0_1;
      end else if (10'h133 == _T_15[9:0]) begin
        image_0_307 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_308 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h134 == _T_37[9:0]) begin
        image_0_308 <= io_pixelVal_in_0_7;
      end else if (10'h134 == _T_34[9:0]) begin
        image_0_308 <= io_pixelVal_in_0_6;
      end else if (10'h134 == _T_31[9:0]) begin
        image_0_308 <= io_pixelVal_in_0_5;
      end else if (10'h134 == _T_28[9:0]) begin
        image_0_308 <= io_pixelVal_in_0_4;
      end else if (10'h134 == _T_25[9:0]) begin
        image_0_308 <= io_pixelVal_in_0_3;
      end else if (10'h134 == _T_22[9:0]) begin
        image_0_308 <= io_pixelVal_in_0_2;
      end else if (10'h134 == _T_19[9:0]) begin
        image_0_308 <= io_pixelVal_in_0_1;
      end else if (10'h134 == _T_15[9:0]) begin
        image_0_308 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_309 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h135 == _T_37[9:0]) begin
        image_0_309 <= io_pixelVal_in_0_7;
      end else if (10'h135 == _T_34[9:0]) begin
        image_0_309 <= io_pixelVal_in_0_6;
      end else if (10'h135 == _T_31[9:0]) begin
        image_0_309 <= io_pixelVal_in_0_5;
      end else if (10'h135 == _T_28[9:0]) begin
        image_0_309 <= io_pixelVal_in_0_4;
      end else if (10'h135 == _T_25[9:0]) begin
        image_0_309 <= io_pixelVal_in_0_3;
      end else if (10'h135 == _T_22[9:0]) begin
        image_0_309 <= io_pixelVal_in_0_2;
      end else if (10'h135 == _T_19[9:0]) begin
        image_0_309 <= io_pixelVal_in_0_1;
      end else if (10'h135 == _T_15[9:0]) begin
        image_0_309 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_310 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h136 == _T_37[9:0]) begin
        image_0_310 <= io_pixelVal_in_0_7;
      end else if (10'h136 == _T_34[9:0]) begin
        image_0_310 <= io_pixelVal_in_0_6;
      end else if (10'h136 == _T_31[9:0]) begin
        image_0_310 <= io_pixelVal_in_0_5;
      end else if (10'h136 == _T_28[9:0]) begin
        image_0_310 <= io_pixelVal_in_0_4;
      end else if (10'h136 == _T_25[9:0]) begin
        image_0_310 <= io_pixelVal_in_0_3;
      end else if (10'h136 == _T_22[9:0]) begin
        image_0_310 <= io_pixelVal_in_0_2;
      end else if (10'h136 == _T_19[9:0]) begin
        image_0_310 <= io_pixelVal_in_0_1;
      end else if (10'h136 == _T_15[9:0]) begin
        image_0_310 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_311 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h137 == _T_37[9:0]) begin
        image_0_311 <= io_pixelVal_in_0_7;
      end else if (10'h137 == _T_34[9:0]) begin
        image_0_311 <= io_pixelVal_in_0_6;
      end else if (10'h137 == _T_31[9:0]) begin
        image_0_311 <= io_pixelVal_in_0_5;
      end else if (10'h137 == _T_28[9:0]) begin
        image_0_311 <= io_pixelVal_in_0_4;
      end else if (10'h137 == _T_25[9:0]) begin
        image_0_311 <= io_pixelVal_in_0_3;
      end else if (10'h137 == _T_22[9:0]) begin
        image_0_311 <= io_pixelVal_in_0_2;
      end else if (10'h137 == _T_19[9:0]) begin
        image_0_311 <= io_pixelVal_in_0_1;
      end else if (10'h137 == _T_15[9:0]) begin
        image_0_311 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_312 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h138 == _T_37[9:0]) begin
        image_0_312 <= io_pixelVal_in_0_7;
      end else if (10'h138 == _T_34[9:0]) begin
        image_0_312 <= io_pixelVal_in_0_6;
      end else if (10'h138 == _T_31[9:0]) begin
        image_0_312 <= io_pixelVal_in_0_5;
      end else if (10'h138 == _T_28[9:0]) begin
        image_0_312 <= io_pixelVal_in_0_4;
      end else if (10'h138 == _T_25[9:0]) begin
        image_0_312 <= io_pixelVal_in_0_3;
      end else if (10'h138 == _T_22[9:0]) begin
        image_0_312 <= io_pixelVal_in_0_2;
      end else if (10'h138 == _T_19[9:0]) begin
        image_0_312 <= io_pixelVal_in_0_1;
      end else if (10'h138 == _T_15[9:0]) begin
        image_0_312 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_313 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h139 == _T_37[9:0]) begin
        image_0_313 <= io_pixelVal_in_0_7;
      end else if (10'h139 == _T_34[9:0]) begin
        image_0_313 <= io_pixelVal_in_0_6;
      end else if (10'h139 == _T_31[9:0]) begin
        image_0_313 <= io_pixelVal_in_0_5;
      end else if (10'h139 == _T_28[9:0]) begin
        image_0_313 <= io_pixelVal_in_0_4;
      end else if (10'h139 == _T_25[9:0]) begin
        image_0_313 <= io_pixelVal_in_0_3;
      end else if (10'h139 == _T_22[9:0]) begin
        image_0_313 <= io_pixelVal_in_0_2;
      end else if (10'h139 == _T_19[9:0]) begin
        image_0_313 <= io_pixelVal_in_0_1;
      end else if (10'h139 == _T_15[9:0]) begin
        image_0_313 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_314 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h13a == _T_37[9:0]) begin
        image_0_314 <= io_pixelVal_in_0_7;
      end else if (10'h13a == _T_34[9:0]) begin
        image_0_314 <= io_pixelVal_in_0_6;
      end else if (10'h13a == _T_31[9:0]) begin
        image_0_314 <= io_pixelVal_in_0_5;
      end else if (10'h13a == _T_28[9:0]) begin
        image_0_314 <= io_pixelVal_in_0_4;
      end else if (10'h13a == _T_25[9:0]) begin
        image_0_314 <= io_pixelVal_in_0_3;
      end else if (10'h13a == _T_22[9:0]) begin
        image_0_314 <= io_pixelVal_in_0_2;
      end else if (10'h13a == _T_19[9:0]) begin
        image_0_314 <= io_pixelVal_in_0_1;
      end else if (10'h13a == _T_15[9:0]) begin
        image_0_314 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_315 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h13b == _T_37[9:0]) begin
        image_0_315 <= io_pixelVal_in_0_7;
      end else if (10'h13b == _T_34[9:0]) begin
        image_0_315 <= io_pixelVal_in_0_6;
      end else if (10'h13b == _T_31[9:0]) begin
        image_0_315 <= io_pixelVal_in_0_5;
      end else if (10'h13b == _T_28[9:0]) begin
        image_0_315 <= io_pixelVal_in_0_4;
      end else if (10'h13b == _T_25[9:0]) begin
        image_0_315 <= io_pixelVal_in_0_3;
      end else if (10'h13b == _T_22[9:0]) begin
        image_0_315 <= io_pixelVal_in_0_2;
      end else if (10'h13b == _T_19[9:0]) begin
        image_0_315 <= io_pixelVal_in_0_1;
      end else if (10'h13b == _T_15[9:0]) begin
        image_0_315 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_316 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h13c == _T_37[9:0]) begin
        image_0_316 <= io_pixelVal_in_0_7;
      end else if (10'h13c == _T_34[9:0]) begin
        image_0_316 <= io_pixelVal_in_0_6;
      end else if (10'h13c == _T_31[9:0]) begin
        image_0_316 <= io_pixelVal_in_0_5;
      end else if (10'h13c == _T_28[9:0]) begin
        image_0_316 <= io_pixelVal_in_0_4;
      end else if (10'h13c == _T_25[9:0]) begin
        image_0_316 <= io_pixelVal_in_0_3;
      end else if (10'h13c == _T_22[9:0]) begin
        image_0_316 <= io_pixelVal_in_0_2;
      end else if (10'h13c == _T_19[9:0]) begin
        image_0_316 <= io_pixelVal_in_0_1;
      end else if (10'h13c == _T_15[9:0]) begin
        image_0_316 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_317 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h13d == _T_37[9:0]) begin
        image_0_317 <= io_pixelVal_in_0_7;
      end else if (10'h13d == _T_34[9:0]) begin
        image_0_317 <= io_pixelVal_in_0_6;
      end else if (10'h13d == _T_31[9:0]) begin
        image_0_317 <= io_pixelVal_in_0_5;
      end else if (10'h13d == _T_28[9:0]) begin
        image_0_317 <= io_pixelVal_in_0_4;
      end else if (10'h13d == _T_25[9:0]) begin
        image_0_317 <= io_pixelVal_in_0_3;
      end else if (10'h13d == _T_22[9:0]) begin
        image_0_317 <= io_pixelVal_in_0_2;
      end else if (10'h13d == _T_19[9:0]) begin
        image_0_317 <= io_pixelVal_in_0_1;
      end else if (10'h13d == _T_15[9:0]) begin
        image_0_317 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_318 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h13e == _T_37[9:0]) begin
        image_0_318 <= io_pixelVal_in_0_7;
      end else if (10'h13e == _T_34[9:0]) begin
        image_0_318 <= io_pixelVal_in_0_6;
      end else if (10'h13e == _T_31[9:0]) begin
        image_0_318 <= io_pixelVal_in_0_5;
      end else if (10'h13e == _T_28[9:0]) begin
        image_0_318 <= io_pixelVal_in_0_4;
      end else if (10'h13e == _T_25[9:0]) begin
        image_0_318 <= io_pixelVal_in_0_3;
      end else if (10'h13e == _T_22[9:0]) begin
        image_0_318 <= io_pixelVal_in_0_2;
      end else if (10'h13e == _T_19[9:0]) begin
        image_0_318 <= io_pixelVal_in_0_1;
      end else if (10'h13e == _T_15[9:0]) begin
        image_0_318 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_319 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h13f == _T_37[9:0]) begin
        image_0_319 <= io_pixelVal_in_0_7;
      end else if (10'h13f == _T_34[9:0]) begin
        image_0_319 <= io_pixelVal_in_0_6;
      end else if (10'h13f == _T_31[9:0]) begin
        image_0_319 <= io_pixelVal_in_0_5;
      end else if (10'h13f == _T_28[9:0]) begin
        image_0_319 <= io_pixelVal_in_0_4;
      end else if (10'h13f == _T_25[9:0]) begin
        image_0_319 <= io_pixelVal_in_0_3;
      end else if (10'h13f == _T_22[9:0]) begin
        image_0_319 <= io_pixelVal_in_0_2;
      end else if (10'h13f == _T_19[9:0]) begin
        image_0_319 <= io_pixelVal_in_0_1;
      end else if (10'h13f == _T_15[9:0]) begin
        image_0_319 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_320 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h140 == _T_37[9:0]) begin
        image_0_320 <= io_pixelVal_in_0_7;
      end else if (10'h140 == _T_34[9:0]) begin
        image_0_320 <= io_pixelVal_in_0_6;
      end else if (10'h140 == _T_31[9:0]) begin
        image_0_320 <= io_pixelVal_in_0_5;
      end else if (10'h140 == _T_28[9:0]) begin
        image_0_320 <= io_pixelVal_in_0_4;
      end else if (10'h140 == _T_25[9:0]) begin
        image_0_320 <= io_pixelVal_in_0_3;
      end else if (10'h140 == _T_22[9:0]) begin
        image_0_320 <= io_pixelVal_in_0_2;
      end else if (10'h140 == _T_19[9:0]) begin
        image_0_320 <= io_pixelVal_in_0_1;
      end else if (10'h140 == _T_15[9:0]) begin
        image_0_320 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_321 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h141 == _T_37[9:0]) begin
        image_0_321 <= io_pixelVal_in_0_7;
      end else if (10'h141 == _T_34[9:0]) begin
        image_0_321 <= io_pixelVal_in_0_6;
      end else if (10'h141 == _T_31[9:0]) begin
        image_0_321 <= io_pixelVal_in_0_5;
      end else if (10'h141 == _T_28[9:0]) begin
        image_0_321 <= io_pixelVal_in_0_4;
      end else if (10'h141 == _T_25[9:0]) begin
        image_0_321 <= io_pixelVal_in_0_3;
      end else if (10'h141 == _T_22[9:0]) begin
        image_0_321 <= io_pixelVal_in_0_2;
      end else if (10'h141 == _T_19[9:0]) begin
        image_0_321 <= io_pixelVal_in_0_1;
      end else if (10'h141 == _T_15[9:0]) begin
        image_0_321 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_322 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h142 == _T_37[9:0]) begin
        image_0_322 <= io_pixelVal_in_0_7;
      end else if (10'h142 == _T_34[9:0]) begin
        image_0_322 <= io_pixelVal_in_0_6;
      end else if (10'h142 == _T_31[9:0]) begin
        image_0_322 <= io_pixelVal_in_0_5;
      end else if (10'h142 == _T_28[9:0]) begin
        image_0_322 <= io_pixelVal_in_0_4;
      end else if (10'h142 == _T_25[9:0]) begin
        image_0_322 <= io_pixelVal_in_0_3;
      end else if (10'h142 == _T_22[9:0]) begin
        image_0_322 <= io_pixelVal_in_0_2;
      end else if (10'h142 == _T_19[9:0]) begin
        image_0_322 <= io_pixelVal_in_0_1;
      end else if (10'h142 == _T_15[9:0]) begin
        image_0_322 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_323 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h143 == _T_37[9:0]) begin
        image_0_323 <= io_pixelVal_in_0_7;
      end else if (10'h143 == _T_34[9:0]) begin
        image_0_323 <= io_pixelVal_in_0_6;
      end else if (10'h143 == _T_31[9:0]) begin
        image_0_323 <= io_pixelVal_in_0_5;
      end else if (10'h143 == _T_28[9:0]) begin
        image_0_323 <= io_pixelVal_in_0_4;
      end else if (10'h143 == _T_25[9:0]) begin
        image_0_323 <= io_pixelVal_in_0_3;
      end else if (10'h143 == _T_22[9:0]) begin
        image_0_323 <= io_pixelVal_in_0_2;
      end else if (10'h143 == _T_19[9:0]) begin
        image_0_323 <= io_pixelVal_in_0_1;
      end else if (10'h143 == _T_15[9:0]) begin
        image_0_323 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_324 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h144 == _T_37[9:0]) begin
        image_0_324 <= io_pixelVal_in_0_7;
      end else if (10'h144 == _T_34[9:0]) begin
        image_0_324 <= io_pixelVal_in_0_6;
      end else if (10'h144 == _T_31[9:0]) begin
        image_0_324 <= io_pixelVal_in_0_5;
      end else if (10'h144 == _T_28[9:0]) begin
        image_0_324 <= io_pixelVal_in_0_4;
      end else if (10'h144 == _T_25[9:0]) begin
        image_0_324 <= io_pixelVal_in_0_3;
      end else if (10'h144 == _T_22[9:0]) begin
        image_0_324 <= io_pixelVal_in_0_2;
      end else if (10'h144 == _T_19[9:0]) begin
        image_0_324 <= io_pixelVal_in_0_1;
      end else if (10'h144 == _T_15[9:0]) begin
        image_0_324 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_325 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h145 == _T_37[9:0]) begin
        image_0_325 <= io_pixelVal_in_0_7;
      end else if (10'h145 == _T_34[9:0]) begin
        image_0_325 <= io_pixelVal_in_0_6;
      end else if (10'h145 == _T_31[9:0]) begin
        image_0_325 <= io_pixelVal_in_0_5;
      end else if (10'h145 == _T_28[9:0]) begin
        image_0_325 <= io_pixelVal_in_0_4;
      end else if (10'h145 == _T_25[9:0]) begin
        image_0_325 <= io_pixelVal_in_0_3;
      end else if (10'h145 == _T_22[9:0]) begin
        image_0_325 <= io_pixelVal_in_0_2;
      end else if (10'h145 == _T_19[9:0]) begin
        image_0_325 <= io_pixelVal_in_0_1;
      end else if (10'h145 == _T_15[9:0]) begin
        image_0_325 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_326 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h146 == _T_37[9:0]) begin
        image_0_326 <= io_pixelVal_in_0_7;
      end else if (10'h146 == _T_34[9:0]) begin
        image_0_326 <= io_pixelVal_in_0_6;
      end else if (10'h146 == _T_31[9:0]) begin
        image_0_326 <= io_pixelVal_in_0_5;
      end else if (10'h146 == _T_28[9:0]) begin
        image_0_326 <= io_pixelVal_in_0_4;
      end else if (10'h146 == _T_25[9:0]) begin
        image_0_326 <= io_pixelVal_in_0_3;
      end else if (10'h146 == _T_22[9:0]) begin
        image_0_326 <= io_pixelVal_in_0_2;
      end else if (10'h146 == _T_19[9:0]) begin
        image_0_326 <= io_pixelVal_in_0_1;
      end else if (10'h146 == _T_15[9:0]) begin
        image_0_326 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_327 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h147 == _T_37[9:0]) begin
        image_0_327 <= io_pixelVal_in_0_7;
      end else if (10'h147 == _T_34[9:0]) begin
        image_0_327 <= io_pixelVal_in_0_6;
      end else if (10'h147 == _T_31[9:0]) begin
        image_0_327 <= io_pixelVal_in_0_5;
      end else if (10'h147 == _T_28[9:0]) begin
        image_0_327 <= io_pixelVal_in_0_4;
      end else if (10'h147 == _T_25[9:0]) begin
        image_0_327 <= io_pixelVal_in_0_3;
      end else if (10'h147 == _T_22[9:0]) begin
        image_0_327 <= io_pixelVal_in_0_2;
      end else if (10'h147 == _T_19[9:0]) begin
        image_0_327 <= io_pixelVal_in_0_1;
      end else if (10'h147 == _T_15[9:0]) begin
        image_0_327 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_328 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h148 == _T_37[9:0]) begin
        image_0_328 <= io_pixelVal_in_0_7;
      end else if (10'h148 == _T_34[9:0]) begin
        image_0_328 <= io_pixelVal_in_0_6;
      end else if (10'h148 == _T_31[9:0]) begin
        image_0_328 <= io_pixelVal_in_0_5;
      end else if (10'h148 == _T_28[9:0]) begin
        image_0_328 <= io_pixelVal_in_0_4;
      end else if (10'h148 == _T_25[9:0]) begin
        image_0_328 <= io_pixelVal_in_0_3;
      end else if (10'h148 == _T_22[9:0]) begin
        image_0_328 <= io_pixelVal_in_0_2;
      end else if (10'h148 == _T_19[9:0]) begin
        image_0_328 <= io_pixelVal_in_0_1;
      end else if (10'h148 == _T_15[9:0]) begin
        image_0_328 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_329 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h149 == _T_37[9:0]) begin
        image_0_329 <= io_pixelVal_in_0_7;
      end else if (10'h149 == _T_34[9:0]) begin
        image_0_329 <= io_pixelVal_in_0_6;
      end else if (10'h149 == _T_31[9:0]) begin
        image_0_329 <= io_pixelVal_in_0_5;
      end else if (10'h149 == _T_28[9:0]) begin
        image_0_329 <= io_pixelVal_in_0_4;
      end else if (10'h149 == _T_25[9:0]) begin
        image_0_329 <= io_pixelVal_in_0_3;
      end else if (10'h149 == _T_22[9:0]) begin
        image_0_329 <= io_pixelVal_in_0_2;
      end else if (10'h149 == _T_19[9:0]) begin
        image_0_329 <= io_pixelVal_in_0_1;
      end else if (10'h149 == _T_15[9:0]) begin
        image_0_329 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_330 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h14a == _T_37[9:0]) begin
        image_0_330 <= io_pixelVal_in_0_7;
      end else if (10'h14a == _T_34[9:0]) begin
        image_0_330 <= io_pixelVal_in_0_6;
      end else if (10'h14a == _T_31[9:0]) begin
        image_0_330 <= io_pixelVal_in_0_5;
      end else if (10'h14a == _T_28[9:0]) begin
        image_0_330 <= io_pixelVal_in_0_4;
      end else if (10'h14a == _T_25[9:0]) begin
        image_0_330 <= io_pixelVal_in_0_3;
      end else if (10'h14a == _T_22[9:0]) begin
        image_0_330 <= io_pixelVal_in_0_2;
      end else if (10'h14a == _T_19[9:0]) begin
        image_0_330 <= io_pixelVal_in_0_1;
      end else if (10'h14a == _T_15[9:0]) begin
        image_0_330 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_331 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h14b == _T_37[9:0]) begin
        image_0_331 <= io_pixelVal_in_0_7;
      end else if (10'h14b == _T_34[9:0]) begin
        image_0_331 <= io_pixelVal_in_0_6;
      end else if (10'h14b == _T_31[9:0]) begin
        image_0_331 <= io_pixelVal_in_0_5;
      end else if (10'h14b == _T_28[9:0]) begin
        image_0_331 <= io_pixelVal_in_0_4;
      end else if (10'h14b == _T_25[9:0]) begin
        image_0_331 <= io_pixelVal_in_0_3;
      end else if (10'h14b == _T_22[9:0]) begin
        image_0_331 <= io_pixelVal_in_0_2;
      end else if (10'h14b == _T_19[9:0]) begin
        image_0_331 <= io_pixelVal_in_0_1;
      end else if (10'h14b == _T_15[9:0]) begin
        image_0_331 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_332 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h14c == _T_37[9:0]) begin
        image_0_332 <= io_pixelVal_in_0_7;
      end else if (10'h14c == _T_34[9:0]) begin
        image_0_332 <= io_pixelVal_in_0_6;
      end else if (10'h14c == _T_31[9:0]) begin
        image_0_332 <= io_pixelVal_in_0_5;
      end else if (10'h14c == _T_28[9:0]) begin
        image_0_332 <= io_pixelVal_in_0_4;
      end else if (10'h14c == _T_25[9:0]) begin
        image_0_332 <= io_pixelVal_in_0_3;
      end else if (10'h14c == _T_22[9:0]) begin
        image_0_332 <= io_pixelVal_in_0_2;
      end else if (10'h14c == _T_19[9:0]) begin
        image_0_332 <= io_pixelVal_in_0_1;
      end else if (10'h14c == _T_15[9:0]) begin
        image_0_332 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_333 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h14d == _T_37[9:0]) begin
        image_0_333 <= io_pixelVal_in_0_7;
      end else if (10'h14d == _T_34[9:0]) begin
        image_0_333 <= io_pixelVal_in_0_6;
      end else if (10'h14d == _T_31[9:0]) begin
        image_0_333 <= io_pixelVal_in_0_5;
      end else if (10'h14d == _T_28[9:0]) begin
        image_0_333 <= io_pixelVal_in_0_4;
      end else if (10'h14d == _T_25[9:0]) begin
        image_0_333 <= io_pixelVal_in_0_3;
      end else if (10'h14d == _T_22[9:0]) begin
        image_0_333 <= io_pixelVal_in_0_2;
      end else if (10'h14d == _T_19[9:0]) begin
        image_0_333 <= io_pixelVal_in_0_1;
      end else if (10'h14d == _T_15[9:0]) begin
        image_0_333 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_334 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h14e == _T_37[9:0]) begin
        image_0_334 <= io_pixelVal_in_0_7;
      end else if (10'h14e == _T_34[9:0]) begin
        image_0_334 <= io_pixelVal_in_0_6;
      end else if (10'h14e == _T_31[9:0]) begin
        image_0_334 <= io_pixelVal_in_0_5;
      end else if (10'h14e == _T_28[9:0]) begin
        image_0_334 <= io_pixelVal_in_0_4;
      end else if (10'h14e == _T_25[9:0]) begin
        image_0_334 <= io_pixelVal_in_0_3;
      end else if (10'h14e == _T_22[9:0]) begin
        image_0_334 <= io_pixelVal_in_0_2;
      end else if (10'h14e == _T_19[9:0]) begin
        image_0_334 <= io_pixelVal_in_0_1;
      end else if (10'h14e == _T_15[9:0]) begin
        image_0_334 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_335 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h14f == _T_37[9:0]) begin
        image_0_335 <= io_pixelVal_in_0_7;
      end else if (10'h14f == _T_34[9:0]) begin
        image_0_335 <= io_pixelVal_in_0_6;
      end else if (10'h14f == _T_31[9:0]) begin
        image_0_335 <= io_pixelVal_in_0_5;
      end else if (10'h14f == _T_28[9:0]) begin
        image_0_335 <= io_pixelVal_in_0_4;
      end else if (10'h14f == _T_25[9:0]) begin
        image_0_335 <= io_pixelVal_in_0_3;
      end else if (10'h14f == _T_22[9:0]) begin
        image_0_335 <= io_pixelVal_in_0_2;
      end else if (10'h14f == _T_19[9:0]) begin
        image_0_335 <= io_pixelVal_in_0_1;
      end else if (10'h14f == _T_15[9:0]) begin
        image_0_335 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_336 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h150 == _T_37[9:0]) begin
        image_0_336 <= io_pixelVal_in_0_7;
      end else if (10'h150 == _T_34[9:0]) begin
        image_0_336 <= io_pixelVal_in_0_6;
      end else if (10'h150 == _T_31[9:0]) begin
        image_0_336 <= io_pixelVal_in_0_5;
      end else if (10'h150 == _T_28[9:0]) begin
        image_0_336 <= io_pixelVal_in_0_4;
      end else if (10'h150 == _T_25[9:0]) begin
        image_0_336 <= io_pixelVal_in_0_3;
      end else if (10'h150 == _T_22[9:0]) begin
        image_0_336 <= io_pixelVal_in_0_2;
      end else if (10'h150 == _T_19[9:0]) begin
        image_0_336 <= io_pixelVal_in_0_1;
      end else if (10'h150 == _T_15[9:0]) begin
        image_0_336 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_337 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h151 == _T_37[9:0]) begin
        image_0_337 <= io_pixelVal_in_0_7;
      end else if (10'h151 == _T_34[9:0]) begin
        image_0_337 <= io_pixelVal_in_0_6;
      end else if (10'h151 == _T_31[9:0]) begin
        image_0_337 <= io_pixelVal_in_0_5;
      end else if (10'h151 == _T_28[9:0]) begin
        image_0_337 <= io_pixelVal_in_0_4;
      end else if (10'h151 == _T_25[9:0]) begin
        image_0_337 <= io_pixelVal_in_0_3;
      end else if (10'h151 == _T_22[9:0]) begin
        image_0_337 <= io_pixelVal_in_0_2;
      end else if (10'h151 == _T_19[9:0]) begin
        image_0_337 <= io_pixelVal_in_0_1;
      end else if (10'h151 == _T_15[9:0]) begin
        image_0_337 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_338 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h152 == _T_37[9:0]) begin
        image_0_338 <= io_pixelVal_in_0_7;
      end else if (10'h152 == _T_34[9:0]) begin
        image_0_338 <= io_pixelVal_in_0_6;
      end else if (10'h152 == _T_31[9:0]) begin
        image_0_338 <= io_pixelVal_in_0_5;
      end else if (10'h152 == _T_28[9:0]) begin
        image_0_338 <= io_pixelVal_in_0_4;
      end else if (10'h152 == _T_25[9:0]) begin
        image_0_338 <= io_pixelVal_in_0_3;
      end else if (10'h152 == _T_22[9:0]) begin
        image_0_338 <= io_pixelVal_in_0_2;
      end else if (10'h152 == _T_19[9:0]) begin
        image_0_338 <= io_pixelVal_in_0_1;
      end else if (10'h152 == _T_15[9:0]) begin
        image_0_338 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_339 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h153 == _T_37[9:0]) begin
        image_0_339 <= io_pixelVal_in_0_7;
      end else if (10'h153 == _T_34[9:0]) begin
        image_0_339 <= io_pixelVal_in_0_6;
      end else if (10'h153 == _T_31[9:0]) begin
        image_0_339 <= io_pixelVal_in_0_5;
      end else if (10'h153 == _T_28[9:0]) begin
        image_0_339 <= io_pixelVal_in_0_4;
      end else if (10'h153 == _T_25[9:0]) begin
        image_0_339 <= io_pixelVal_in_0_3;
      end else if (10'h153 == _T_22[9:0]) begin
        image_0_339 <= io_pixelVal_in_0_2;
      end else if (10'h153 == _T_19[9:0]) begin
        image_0_339 <= io_pixelVal_in_0_1;
      end else if (10'h153 == _T_15[9:0]) begin
        image_0_339 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_340 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h154 == _T_37[9:0]) begin
        image_0_340 <= io_pixelVal_in_0_7;
      end else if (10'h154 == _T_34[9:0]) begin
        image_0_340 <= io_pixelVal_in_0_6;
      end else if (10'h154 == _T_31[9:0]) begin
        image_0_340 <= io_pixelVal_in_0_5;
      end else if (10'h154 == _T_28[9:0]) begin
        image_0_340 <= io_pixelVal_in_0_4;
      end else if (10'h154 == _T_25[9:0]) begin
        image_0_340 <= io_pixelVal_in_0_3;
      end else if (10'h154 == _T_22[9:0]) begin
        image_0_340 <= io_pixelVal_in_0_2;
      end else if (10'h154 == _T_19[9:0]) begin
        image_0_340 <= io_pixelVal_in_0_1;
      end else if (10'h154 == _T_15[9:0]) begin
        image_0_340 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_341 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h155 == _T_37[9:0]) begin
        image_0_341 <= io_pixelVal_in_0_7;
      end else if (10'h155 == _T_34[9:0]) begin
        image_0_341 <= io_pixelVal_in_0_6;
      end else if (10'h155 == _T_31[9:0]) begin
        image_0_341 <= io_pixelVal_in_0_5;
      end else if (10'h155 == _T_28[9:0]) begin
        image_0_341 <= io_pixelVal_in_0_4;
      end else if (10'h155 == _T_25[9:0]) begin
        image_0_341 <= io_pixelVal_in_0_3;
      end else if (10'h155 == _T_22[9:0]) begin
        image_0_341 <= io_pixelVal_in_0_2;
      end else if (10'h155 == _T_19[9:0]) begin
        image_0_341 <= io_pixelVal_in_0_1;
      end else if (10'h155 == _T_15[9:0]) begin
        image_0_341 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_342 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h156 == _T_37[9:0]) begin
        image_0_342 <= io_pixelVal_in_0_7;
      end else if (10'h156 == _T_34[9:0]) begin
        image_0_342 <= io_pixelVal_in_0_6;
      end else if (10'h156 == _T_31[9:0]) begin
        image_0_342 <= io_pixelVal_in_0_5;
      end else if (10'h156 == _T_28[9:0]) begin
        image_0_342 <= io_pixelVal_in_0_4;
      end else if (10'h156 == _T_25[9:0]) begin
        image_0_342 <= io_pixelVal_in_0_3;
      end else if (10'h156 == _T_22[9:0]) begin
        image_0_342 <= io_pixelVal_in_0_2;
      end else if (10'h156 == _T_19[9:0]) begin
        image_0_342 <= io_pixelVal_in_0_1;
      end else if (10'h156 == _T_15[9:0]) begin
        image_0_342 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_343 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h157 == _T_37[9:0]) begin
        image_0_343 <= io_pixelVal_in_0_7;
      end else if (10'h157 == _T_34[9:0]) begin
        image_0_343 <= io_pixelVal_in_0_6;
      end else if (10'h157 == _T_31[9:0]) begin
        image_0_343 <= io_pixelVal_in_0_5;
      end else if (10'h157 == _T_28[9:0]) begin
        image_0_343 <= io_pixelVal_in_0_4;
      end else if (10'h157 == _T_25[9:0]) begin
        image_0_343 <= io_pixelVal_in_0_3;
      end else if (10'h157 == _T_22[9:0]) begin
        image_0_343 <= io_pixelVal_in_0_2;
      end else if (10'h157 == _T_19[9:0]) begin
        image_0_343 <= io_pixelVal_in_0_1;
      end else if (10'h157 == _T_15[9:0]) begin
        image_0_343 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_344 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h158 == _T_37[9:0]) begin
        image_0_344 <= io_pixelVal_in_0_7;
      end else if (10'h158 == _T_34[9:0]) begin
        image_0_344 <= io_pixelVal_in_0_6;
      end else if (10'h158 == _T_31[9:0]) begin
        image_0_344 <= io_pixelVal_in_0_5;
      end else if (10'h158 == _T_28[9:0]) begin
        image_0_344 <= io_pixelVal_in_0_4;
      end else if (10'h158 == _T_25[9:0]) begin
        image_0_344 <= io_pixelVal_in_0_3;
      end else if (10'h158 == _T_22[9:0]) begin
        image_0_344 <= io_pixelVal_in_0_2;
      end else if (10'h158 == _T_19[9:0]) begin
        image_0_344 <= io_pixelVal_in_0_1;
      end else if (10'h158 == _T_15[9:0]) begin
        image_0_344 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_345 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h159 == _T_37[9:0]) begin
        image_0_345 <= io_pixelVal_in_0_7;
      end else if (10'h159 == _T_34[9:0]) begin
        image_0_345 <= io_pixelVal_in_0_6;
      end else if (10'h159 == _T_31[9:0]) begin
        image_0_345 <= io_pixelVal_in_0_5;
      end else if (10'h159 == _T_28[9:0]) begin
        image_0_345 <= io_pixelVal_in_0_4;
      end else if (10'h159 == _T_25[9:0]) begin
        image_0_345 <= io_pixelVal_in_0_3;
      end else if (10'h159 == _T_22[9:0]) begin
        image_0_345 <= io_pixelVal_in_0_2;
      end else if (10'h159 == _T_19[9:0]) begin
        image_0_345 <= io_pixelVal_in_0_1;
      end else if (10'h159 == _T_15[9:0]) begin
        image_0_345 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_346 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h15a == _T_37[9:0]) begin
        image_0_346 <= io_pixelVal_in_0_7;
      end else if (10'h15a == _T_34[9:0]) begin
        image_0_346 <= io_pixelVal_in_0_6;
      end else if (10'h15a == _T_31[9:0]) begin
        image_0_346 <= io_pixelVal_in_0_5;
      end else if (10'h15a == _T_28[9:0]) begin
        image_0_346 <= io_pixelVal_in_0_4;
      end else if (10'h15a == _T_25[9:0]) begin
        image_0_346 <= io_pixelVal_in_0_3;
      end else if (10'h15a == _T_22[9:0]) begin
        image_0_346 <= io_pixelVal_in_0_2;
      end else if (10'h15a == _T_19[9:0]) begin
        image_0_346 <= io_pixelVal_in_0_1;
      end else if (10'h15a == _T_15[9:0]) begin
        image_0_346 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_347 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h15b == _T_37[9:0]) begin
        image_0_347 <= io_pixelVal_in_0_7;
      end else if (10'h15b == _T_34[9:0]) begin
        image_0_347 <= io_pixelVal_in_0_6;
      end else if (10'h15b == _T_31[9:0]) begin
        image_0_347 <= io_pixelVal_in_0_5;
      end else if (10'h15b == _T_28[9:0]) begin
        image_0_347 <= io_pixelVal_in_0_4;
      end else if (10'h15b == _T_25[9:0]) begin
        image_0_347 <= io_pixelVal_in_0_3;
      end else if (10'h15b == _T_22[9:0]) begin
        image_0_347 <= io_pixelVal_in_0_2;
      end else if (10'h15b == _T_19[9:0]) begin
        image_0_347 <= io_pixelVal_in_0_1;
      end else if (10'h15b == _T_15[9:0]) begin
        image_0_347 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_348 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h15c == _T_37[9:0]) begin
        image_0_348 <= io_pixelVal_in_0_7;
      end else if (10'h15c == _T_34[9:0]) begin
        image_0_348 <= io_pixelVal_in_0_6;
      end else if (10'h15c == _T_31[9:0]) begin
        image_0_348 <= io_pixelVal_in_0_5;
      end else if (10'h15c == _T_28[9:0]) begin
        image_0_348 <= io_pixelVal_in_0_4;
      end else if (10'h15c == _T_25[9:0]) begin
        image_0_348 <= io_pixelVal_in_0_3;
      end else if (10'h15c == _T_22[9:0]) begin
        image_0_348 <= io_pixelVal_in_0_2;
      end else if (10'h15c == _T_19[9:0]) begin
        image_0_348 <= io_pixelVal_in_0_1;
      end else if (10'h15c == _T_15[9:0]) begin
        image_0_348 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_349 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h15d == _T_37[9:0]) begin
        image_0_349 <= io_pixelVal_in_0_7;
      end else if (10'h15d == _T_34[9:0]) begin
        image_0_349 <= io_pixelVal_in_0_6;
      end else if (10'h15d == _T_31[9:0]) begin
        image_0_349 <= io_pixelVal_in_0_5;
      end else if (10'h15d == _T_28[9:0]) begin
        image_0_349 <= io_pixelVal_in_0_4;
      end else if (10'h15d == _T_25[9:0]) begin
        image_0_349 <= io_pixelVal_in_0_3;
      end else if (10'h15d == _T_22[9:0]) begin
        image_0_349 <= io_pixelVal_in_0_2;
      end else if (10'h15d == _T_19[9:0]) begin
        image_0_349 <= io_pixelVal_in_0_1;
      end else if (10'h15d == _T_15[9:0]) begin
        image_0_349 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_350 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h15e == _T_37[9:0]) begin
        image_0_350 <= io_pixelVal_in_0_7;
      end else if (10'h15e == _T_34[9:0]) begin
        image_0_350 <= io_pixelVal_in_0_6;
      end else if (10'h15e == _T_31[9:0]) begin
        image_0_350 <= io_pixelVal_in_0_5;
      end else if (10'h15e == _T_28[9:0]) begin
        image_0_350 <= io_pixelVal_in_0_4;
      end else if (10'h15e == _T_25[9:0]) begin
        image_0_350 <= io_pixelVal_in_0_3;
      end else if (10'h15e == _T_22[9:0]) begin
        image_0_350 <= io_pixelVal_in_0_2;
      end else if (10'h15e == _T_19[9:0]) begin
        image_0_350 <= io_pixelVal_in_0_1;
      end else if (10'h15e == _T_15[9:0]) begin
        image_0_350 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_351 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h15f == _T_37[9:0]) begin
        image_0_351 <= io_pixelVal_in_0_7;
      end else if (10'h15f == _T_34[9:0]) begin
        image_0_351 <= io_pixelVal_in_0_6;
      end else if (10'h15f == _T_31[9:0]) begin
        image_0_351 <= io_pixelVal_in_0_5;
      end else if (10'h15f == _T_28[9:0]) begin
        image_0_351 <= io_pixelVal_in_0_4;
      end else if (10'h15f == _T_25[9:0]) begin
        image_0_351 <= io_pixelVal_in_0_3;
      end else if (10'h15f == _T_22[9:0]) begin
        image_0_351 <= io_pixelVal_in_0_2;
      end else if (10'h15f == _T_19[9:0]) begin
        image_0_351 <= io_pixelVal_in_0_1;
      end else if (10'h15f == _T_15[9:0]) begin
        image_0_351 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_352 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h160 == _T_37[9:0]) begin
        image_0_352 <= io_pixelVal_in_0_7;
      end else if (10'h160 == _T_34[9:0]) begin
        image_0_352 <= io_pixelVal_in_0_6;
      end else if (10'h160 == _T_31[9:0]) begin
        image_0_352 <= io_pixelVal_in_0_5;
      end else if (10'h160 == _T_28[9:0]) begin
        image_0_352 <= io_pixelVal_in_0_4;
      end else if (10'h160 == _T_25[9:0]) begin
        image_0_352 <= io_pixelVal_in_0_3;
      end else if (10'h160 == _T_22[9:0]) begin
        image_0_352 <= io_pixelVal_in_0_2;
      end else if (10'h160 == _T_19[9:0]) begin
        image_0_352 <= io_pixelVal_in_0_1;
      end else if (10'h160 == _T_15[9:0]) begin
        image_0_352 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_353 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h161 == _T_37[9:0]) begin
        image_0_353 <= io_pixelVal_in_0_7;
      end else if (10'h161 == _T_34[9:0]) begin
        image_0_353 <= io_pixelVal_in_0_6;
      end else if (10'h161 == _T_31[9:0]) begin
        image_0_353 <= io_pixelVal_in_0_5;
      end else if (10'h161 == _T_28[9:0]) begin
        image_0_353 <= io_pixelVal_in_0_4;
      end else if (10'h161 == _T_25[9:0]) begin
        image_0_353 <= io_pixelVal_in_0_3;
      end else if (10'h161 == _T_22[9:0]) begin
        image_0_353 <= io_pixelVal_in_0_2;
      end else if (10'h161 == _T_19[9:0]) begin
        image_0_353 <= io_pixelVal_in_0_1;
      end else if (10'h161 == _T_15[9:0]) begin
        image_0_353 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_354 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h162 == _T_37[9:0]) begin
        image_0_354 <= io_pixelVal_in_0_7;
      end else if (10'h162 == _T_34[9:0]) begin
        image_0_354 <= io_pixelVal_in_0_6;
      end else if (10'h162 == _T_31[9:0]) begin
        image_0_354 <= io_pixelVal_in_0_5;
      end else if (10'h162 == _T_28[9:0]) begin
        image_0_354 <= io_pixelVal_in_0_4;
      end else if (10'h162 == _T_25[9:0]) begin
        image_0_354 <= io_pixelVal_in_0_3;
      end else if (10'h162 == _T_22[9:0]) begin
        image_0_354 <= io_pixelVal_in_0_2;
      end else if (10'h162 == _T_19[9:0]) begin
        image_0_354 <= io_pixelVal_in_0_1;
      end else if (10'h162 == _T_15[9:0]) begin
        image_0_354 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_355 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h163 == _T_37[9:0]) begin
        image_0_355 <= io_pixelVal_in_0_7;
      end else if (10'h163 == _T_34[9:0]) begin
        image_0_355 <= io_pixelVal_in_0_6;
      end else if (10'h163 == _T_31[9:0]) begin
        image_0_355 <= io_pixelVal_in_0_5;
      end else if (10'h163 == _T_28[9:0]) begin
        image_0_355 <= io_pixelVal_in_0_4;
      end else if (10'h163 == _T_25[9:0]) begin
        image_0_355 <= io_pixelVal_in_0_3;
      end else if (10'h163 == _T_22[9:0]) begin
        image_0_355 <= io_pixelVal_in_0_2;
      end else if (10'h163 == _T_19[9:0]) begin
        image_0_355 <= io_pixelVal_in_0_1;
      end else if (10'h163 == _T_15[9:0]) begin
        image_0_355 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_356 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h164 == _T_37[9:0]) begin
        image_0_356 <= io_pixelVal_in_0_7;
      end else if (10'h164 == _T_34[9:0]) begin
        image_0_356 <= io_pixelVal_in_0_6;
      end else if (10'h164 == _T_31[9:0]) begin
        image_0_356 <= io_pixelVal_in_0_5;
      end else if (10'h164 == _T_28[9:0]) begin
        image_0_356 <= io_pixelVal_in_0_4;
      end else if (10'h164 == _T_25[9:0]) begin
        image_0_356 <= io_pixelVal_in_0_3;
      end else if (10'h164 == _T_22[9:0]) begin
        image_0_356 <= io_pixelVal_in_0_2;
      end else if (10'h164 == _T_19[9:0]) begin
        image_0_356 <= io_pixelVal_in_0_1;
      end else if (10'h164 == _T_15[9:0]) begin
        image_0_356 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_357 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h165 == _T_37[9:0]) begin
        image_0_357 <= io_pixelVal_in_0_7;
      end else if (10'h165 == _T_34[9:0]) begin
        image_0_357 <= io_pixelVal_in_0_6;
      end else if (10'h165 == _T_31[9:0]) begin
        image_0_357 <= io_pixelVal_in_0_5;
      end else if (10'h165 == _T_28[9:0]) begin
        image_0_357 <= io_pixelVal_in_0_4;
      end else if (10'h165 == _T_25[9:0]) begin
        image_0_357 <= io_pixelVal_in_0_3;
      end else if (10'h165 == _T_22[9:0]) begin
        image_0_357 <= io_pixelVal_in_0_2;
      end else if (10'h165 == _T_19[9:0]) begin
        image_0_357 <= io_pixelVal_in_0_1;
      end else if (10'h165 == _T_15[9:0]) begin
        image_0_357 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_358 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h166 == _T_37[9:0]) begin
        image_0_358 <= io_pixelVal_in_0_7;
      end else if (10'h166 == _T_34[9:0]) begin
        image_0_358 <= io_pixelVal_in_0_6;
      end else if (10'h166 == _T_31[9:0]) begin
        image_0_358 <= io_pixelVal_in_0_5;
      end else if (10'h166 == _T_28[9:0]) begin
        image_0_358 <= io_pixelVal_in_0_4;
      end else if (10'h166 == _T_25[9:0]) begin
        image_0_358 <= io_pixelVal_in_0_3;
      end else if (10'h166 == _T_22[9:0]) begin
        image_0_358 <= io_pixelVal_in_0_2;
      end else if (10'h166 == _T_19[9:0]) begin
        image_0_358 <= io_pixelVal_in_0_1;
      end else if (10'h166 == _T_15[9:0]) begin
        image_0_358 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_359 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h167 == _T_37[9:0]) begin
        image_0_359 <= io_pixelVal_in_0_7;
      end else if (10'h167 == _T_34[9:0]) begin
        image_0_359 <= io_pixelVal_in_0_6;
      end else if (10'h167 == _T_31[9:0]) begin
        image_0_359 <= io_pixelVal_in_0_5;
      end else if (10'h167 == _T_28[9:0]) begin
        image_0_359 <= io_pixelVal_in_0_4;
      end else if (10'h167 == _T_25[9:0]) begin
        image_0_359 <= io_pixelVal_in_0_3;
      end else if (10'h167 == _T_22[9:0]) begin
        image_0_359 <= io_pixelVal_in_0_2;
      end else if (10'h167 == _T_19[9:0]) begin
        image_0_359 <= io_pixelVal_in_0_1;
      end else if (10'h167 == _T_15[9:0]) begin
        image_0_359 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_360 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h168 == _T_37[9:0]) begin
        image_0_360 <= io_pixelVal_in_0_7;
      end else if (10'h168 == _T_34[9:0]) begin
        image_0_360 <= io_pixelVal_in_0_6;
      end else if (10'h168 == _T_31[9:0]) begin
        image_0_360 <= io_pixelVal_in_0_5;
      end else if (10'h168 == _T_28[9:0]) begin
        image_0_360 <= io_pixelVal_in_0_4;
      end else if (10'h168 == _T_25[9:0]) begin
        image_0_360 <= io_pixelVal_in_0_3;
      end else if (10'h168 == _T_22[9:0]) begin
        image_0_360 <= io_pixelVal_in_0_2;
      end else if (10'h168 == _T_19[9:0]) begin
        image_0_360 <= io_pixelVal_in_0_1;
      end else if (10'h168 == _T_15[9:0]) begin
        image_0_360 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_361 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h169 == _T_37[9:0]) begin
        image_0_361 <= io_pixelVal_in_0_7;
      end else if (10'h169 == _T_34[9:0]) begin
        image_0_361 <= io_pixelVal_in_0_6;
      end else if (10'h169 == _T_31[9:0]) begin
        image_0_361 <= io_pixelVal_in_0_5;
      end else if (10'h169 == _T_28[9:0]) begin
        image_0_361 <= io_pixelVal_in_0_4;
      end else if (10'h169 == _T_25[9:0]) begin
        image_0_361 <= io_pixelVal_in_0_3;
      end else if (10'h169 == _T_22[9:0]) begin
        image_0_361 <= io_pixelVal_in_0_2;
      end else if (10'h169 == _T_19[9:0]) begin
        image_0_361 <= io_pixelVal_in_0_1;
      end else if (10'h169 == _T_15[9:0]) begin
        image_0_361 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_362 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h16a == _T_37[9:0]) begin
        image_0_362 <= io_pixelVal_in_0_7;
      end else if (10'h16a == _T_34[9:0]) begin
        image_0_362 <= io_pixelVal_in_0_6;
      end else if (10'h16a == _T_31[9:0]) begin
        image_0_362 <= io_pixelVal_in_0_5;
      end else if (10'h16a == _T_28[9:0]) begin
        image_0_362 <= io_pixelVal_in_0_4;
      end else if (10'h16a == _T_25[9:0]) begin
        image_0_362 <= io_pixelVal_in_0_3;
      end else if (10'h16a == _T_22[9:0]) begin
        image_0_362 <= io_pixelVal_in_0_2;
      end else if (10'h16a == _T_19[9:0]) begin
        image_0_362 <= io_pixelVal_in_0_1;
      end else if (10'h16a == _T_15[9:0]) begin
        image_0_362 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_363 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h16b == _T_37[9:0]) begin
        image_0_363 <= io_pixelVal_in_0_7;
      end else if (10'h16b == _T_34[9:0]) begin
        image_0_363 <= io_pixelVal_in_0_6;
      end else if (10'h16b == _T_31[9:0]) begin
        image_0_363 <= io_pixelVal_in_0_5;
      end else if (10'h16b == _T_28[9:0]) begin
        image_0_363 <= io_pixelVal_in_0_4;
      end else if (10'h16b == _T_25[9:0]) begin
        image_0_363 <= io_pixelVal_in_0_3;
      end else if (10'h16b == _T_22[9:0]) begin
        image_0_363 <= io_pixelVal_in_0_2;
      end else if (10'h16b == _T_19[9:0]) begin
        image_0_363 <= io_pixelVal_in_0_1;
      end else if (10'h16b == _T_15[9:0]) begin
        image_0_363 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_364 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h16c == _T_37[9:0]) begin
        image_0_364 <= io_pixelVal_in_0_7;
      end else if (10'h16c == _T_34[9:0]) begin
        image_0_364 <= io_pixelVal_in_0_6;
      end else if (10'h16c == _T_31[9:0]) begin
        image_0_364 <= io_pixelVal_in_0_5;
      end else if (10'h16c == _T_28[9:0]) begin
        image_0_364 <= io_pixelVal_in_0_4;
      end else if (10'h16c == _T_25[9:0]) begin
        image_0_364 <= io_pixelVal_in_0_3;
      end else if (10'h16c == _T_22[9:0]) begin
        image_0_364 <= io_pixelVal_in_0_2;
      end else if (10'h16c == _T_19[9:0]) begin
        image_0_364 <= io_pixelVal_in_0_1;
      end else if (10'h16c == _T_15[9:0]) begin
        image_0_364 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_365 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h16d == _T_37[9:0]) begin
        image_0_365 <= io_pixelVal_in_0_7;
      end else if (10'h16d == _T_34[9:0]) begin
        image_0_365 <= io_pixelVal_in_0_6;
      end else if (10'h16d == _T_31[9:0]) begin
        image_0_365 <= io_pixelVal_in_0_5;
      end else if (10'h16d == _T_28[9:0]) begin
        image_0_365 <= io_pixelVal_in_0_4;
      end else if (10'h16d == _T_25[9:0]) begin
        image_0_365 <= io_pixelVal_in_0_3;
      end else if (10'h16d == _T_22[9:0]) begin
        image_0_365 <= io_pixelVal_in_0_2;
      end else if (10'h16d == _T_19[9:0]) begin
        image_0_365 <= io_pixelVal_in_0_1;
      end else if (10'h16d == _T_15[9:0]) begin
        image_0_365 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_366 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h16e == _T_37[9:0]) begin
        image_0_366 <= io_pixelVal_in_0_7;
      end else if (10'h16e == _T_34[9:0]) begin
        image_0_366 <= io_pixelVal_in_0_6;
      end else if (10'h16e == _T_31[9:0]) begin
        image_0_366 <= io_pixelVal_in_0_5;
      end else if (10'h16e == _T_28[9:0]) begin
        image_0_366 <= io_pixelVal_in_0_4;
      end else if (10'h16e == _T_25[9:0]) begin
        image_0_366 <= io_pixelVal_in_0_3;
      end else if (10'h16e == _T_22[9:0]) begin
        image_0_366 <= io_pixelVal_in_0_2;
      end else if (10'h16e == _T_19[9:0]) begin
        image_0_366 <= io_pixelVal_in_0_1;
      end else if (10'h16e == _T_15[9:0]) begin
        image_0_366 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_367 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h16f == _T_37[9:0]) begin
        image_0_367 <= io_pixelVal_in_0_7;
      end else if (10'h16f == _T_34[9:0]) begin
        image_0_367 <= io_pixelVal_in_0_6;
      end else if (10'h16f == _T_31[9:0]) begin
        image_0_367 <= io_pixelVal_in_0_5;
      end else if (10'h16f == _T_28[9:0]) begin
        image_0_367 <= io_pixelVal_in_0_4;
      end else if (10'h16f == _T_25[9:0]) begin
        image_0_367 <= io_pixelVal_in_0_3;
      end else if (10'h16f == _T_22[9:0]) begin
        image_0_367 <= io_pixelVal_in_0_2;
      end else if (10'h16f == _T_19[9:0]) begin
        image_0_367 <= io_pixelVal_in_0_1;
      end else if (10'h16f == _T_15[9:0]) begin
        image_0_367 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_368 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h170 == _T_37[9:0]) begin
        image_0_368 <= io_pixelVal_in_0_7;
      end else if (10'h170 == _T_34[9:0]) begin
        image_0_368 <= io_pixelVal_in_0_6;
      end else if (10'h170 == _T_31[9:0]) begin
        image_0_368 <= io_pixelVal_in_0_5;
      end else if (10'h170 == _T_28[9:0]) begin
        image_0_368 <= io_pixelVal_in_0_4;
      end else if (10'h170 == _T_25[9:0]) begin
        image_0_368 <= io_pixelVal_in_0_3;
      end else if (10'h170 == _T_22[9:0]) begin
        image_0_368 <= io_pixelVal_in_0_2;
      end else if (10'h170 == _T_19[9:0]) begin
        image_0_368 <= io_pixelVal_in_0_1;
      end else if (10'h170 == _T_15[9:0]) begin
        image_0_368 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_369 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h171 == _T_37[9:0]) begin
        image_0_369 <= io_pixelVal_in_0_7;
      end else if (10'h171 == _T_34[9:0]) begin
        image_0_369 <= io_pixelVal_in_0_6;
      end else if (10'h171 == _T_31[9:0]) begin
        image_0_369 <= io_pixelVal_in_0_5;
      end else if (10'h171 == _T_28[9:0]) begin
        image_0_369 <= io_pixelVal_in_0_4;
      end else if (10'h171 == _T_25[9:0]) begin
        image_0_369 <= io_pixelVal_in_0_3;
      end else if (10'h171 == _T_22[9:0]) begin
        image_0_369 <= io_pixelVal_in_0_2;
      end else if (10'h171 == _T_19[9:0]) begin
        image_0_369 <= io_pixelVal_in_0_1;
      end else if (10'h171 == _T_15[9:0]) begin
        image_0_369 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_370 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h172 == _T_37[9:0]) begin
        image_0_370 <= io_pixelVal_in_0_7;
      end else if (10'h172 == _T_34[9:0]) begin
        image_0_370 <= io_pixelVal_in_0_6;
      end else if (10'h172 == _T_31[9:0]) begin
        image_0_370 <= io_pixelVal_in_0_5;
      end else if (10'h172 == _T_28[9:0]) begin
        image_0_370 <= io_pixelVal_in_0_4;
      end else if (10'h172 == _T_25[9:0]) begin
        image_0_370 <= io_pixelVal_in_0_3;
      end else if (10'h172 == _T_22[9:0]) begin
        image_0_370 <= io_pixelVal_in_0_2;
      end else if (10'h172 == _T_19[9:0]) begin
        image_0_370 <= io_pixelVal_in_0_1;
      end else if (10'h172 == _T_15[9:0]) begin
        image_0_370 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_371 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h173 == _T_37[9:0]) begin
        image_0_371 <= io_pixelVal_in_0_7;
      end else if (10'h173 == _T_34[9:0]) begin
        image_0_371 <= io_pixelVal_in_0_6;
      end else if (10'h173 == _T_31[9:0]) begin
        image_0_371 <= io_pixelVal_in_0_5;
      end else if (10'h173 == _T_28[9:0]) begin
        image_0_371 <= io_pixelVal_in_0_4;
      end else if (10'h173 == _T_25[9:0]) begin
        image_0_371 <= io_pixelVal_in_0_3;
      end else if (10'h173 == _T_22[9:0]) begin
        image_0_371 <= io_pixelVal_in_0_2;
      end else if (10'h173 == _T_19[9:0]) begin
        image_0_371 <= io_pixelVal_in_0_1;
      end else if (10'h173 == _T_15[9:0]) begin
        image_0_371 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_372 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h174 == _T_37[9:0]) begin
        image_0_372 <= io_pixelVal_in_0_7;
      end else if (10'h174 == _T_34[9:0]) begin
        image_0_372 <= io_pixelVal_in_0_6;
      end else if (10'h174 == _T_31[9:0]) begin
        image_0_372 <= io_pixelVal_in_0_5;
      end else if (10'h174 == _T_28[9:0]) begin
        image_0_372 <= io_pixelVal_in_0_4;
      end else if (10'h174 == _T_25[9:0]) begin
        image_0_372 <= io_pixelVal_in_0_3;
      end else if (10'h174 == _T_22[9:0]) begin
        image_0_372 <= io_pixelVal_in_0_2;
      end else if (10'h174 == _T_19[9:0]) begin
        image_0_372 <= io_pixelVal_in_0_1;
      end else if (10'h174 == _T_15[9:0]) begin
        image_0_372 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_373 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h175 == _T_37[9:0]) begin
        image_0_373 <= io_pixelVal_in_0_7;
      end else if (10'h175 == _T_34[9:0]) begin
        image_0_373 <= io_pixelVal_in_0_6;
      end else if (10'h175 == _T_31[9:0]) begin
        image_0_373 <= io_pixelVal_in_0_5;
      end else if (10'h175 == _T_28[9:0]) begin
        image_0_373 <= io_pixelVal_in_0_4;
      end else if (10'h175 == _T_25[9:0]) begin
        image_0_373 <= io_pixelVal_in_0_3;
      end else if (10'h175 == _T_22[9:0]) begin
        image_0_373 <= io_pixelVal_in_0_2;
      end else if (10'h175 == _T_19[9:0]) begin
        image_0_373 <= io_pixelVal_in_0_1;
      end else if (10'h175 == _T_15[9:0]) begin
        image_0_373 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_374 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h176 == _T_37[9:0]) begin
        image_0_374 <= io_pixelVal_in_0_7;
      end else if (10'h176 == _T_34[9:0]) begin
        image_0_374 <= io_pixelVal_in_0_6;
      end else if (10'h176 == _T_31[9:0]) begin
        image_0_374 <= io_pixelVal_in_0_5;
      end else if (10'h176 == _T_28[9:0]) begin
        image_0_374 <= io_pixelVal_in_0_4;
      end else if (10'h176 == _T_25[9:0]) begin
        image_0_374 <= io_pixelVal_in_0_3;
      end else if (10'h176 == _T_22[9:0]) begin
        image_0_374 <= io_pixelVal_in_0_2;
      end else if (10'h176 == _T_19[9:0]) begin
        image_0_374 <= io_pixelVal_in_0_1;
      end else if (10'h176 == _T_15[9:0]) begin
        image_0_374 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_375 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h177 == _T_37[9:0]) begin
        image_0_375 <= io_pixelVal_in_0_7;
      end else if (10'h177 == _T_34[9:0]) begin
        image_0_375 <= io_pixelVal_in_0_6;
      end else if (10'h177 == _T_31[9:0]) begin
        image_0_375 <= io_pixelVal_in_0_5;
      end else if (10'h177 == _T_28[9:0]) begin
        image_0_375 <= io_pixelVal_in_0_4;
      end else if (10'h177 == _T_25[9:0]) begin
        image_0_375 <= io_pixelVal_in_0_3;
      end else if (10'h177 == _T_22[9:0]) begin
        image_0_375 <= io_pixelVal_in_0_2;
      end else if (10'h177 == _T_19[9:0]) begin
        image_0_375 <= io_pixelVal_in_0_1;
      end else if (10'h177 == _T_15[9:0]) begin
        image_0_375 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_376 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h178 == _T_37[9:0]) begin
        image_0_376 <= io_pixelVal_in_0_7;
      end else if (10'h178 == _T_34[9:0]) begin
        image_0_376 <= io_pixelVal_in_0_6;
      end else if (10'h178 == _T_31[9:0]) begin
        image_0_376 <= io_pixelVal_in_0_5;
      end else if (10'h178 == _T_28[9:0]) begin
        image_0_376 <= io_pixelVal_in_0_4;
      end else if (10'h178 == _T_25[9:0]) begin
        image_0_376 <= io_pixelVal_in_0_3;
      end else if (10'h178 == _T_22[9:0]) begin
        image_0_376 <= io_pixelVal_in_0_2;
      end else if (10'h178 == _T_19[9:0]) begin
        image_0_376 <= io_pixelVal_in_0_1;
      end else if (10'h178 == _T_15[9:0]) begin
        image_0_376 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_377 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h179 == _T_37[9:0]) begin
        image_0_377 <= io_pixelVal_in_0_7;
      end else if (10'h179 == _T_34[9:0]) begin
        image_0_377 <= io_pixelVal_in_0_6;
      end else if (10'h179 == _T_31[9:0]) begin
        image_0_377 <= io_pixelVal_in_0_5;
      end else if (10'h179 == _T_28[9:0]) begin
        image_0_377 <= io_pixelVal_in_0_4;
      end else if (10'h179 == _T_25[9:0]) begin
        image_0_377 <= io_pixelVal_in_0_3;
      end else if (10'h179 == _T_22[9:0]) begin
        image_0_377 <= io_pixelVal_in_0_2;
      end else if (10'h179 == _T_19[9:0]) begin
        image_0_377 <= io_pixelVal_in_0_1;
      end else if (10'h179 == _T_15[9:0]) begin
        image_0_377 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_378 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h17a == _T_37[9:0]) begin
        image_0_378 <= io_pixelVal_in_0_7;
      end else if (10'h17a == _T_34[9:0]) begin
        image_0_378 <= io_pixelVal_in_0_6;
      end else if (10'h17a == _T_31[9:0]) begin
        image_0_378 <= io_pixelVal_in_0_5;
      end else if (10'h17a == _T_28[9:0]) begin
        image_0_378 <= io_pixelVal_in_0_4;
      end else if (10'h17a == _T_25[9:0]) begin
        image_0_378 <= io_pixelVal_in_0_3;
      end else if (10'h17a == _T_22[9:0]) begin
        image_0_378 <= io_pixelVal_in_0_2;
      end else if (10'h17a == _T_19[9:0]) begin
        image_0_378 <= io_pixelVal_in_0_1;
      end else if (10'h17a == _T_15[9:0]) begin
        image_0_378 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_379 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h17b == _T_37[9:0]) begin
        image_0_379 <= io_pixelVal_in_0_7;
      end else if (10'h17b == _T_34[9:0]) begin
        image_0_379 <= io_pixelVal_in_0_6;
      end else if (10'h17b == _T_31[9:0]) begin
        image_0_379 <= io_pixelVal_in_0_5;
      end else if (10'h17b == _T_28[9:0]) begin
        image_0_379 <= io_pixelVal_in_0_4;
      end else if (10'h17b == _T_25[9:0]) begin
        image_0_379 <= io_pixelVal_in_0_3;
      end else if (10'h17b == _T_22[9:0]) begin
        image_0_379 <= io_pixelVal_in_0_2;
      end else if (10'h17b == _T_19[9:0]) begin
        image_0_379 <= io_pixelVal_in_0_1;
      end else if (10'h17b == _T_15[9:0]) begin
        image_0_379 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_380 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h17c == _T_37[9:0]) begin
        image_0_380 <= io_pixelVal_in_0_7;
      end else if (10'h17c == _T_34[9:0]) begin
        image_0_380 <= io_pixelVal_in_0_6;
      end else if (10'h17c == _T_31[9:0]) begin
        image_0_380 <= io_pixelVal_in_0_5;
      end else if (10'h17c == _T_28[9:0]) begin
        image_0_380 <= io_pixelVal_in_0_4;
      end else if (10'h17c == _T_25[9:0]) begin
        image_0_380 <= io_pixelVal_in_0_3;
      end else if (10'h17c == _T_22[9:0]) begin
        image_0_380 <= io_pixelVal_in_0_2;
      end else if (10'h17c == _T_19[9:0]) begin
        image_0_380 <= io_pixelVal_in_0_1;
      end else if (10'h17c == _T_15[9:0]) begin
        image_0_380 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_381 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h17d == _T_37[9:0]) begin
        image_0_381 <= io_pixelVal_in_0_7;
      end else if (10'h17d == _T_34[9:0]) begin
        image_0_381 <= io_pixelVal_in_0_6;
      end else if (10'h17d == _T_31[9:0]) begin
        image_0_381 <= io_pixelVal_in_0_5;
      end else if (10'h17d == _T_28[9:0]) begin
        image_0_381 <= io_pixelVal_in_0_4;
      end else if (10'h17d == _T_25[9:0]) begin
        image_0_381 <= io_pixelVal_in_0_3;
      end else if (10'h17d == _T_22[9:0]) begin
        image_0_381 <= io_pixelVal_in_0_2;
      end else if (10'h17d == _T_19[9:0]) begin
        image_0_381 <= io_pixelVal_in_0_1;
      end else if (10'h17d == _T_15[9:0]) begin
        image_0_381 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_382 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h17e == _T_37[9:0]) begin
        image_0_382 <= io_pixelVal_in_0_7;
      end else if (10'h17e == _T_34[9:0]) begin
        image_0_382 <= io_pixelVal_in_0_6;
      end else if (10'h17e == _T_31[9:0]) begin
        image_0_382 <= io_pixelVal_in_0_5;
      end else if (10'h17e == _T_28[9:0]) begin
        image_0_382 <= io_pixelVal_in_0_4;
      end else if (10'h17e == _T_25[9:0]) begin
        image_0_382 <= io_pixelVal_in_0_3;
      end else if (10'h17e == _T_22[9:0]) begin
        image_0_382 <= io_pixelVal_in_0_2;
      end else if (10'h17e == _T_19[9:0]) begin
        image_0_382 <= io_pixelVal_in_0_1;
      end else if (10'h17e == _T_15[9:0]) begin
        image_0_382 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_383 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h17f == _T_37[9:0]) begin
        image_0_383 <= io_pixelVal_in_0_7;
      end else if (10'h17f == _T_34[9:0]) begin
        image_0_383 <= io_pixelVal_in_0_6;
      end else if (10'h17f == _T_31[9:0]) begin
        image_0_383 <= io_pixelVal_in_0_5;
      end else if (10'h17f == _T_28[9:0]) begin
        image_0_383 <= io_pixelVal_in_0_4;
      end else if (10'h17f == _T_25[9:0]) begin
        image_0_383 <= io_pixelVal_in_0_3;
      end else if (10'h17f == _T_22[9:0]) begin
        image_0_383 <= io_pixelVal_in_0_2;
      end else if (10'h17f == _T_19[9:0]) begin
        image_0_383 <= io_pixelVal_in_0_1;
      end else if (10'h17f == _T_15[9:0]) begin
        image_0_383 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_384 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h180 == _T_37[9:0]) begin
        image_0_384 <= io_pixelVal_in_0_7;
      end else if (10'h180 == _T_34[9:0]) begin
        image_0_384 <= io_pixelVal_in_0_6;
      end else if (10'h180 == _T_31[9:0]) begin
        image_0_384 <= io_pixelVal_in_0_5;
      end else if (10'h180 == _T_28[9:0]) begin
        image_0_384 <= io_pixelVal_in_0_4;
      end else if (10'h180 == _T_25[9:0]) begin
        image_0_384 <= io_pixelVal_in_0_3;
      end else if (10'h180 == _T_22[9:0]) begin
        image_0_384 <= io_pixelVal_in_0_2;
      end else if (10'h180 == _T_19[9:0]) begin
        image_0_384 <= io_pixelVal_in_0_1;
      end else if (10'h180 == _T_15[9:0]) begin
        image_0_384 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_385 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h181 == _T_37[9:0]) begin
        image_0_385 <= io_pixelVal_in_0_7;
      end else if (10'h181 == _T_34[9:0]) begin
        image_0_385 <= io_pixelVal_in_0_6;
      end else if (10'h181 == _T_31[9:0]) begin
        image_0_385 <= io_pixelVal_in_0_5;
      end else if (10'h181 == _T_28[9:0]) begin
        image_0_385 <= io_pixelVal_in_0_4;
      end else if (10'h181 == _T_25[9:0]) begin
        image_0_385 <= io_pixelVal_in_0_3;
      end else if (10'h181 == _T_22[9:0]) begin
        image_0_385 <= io_pixelVal_in_0_2;
      end else if (10'h181 == _T_19[9:0]) begin
        image_0_385 <= io_pixelVal_in_0_1;
      end else if (10'h181 == _T_15[9:0]) begin
        image_0_385 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_386 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h182 == _T_37[9:0]) begin
        image_0_386 <= io_pixelVal_in_0_7;
      end else if (10'h182 == _T_34[9:0]) begin
        image_0_386 <= io_pixelVal_in_0_6;
      end else if (10'h182 == _T_31[9:0]) begin
        image_0_386 <= io_pixelVal_in_0_5;
      end else if (10'h182 == _T_28[9:0]) begin
        image_0_386 <= io_pixelVal_in_0_4;
      end else if (10'h182 == _T_25[9:0]) begin
        image_0_386 <= io_pixelVal_in_0_3;
      end else if (10'h182 == _T_22[9:0]) begin
        image_0_386 <= io_pixelVal_in_0_2;
      end else if (10'h182 == _T_19[9:0]) begin
        image_0_386 <= io_pixelVal_in_0_1;
      end else if (10'h182 == _T_15[9:0]) begin
        image_0_386 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_387 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h183 == _T_37[9:0]) begin
        image_0_387 <= io_pixelVal_in_0_7;
      end else if (10'h183 == _T_34[9:0]) begin
        image_0_387 <= io_pixelVal_in_0_6;
      end else if (10'h183 == _T_31[9:0]) begin
        image_0_387 <= io_pixelVal_in_0_5;
      end else if (10'h183 == _T_28[9:0]) begin
        image_0_387 <= io_pixelVal_in_0_4;
      end else if (10'h183 == _T_25[9:0]) begin
        image_0_387 <= io_pixelVal_in_0_3;
      end else if (10'h183 == _T_22[9:0]) begin
        image_0_387 <= io_pixelVal_in_0_2;
      end else if (10'h183 == _T_19[9:0]) begin
        image_0_387 <= io_pixelVal_in_0_1;
      end else if (10'h183 == _T_15[9:0]) begin
        image_0_387 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_388 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h184 == _T_37[9:0]) begin
        image_0_388 <= io_pixelVal_in_0_7;
      end else if (10'h184 == _T_34[9:0]) begin
        image_0_388 <= io_pixelVal_in_0_6;
      end else if (10'h184 == _T_31[9:0]) begin
        image_0_388 <= io_pixelVal_in_0_5;
      end else if (10'h184 == _T_28[9:0]) begin
        image_0_388 <= io_pixelVal_in_0_4;
      end else if (10'h184 == _T_25[9:0]) begin
        image_0_388 <= io_pixelVal_in_0_3;
      end else if (10'h184 == _T_22[9:0]) begin
        image_0_388 <= io_pixelVal_in_0_2;
      end else if (10'h184 == _T_19[9:0]) begin
        image_0_388 <= io_pixelVal_in_0_1;
      end else if (10'h184 == _T_15[9:0]) begin
        image_0_388 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_389 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h185 == _T_37[9:0]) begin
        image_0_389 <= io_pixelVal_in_0_7;
      end else if (10'h185 == _T_34[9:0]) begin
        image_0_389 <= io_pixelVal_in_0_6;
      end else if (10'h185 == _T_31[9:0]) begin
        image_0_389 <= io_pixelVal_in_0_5;
      end else if (10'h185 == _T_28[9:0]) begin
        image_0_389 <= io_pixelVal_in_0_4;
      end else if (10'h185 == _T_25[9:0]) begin
        image_0_389 <= io_pixelVal_in_0_3;
      end else if (10'h185 == _T_22[9:0]) begin
        image_0_389 <= io_pixelVal_in_0_2;
      end else if (10'h185 == _T_19[9:0]) begin
        image_0_389 <= io_pixelVal_in_0_1;
      end else if (10'h185 == _T_15[9:0]) begin
        image_0_389 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_390 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h186 == _T_37[9:0]) begin
        image_0_390 <= io_pixelVal_in_0_7;
      end else if (10'h186 == _T_34[9:0]) begin
        image_0_390 <= io_pixelVal_in_0_6;
      end else if (10'h186 == _T_31[9:0]) begin
        image_0_390 <= io_pixelVal_in_0_5;
      end else if (10'h186 == _T_28[9:0]) begin
        image_0_390 <= io_pixelVal_in_0_4;
      end else if (10'h186 == _T_25[9:0]) begin
        image_0_390 <= io_pixelVal_in_0_3;
      end else if (10'h186 == _T_22[9:0]) begin
        image_0_390 <= io_pixelVal_in_0_2;
      end else if (10'h186 == _T_19[9:0]) begin
        image_0_390 <= io_pixelVal_in_0_1;
      end else if (10'h186 == _T_15[9:0]) begin
        image_0_390 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_391 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h187 == _T_37[9:0]) begin
        image_0_391 <= io_pixelVal_in_0_7;
      end else if (10'h187 == _T_34[9:0]) begin
        image_0_391 <= io_pixelVal_in_0_6;
      end else if (10'h187 == _T_31[9:0]) begin
        image_0_391 <= io_pixelVal_in_0_5;
      end else if (10'h187 == _T_28[9:0]) begin
        image_0_391 <= io_pixelVal_in_0_4;
      end else if (10'h187 == _T_25[9:0]) begin
        image_0_391 <= io_pixelVal_in_0_3;
      end else if (10'h187 == _T_22[9:0]) begin
        image_0_391 <= io_pixelVal_in_0_2;
      end else if (10'h187 == _T_19[9:0]) begin
        image_0_391 <= io_pixelVal_in_0_1;
      end else if (10'h187 == _T_15[9:0]) begin
        image_0_391 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_392 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h188 == _T_37[9:0]) begin
        image_0_392 <= io_pixelVal_in_0_7;
      end else if (10'h188 == _T_34[9:0]) begin
        image_0_392 <= io_pixelVal_in_0_6;
      end else if (10'h188 == _T_31[9:0]) begin
        image_0_392 <= io_pixelVal_in_0_5;
      end else if (10'h188 == _T_28[9:0]) begin
        image_0_392 <= io_pixelVal_in_0_4;
      end else if (10'h188 == _T_25[9:0]) begin
        image_0_392 <= io_pixelVal_in_0_3;
      end else if (10'h188 == _T_22[9:0]) begin
        image_0_392 <= io_pixelVal_in_0_2;
      end else if (10'h188 == _T_19[9:0]) begin
        image_0_392 <= io_pixelVal_in_0_1;
      end else if (10'h188 == _T_15[9:0]) begin
        image_0_392 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_393 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h189 == _T_37[9:0]) begin
        image_0_393 <= io_pixelVal_in_0_7;
      end else if (10'h189 == _T_34[9:0]) begin
        image_0_393 <= io_pixelVal_in_0_6;
      end else if (10'h189 == _T_31[9:0]) begin
        image_0_393 <= io_pixelVal_in_0_5;
      end else if (10'h189 == _T_28[9:0]) begin
        image_0_393 <= io_pixelVal_in_0_4;
      end else if (10'h189 == _T_25[9:0]) begin
        image_0_393 <= io_pixelVal_in_0_3;
      end else if (10'h189 == _T_22[9:0]) begin
        image_0_393 <= io_pixelVal_in_0_2;
      end else if (10'h189 == _T_19[9:0]) begin
        image_0_393 <= io_pixelVal_in_0_1;
      end else if (10'h189 == _T_15[9:0]) begin
        image_0_393 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_394 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h18a == _T_37[9:0]) begin
        image_0_394 <= io_pixelVal_in_0_7;
      end else if (10'h18a == _T_34[9:0]) begin
        image_0_394 <= io_pixelVal_in_0_6;
      end else if (10'h18a == _T_31[9:0]) begin
        image_0_394 <= io_pixelVal_in_0_5;
      end else if (10'h18a == _T_28[9:0]) begin
        image_0_394 <= io_pixelVal_in_0_4;
      end else if (10'h18a == _T_25[9:0]) begin
        image_0_394 <= io_pixelVal_in_0_3;
      end else if (10'h18a == _T_22[9:0]) begin
        image_0_394 <= io_pixelVal_in_0_2;
      end else if (10'h18a == _T_19[9:0]) begin
        image_0_394 <= io_pixelVal_in_0_1;
      end else if (10'h18a == _T_15[9:0]) begin
        image_0_394 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_395 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h18b == _T_37[9:0]) begin
        image_0_395 <= io_pixelVal_in_0_7;
      end else if (10'h18b == _T_34[9:0]) begin
        image_0_395 <= io_pixelVal_in_0_6;
      end else if (10'h18b == _T_31[9:0]) begin
        image_0_395 <= io_pixelVal_in_0_5;
      end else if (10'h18b == _T_28[9:0]) begin
        image_0_395 <= io_pixelVal_in_0_4;
      end else if (10'h18b == _T_25[9:0]) begin
        image_0_395 <= io_pixelVal_in_0_3;
      end else if (10'h18b == _T_22[9:0]) begin
        image_0_395 <= io_pixelVal_in_0_2;
      end else if (10'h18b == _T_19[9:0]) begin
        image_0_395 <= io_pixelVal_in_0_1;
      end else if (10'h18b == _T_15[9:0]) begin
        image_0_395 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_396 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h18c == _T_37[9:0]) begin
        image_0_396 <= io_pixelVal_in_0_7;
      end else if (10'h18c == _T_34[9:0]) begin
        image_0_396 <= io_pixelVal_in_0_6;
      end else if (10'h18c == _T_31[9:0]) begin
        image_0_396 <= io_pixelVal_in_0_5;
      end else if (10'h18c == _T_28[9:0]) begin
        image_0_396 <= io_pixelVal_in_0_4;
      end else if (10'h18c == _T_25[9:0]) begin
        image_0_396 <= io_pixelVal_in_0_3;
      end else if (10'h18c == _T_22[9:0]) begin
        image_0_396 <= io_pixelVal_in_0_2;
      end else if (10'h18c == _T_19[9:0]) begin
        image_0_396 <= io_pixelVal_in_0_1;
      end else if (10'h18c == _T_15[9:0]) begin
        image_0_396 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_397 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h18d == _T_37[9:0]) begin
        image_0_397 <= io_pixelVal_in_0_7;
      end else if (10'h18d == _T_34[9:0]) begin
        image_0_397 <= io_pixelVal_in_0_6;
      end else if (10'h18d == _T_31[9:0]) begin
        image_0_397 <= io_pixelVal_in_0_5;
      end else if (10'h18d == _T_28[9:0]) begin
        image_0_397 <= io_pixelVal_in_0_4;
      end else if (10'h18d == _T_25[9:0]) begin
        image_0_397 <= io_pixelVal_in_0_3;
      end else if (10'h18d == _T_22[9:0]) begin
        image_0_397 <= io_pixelVal_in_0_2;
      end else if (10'h18d == _T_19[9:0]) begin
        image_0_397 <= io_pixelVal_in_0_1;
      end else if (10'h18d == _T_15[9:0]) begin
        image_0_397 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_398 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h18e == _T_37[9:0]) begin
        image_0_398 <= io_pixelVal_in_0_7;
      end else if (10'h18e == _T_34[9:0]) begin
        image_0_398 <= io_pixelVal_in_0_6;
      end else if (10'h18e == _T_31[9:0]) begin
        image_0_398 <= io_pixelVal_in_0_5;
      end else if (10'h18e == _T_28[9:0]) begin
        image_0_398 <= io_pixelVal_in_0_4;
      end else if (10'h18e == _T_25[9:0]) begin
        image_0_398 <= io_pixelVal_in_0_3;
      end else if (10'h18e == _T_22[9:0]) begin
        image_0_398 <= io_pixelVal_in_0_2;
      end else if (10'h18e == _T_19[9:0]) begin
        image_0_398 <= io_pixelVal_in_0_1;
      end else if (10'h18e == _T_15[9:0]) begin
        image_0_398 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_399 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h18f == _T_37[9:0]) begin
        image_0_399 <= io_pixelVal_in_0_7;
      end else if (10'h18f == _T_34[9:0]) begin
        image_0_399 <= io_pixelVal_in_0_6;
      end else if (10'h18f == _T_31[9:0]) begin
        image_0_399 <= io_pixelVal_in_0_5;
      end else if (10'h18f == _T_28[9:0]) begin
        image_0_399 <= io_pixelVal_in_0_4;
      end else if (10'h18f == _T_25[9:0]) begin
        image_0_399 <= io_pixelVal_in_0_3;
      end else if (10'h18f == _T_22[9:0]) begin
        image_0_399 <= io_pixelVal_in_0_2;
      end else if (10'h18f == _T_19[9:0]) begin
        image_0_399 <= io_pixelVal_in_0_1;
      end else if (10'h18f == _T_15[9:0]) begin
        image_0_399 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_400 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h190 == _T_37[9:0]) begin
        image_0_400 <= io_pixelVal_in_0_7;
      end else if (10'h190 == _T_34[9:0]) begin
        image_0_400 <= io_pixelVal_in_0_6;
      end else if (10'h190 == _T_31[9:0]) begin
        image_0_400 <= io_pixelVal_in_0_5;
      end else if (10'h190 == _T_28[9:0]) begin
        image_0_400 <= io_pixelVal_in_0_4;
      end else if (10'h190 == _T_25[9:0]) begin
        image_0_400 <= io_pixelVal_in_0_3;
      end else if (10'h190 == _T_22[9:0]) begin
        image_0_400 <= io_pixelVal_in_0_2;
      end else if (10'h190 == _T_19[9:0]) begin
        image_0_400 <= io_pixelVal_in_0_1;
      end else if (10'h190 == _T_15[9:0]) begin
        image_0_400 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_401 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h191 == _T_37[9:0]) begin
        image_0_401 <= io_pixelVal_in_0_7;
      end else if (10'h191 == _T_34[9:0]) begin
        image_0_401 <= io_pixelVal_in_0_6;
      end else if (10'h191 == _T_31[9:0]) begin
        image_0_401 <= io_pixelVal_in_0_5;
      end else if (10'h191 == _T_28[9:0]) begin
        image_0_401 <= io_pixelVal_in_0_4;
      end else if (10'h191 == _T_25[9:0]) begin
        image_0_401 <= io_pixelVal_in_0_3;
      end else if (10'h191 == _T_22[9:0]) begin
        image_0_401 <= io_pixelVal_in_0_2;
      end else if (10'h191 == _T_19[9:0]) begin
        image_0_401 <= io_pixelVal_in_0_1;
      end else if (10'h191 == _T_15[9:0]) begin
        image_0_401 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_402 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h192 == _T_37[9:0]) begin
        image_0_402 <= io_pixelVal_in_0_7;
      end else if (10'h192 == _T_34[9:0]) begin
        image_0_402 <= io_pixelVal_in_0_6;
      end else if (10'h192 == _T_31[9:0]) begin
        image_0_402 <= io_pixelVal_in_0_5;
      end else if (10'h192 == _T_28[9:0]) begin
        image_0_402 <= io_pixelVal_in_0_4;
      end else if (10'h192 == _T_25[9:0]) begin
        image_0_402 <= io_pixelVal_in_0_3;
      end else if (10'h192 == _T_22[9:0]) begin
        image_0_402 <= io_pixelVal_in_0_2;
      end else if (10'h192 == _T_19[9:0]) begin
        image_0_402 <= io_pixelVal_in_0_1;
      end else if (10'h192 == _T_15[9:0]) begin
        image_0_402 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_403 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h193 == _T_37[9:0]) begin
        image_0_403 <= io_pixelVal_in_0_7;
      end else if (10'h193 == _T_34[9:0]) begin
        image_0_403 <= io_pixelVal_in_0_6;
      end else if (10'h193 == _T_31[9:0]) begin
        image_0_403 <= io_pixelVal_in_0_5;
      end else if (10'h193 == _T_28[9:0]) begin
        image_0_403 <= io_pixelVal_in_0_4;
      end else if (10'h193 == _T_25[9:0]) begin
        image_0_403 <= io_pixelVal_in_0_3;
      end else if (10'h193 == _T_22[9:0]) begin
        image_0_403 <= io_pixelVal_in_0_2;
      end else if (10'h193 == _T_19[9:0]) begin
        image_0_403 <= io_pixelVal_in_0_1;
      end else if (10'h193 == _T_15[9:0]) begin
        image_0_403 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_404 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h194 == _T_37[9:0]) begin
        image_0_404 <= io_pixelVal_in_0_7;
      end else if (10'h194 == _T_34[9:0]) begin
        image_0_404 <= io_pixelVal_in_0_6;
      end else if (10'h194 == _T_31[9:0]) begin
        image_0_404 <= io_pixelVal_in_0_5;
      end else if (10'h194 == _T_28[9:0]) begin
        image_0_404 <= io_pixelVal_in_0_4;
      end else if (10'h194 == _T_25[9:0]) begin
        image_0_404 <= io_pixelVal_in_0_3;
      end else if (10'h194 == _T_22[9:0]) begin
        image_0_404 <= io_pixelVal_in_0_2;
      end else if (10'h194 == _T_19[9:0]) begin
        image_0_404 <= io_pixelVal_in_0_1;
      end else if (10'h194 == _T_15[9:0]) begin
        image_0_404 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_405 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h195 == _T_37[9:0]) begin
        image_0_405 <= io_pixelVal_in_0_7;
      end else if (10'h195 == _T_34[9:0]) begin
        image_0_405 <= io_pixelVal_in_0_6;
      end else if (10'h195 == _T_31[9:0]) begin
        image_0_405 <= io_pixelVal_in_0_5;
      end else if (10'h195 == _T_28[9:0]) begin
        image_0_405 <= io_pixelVal_in_0_4;
      end else if (10'h195 == _T_25[9:0]) begin
        image_0_405 <= io_pixelVal_in_0_3;
      end else if (10'h195 == _T_22[9:0]) begin
        image_0_405 <= io_pixelVal_in_0_2;
      end else if (10'h195 == _T_19[9:0]) begin
        image_0_405 <= io_pixelVal_in_0_1;
      end else if (10'h195 == _T_15[9:0]) begin
        image_0_405 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_406 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h196 == _T_37[9:0]) begin
        image_0_406 <= io_pixelVal_in_0_7;
      end else if (10'h196 == _T_34[9:0]) begin
        image_0_406 <= io_pixelVal_in_0_6;
      end else if (10'h196 == _T_31[9:0]) begin
        image_0_406 <= io_pixelVal_in_0_5;
      end else if (10'h196 == _T_28[9:0]) begin
        image_0_406 <= io_pixelVal_in_0_4;
      end else if (10'h196 == _T_25[9:0]) begin
        image_0_406 <= io_pixelVal_in_0_3;
      end else if (10'h196 == _T_22[9:0]) begin
        image_0_406 <= io_pixelVal_in_0_2;
      end else if (10'h196 == _T_19[9:0]) begin
        image_0_406 <= io_pixelVal_in_0_1;
      end else if (10'h196 == _T_15[9:0]) begin
        image_0_406 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_407 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h197 == _T_37[9:0]) begin
        image_0_407 <= io_pixelVal_in_0_7;
      end else if (10'h197 == _T_34[9:0]) begin
        image_0_407 <= io_pixelVal_in_0_6;
      end else if (10'h197 == _T_31[9:0]) begin
        image_0_407 <= io_pixelVal_in_0_5;
      end else if (10'h197 == _T_28[9:0]) begin
        image_0_407 <= io_pixelVal_in_0_4;
      end else if (10'h197 == _T_25[9:0]) begin
        image_0_407 <= io_pixelVal_in_0_3;
      end else if (10'h197 == _T_22[9:0]) begin
        image_0_407 <= io_pixelVal_in_0_2;
      end else if (10'h197 == _T_19[9:0]) begin
        image_0_407 <= io_pixelVal_in_0_1;
      end else if (10'h197 == _T_15[9:0]) begin
        image_0_407 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_408 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h198 == _T_37[9:0]) begin
        image_0_408 <= io_pixelVal_in_0_7;
      end else if (10'h198 == _T_34[9:0]) begin
        image_0_408 <= io_pixelVal_in_0_6;
      end else if (10'h198 == _T_31[9:0]) begin
        image_0_408 <= io_pixelVal_in_0_5;
      end else if (10'h198 == _T_28[9:0]) begin
        image_0_408 <= io_pixelVal_in_0_4;
      end else if (10'h198 == _T_25[9:0]) begin
        image_0_408 <= io_pixelVal_in_0_3;
      end else if (10'h198 == _T_22[9:0]) begin
        image_0_408 <= io_pixelVal_in_0_2;
      end else if (10'h198 == _T_19[9:0]) begin
        image_0_408 <= io_pixelVal_in_0_1;
      end else if (10'h198 == _T_15[9:0]) begin
        image_0_408 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_409 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h199 == _T_37[9:0]) begin
        image_0_409 <= io_pixelVal_in_0_7;
      end else if (10'h199 == _T_34[9:0]) begin
        image_0_409 <= io_pixelVal_in_0_6;
      end else if (10'h199 == _T_31[9:0]) begin
        image_0_409 <= io_pixelVal_in_0_5;
      end else if (10'h199 == _T_28[9:0]) begin
        image_0_409 <= io_pixelVal_in_0_4;
      end else if (10'h199 == _T_25[9:0]) begin
        image_0_409 <= io_pixelVal_in_0_3;
      end else if (10'h199 == _T_22[9:0]) begin
        image_0_409 <= io_pixelVal_in_0_2;
      end else if (10'h199 == _T_19[9:0]) begin
        image_0_409 <= io_pixelVal_in_0_1;
      end else if (10'h199 == _T_15[9:0]) begin
        image_0_409 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_410 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h19a == _T_37[9:0]) begin
        image_0_410 <= io_pixelVal_in_0_7;
      end else if (10'h19a == _T_34[9:0]) begin
        image_0_410 <= io_pixelVal_in_0_6;
      end else if (10'h19a == _T_31[9:0]) begin
        image_0_410 <= io_pixelVal_in_0_5;
      end else if (10'h19a == _T_28[9:0]) begin
        image_0_410 <= io_pixelVal_in_0_4;
      end else if (10'h19a == _T_25[9:0]) begin
        image_0_410 <= io_pixelVal_in_0_3;
      end else if (10'h19a == _T_22[9:0]) begin
        image_0_410 <= io_pixelVal_in_0_2;
      end else if (10'h19a == _T_19[9:0]) begin
        image_0_410 <= io_pixelVal_in_0_1;
      end else if (10'h19a == _T_15[9:0]) begin
        image_0_410 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_411 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h19b == _T_37[9:0]) begin
        image_0_411 <= io_pixelVal_in_0_7;
      end else if (10'h19b == _T_34[9:0]) begin
        image_0_411 <= io_pixelVal_in_0_6;
      end else if (10'h19b == _T_31[9:0]) begin
        image_0_411 <= io_pixelVal_in_0_5;
      end else if (10'h19b == _T_28[9:0]) begin
        image_0_411 <= io_pixelVal_in_0_4;
      end else if (10'h19b == _T_25[9:0]) begin
        image_0_411 <= io_pixelVal_in_0_3;
      end else if (10'h19b == _T_22[9:0]) begin
        image_0_411 <= io_pixelVal_in_0_2;
      end else if (10'h19b == _T_19[9:0]) begin
        image_0_411 <= io_pixelVal_in_0_1;
      end else if (10'h19b == _T_15[9:0]) begin
        image_0_411 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_412 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h19c == _T_37[9:0]) begin
        image_0_412 <= io_pixelVal_in_0_7;
      end else if (10'h19c == _T_34[9:0]) begin
        image_0_412 <= io_pixelVal_in_0_6;
      end else if (10'h19c == _T_31[9:0]) begin
        image_0_412 <= io_pixelVal_in_0_5;
      end else if (10'h19c == _T_28[9:0]) begin
        image_0_412 <= io_pixelVal_in_0_4;
      end else if (10'h19c == _T_25[9:0]) begin
        image_0_412 <= io_pixelVal_in_0_3;
      end else if (10'h19c == _T_22[9:0]) begin
        image_0_412 <= io_pixelVal_in_0_2;
      end else if (10'h19c == _T_19[9:0]) begin
        image_0_412 <= io_pixelVal_in_0_1;
      end else if (10'h19c == _T_15[9:0]) begin
        image_0_412 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_413 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h19d == _T_37[9:0]) begin
        image_0_413 <= io_pixelVal_in_0_7;
      end else if (10'h19d == _T_34[9:0]) begin
        image_0_413 <= io_pixelVal_in_0_6;
      end else if (10'h19d == _T_31[9:0]) begin
        image_0_413 <= io_pixelVal_in_0_5;
      end else if (10'h19d == _T_28[9:0]) begin
        image_0_413 <= io_pixelVal_in_0_4;
      end else if (10'h19d == _T_25[9:0]) begin
        image_0_413 <= io_pixelVal_in_0_3;
      end else if (10'h19d == _T_22[9:0]) begin
        image_0_413 <= io_pixelVal_in_0_2;
      end else if (10'h19d == _T_19[9:0]) begin
        image_0_413 <= io_pixelVal_in_0_1;
      end else if (10'h19d == _T_15[9:0]) begin
        image_0_413 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_414 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h19e == _T_37[9:0]) begin
        image_0_414 <= io_pixelVal_in_0_7;
      end else if (10'h19e == _T_34[9:0]) begin
        image_0_414 <= io_pixelVal_in_0_6;
      end else if (10'h19e == _T_31[9:0]) begin
        image_0_414 <= io_pixelVal_in_0_5;
      end else if (10'h19e == _T_28[9:0]) begin
        image_0_414 <= io_pixelVal_in_0_4;
      end else if (10'h19e == _T_25[9:0]) begin
        image_0_414 <= io_pixelVal_in_0_3;
      end else if (10'h19e == _T_22[9:0]) begin
        image_0_414 <= io_pixelVal_in_0_2;
      end else if (10'h19e == _T_19[9:0]) begin
        image_0_414 <= io_pixelVal_in_0_1;
      end else if (10'h19e == _T_15[9:0]) begin
        image_0_414 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_415 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h19f == _T_37[9:0]) begin
        image_0_415 <= io_pixelVal_in_0_7;
      end else if (10'h19f == _T_34[9:0]) begin
        image_0_415 <= io_pixelVal_in_0_6;
      end else if (10'h19f == _T_31[9:0]) begin
        image_0_415 <= io_pixelVal_in_0_5;
      end else if (10'h19f == _T_28[9:0]) begin
        image_0_415 <= io_pixelVal_in_0_4;
      end else if (10'h19f == _T_25[9:0]) begin
        image_0_415 <= io_pixelVal_in_0_3;
      end else if (10'h19f == _T_22[9:0]) begin
        image_0_415 <= io_pixelVal_in_0_2;
      end else if (10'h19f == _T_19[9:0]) begin
        image_0_415 <= io_pixelVal_in_0_1;
      end else if (10'h19f == _T_15[9:0]) begin
        image_0_415 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_416 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1a0 == _T_37[9:0]) begin
        image_0_416 <= io_pixelVal_in_0_7;
      end else if (10'h1a0 == _T_34[9:0]) begin
        image_0_416 <= io_pixelVal_in_0_6;
      end else if (10'h1a0 == _T_31[9:0]) begin
        image_0_416 <= io_pixelVal_in_0_5;
      end else if (10'h1a0 == _T_28[9:0]) begin
        image_0_416 <= io_pixelVal_in_0_4;
      end else if (10'h1a0 == _T_25[9:0]) begin
        image_0_416 <= io_pixelVal_in_0_3;
      end else if (10'h1a0 == _T_22[9:0]) begin
        image_0_416 <= io_pixelVal_in_0_2;
      end else if (10'h1a0 == _T_19[9:0]) begin
        image_0_416 <= io_pixelVal_in_0_1;
      end else if (10'h1a0 == _T_15[9:0]) begin
        image_0_416 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_417 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1a1 == _T_37[9:0]) begin
        image_0_417 <= io_pixelVal_in_0_7;
      end else if (10'h1a1 == _T_34[9:0]) begin
        image_0_417 <= io_pixelVal_in_0_6;
      end else if (10'h1a1 == _T_31[9:0]) begin
        image_0_417 <= io_pixelVal_in_0_5;
      end else if (10'h1a1 == _T_28[9:0]) begin
        image_0_417 <= io_pixelVal_in_0_4;
      end else if (10'h1a1 == _T_25[9:0]) begin
        image_0_417 <= io_pixelVal_in_0_3;
      end else if (10'h1a1 == _T_22[9:0]) begin
        image_0_417 <= io_pixelVal_in_0_2;
      end else if (10'h1a1 == _T_19[9:0]) begin
        image_0_417 <= io_pixelVal_in_0_1;
      end else if (10'h1a1 == _T_15[9:0]) begin
        image_0_417 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_418 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1a2 == _T_37[9:0]) begin
        image_0_418 <= io_pixelVal_in_0_7;
      end else if (10'h1a2 == _T_34[9:0]) begin
        image_0_418 <= io_pixelVal_in_0_6;
      end else if (10'h1a2 == _T_31[9:0]) begin
        image_0_418 <= io_pixelVal_in_0_5;
      end else if (10'h1a2 == _T_28[9:0]) begin
        image_0_418 <= io_pixelVal_in_0_4;
      end else if (10'h1a2 == _T_25[9:0]) begin
        image_0_418 <= io_pixelVal_in_0_3;
      end else if (10'h1a2 == _T_22[9:0]) begin
        image_0_418 <= io_pixelVal_in_0_2;
      end else if (10'h1a2 == _T_19[9:0]) begin
        image_0_418 <= io_pixelVal_in_0_1;
      end else if (10'h1a2 == _T_15[9:0]) begin
        image_0_418 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_419 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1a3 == _T_37[9:0]) begin
        image_0_419 <= io_pixelVal_in_0_7;
      end else if (10'h1a3 == _T_34[9:0]) begin
        image_0_419 <= io_pixelVal_in_0_6;
      end else if (10'h1a3 == _T_31[9:0]) begin
        image_0_419 <= io_pixelVal_in_0_5;
      end else if (10'h1a3 == _T_28[9:0]) begin
        image_0_419 <= io_pixelVal_in_0_4;
      end else if (10'h1a3 == _T_25[9:0]) begin
        image_0_419 <= io_pixelVal_in_0_3;
      end else if (10'h1a3 == _T_22[9:0]) begin
        image_0_419 <= io_pixelVal_in_0_2;
      end else if (10'h1a3 == _T_19[9:0]) begin
        image_0_419 <= io_pixelVal_in_0_1;
      end else if (10'h1a3 == _T_15[9:0]) begin
        image_0_419 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_420 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1a4 == _T_37[9:0]) begin
        image_0_420 <= io_pixelVal_in_0_7;
      end else if (10'h1a4 == _T_34[9:0]) begin
        image_0_420 <= io_pixelVal_in_0_6;
      end else if (10'h1a4 == _T_31[9:0]) begin
        image_0_420 <= io_pixelVal_in_0_5;
      end else if (10'h1a4 == _T_28[9:0]) begin
        image_0_420 <= io_pixelVal_in_0_4;
      end else if (10'h1a4 == _T_25[9:0]) begin
        image_0_420 <= io_pixelVal_in_0_3;
      end else if (10'h1a4 == _T_22[9:0]) begin
        image_0_420 <= io_pixelVal_in_0_2;
      end else if (10'h1a4 == _T_19[9:0]) begin
        image_0_420 <= io_pixelVal_in_0_1;
      end else if (10'h1a4 == _T_15[9:0]) begin
        image_0_420 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_421 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1a5 == _T_37[9:0]) begin
        image_0_421 <= io_pixelVal_in_0_7;
      end else if (10'h1a5 == _T_34[9:0]) begin
        image_0_421 <= io_pixelVal_in_0_6;
      end else if (10'h1a5 == _T_31[9:0]) begin
        image_0_421 <= io_pixelVal_in_0_5;
      end else if (10'h1a5 == _T_28[9:0]) begin
        image_0_421 <= io_pixelVal_in_0_4;
      end else if (10'h1a5 == _T_25[9:0]) begin
        image_0_421 <= io_pixelVal_in_0_3;
      end else if (10'h1a5 == _T_22[9:0]) begin
        image_0_421 <= io_pixelVal_in_0_2;
      end else if (10'h1a5 == _T_19[9:0]) begin
        image_0_421 <= io_pixelVal_in_0_1;
      end else if (10'h1a5 == _T_15[9:0]) begin
        image_0_421 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_422 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1a6 == _T_37[9:0]) begin
        image_0_422 <= io_pixelVal_in_0_7;
      end else if (10'h1a6 == _T_34[9:0]) begin
        image_0_422 <= io_pixelVal_in_0_6;
      end else if (10'h1a6 == _T_31[9:0]) begin
        image_0_422 <= io_pixelVal_in_0_5;
      end else if (10'h1a6 == _T_28[9:0]) begin
        image_0_422 <= io_pixelVal_in_0_4;
      end else if (10'h1a6 == _T_25[9:0]) begin
        image_0_422 <= io_pixelVal_in_0_3;
      end else if (10'h1a6 == _T_22[9:0]) begin
        image_0_422 <= io_pixelVal_in_0_2;
      end else if (10'h1a6 == _T_19[9:0]) begin
        image_0_422 <= io_pixelVal_in_0_1;
      end else if (10'h1a6 == _T_15[9:0]) begin
        image_0_422 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_423 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1a7 == _T_37[9:0]) begin
        image_0_423 <= io_pixelVal_in_0_7;
      end else if (10'h1a7 == _T_34[9:0]) begin
        image_0_423 <= io_pixelVal_in_0_6;
      end else if (10'h1a7 == _T_31[9:0]) begin
        image_0_423 <= io_pixelVal_in_0_5;
      end else if (10'h1a7 == _T_28[9:0]) begin
        image_0_423 <= io_pixelVal_in_0_4;
      end else if (10'h1a7 == _T_25[9:0]) begin
        image_0_423 <= io_pixelVal_in_0_3;
      end else if (10'h1a7 == _T_22[9:0]) begin
        image_0_423 <= io_pixelVal_in_0_2;
      end else if (10'h1a7 == _T_19[9:0]) begin
        image_0_423 <= io_pixelVal_in_0_1;
      end else if (10'h1a7 == _T_15[9:0]) begin
        image_0_423 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_424 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1a8 == _T_37[9:0]) begin
        image_0_424 <= io_pixelVal_in_0_7;
      end else if (10'h1a8 == _T_34[9:0]) begin
        image_0_424 <= io_pixelVal_in_0_6;
      end else if (10'h1a8 == _T_31[9:0]) begin
        image_0_424 <= io_pixelVal_in_0_5;
      end else if (10'h1a8 == _T_28[9:0]) begin
        image_0_424 <= io_pixelVal_in_0_4;
      end else if (10'h1a8 == _T_25[9:0]) begin
        image_0_424 <= io_pixelVal_in_0_3;
      end else if (10'h1a8 == _T_22[9:0]) begin
        image_0_424 <= io_pixelVal_in_0_2;
      end else if (10'h1a8 == _T_19[9:0]) begin
        image_0_424 <= io_pixelVal_in_0_1;
      end else if (10'h1a8 == _T_15[9:0]) begin
        image_0_424 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_425 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1a9 == _T_37[9:0]) begin
        image_0_425 <= io_pixelVal_in_0_7;
      end else if (10'h1a9 == _T_34[9:0]) begin
        image_0_425 <= io_pixelVal_in_0_6;
      end else if (10'h1a9 == _T_31[9:0]) begin
        image_0_425 <= io_pixelVal_in_0_5;
      end else if (10'h1a9 == _T_28[9:0]) begin
        image_0_425 <= io_pixelVal_in_0_4;
      end else if (10'h1a9 == _T_25[9:0]) begin
        image_0_425 <= io_pixelVal_in_0_3;
      end else if (10'h1a9 == _T_22[9:0]) begin
        image_0_425 <= io_pixelVal_in_0_2;
      end else if (10'h1a9 == _T_19[9:0]) begin
        image_0_425 <= io_pixelVal_in_0_1;
      end else if (10'h1a9 == _T_15[9:0]) begin
        image_0_425 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_426 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1aa == _T_37[9:0]) begin
        image_0_426 <= io_pixelVal_in_0_7;
      end else if (10'h1aa == _T_34[9:0]) begin
        image_0_426 <= io_pixelVal_in_0_6;
      end else if (10'h1aa == _T_31[9:0]) begin
        image_0_426 <= io_pixelVal_in_0_5;
      end else if (10'h1aa == _T_28[9:0]) begin
        image_0_426 <= io_pixelVal_in_0_4;
      end else if (10'h1aa == _T_25[9:0]) begin
        image_0_426 <= io_pixelVal_in_0_3;
      end else if (10'h1aa == _T_22[9:0]) begin
        image_0_426 <= io_pixelVal_in_0_2;
      end else if (10'h1aa == _T_19[9:0]) begin
        image_0_426 <= io_pixelVal_in_0_1;
      end else if (10'h1aa == _T_15[9:0]) begin
        image_0_426 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_427 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1ab == _T_37[9:0]) begin
        image_0_427 <= io_pixelVal_in_0_7;
      end else if (10'h1ab == _T_34[9:0]) begin
        image_0_427 <= io_pixelVal_in_0_6;
      end else if (10'h1ab == _T_31[9:0]) begin
        image_0_427 <= io_pixelVal_in_0_5;
      end else if (10'h1ab == _T_28[9:0]) begin
        image_0_427 <= io_pixelVal_in_0_4;
      end else if (10'h1ab == _T_25[9:0]) begin
        image_0_427 <= io_pixelVal_in_0_3;
      end else if (10'h1ab == _T_22[9:0]) begin
        image_0_427 <= io_pixelVal_in_0_2;
      end else if (10'h1ab == _T_19[9:0]) begin
        image_0_427 <= io_pixelVal_in_0_1;
      end else if (10'h1ab == _T_15[9:0]) begin
        image_0_427 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_428 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1ac == _T_37[9:0]) begin
        image_0_428 <= io_pixelVal_in_0_7;
      end else if (10'h1ac == _T_34[9:0]) begin
        image_0_428 <= io_pixelVal_in_0_6;
      end else if (10'h1ac == _T_31[9:0]) begin
        image_0_428 <= io_pixelVal_in_0_5;
      end else if (10'h1ac == _T_28[9:0]) begin
        image_0_428 <= io_pixelVal_in_0_4;
      end else if (10'h1ac == _T_25[9:0]) begin
        image_0_428 <= io_pixelVal_in_0_3;
      end else if (10'h1ac == _T_22[9:0]) begin
        image_0_428 <= io_pixelVal_in_0_2;
      end else if (10'h1ac == _T_19[9:0]) begin
        image_0_428 <= io_pixelVal_in_0_1;
      end else if (10'h1ac == _T_15[9:0]) begin
        image_0_428 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_429 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1ad == _T_37[9:0]) begin
        image_0_429 <= io_pixelVal_in_0_7;
      end else if (10'h1ad == _T_34[9:0]) begin
        image_0_429 <= io_pixelVal_in_0_6;
      end else if (10'h1ad == _T_31[9:0]) begin
        image_0_429 <= io_pixelVal_in_0_5;
      end else if (10'h1ad == _T_28[9:0]) begin
        image_0_429 <= io_pixelVal_in_0_4;
      end else if (10'h1ad == _T_25[9:0]) begin
        image_0_429 <= io_pixelVal_in_0_3;
      end else if (10'h1ad == _T_22[9:0]) begin
        image_0_429 <= io_pixelVal_in_0_2;
      end else if (10'h1ad == _T_19[9:0]) begin
        image_0_429 <= io_pixelVal_in_0_1;
      end else if (10'h1ad == _T_15[9:0]) begin
        image_0_429 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_430 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1ae == _T_37[9:0]) begin
        image_0_430 <= io_pixelVal_in_0_7;
      end else if (10'h1ae == _T_34[9:0]) begin
        image_0_430 <= io_pixelVal_in_0_6;
      end else if (10'h1ae == _T_31[9:0]) begin
        image_0_430 <= io_pixelVal_in_0_5;
      end else if (10'h1ae == _T_28[9:0]) begin
        image_0_430 <= io_pixelVal_in_0_4;
      end else if (10'h1ae == _T_25[9:0]) begin
        image_0_430 <= io_pixelVal_in_0_3;
      end else if (10'h1ae == _T_22[9:0]) begin
        image_0_430 <= io_pixelVal_in_0_2;
      end else if (10'h1ae == _T_19[9:0]) begin
        image_0_430 <= io_pixelVal_in_0_1;
      end else if (10'h1ae == _T_15[9:0]) begin
        image_0_430 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_431 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1af == _T_37[9:0]) begin
        image_0_431 <= io_pixelVal_in_0_7;
      end else if (10'h1af == _T_34[9:0]) begin
        image_0_431 <= io_pixelVal_in_0_6;
      end else if (10'h1af == _T_31[9:0]) begin
        image_0_431 <= io_pixelVal_in_0_5;
      end else if (10'h1af == _T_28[9:0]) begin
        image_0_431 <= io_pixelVal_in_0_4;
      end else if (10'h1af == _T_25[9:0]) begin
        image_0_431 <= io_pixelVal_in_0_3;
      end else if (10'h1af == _T_22[9:0]) begin
        image_0_431 <= io_pixelVal_in_0_2;
      end else if (10'h1af == _T_19[9:0]) begin
        image_0_431 <= io_pixelVal_in_0_1;
      end else if (10'h1af == _T_15[9:0]) begin
        image_0_431 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_432 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1b0 == _T_37[9:0]) begin
        image_0_432 <= io_pixelVal_in_0_7;
      end else if (10'h1b0 == _T_34[9:0]) begin
        image_0_432 <= io_pixelVal_in_0_6;
      end else if (10'h1b0 == _T_31[9:0]) begin
        image_0_432 <= io_pixelVal_in_0_5;
      end else if (10'h1b0 == _T_28[9:0]) begin
        image_0_432 <= io_pixelVal_in_0_4;
      end else if (10'h1b0 == _T_25[9:0]) begin
        image_0_432 <= io_pixelVal_in_0_3;
      end else if (10'h1b0 == _T_22[9:0]) begin
        image_0_432 <= io_pixelVal_in_0_2;
      end else if (10'h1b0 == _T_19[9:0]) begin
        image_0_432 <= io_pixelVal_in_0_1;
      end else if (10'h1b0 == _T_15[9:0]) begin
        image_0_432 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_433 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1b1 == _T_37[9:0]) begin
        image_0_433 <= io_pixelVal_in_0_7;
      end else if (10'h1b1 == _T_34[9:0]) begin
        image_0_433 <= io_pixelVal_in_0_6;
      end else if (10'h1b1 == _T_31[9:0]) begin
        image_0_433 <= io_pixelVal_in_0_5;
      end else if (10'h1b1 == _T_28[9:0]) begin
        image_0_433 <= io_pixelVal_in_0_4;
      end else if (10'h1b1 == _T_25[9:0]) begin
        image_0_433 <= io_pixelVal_in_0_3;
      end else if (10'h1b1 == _T_22[9:0]) begin
        image_0_433 <= io_pixelVal_in_0_2;
      end else if (10'h1b1 == _T_19[9:0]) begin
        image_0_433 <= io_pixelVal_in_0_1;
      end else if (10'h1b1 == _T_15[9:0]) begin
        image_0_433 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_434 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1b2 == _T_37[9:0]) begin
        image_0_434 <= io_pixelVal_in_0_7;
      end else if (10'h1b2 == _T_34[9:0]) begin
        image_0_434 <= io_pixelVal_in_0_6;
      end else if (10'h1b2 == _T_31[9:0]) begin
        image_0_434 <= io_pixelVal_in_0_5;
      end else if (10'h1b2 == _T_28[9:0]) begin
        image_0_434 <= io_pixelVal_in_0_4;
      end else if (10'h1b2 == _T_25[9:0]) begin
        image_0_434 <= io_pixelVal_in_0_3;
      end else if (10'h1b2 == _T_22[9:0]) begin
        image_0_434 <= io_pixelVal_in_0_2;
      end else if (10'h1b2 == _T_19[9:0]) begin
        image_0_434 <= io_pixelVal_in_0_1;
      end else if (10'h1b2 == _T_15[9:0]) begin
        image_0_434 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_435 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1b3 == _T_37[9:0]) begin
        image_0_435 <= io_pixelVal_in_0_7;
      end else if (10'h1b3 == _T_34[9:0]) begin
        image_0_435 <= io_pixelVal_in_0_6;
      end else if (10'h1b3 == _T_31[9:0]) begin
        image_0_435 <= io_pixelVal_in_0_5;
      end else if (10'h1b3 == _T_28[9:0]) begin
        image_0_435 <= io_pixelVal_in_0_4;
      end else if (10'h1b3 == _T_25[9:0]) begin
        image_0_435 <= io_pixelVal_in_0_3;
      end else if (10'h1b3 == _T_22[9:0]) begin
        image_0_435 <= io_pixelVal_in_0_2;
      end else if (10'h1b3 == _T_19[9:0]) begin
        image_0_435 <= io_pixelVal_in_0_1;
      end else if (10'h1b3 == _T_15[9:0]) begin
        image_0_435 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_436 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1b4 == _T_37[9:0]) begin
        image_0_436 <= io_pixelVal_in_0_7;
      end else if (10'h1b4 == _T_34[9:0]) begin
        image_0_436 <= io_pixelVal_in_0_6;
      end else if (10'h1b4 == _T_31[9:0]) begin
        image_0_436 <= io_pixelVal_in_0_5;
      end else if (10'h1b4 == _T_28[9:0]) begin
        image_0_436 <= io_pixelVal_in_0_4;
      end else if (10'h1b4 == _T_25[9:0]) begin
        image_0_436 <= io_pixelVal_in_0_3;
      end else if (10'h1b4 == _T_22[9:0]) begin
        image_0_436 <= io_pixelVal_in_0_2;
      end else if (10'h1b4 == _T_19[9:0]) begin
        image_0_436 <= io_pixelVal_in_0_1;
      end else if (10'h1b4 == _T_15[9:0]) begin
        image_0_436 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_437 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1b5 == _T_37[9:0]) begin
        image_0_437 <= io_pixelVal_in_0_7;
      end else if (10'h1b5 == _T_34[9:0]) begin
        image_0_437 <= io_pixelVal_in_0_6;
      end else if (10'h1b5 == _T_31[9:0]) begin
        image_0_437 <= io_pixelVal_in_0_5;
      end else if (10'h1b5 == _T_28[9:0]) begin
        image_0_437 <= io_pixelVal_in_0_4;
      end else if (10'h1b5 == _T_25[9:0]) begin
        image_0_437 <= io_pixelVal_in_0_3;
      end else if (10'h1b5 == _T_22[9:0]) begin
        image_0_437 <= io_pixelVal_in_0_2;
      end else if (10'h1b5 == _T_19[9:0]) begin
        image_0_437 <= io_pixelVal_in_0_1;
      end else if (10'h1b5 == _T_15[9:0]) begin
        image_0_437 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_438 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1b6 == _T_37[9:0]) begin
        image_0_438 <= io_pixelVal_in_0_7;
      end else if (10'h1b6 == _T_34[9:0]) begin
        image_0_438 <= io_pixelVal_in_0_6;
      end else if (10'h1b6 == _T_31[9:0]) begin
        image_0_438 <= io_pixelVal_in_0_5;
      end else if (10'h1b6 == _T_28[9:0]) begin
        image_0_438 <= io_pixelVal_in_0_4;
      end else if (10'h1b6 == _T_25[9:0]) begin
        image_0_438 <= io_pixelVal_in_0_3;
      end else if (10'h1b6 == _T_22[9:0]) begin
        image_0_438 <= io_pixelVal_in_0_2;
      end else if (10'h1b6 == _T_19[9:0]) begin
        image_0_438 <= io_pixelVal_in_0_1;
      end else if (10'h1b6 == _T_15[9:0]) begin
        image_0_438 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_439 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1b7 == _T_37[9:0]) begin
        image_0_439 <= io_pixelVal_in_0_7;
      end else if (10'h1b7 == _T_34[9:0]) begin
        image_0_439 <= io_pixelVal_in_0_6;
      end else if (10'h1b7 == _T_31[9:0]) begin
        image_0_439 <= io_pixelVal_in_0_5;
      end else if (10'h1b7 == _T_28[9:0]) begin
        image_0_439 <= io_pixelVal_in_0_4;
      end else if (10'h1b7 == _T_25[9:0]) begin
        image_0_439 <= io_pixelVal_in_0_3;
      end else if (10'h1b7 == _T_22[9:0]) begin
        image_0_439 <= io_pixelVal_in_0_2;
      end else if (10'h1b7 == _T_19[9:0]) begin
        image_0_439 <= io_pixelVal_in_0_1;
      end else if (10'h1b7 == _T_15[9:0]) begin
        image_0_439 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_440 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1b8 == _T_37[9:0]) begin
        image_0_440 <= io_pixelVal_in_0_7;
      end else if (10'h1b8 == _T_34[9:0]) begin
        image_0_440 <= io_pixelVal_in_0_6;
      end else if (10'h1b8 == _T_31[9:0]) begin
        image_0_440 <= io_pixelVal_in_0_5;
      end else if (10'h1b8 == _T_28[9:0]) begin
        image_0_440 <= io_pixelVal_in_0_4;
      end else if (10'h1b8 == _T_25[9:0]) begin
        image_0_440 <= io_pixelVal_in_0_3;
      end else if (10'h1b8 == _T_22[9:0]) begin
        image_0_440 <= io_pixelVal_in_0_2;
      end else if (10'h1b8 == _T_19[9:0]) begin
        image_0_440 <= io_pixelVal_in_0_1;
      end else if (10'h1b8 == _T_15[9:0]) begin
        image_0_440 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_441 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1b9 == _T_37[9:0]) begin
        image_0_441 <= io_pixelVal_in_0_7;
      end else if (10'h1b9 == _T_34[9:0]) begin
        image_0_441 <= io_pixelVal_in_0_6;
      end else if (10'h1b9 == _T_31[9:0]) begin
        image_0_441 <= io_pixelVal_in_0_5;
      end else if (10'h1b9 == _T_28[9:0]) begin
        image_0_441 <= io_pixelVal_in_0_4;
      end else if (10'h1b9 == _T_25[9:0]) begin
        image_0_441 <= io_pixelVal_in_0_3;
      end else if (10'h1b9 == _T_22[9:0]) begin
        image_0_441 <= io_pixelVal_in_0_2;
      end else if (10'h1b9 == _T_19[9:0]) begin
        image_0_441 <= io_pixelVal_in_0_1;
      end else if (10'h1b9 == _T_15[9:0]) begin
        image_0_441 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_442 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1ba == _T_37[9:0]) begin
        image_0_442 <= io_pixelVal_in_0_7;
      end else if (10'h1ba == _T_34[9:0]) begin
        image_0_442 <= io_pixelVal_in_0_6;
      end else if (10'h1ba == _T_31[9:0]) begin
        image_0_442 <= io_pixelVal_in_0_5;
      end else if (10'h1ba == _T_28[9:0]) begin
        image_0_442 <= io_pixelVal_in_0_4;
      end else if (10'h1ba == _T_25[9:0]) begin
        image_0_442 <= io_pixelVal_in_0_3;
      end else if (10'h1ba == _T_22[9:0]) begin
        image_0_442 <= io_pixelVal_in_0_2;
      end else if (10'h1ba == _T_19[9:0]) begin
        image_0_442 <= io_pixelVal_in_0_1;
      end else if (10'h1ba == _T_15[9:0]) begin
        image_0_442 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_443 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1bb == _T_37[9:0]) begin
        image_0_443 <= io_pixelVal_in_0_7;
      end else if (10'h1bb == _T_34[9:0]) begin
        image_0_443 <= io_pixelVal_in_0_6;
      end else if (10'h1bb == _T_31[9:0]) begin
        image_0_443 <= io_pixelVal_in_0_5;
      end else if (10'h1bb == _T_28[9:0]) begin
        image_0_443 <= io_pixelVal_in_0_4;
      end else if (10'h1bb == _T_25[9:0]) begin
        image_0_443 <= io_pixelVal_in_0_3;
      end else if (10'h1bb == _T_22[9:0]) begin
        image_0_443 <= io_pixelVal_in_0_2;
      end else if (10'h1bb == _T_19[9:0]) begin
        image_0_443 <= io_pixelVal_in_0_1;
      end else if (10'h1bb == _T_15[9:0]) begin
        image_0_443 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_444 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1bc == _T_37[9:0]) begin
        image_0_444 <= io_pixelVal_in_0_7;
      end else if (10'h1bc == _T_34[9:0]) begin
        image_0_444 <= io_pixelVal_in_0_6;
      end else if (10'h1bc == _T_31[9:0]) begin
        image_0_444 <= io_pixelVal_in_0_5;
      end else if (10'h1bc == _T_28[9:0]) begin
        image_0_444 <= io_pixelVal_in_0_4;
      end else if (10'h1bc == _T_25[9:0]) begin
        image_0_444 <= io_pixelVal_in_0_3;
      end else if (10'h1bc == _T_22[9:0]) begin
        image_0_444 <= io_pixelVal_in_0_2;
      end else if (10'h1bc == _T_19[9:0]) begin
        image_0_444 <= io_pixelVal_in_0_1;
      end else if (10'h1bc == _T_15[9:0]) begin
        image_0_444 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_445 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1bd == _T_37[9:0]) begin
        image_0_445 <= io_pixelVal_in_0_7;
      end else if (10'h1bd == _T_34[9:0]) begin
        image_0_445 <= io_pixelVal_in_0_6;
      end else if (10'h1bd == _T_31[9:0]) begin
        image_0_445 <= io_pixelVal_in_0_5;
      end else if (10'h1bd == _T_28[9:0]) begin
        image_0_445 <= io_pixelVal_in_0_4;
      end else if (10'h1bd == _T_25[9:0]) begin
        image_0_445 <= io_pixelVal_in_0_3;
      end else if (10'h1bd == _T_22[9:0]) begin
        image_0_445 <= io_pixelVal_in_0_2;
      end else if (10'h1bd == _T_19[9:0]) begin
        image_0_445 <= io_pixelVal_in_0_1;
      end else if (10'h1bd == _T_15[9:0]) begin
        image_0_445 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_446 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1be == _T_37[9:0]) begin
        image_0_446 <= io_pixelVal_in_0_7;
      end else if (10'h1be == _T_34[9:0]) begin
        image_0_446 <= io_pixelVal_in_0_6;
      end else if (10'h1be == _T_31[9:0]) begin
        image_0_446 <= io_pixelVal_in_0_5;
      end else if (10'h1be == _T_28[9:0]) begin
        image_0_446 <= io_pixelVal_in_0_4;
      end else if (10'h1be == _T_25[9:0]) begin
        image_0_446 <= io_pixelVal_in_0_3;
      end else if (10'h1be == _T_22[9:0]) begin
        image_0_446 <= io_pixelVal_in_0_2;
      end else if (10'h1be == _T_19[9:0]) begin
        image_0_446 <= io_pixelVal_in_0_1;
      end else if (10'h1be == _T_15[9:0]) begin
        image_0_446 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_447 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1bf == _T_37[9:0]) begin
        image_0_447 <= io_pixelVal_in_0_7;
      end else if (10'h1bf == _T_34[9:0]) begin
        image_0_447 <= io_pixelVal_in_0_6;
      end else if (10'h1bf == _T_31[9:0]) begin
        image_0_447 <= io_pixelVal_in_0_5;
      end else if (10'h1bf == _T_28[9:0]) begin
        image_0_447 <= io_pixelVal_in_0_4;
      end else if (10'h1bf == _T_25[9:0]) begin
        image_0_447 <= io_pixelVal_in_0_3;
      end else if (10'h1bf == _T_22[9:0]) begin
        image_0_447 <= io_pixelVal_in_0_2;
      end else if (10'h1bf == _T_19[9:0]) begin
        image_0_447 <= io_pixelVal_in_0_1;
      end else if (10'h1bf == _T_15[9:0]) begin
        image_0_447 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_448 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1c0 == _T_37[9:0]) begin
        image_0_448 <= io_pixelVal_in_0_7;
      end else if (10'h1c0 == _T_34[9:0]) begin
        image_0_448 <= io_pixelVal_in_0_6;
      end else if (10'h1c0 == _T_31[9:0]) begin
        image_0_448 <= io_pixelVal_in_0_5;
      end else if (10'h1c0 == _T_28[9:0]) begin
        image_0_448 <= io_pixelVal_in_0_4;
      end else if (10'h1c0 == _T_25[9:0]) begin
        image_0_448 <= io_pixelVal_in_0_3;
      end else if (10'h1c0 == _T_22[9:0]) begin
        image_0_448 <= io_pixelVal_in_0_2;
      end else if (10'h1c0 == _T_19[9:0]) begin
        image_0_448 <= io_pixelVal_in_0_1;
      end else if (10'h1c0 == _T_15[9:0]) begin
        image_0_448 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_449 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1c1 == _T_37[9:0]) begin
        image_0_449 <= io_pixelVal_in_0_7;
      end else if (10'h1c1 == _T_34[9:0]) begin
        image_0_449 <= io_pixelVal_in_0_6;
      end else if (10'h1c1 == _T_31[9:0]) begin
        image_0_449 <= io_pixelVal_in_0_5;
      end else if (10'h1c1 == _T_28[9:0]) begin
        image_0_449 <= io_pixelVal_in_0_4;
      end else if (10'h1c1 == _T_25[9:0]) begin
        image_0_449 <= io_pixelVal_in_0_3;
      end else if (10'h1c1 == _T_22[9:0]) begin
        image_0_449 <= io_pixelVal_in_0_2;
      end else if (10'h1c1 == _T_19[9:0]) begin
        image_0_449 <= io_pixelVal_in_0_1;
      end else if (10'h1c1 == _T_15[9:0]) begin
        image_0_449 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_450 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1c2 == _T_37[9:0]) begin
        image_0_450 <= io_pixelVal_in_0_7;
      end else if (10'h1c2 == _T_34[9:0]) begin
        image_0_450 <= io_pixelVal_in_0_6;
      end else if (10'h1c2 == _T_31[9:0]) begin
        image_0_450 <= io_pixelVal_in_0_5;
      end else if (10'h1c2 == _T_28[9:0]) begin
        image_0_450 <= io_pixelVal_in_0_4;
      end else if (10'h1c2 == _T_25[9:0]) begin
        image_0_450 <= io_pixelVal_in_0_3;
      end else if (10'h1c2 == _T_22[9:0]) begin
        image_0_450 <= io_pixelVal_in_0_2;
      end else if (10'h1c2 == _T_19[9:0]) begin
        image_0_450 <= io_pixelVal_in_0_1;
      end else if (10'h1c2 == _T_15[9:0]) begin
        image_0_450 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_451 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1c3 == _T_37[9:0]) begin
        image_0_451 <= io_pixelVal_in_0_7;
      end else if (10'h1c3 == _T_34[9:0]) begin
        image_0_451 <= io_pixelVal_in_0_6;
      end else if (10'h1c3 == _T_31[9:0]) begin
        image_0_451 <= io_pixelVal_in_0_5;
      end else if (10'h1c3 == _T_28[9:0]) begin
        image_0_451 <= io_pixelVal_in_0_4;
      end else if (10'h1c3 == _T_25[9:0]) begin
        image_0_451 <= io_pixelVal_in_0_3;
      end else if (10'h1c3 == _T_22[9:0]) begin
        image_0_451 <= io_pixelVal_in_0_2;
      end else if (10'h1c3 == _T_19[9:0]) begin
        image_0_451 <= io_pixelVal_in_0_1;
      end else if (10'h1c3 == _T_15[9:0]) begin
        image_0_451 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_452 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1c4 == _T_37[9:0]) begin
        image_0_452 <= io_pixelVal_in_0_7;
      end else if (10'h1c4 == _T_34[9:0]) begin
        image_0_452 <= io_pixelVal_in_0_6;
      end else if (10'h1c4 == _T_31[9:0]) begin
        image_0_452 <= io_pixelVal_in_0_5;
      end else if (10'h1c4 == _T_28[9:0]) begin
        image_0_452 <= io_pixelVal_in_0_4;
      end else if (10'h1c4 == _T_25[9:0]) begin
        image_0_452 <= io_pixelVal_in_0_3;
      end else if (10'h1c4 == _T_22[9:0]) begin
        image_0_452 <= io_pixelVal_in_0_2;
      end else if (10'h1c4 == _T_19[9:0]) begin
        image_0_452 <= io_pixelVal_in_0_1;
      end else if (10'h1c4 == _T_15[9:0]) begin
        image_0_452 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_453 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1c5 == _T_37[9:0]) begin
        image_0_453 <= io_pixelVal_in_0_7;
      end else if (10'h1c5 == _T_34[9:0]) begin
        image_0_453 <= io_pixelVal_in_0_6;
      end else if (10'h1c5 == _T_31[9:0]) begin
        image_0_453 <= io_pixelVal_in_0_5;
      end else if (10'h1c5 == _T_28[9:0]) begin
        image_0_453 <= io_pixelVal_in_0_4;
      end else if (10'h1c5 == _T_25[9:0]) begin
        image_0_453 <= io_pixelVal_in_0_3;
      end else if (10'h1c5 == _T_22[9:0]) begin
        image_0_453 <= io_pixelVal_in_0_2;
      end else if (10'h1c5 == _T_19[9:0]) begin
        image_0_453 <= io_pixelVal_in_0_1;
      end else if (10'h1c5 == _T_15[9:0]) begin
        image_0_453 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_454 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1c6 == _T_37[9:0]) begin
        image_0_454 <= io_pixelVal_in_0_7;
      end else if (10'h1c6 == _T_34[9:0]) begin
        image_0_454 <= io_pixelVal_in_0_6;
      end else if (10'h1c6 == _T_31[9:0]) begin
        image_0_454 <= io_pixelVal_in_0_5;
      end else if (10'h1c6 == _T_28[9:0]) begin
        image_0_454 <= io_pixelVal_in_0_4;
      end else if (10'h1c6 == _T_25[9:0]) begin
        image_0_454 <= io_pixelVal_in_0_3;
      end else if (10'h1c6 == _T_22[9:0]) begin
        image_0_454 <= io_pixelVal_in_0_2;
      end else if (10'h1c6 == _T_19[9:0]) begin
        image_0_454 <= io_pixelVal_in_0_1;
      end else if (10'h1c6 == _T_15[9:0]) begin
        image_0_454 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_455 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1c7 == _T_37[9:0]) begin
        image_0_455 <= io_pixelVal_in_0_7;
      end else if (10'h1c7 == _T_34[9:0]) begin
        image_0_455 <= io_pixelVal_in_0_6;
      end else if (10'h1c7 == _T_31[9:0]) begin
        image_0_455 <= io_pixelVal_in_0_5;
      end else if (10'h1c7 == _T_28[9:0]) begin
        image_0_455 <= io_pixelVal_in_0_4;
      end else if (10'h1c7 == _T_25[9:0]) begin
        image_0_455 <= io_pixelVal_in_0_3;
      end else if (10'h1c7 == _T_22[9:0]) begin
        image_0_455 <= io_pixelVal_in_0_2;
      end else if (10'h1c7 == _T_19[9:0]) begin
        image_0_455 <= io_pixelVal_in_0_1;
      end else if (10'h1c7 == _T_15[9:0]) begin
        image_0_455 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_456 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1c8 == _T_37[9:0]) begin
        image_0_456 <= io_pixelVal_in_0_7;
      end else if (10'h1c8 == _T_34[9:0]) begin
        image_0_456 <= io_pixelVal_in_0_6;
      end else if (10'h1c8 == _T_31[9:0]) begin
        image_0_456 <= io_pixelVal_in_0_5;
      end else if (10'h1c8 == _T_28[9:0]) begin
        image_0_456 <= io_pixelVal_in_0_4;
      end else if (10'h1c8 == _T_25[9:0]) begin
        image_0_456 <= io_pixelVal_in_0_3;
      end else if (10'h1c8 == _T_22[9:0]) begin
        image_0_456 <= io_pixelVal_in_0_2;
      end else if (10'h1c8 == _T_19[9:0]) begin
        image_0_456 <= io_pixelVal_in_0_1;
      end else if (10'h1c8 == _T_15[9:0]) begin
        image_0_456 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_457 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1c9 == _T_37[9:0]) begin
        image_0_457 <= io_pixelVal_in_0_7;
      end else if (10'h1c9 == _T_34[9:0]) begin
        image_0_457 <= io_pixelVal_in_0_6;
      end else if (10'h1c9 == _T_31[9:0]) begin
        image_0_457 <= io_pixelVal_in_0_5;
      end else if (10'h1c9 == _T_28[9:0]) begin
        image_0_457 <= io_pixelVal_in_0_4;
      end else if (10'h1c9 == _T_25[9:0]) begin
        image_0_457 <= io_pixelVal_in_0_3;
      end else if (10'h1c9 == _T_22[9:0]) begin
        image_0_457 <= io_pixelVal_in_0_2;
      end else if (10'h1c9 == _T_19[9:0]) begin
        image_0_457 <= io_pixelVal_in_0_1;
      end else if (10'h1c9 == _T_15[9:0]) begin
        image_0_457 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_458 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1ca == _T_37[9:0]) begin
        image_0_458 <= io_pixelVal_in_0_7;
      end else if (10'h1ca == _T_34[9:0]) begin
        image_0_458 <= io_pixelVal_in_0_6;
      end else if (10'h1ca == _T_31[9:0]) begin
        image_0_458 <= io_pixelVal_in_0_5;
      end else if (10'h1ca == _T_28[9:0]) begin
        image_0_458 <= io_pixelVal_in_0_4;
      end else if (10'h1ca == _T_25[9:0]) begin
        image_0_458 <= io_pixelVal_in_0_3;
      end else if (10'h1ca == _T_22[9:0]) begin
        image_0_458 <= io_pixelVal_in_0_2;
      end else if (10'h1ca == _T_19[9:0]) begin
        image_0_458 <= io_pixelVal_in_0_1;
      end else if (10'h1ca == _T_15[9:0]) begin
        image_0_458 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_459 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1cb == _T_37[9:0]) begin
        image_0_459 <= io_pixelVal_in_0_7;
      end else if (10'h1cb == _T_34[9:0]) begin
        image_0_459 <= io_pixelVal_in_0_6;
      end else if (10'h1cb == _T_31[9:0]) begin
        image_0_459 <= io_pixelVal_in_0_5;
      end else if (10'h1cb == _T_28[9:0]) begin
        image_0_459 <= io_pixelVal_in_0_4;
      end else if (10'h1cb == _T_25[9:0]) begin
        image_0_459 <= io_pixelVal_in_0_3;
      end else if (10'h1cb == _T_22[9:0]) begin
        image_0_459 <= io_pixelVal_in_0_2;
      end else if (10'h1cb == _T_19[9:0]) begin
        image_0_459 <= io_pixelVal_in_0_1;
      end else if (10'h1cb == _T_15[9:0]) begin
        image_0_459 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_460 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1cc == _T_37[9:0]) begin
        image_0_460 <= io_pixelVal_in_0_7;
      end else if (10'h1cc == _T_34[9:0]) begin
        image_0_460 <= io_pixelVal_in_0_6;
      end else if (10'h1cc == _T_31[9:0]) begin
        image_0_460 <= io_pixelVal_in_0_5;
      end else if (10'h1cc == _T_28[9:0]) begin
        image_0_460 <= io_pixelVal_in_0_4;
      end else if (10'h1cc == _T_25[9:0]) begin
        image_0_460 <= io_pixelVal_in_0_3;
      end else if (10'h1cc == _T_22[9:0]) begin
        image_0_460 <= io_pixelVal_in_0_2;
      end else if (10'h1cc == _T_19[9:0]) begin
        image_0_460 <= io_pixelVal_in_0_1;
      end else if (10'h1cc == _T_15[9:0]) begin
        image_0_460 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_461 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1cd == _T_37[9:0]) begin
        image_0_461 <= io_pixelVal_in_0_7;
      end else if (10'h1cd == _T_34[9:0]) begin
        image_0_461 <= io_pixelVal_in_0_6;
      end else if (10'h1cd == _T_31[9:0]) begin
        image_0_461 <= io_pixelVal_in_0_5;
      end else if (10'h1cd == _T_28[9:0]) begin
        image_0_461 <= io_pixelVal_in_0_4;
      end else if (10'h1cd == _T_25[9:0]) begin
        image_0_461 <= io_pixelVal_in_0_3;
      end else if (10'h1cd == _T_22[9:0]) begin
        image_0_461 <= io_pixelVal_in_0_2;
      end else if (10'h1cd == _T_19[9:0]) begin
        image_0_461 <= io_pixelVal_in_0_1;
      end else if (10'h1cd == _T_15[9:0]) begin
        image_0_461 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_462 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1ce == _T_37[9:0]) begin
        image_0_462 <= io_pixelVal_in_0_7;
      end else if (10'h1ce == _T_34[9:0]) begin
        image_0_462 <= io_pixelVal_in_0_6;
      end else if (10'h1ce == _T_31[9:0]) begin
        image_0_462 <= io_pixelVal_in_0_5;
      end else if (10'h1ce == _T_28[9:0]) begin
        image_0_462 <= io_pixelVal_in_0_4;
      end else if (10'h1ce == _T_25[9:0]) begin
        image_0_462 <= io_pixelVal_in_0_3;
      end else if (10'h1ce == _T_22[9:0]) begin
        image_0_462 <= io_pixelVal_in_0_2;
      end else if (10'h1ce == _T_19[9:0]) begin
        image_0_462 <= io_pixelVal_in_0_1;
      end else if (10'h1ce == _T_15[9:0]) begin
        image_0_462 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_463 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1cf == _T_37[9:0]) begin
        image_0_463 <= io_pixelVal_in_0_7;
      end else if (10'h1cf == _T_34[9:0]) begin
        image_0_463 <= io_pixelVal_in_0_6;
      end else if (10'h1cf == _T_31[9:0]) begin
        image_0_463 <= io_pixelVal_in_0_5;
      end else if (10'h1cf == _T_28[9:0]) begin
        image_0_463 <= io_pixelVal_in_0_4;
      end else if (10'h1cf == _T_25[9:0]) begin
        image_0_463 <= io_pixelVal_in_0_3;
      end else if (10'h1cf == _T_22[9:0]) begin
        image_0_463 <= io_pixelVal_in_0_2;
      end else if (10'h1cf == _T_19[9:0]) begin
        image_0_463 <= io_pixelVal_in_0_1;
      end else if (10'h1cf == _T_15[9:0]) begin
        image_0_463 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_464 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1d0 == _T_37[9:0]) begin
        image_0_464 <= io_pixelVal_in_0_7;
      end else if (10'h1d0 == _T_34[9:0]) begin
        image_0_464 <= io_pixelVal_in_0_6;
      end else if (10'h1d0 == _T_31[9:0]) begin
        image_0_464 <= io_pixelVal_in_0_5;
      end else if (10'h1d0 == _T_28[9:0]) begin
        image_0_464 <= io_pixelVal_in_0_4;
      end else if (10'h1d0 == _T_25[9:0]) begin
        image_0_464 <= io_pixelVal_in_0_3;
      end else if (10'h1d0 == _T_22[9:0]) begin
        image_0_464 <= io_pixelVal_in_0_2;
      end else if (10'h1d0 == _T_19[9:0]) begin
        image_0_464 <= io_pixelVal_in_0_1;
      end else if (10'h1d0 == _T_15[9:0]) begin
        image_0_464 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_465 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1d1 == _T_37[9:0]) begin
        image_0_465 <= io_pixelVal_in_0_7;
      end else if (10'h1d1 == _T_34[9:0]) begin
        image_0_465 <= io_pixelVal_in_0_6;
      end else if (10'h1d1 == _T_31[9:0]) begin
        image_0_465 <= io_pixelVal_in_0_5;
      end else if (10'h1d1 == _T_28[9:0]) begin
        image_0_465 <= io_pixelVal_in_0_4;
      end else if (10'h1d1 == _T_25[9:0]) begin
        image_0_465 <= io_pixelVal_in_0_3;
      end else if (10'h1d1 == _T_22[9:0]) begin
        image_0_465 <= io_pixelVal_in_0_2;
      end else if (10'h1d1 == _T_19[9:0]) begin
        image_0_465 <= io_pixelVal_in_0_1;
      end else if (10'h1d1 == _T_15[9:0]) begin
        image_0_465 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_466 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1d2 == _T_37[9:0]) begin
        image_0_466 <= io_pixelVal_in_0_7;
      end else if (10'h1d2 == _T_34[9:0]) begin
        image_0_466 <= io_pixelVal_in_0_6;
      end else if (10'h1d2 == _T_31[9:0]) begin
        image_0_466 <= io_pixelVal_in_0_5;
      end else if (10'h1d2 == _T_28[9:0]) begin
        image_0_466 <= io_pixelVal_in_0_4;
      end else if (10'h1d2 == _T_25[9:0]) begin
        image_0_466 <= io_pixelVal_in_0_3;
      end else if (10'h1d2 == _T_22[9:0]) begin
        image_0_466 <= io_pixelVal_in_0_2;
      end else if (10'h1d2 == _T_19[9:0]) begin
        image_0_466 <= io_pixelVal_in_0_1;
      end else if (10'h1d2 == _T_15[9:0]) begin
        image_0_466 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_467 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1d3 == _T_37[9:0]) begin
        image_0_467 <= io_pixelVal_in_0_7;
      end else if (10'h1d3 == _T_34[9:0]) begin
        image_0_467 <= io_pixelVal_in_0_6;
      end else if (10'h1d3 == _T_31[9:0]) begin
        image_0_467 <= io_pixelVal_in_0_5;
      end else if (10'h1d3 == _T_28[9:0]) begin
        image_0_467 <= io_pixelVal_in_0_4;
      end else if (10'h1d3 == _T_25[9:0]) begin
        image_0_467 <= io_pixelVal_in_0_3;
      end else if (10'h1d3 == _T_22[9:0]) begin
        image_0_467 <= io_pixelVal_in_0_2;
      end else if (10'h1d3 == _T_19[9:0]) begin
        image_0_467 <= io_pixelVal_in_0_1;
      end else if (10'h1d3 == _T_15[9:0]) begin
        image_0_467 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_468 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1d4 == _T_37[9:0]) begin
        image_0_468 <= io_pixelVal_in_0_7;
      end else if (10'h1d4 == _T_34[9:0]) begin
        image_0_468 <= io_pixelVal_in_0_6;
      end else if (10'h1d4 == _T_31[9:0]) begin
        image_0_468 <= io_pixelVal_in_0_5;
      end else if (10'h1d4 == _T_28[9:0]) begin
        image_0_468 <= io_pixelVal_in_0_4;
      end else if (10'h1d4 == _T_25[9:0]) begin
        image_0_468 <= io_pixelVal_in_0_3;
      end else if (10'h1d4 == _T_22[9:0]) begin
        image_0_468 <= io_pixelVal_in_0_2;
      end else if (10'h1d4 == _T_19[9:0]) begin
        image_0_468 <= io_pixelVal_in_0_1;
      end else if (10'h1d4 == _T_15[9:0]) begin
        image_0_468 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_469 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1d5 == _T_37[9:0]) begin
        image_0_469 <= io_pixelVal_in_0_7;
      end else if (10'h1d5 == _T_34[9:0]) begin
        image_0_469 <= io_pixelVal_in_0_6;
      end else if (10'h1d5 == _T_31[9:0]) begin
        image_0_469 <= io_pixelVal_in_0_5;
      end else if (10'h1d5 == _T_28[9:0]) begin
        image_0_469 <= io_pixelVal_in_0_4;
      end else if (10'h1d5 == _T_25[9:0]) begin
        image_0_469 <= io_pixelVal_in_0_3;
      end else if (10'h1d5 == _T_22[9:0]) begin
        image_0_469 <= io_pixelVal_in_0_2;
      end else if (10'h1d5 == _T_19[9:0]) begin
        image_0_469 <= io_pixelVal_in_0_1;
      end else if (10'h1d5 == _T_15[9:0]) begin
        image_0_469 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_470 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1d6 == _T_37[9:0]) begin
        image_0_470 <= io_pixelVal_in_0_7;
      end else if (10'h1d6 == _T_34[9:0]) begin
        image_0_470 <= io_pixelVal_in_0_6;
      end else if (10'h1d6 == _T_31[9:0]) begin
        image_0_470 <= io_pixelVal_in_0_5;
      end else if (10'h1d6 == _T_28[9:0]) begin
        image_0_470 <= io_pixelVal_in_0_4;
      end else if (10'h1d6 == _T_25[9:0]) begin
        image_0_470 <= io_pixelVal_in_0_3;
      end else if (10'h1d6 == _T_22[9:0]) begin
        image_0_470 <= io_pixelVal_in_0_2;
      end else if (10'h1d6 == _T_19[9:0]) begin
        image_0_470 <= io_pixelVal_in_0_1;
      end else if (10'h1d6 == _T_15[9:0]) begin
        image_0_470 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_471 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1d7 == _T_37[9:0]) begin
        image_0_471 <= io_pixelVal_in_0_7;
      end else if (10'h1d7 == _T_34[9:0]) begin
        image_0_471 <= io_pixelVal_in_0_6;
      end else if (10'h1d7 == _T_31[9:0]) begin
        image_0_471 <= io_pixelVal_in_0_5;
      end else if (10'h1d7 == _T_28[9:0]) begin
        image_0_471 <= io_pixelVal_in_0_4;
      end else if (10'h1d7 == _T_25[9:0]) begin
        image_0_471 <= io_pixelVal_in_0_3;
      end else if (10'h1d7 == _T_22[9:0]) begin
        image_0_471 <= io_pixelVal_in_0_2;
      end else if (10'h1d7 == _T_19[9:0]) begin
        image_0_471 <= io_pixelVal_in_0_1;
      end else if (10'h1d7 == _T_15[9:0]) begin
        image_0_471 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_472 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1d8 == _T_37[9:0]) begin
        image_0_472 <= io_pixelVal_in_0_7;
      end else if (10'h1d8 == _T_34[9:0]) begin
        image_0_472 <= io_pixelVal_in_0_6;
      end else if (10'h1d8 == _T_31[9:0]) begin
        image_0_472 <= io_pixelVal_in_0_5;
      end else if (10'h1d8 == _T_28[9:0]) begin
        image_0_472 <= io_pixelVal_in_0_4;
      end else if (10'h1d8 == _T_25[9:0]) begin
        image_0_472 <= io_pixelVal_in_0_3;
      end else if (10'h1d8 == _T_22[9:0]) begin
        image_0_472 <= io_pixelVal_in_0_2;
      end else if (10'h1d8 == _T_19[9:0]) begin
        image_0_472 <= io_pixelVal_in_0_1;
      end else if (10'h1d8 == _T_15[9:0]) begin
        image_0_472 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_473 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1d9 == _T_37[9:0]) begin
        image_0_473 <= io_pixelVal_in_0_7;
      end else if (10'h1d9 == _T_34[9:0]) begin
        image_0_473 <= io_pixelVal_in_0_6;
      end else if (10'h1d9 == _T_31[9:0]) begin
        image_0_473 <= io_pixelVal_in_0_5;
      end else if (10'h1d9 == _T_28[9:0]) begin
        image_0_473 <= io_pixelVal_in_0_4;
      end else if (10'h1d9 == _T_25[9:0]) begin
        image_0_473 <= io_pixelVal_in_0_3;
      end else if (10'h1d9 == _T_22[9:0]) begin
        image_0_473 <= io_pixelVal_in_0_2;
      end else if (10'h1d9 == _T_19[9:0]) begin
        image_0_473 <= io_pixelVal_in_0_1;
      end else if (10'h1d9 == _T_15[9:0]) begin
        image_0_473 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_474 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1da == _T_37[9:0]) begin
        image_0_474 <= io_pixelVal_in_0_7;
      end else if (10'h1da == _T_34[9:0]) begin
        image_0_474 <= io_pixelVal_in_0_6;
      end else if (10'h1da == _T_31[9:0]) begin
        image_0_474 <= io_pixelVal_in_0_5;
      end else if (10'h1da == _T_28[9:0]) begin
        image_0_474 <= io_pixelVal_in_0_4;
      end else if (10'h1da == _T_25[9:0]) begin
        image_0_474 <= io_pixelVal_in_0_3;
      end else if (10'h1da == _T_22[9:0]) begin
        image_0_474 <= io_pixelVal_in_0_2;
      end else if (10'h1da == _T_19[9:0]) begin
        image_0_474 <= io_pixelVal_in_0_1;
      end else if (10'h1da == _T_15[9:0]) begin
        image_0_474 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_475 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1db == _T_37[9:0]) begin
        image_0_475 <= io_pixelVal_in_0_7;
      end else if (10'h1db == _T_34[9:0]) begin
        image_0_475 <= io_pixelVal_in_0_6;
      end else if (10'h1db == _T_31[9:0]) begin
        image_0_475 <= io_pixelVal_in_0_5;
      end else if (10'h1db == _T_28[9:0]) begin
        image_0_475 <= io_pixelVal_in_0_4;
      end else if (10'h1db == _T_25[9:0]) begin
        image_0_475 <= io_pixelVal_in_0_3;
      end else if (10'h1db == _T_22[9:0]) begin
        image_0_475 <= io_pixelVal_in_0_2;
      end else if (10'h1db == _T_19[9:0]) begin
        image_0_475 <= io_pixelVal_in_0_1;
      end else if (10'h1db == _T_15[9:0]) begin
        image_0_475 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_476 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1dc == _T_37[9:0]) begin
        image_0_476 <= io_pixelVal_in_0_7;
      end else if (10'h1dc == _T_34[9:0]) begin
        image_0_476 <= io_pixelVal_in_0_6;
      end else if (10'h1dc == _T_31[9:0]) begin
        image_0_476 <= io_pixelVal_in_0_5;
      end else if (10'h1dc == _T_28[9:0]) begin
        image_0_476 <= io_pixelVal_in_0_4;
      end else if (10'h1dc == _T_25[9:0]) begin
        image_0_476 <= io_pixelVal_in_0_3;
      end else if (10'h1dc == _T_22[9:0]) begin
        image_0_476 <= io_pixelVal_in_0_2;
      end else if (10'h1dc == _T_19[9:0]) begin
        image_0_476 <= io_pixelVal_in_0_1;
      end else if (10'h1dc == _T_15[9:0]) begin
        image_0_476 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_477 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1dd == _T_37[9:0]) begin
        image_0_477 <= io_pixelVal_in_0_7;
      end else if (10'h1dd == _T_34[9:0]) begin
        image_0_477 <= io_pixelVal_in_0_6;
      end else if (10'h1dd == _T_31[9:0]) begin
        image_0_477 <= io_pixelVal_in_0_5;
      end else if (10'h1dd == _T_28[9:0]) begin
        image_0_477 <= io_pixelVal_in_0_4;
      end else if (10'h1dd == _T_25[9:0]) begin
        image_0_477 <= io_pixelVal_in_0_3;
      end else if (10'h1dd == _T_22[9:0]) begin
        image_0_477 <= io_pixelVal_in_0_2;
      end else if (10'h1dd == _T_19[9:0]) begin
        image_0_477 <= io_pixelVal_in_0_1;
      end else if (10'h1dd == _T_15[9:0]) begin
        image_0_477 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_478 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1de == _T_37[9:0]) begin
        image_0_478 <= io_pixelVal_in_0_7;
      end else if (10'h1de == _T_34[9:0]) begin
        image_0_478 <= io_pixelVal_in_0_6;
      end else if (10'h1de == _T_31[9:0]) begin
        image_0_478 <= io_pixelVal_in_0_5;
      end else if (10'h1de == _T_28[9:0]) begin
        image_0_478 <= io_pixelVal_in_0_4;
      end else if (10'h1de == _T_25[9:0]) begin
        image_0_478 <= io_pixelVal_in_0_3;
      end else if (10'h1de == _T_22[9:0]) begin
        image_0_478 <= io_pixelVal_in_0_2;
      end else if (10'h1de == _T_19[9:0]) begin
        image_0_478 <= io_pixelVal_in_0_1;
      end else if (10'h1de == _T_15[9:0]) begin
        image_0_478 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_479 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1df == _T_37[9:0]) begin
        image_0_479 <= io_pixelVal_in_0_7;
      end else if (10'h1df == _T_34[9:0]) begin
        image_0_479 <= io_pixelVal_in_0_6;
      end else if (10'h1df == _T_31[9:0]) begin
        image_0_479 <= io_pixelVal_in_0_5;
      end else if (10'h1df == _T_28[9:0]) begin
        image_0_479 <= io_pixelVal_in_0_4;
      end else if (10'h1df == _T_25[9:0]) begin
        image_0_479 <= io_pixelVal_in_0_3;
      end else if (10'h1df == _T_22[9:0]) begin
        image_0_479 <= io_pixelVal_in_0_2;
      end else if (10'h1df == _T_19[9:0]) begin
        image_0_479 <= io_pixelVal_in_0_1;
      end else if (10'h1df == _T_15[9:0]) begin
        image_0_479 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_480 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1e0 == _T_37[9:0]) begin
        image_0_480 <= io_pixelVal_in_0_7;
      end else if (10'h1e0 == _T_34[9:0]) begin
        image_0_480 <= io_pixelVal_in_0_6;
      end else if (10'h1e0 == _T_31[9:0]) begin
        image_0_480 <= io_pixelVal_in_0_5;
      end else if (10'h1e0 == _T_28[9:0]) begin
        image_0_480 <= io_pixelVal_in_0_4;
      end else if (10'h1e0 == _T_25[9:0]) begin
        image_0_480 <= io_pixelVal_in_0_3;
      end else if (10'h1e0 == _T_22[9:0]) begin
        image_0_480 <= io_pixelVal_in_0_2;
      end else if (10'h1e0 == _T_19[9:0]) begin
        image_0_480 <= io_pixelVal_in_0_1;
      end else if (10'h1e0 == _T_15[9:0]) begin
        image_0_480 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_481 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1e1 == _T_37[9:0]) begin
        image_0_481 <= io_pixelVal_in_0_7;
      end else if (10'h1e1 == _T_34[9:0]) begin
        image_0_481 <= io_pixelVal_in_0_6;
      end else if (10'h1e1 == _T_31[9:0]) begin
        image_0_481 <= io_pixelVal_in_0_5;
      end else if (10'h1e1 == _T_28[9:0]) begin
        image_0_481 <= io_pixelVal_in_0_4;
      end else if (10'h1e1 == _T_25[9:0]) begin
        image_0_481 <= io_pixelVal_in_0_3;
      end else if (10'h1e1 == _T_22[9:0]) begin
        image_0_481 <= io_pixelVal_in_0_2;
      end else if (10'h1e1 == _T_19[9:0]) begin
        image_0_481 <= io_pixelVal_in_0_1;
      end else if (10'h1e1 == _T_15[9:0]) begin
        image_0_481 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_482 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1e2 == _T_37[9:0]) begin
        image_0_482 <= io_pixelVal_in_0_7;
      end else if (10'h1e2 == _T_34[9:0]) begin
        image_0_482 <= io_pixelVal_in_0_6;
      end else if (10'h1e2 == _T_31[9:0]) begin
        image_0_482 <= io_pixelVal_in_0_5;
      end else if (10'h1e2 == _T_28[9:0]) begin
        image_0_482 <= io_pixelVal_in_0_4;
      end else if (10'h1e2 == _T_25[9:0]) begin
        image_0_482 <= io_pixelVal_in_0_3;
      end else if (10'h1e2 == _T_22[9:0]) begin
        image_0_482 <= io_pixelVal_in_0_2;
      end else if (10'h1e2 == _T_19[9:0]) begin
        image_0_482 <= io_pixelVal_in_0_1;
      end else if (10'h1e2 == _T_15[9:0]) begin
        image_0_482 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_483 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1e3 == _T_37[9:0]) begin
        image_0_483 <= io_pixelVal_in_0_7;
      end else if (10'h1e3 == _T_34[9:0]) begin
        image_0_483 <= io_pixelVal_in_0_6;
      end else if (10'h1e3 == _T_31[9:0]) begin
        image_0_483 <= io_pixelVal_in_0_5;
      end else if (10'h1e3 == _T_28[9:0]) begin
        image_0_483 <= io_pixelVal_in_0_4;
      end else if (10'h1e3 == _T_25[9:0]) begin
        image_0_483 <= io_pixelVal_in_0_3;
      end else if (10'h1e3 == _T_22[9:0]) begin
        image_0_483 <= io_pixelVal_in_0_2;
      end else if (10'h1e3 == _T_19[9:0]) begin
        image_0_483 <= io_pixelVal_in_0_1;
      end else if (10'h1e3 == _T_15[9:0]) begin
        image_0_483 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_484 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1e4 == _T_37[9:0]) begin
        image_0_484 <= io_pixelVal_in_0_7;
      end else if (10'h1e4 == _T_34[9:0]) begin
        image_0_484 <= io_pixelVal_in_0_6;
      end else if (10'h1e4 == _T_31[9:0]) begin
        image_0_484 <= io_pixelVal_in_0_5;
      end else if (10'h1e4 == _T_28[9:0]) begin
        image_0_484 <= io_pixelVal_in_0_4;
      end else if (10'h1e4 == _T_25[9:0]) begin
        image_0_484 <= io_pixelVal_in_0_3;
      end else if (10'h1e4 == _T_22[9:0]) begin
        image_0_484 <= io_pixelVal_in_0_2;
      end else if (10'h1e4 == _T_19[9:0]) begin
        image_0_484 <= io_pixelVal_in_0_1;
      end else if (10'h1e4 == _T_15[9:0]) begin
        image_0_484 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_485 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1e5 == _T_37[9:0]) begin
        image_0_485 <= io_pixelVal_in_0_7;
      end else if (10'h1e5 == _T_34[9:0]) begin
        image_0_485 <= io_pixelVal_in_0_6;
      end else if (10'h1e5 == _T_31[9:0]) begin
        image_0_485 <= io_pixelVal_in_0_5;
      end else if (10'h1e5 == _T_28[9:0]) begin
        image_0_485 <= io_pixelVal_in_0_4;
      end else if (10'h1e5 == _T_25[9:0]) begin
        image_0_485 <= io_pixelVal_in_0_3;
      end else if (10'h1e5 == _T_22[9:0]) begin
        image_0_485 <= io_pixelVal_in_0_2;
      end else if (10'h1e5 == _T_19[9:0]) begin
        image_0_485 <= io_pixelVal_in_0_1;
      end else if (10'h1e5 == _T_15[9:0]) begin
        image_0_485 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_486 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1e6 == _T_37[9:0]) begin
        image_0_486 <= io_pixelVal_in_0_7;
      end else if (10'h1e6 == _T_34[9:0]) begin
        image_0_486 <= io_pixelVal_in_0_6;
      end else if (10'h1e6 == _T_31[9:0]) begin
        image_0_486 <= io_pixelVal_in_0_5;
      end else if (10'h1e6 == _T_28[9:0]) begin
        image_0_486 <= io_pixelVal_in_0_4;
      end else if (10'h1e6 == _T_25[9:0]) begin
        image_0_486 <= io_pixelVal_in_0_3;
      end else if (10'h1e6 == _T_22[9:0]) begin
        image_0_486 <= io_pixelVal_in_0_2;
      end else if (10'h1e6 == _T_19[9:0]) begin
        image_0_486 <= io_pixelVal_in_0_1;
      end else if (10'h1e6 == _T_15[9:0]) begin
        image_0_486 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_487 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1e7 == _T_37[9:0]) begin
        image_0_487 <= io_pixelVal_in_0_7;
      end else if (10'h1e7 == _T_34[9:0]) begin
        image_0_487 <= io_pixelVal_in_0_6;
      end else if (10'h1e7 == _T_31[9:0]) begin
        image_0_487 <= io_pixelVal_in_0_5;
      end else if (10'h1e7 == _T_28[9:0]) begin
        image_0_487 <= io_pixelVal_in_0_4;
      end else if (10'h1e7 == _T_25[9:0]) begin
        image_0_487 <= io_pixelVal_in_0_3;
      end else if (10'h1e7 == _T_22[9:0]) begin
        image_0_487 <= io_pixelVal_in_0_2;
      end else if (10'h1e7 == _T_19[9:0]) begin
        image_0_487 <= io_pixelVal_in_0_1;
      end else if (10'h1e7 == _T_15[9:0]) begin
        image_0_487 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_488 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1e8 == _T_37[9:0]) begin
        image_0_488 <= io_pixelVal_in_0_7;
      end else if (10'h1e8 == _T_34[9:0]) begin
        image_0_488 <= io_pixelVal_in_0_6;
      end else if (10'h1e8 == _T_31[9:0]) begin
        image_0_488 <= io_pixelVal_in_0_5;
      end else if (10'h1e8 == _T_28[9:0]) begin
        image_0_488 <= io_pixelVal_in_0_4;
      end else if (10'h1e8 == _T_25[9:0]) begin
        image_0_488 <= io_pixelVal_in_0_3;
      end else if (10'h1e8 == _T_22[9:0]) begin
        image_0_488 <= io_pixelVal_in_0_2;
      end else if (10'h1e8 == _T_19[9:0]) begin
        image_0_488 <= io_pixelVal_in_0_1;
      end else if (10'h1e8 == _T_15[9:0]) begin
        image_0_488 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_489 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1e9 == _T_37[9:0]) begin
        image_0_489 <= io_pixelVal_in_0_7;
      end else if (10'h1e9 == _T_34[9:0]) begin
        image_0_489 <= io_pixelVal_in_0_6;
      end else if (10'h1e9 == _T_31[9:0]) begin
        image_0_489 <= io_pixelVal_in_0_5;
      end else if (10'h1e9 == _T_28[9:0]) begin
        image_0_489 <= io_pixelVal_in_0_4;
      end else if (10'h1e9 == _T_25[9:0]) begin
        image_0_489 <= io_pixelVal_in_0_3;
      end else if (10'h1e9 == _T_22[9:0]) begin
        image_0_489 <= io_pixelVal_in_0_2;
      end else if (10'h1e9 == _T_19[9:0]) begin
        image_0_489 <= io_pixelVal_in_0_1;
      end else if (10'h1e9 == _T_15[9:0]) begin
        image_0_489 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_490 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1ea == _T_37[9:0]) begin
        image_0_490 <= io_pixelVal_in_0_7;
      end else if (10'h1ea == _T_34[9:0]) begin
        image_0_490 <= io_pixelVal_in_0_6;
      end else if (10'h1ea == _T_31[9:0]) begin
        image_0_490 <= io_pixelVal_in_0_5;
      end else if (10'h1ea == _T_28[9:0]) begin
        image_0_490 <= io_pixelVal_in_0_4;
      end else if (10'h1ea == _T_25[9:0]) begin
        image_0_490 <= io_pixelVal_in_0_3;
      end else if (10'h1ea == _T_22[9:0]) begin
        image_0_490 <= io_pixelVal_in_0_2;
      end else if (10'h1ea == _T_19[9:0]) begin
        image_0_490 <= io_pixelVal_in_0_1;
      end else if (10'h1ea == _T_15[9:0]) begin
        image_0_490 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_491 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1eb == _T_37[9:0]) begin
        image_0_491 <= io_pixelVal_in_0_7;
      end else if (10'h1eb == _T_34[9:0]) begin
        image_0_491 <= io_pixelVal_in_0_6;
      end else if (10'h1eb == _T_31[9:0]) begin
        image_0_491 <= io_pixelVal_in_0_5;
      end else if (10'h1eb == _T_28[9:0]) begin
        image_0_491 <= io_pixelVal_in_0_4;
      end else if (10'h1eb == _T_25[9:0]) begin
        image_0_491 <= io_pixelVal_in_0_3;
      end else if (10'h1eb == _T_22[9:0]) begin
        image_0_491 <= io_pixelVal_in_0_2;
      end else if (10'h1eb == _T_19[9:0]) begin
        image_0_491 <= io_pixelVal_in_0_1;
      end else if (10'h1eb == _T_15[9:0]) begin
        image_0_491 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_492 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1ec == _T_37[9:0]) begin
        image_0_492 <= io_pixelVal_in_0_7;
      end else if (10'h1ec == _T_34[9:0]) begin
        image_0_492 <= io_pixelVal_in_0_6;
      end else if (10'h1ec == _T_31[9:0]) begin
        image_0_492 <= io_pixelVal_in_0_5;
      end else if (10'h1ec == _T_28[9:0]) begin
        image_0_492 <= io_pixelVal_in_0_4;
      end else if (10'h1ec == _T_25[9:0]) begin
        image_0_492 <= io_pixelVal_in_0_3;
      end else if (10'h1ec == _T_22[9:0]) begin
        image_0_492 <= io_pixelVal_in_0_2;
      end else if (10'h1ec == _T_19[9:0]) begin
        image_0_492 <= io_pixelVal_in_0_1;
      end else if (10'h1ec == _T_15[9:0]) begin
        image_0_492 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_493 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1ed == _T_37[9:0]) begin
        image_0_493 <= io_pixelVal_in_0_7;
      end else if (10'h1ed == _T_34[9:0]) begin
        image_0_493 <= io_pixelVal_in_0_6;
      end else if (10'h1ed == _T_31[9:0]) begin
        image_0_493 <= io_pixelVal_in_0_5;
      end else if (10'h1ed == _T_28[9:0]) begin
        image_0_493 <= io_pixelVal_in_0_4;
      end else if (10'h1ed == _T_25[9:0]) begin
        image_0_493 <= io_pixelVal_in_0_3;
      end else if (10'h1ed == _T_22[9:0]) begin
        image_0_493 <= io_pixelVal_in_0_2;
      end else if (10'h1ed == _T_19[9:0]) begin
        image_0_493 <= io_pixelVal_in_0_1;
      end else if (10'h1ed == _T_15[9:0]) begin
        image_0_493 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_494 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1ee == _T_37[9:0]) begin
        image_0_494 <= io_pixelVal_in_0_7;
      end else if (10'h1ee == _T_34[9:0]) begin
        image_0_494 <= io_pixelVal_in_0_6;
      end else if (10'h1ee == _T_31[9:0]) begin
        image_0_494 <= io_pixelVal_in_0_5;
      end else if (10'h1ee == _T_28[9:0]) begin
        image_0_494 <= io_pixelVal_in_0_4;
      end else if (10'h1ee == _T_25[9:0]) begin
        image_0_494 <= io_pixelVal_in_0_3;
      end else if (10'h1ee == _T_22[9:0]) begin
        image_0_494 <= io_pixelVal_in_0_2;
      end else if (10'h1ee == _T_19[9:0]) begin
        image_0_494 <= io_pixelVal_in_0_1;
      end else if (10'h1ee == _T_15[9:0]) begin
        image_0_494 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_495 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1ef == _T_37[9:0]) begin
        image_0_495 <= io_pixelVal_in_0_7;
      end else if (10'h1ef == _T_34[9:0]) begin
        image_0_495 <= io_pixelVal_in_0_6;
      end else if (10'h1ef == _T_31[9:0]) begin
        image_0_495 <= io_pixelVal_in_0_5;
      end else if (10'h1ef == _T_28[9:0]) begin
        image_0_495 <= io_pixelVal_in_0_4;
      end else if (10'h1ef == _T_25[9:0]) begin
        image_0_495 <= io_pixelVal_in_0_3;
      end else if (10'h1ef == _T_22[9:0]) begin
        image_0_495 <= io_pixelVal_in_0_2;
      end else if (10'h1ef == _T_19[9:0]) begin
        image_0_495 <= io_pixelVal_in_0_1;
      end else if (10'h1ef == _T_15[9:0]) begin
        image_0_495 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_496 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1f0 == _T_37[9:0]) begin
        image_0_496 <= io_pixelVal_in_0_7;
      end else if (10'h1f0 == _T_34[9:0]) begin
        image_0_496 <= io_pixelVal_in_0_6;
      end else if (10'h1f0 == _T_31[9:0]) begin
        image_0_496 <= io_pixelVal_in_0_5;
      end else if (10'h1f0 == _T_28[9:0]) begin
        image_0_496 <= io_pixelVal_in_0_4;
      end else if (10'h1f0 == _T_25[9:0]) begin
        image_0_496 <= io_pixelVal_in_0_3;
      end else if (10'h1f0 == _T_22[9:0]) begin
        image_0_496 <= io_pixelVal_in_0_2;
      end else if (10'h1f0 == _T_19[9:0]) begin
        image_0_496 <= io_pixelVal_in_0_1;
      end else if (10'h1f0 == _T_15[9:0]) begin
        image_0_496 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_497 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1f1 == _T_37[9:0]) begin
        image_0_497 <= io_pixelVal_in_0_7;
      end else if (10'h1f1 == _T_34[9:0]) begin
        image_0_497 <= io_pixelVal_in_0_6;
      end else if (10'h1f1 == _T_31[9:0]) begin
        image_0_497 <= io_pixelVal_in_0_5;
      end else if (10'h1f1 == _T_28[9:0]) begin
        image_0_497 <= io_pixelVal_in_0_4;
      end else if (10'h1f1 == _T_25[9:0]) begin
        image_0_497 <= io_pixelVal_in_0_3;
      end else if (10'h1f1 == _T_22[9:0]) begin
        image_0_497 <= io_pixelVal_in_0_2;
      end else if (10'h1f1 == _T_19[9:0]) begin
        image_0_497 <= io_pixelVal_in_0_1;
      end else if (10'h1f1 == _T_15[9:0]) begin
        image_0_497 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_498 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1f2 == _T_37[9:0]) begin
        image_0_498 <= io_pixelVal_in_0_7;
      end else if (10'h1f2 == _T_34[9:0]) begin
        image_0_498 <= io_pixelVal_in_0_6;
      end else if (10'h1f2 == _T_31[9:0]) begin
        image_0_498 <= io_pixelVal_in_0_5;
      end else if (10'h1f2 == _T_28[9:0]) begin
        image_0_498 <= io_pixelVal_in_0_4;
      end else if (10'h1f2 == _T_25[9:0]) begin
        image_0_498 <= io_pixelVal_in_0_3;
      end else if (10'h1f2 == _T_22[9:0]) begin
        image_0_498 <= io_pixelVal_in_0_2;
      end else if (10'h1f2 == _T_19[9:0]) begin
        image_0_498 <= io_pixelVal_in_0_1;
      end else if (10'h1f2 == _T_15[9:0]) begin
        image_0_498 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_499 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1f3 == _T_37[9:0]) begin
        image_0_499 <= io_pixelVal_in_0_7;
      end else if (10'h1f3 == _T_34[9:0]) begin
        image_0_499 <= io_pixelVal_in_0_6;
      end else if (10'h1f3 == _T_31[9:0]) begin
        image_0_499 <= io_pixelVal_in_0_5;
      end else if (10'h1f3 == _T_28[9:0]) begin
        image_0_499 <= io_pixelVal_in_0_4;
      end else if (10'h1f3 == _T_25[9:0]) begin
        image_0_499 <= io_pixelVal_in_0_3;
      end else if (10'h1f3 == _T_22[9:0]) begin
        image_0_499 <= io_pixelVal_in_0_2;
      end else if (10'h1f3 == _T_19[9:0]) begin
        image_0_499 <= io_pixelVal_in_0_1;
      end else if (10'h1f3 == _T_15[9:0]) begin
        image_0_499 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_500 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1f4 == _T_37[9:0]) begin
        image_0_500 <= io_pixelVal_in_0_7;
      end else if (10'h1f4 == _T_34[9:0]) begin
        image_0_500 <= io_pixelVal_in_0_6;
      end else if (10'h1f4 == _T_31[9:0]) begin
        image_0_500 <= io_pixelVal_in_0_5;
      end else if (10'h1f4 == _T_28[9:0]) begin
        image_0_500 <= io_pixelVal_in_0_4;
      end else if (10'h1f4 == _T_25[9:0]) begin
        image_0_500 <= io_pixelVal_in_0_3;
      end else if (10'h1f4 == _T_22[9:0]) begin
        image_0_500 <= io_pixelVal_in_0_2;
      end else if (10'h1f4 == _T_19[9:0]) begin
        image_0_500 <= io_pixelVal_in_0_1;
      end else if (10'h1f4 == _T_15[9:0]) begin
        image_0_500 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_501 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1f5 == _T_37[9:0]) begin
        image_0_501 <= io_pixelVal_in_0_7;
      end else if (10'h1f5 == _T_34[9:0]) begin
        image_0_501 <= io_pixelVal_in_0_6;
      end else if (10'h1f5 == _T_31[9:0]) begin
        image_0_501 <= io_pixelVal_in_0_5;
      end else if (10'h1f5 == _T_28[9:0]) begin
        image_0_501 <= io_pixelVal_in_0_4;
      end else if (10'h1f5 == _T_25[9:0]) begin
        image_0_501 <= io_pixelVal_in_0_3;
      end else if (10'h1f5 == _T_22[9:0]) begin
        image_0_501 <= io_pixelVal_in_0_2;
      end else if (10'h1f5 == _T_19[9:0]) begin
        image_0_501 <= io_pixelVal_in_0_1;
      end else if (10'h1f5 == _T_15[9:0]) begin
        image_0_501 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_502 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1f6 == _T_37[9:0]) begin
        image_0_502 <= io_pixelVal_in_0_7;
      end else if (10'h1f6 == _T_34[9:0]) begin
        image_0_502 <= io_pixelVal_in_0_6;
      end else if (10'h1f6 == _T_31[9:0]) begin
        image_0_502 <= io_pixelVal_in_0_5;
      end else if (10'h1f6 == _T_28[9:0]) begin
        image_0_502 <= io_pixelVal_in_0_4;
      end else if (10'h1f6 == _T_25[9:0]) begin
        image_0_502 <= io_pixelVal_in_0_3;
      end else if (10'h1f6 == _T_22[9:0]) begin
        image_0_502 <= io_pixelVal_in_0_2;
      end else if (10'h1f6 == _T_19[9:0]) begin
        image_0_502 <= io_pixelVal_in_0_1;
      end else if (10'h1f6 == _T_15[9:0]) begin
        image_0_502 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_503 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1f7 == _T_37[9:0]) begin
        image_0_503 <= io_pixelVal_in_0_7;
      end else if (10'h1f7 == _T_34[9:0]) begin
        image_0_503 <= io_pixelVal_in_0_6;
      end else if (10'h1f7 == _T_31[9:0]) begin
        image_0_503 <= io_pixelVal_in_0_5;
      end else if (10'h1f7 == _T_28[9:0]) begin
        image_0_503 <= io_pixelVal_in_0_4;
      end else if (10'h1f7 == _T_25[9:0]) begin
        image_0_503 <= io_pixelVal_in_0_3;
      end else if (10'h1f7 == _T_22[9:0]) begin
        image_0_503 <= io_pixelVal_in_0_2;
      end else if (10'h1f7 == _T_19[9:0]) begin
        image_0_503 <= io_pixelVal_in_0_1;
      end else if (10'h1f7 == _T_15[9:0]) begin
        image_0_503 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_504 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1f8 == _T_37[9:0]) begin
        image_0_504 <= io_pixelVal_in_0_7;
      end else if (10'h1f8 == _T_34[9:0]) begin
        image_0_504 <= io_pixelVal_in_0_6;
      end else if (10'h1f8 == _T_31[9:0]) begin
        image_0_504 <= io_pixelVal_in_0_5;
      end else if (10'h1f8 == _T_28[9:0]) begin
        image_0_504 <= io_pixelVal_in_0_4;
      end else if (10'h1f8 == _T_25[9:0]) begin
        image_0_504 <= io_pixelVal_in_0_3;
      end else if (10'h1f8 == _T_22[9:0]) begin
        image_0_504 <= io_pixelVal_in_0_2;
      end else if (10'h1f8 == _T_19[9:0]) begin
        image_0_504 <= io_pixelVal_in_0_1;
      end else if (10'h1f8 == _T_15[9:0]) begin
        image_0_504 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_505 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1f9 == _T_37[9:0]) begin
        image_0_505 <= io_pixelVal_in_0_7;
      end else if (10'h1f9 == _T_34[9:0]) begin
        image_0_505 <= io_pixelVal_in_0_6;
      end else if (10'h1f9 == _T_31[9:0]) begin
        image_0_505 <= io_pixelVal_in_0_5;
      end else if (10'h1f9 == _T_28[9:0]) begin
        image_0_505 <= io_pixelVal_in_0_4;
      end else if (10'h1f9 == _T_25[9:0]) begin
        image_0_505 <= io_pixelVal_in_0_3;
      end else if (10'h1f9 == _T_22[9:0]) begin
        image_0_505 <= io_pixelVal_in_0_2;
      end else if (10'h1f9 == _T_19[9:0]) begin
        image_0_505 <= io_pixelVal_in_0_1;
      end else if (10'h1f9 == _T_15[9:0]) begin
        image_0_505 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_506 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1fa == _T_37[9:0]) begin
        image_0_506 <= io_pixelVal_in_0_7;
      end else if (10'h1fa == _T_34[9:0]) begin
        image_0_506 <= io_pixelVal_in_0_6;
      end else if (10'h1fa == _T_31[9:0]) begin
        image_0_506 <= io_pixelVal_in_0_5;
      end else if (10'h1fa == _T_28[9:0]) begin
        image_0_506 <= io_pixelVal_in_0_4;
      end else if (10'h1fa == _T_25[9:0]) begin
        image_0_506 <= io_pixelVal_in_0_3;
      end else if (10'h1fa == _T_22[9:0]) begin
        image_0_506 <= io_pixelVal_in_0_2;
      end else if (10'h1fa == _T_19[9:0]) begin
        image_0_506 <= io_pixelVal_in_0_1;
      end else if (10'h1fa == _T_15[9:0]) begin
        image_0_506 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_507 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1fb == _T_37[9:0]) begin
        image_0_507 <= io_pixelVal_in_0_7;
      end else if (10'h1fb == _T_34[9:0]) begin
        image_0_507 <= io_pixelVal_in_0_6;
      end else if (10'h1fb == _T_31[9:0]) begin
        image_0_507 <= io_pixelVal_in_0_5;
      end else if (10'h1fb == _T_28[9:0]) begin
        image_0_507 <= io_pixelVal_in_0_4;
      end else if (10'h1fb == _T_25[9:0]) begin
        image_0_507 <= io_pixelVal_in_0_3;
      end else if (10'h1fb == _T_22[9:0]) begin
        image_0_507 <= io_pixelVal_in_0_2;
      end else if (10'h1fb == _T_19[9:0]) begin
        image_0_507 <= io_pixelVal_in_0_1;
      end else if (10'h1fb == _T_15[9:0]) begin
        image_0_507 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_508 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1fc == _T_37[9:0]) begin
        image_0_508 <= io_pixelVal_in_0_7;
      end else if (10'h1fc == _T_34[9:0]) begin
        image_0_508 <= io_pixelVal_in_0_6;
      end else if (10'h1fc == _T_31[9:0]) begin
        image_0_508 <= io_pixelVal_in_0_5;
      end else if (10'h1fc == _T_28[9:0]) begin
        image_0_508 <= io_pixelVal_in_0_4;
      end else if (10'h1fc == _T_25[9:0]) begin
        image_0_508 <= io_pixelVal_in_0_3;
      end else if (10'h1fc == _T_22[9:0]) begin
        image_0_508 <= io_pixelVal_in_0_2;
      end else if (10'h1fc == _T_19[9:0]) begin
        image_0_508 <= io_pixelVal_in_0_1;
      end else if (10'h1fc == _T_15[9:0]) begin
        image_0_508 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_509 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1fd == _T_37[9:0]) begin
        image_0_509 <= io_pixelVal_in_0_7;
      end else if (10'h1fd == _T_34[9:0]) begin
        image_0_509 <= io_pixelVal_in_0_6;
      end else if (10'h1fd == _T_31[9:0]) begin
        image_0_509 <= io_pixelVal_in_0_5;
      end else if (10'h1fd == _T_28[9:0]) begin
        image_0_509 <= io_pixelVal_in_0_4;
      end else if (10'h1fd == _T_25[9:0]) begin
        image_0_509 <= io_pixelVal_in_0_3;
      end else if (10'h1fd == _T_22[9:0]) begin
        image_0_509 <= io_pixelVal_in_0_2;
      end else if (10'h1fd == _T_19[9:0]) begin
        image_0_509 <= io_pixelVal_in_0_1;
      end else if (10'h1fd == _T_15[9:0]) begin
        image_0_509 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_510 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1fe == _T_37[9:0]) begin
        image_0_510 <= io_pixelVal_in_0_7;
      end else if (10'h1fe == _T_34[9:0]) begin
        image_0_510 <= io_pixelVal_in_0_6;
      end else if (10'h1fe == _T_31[9:0]) begin
        image_0_510 <= io_pixelVal_in_0_5;
      end else if (10'h1fe == _T_28[9:0]) begin
        image_0_510 <= io_pixelVal_in_0_4;
      end else if (10'h1fe == _T_25[9:0]) begin
        image_0_510 <= io_pixelVal_in_0_3;
      end else if (10'h1fe == _T_22[9:0]) begin
        image_0_510 <= io_pixelVal_in_0_2;
      end else if (10'h1fe == _T_19[9:0]) begin
        image_0_510 <= io_pixelVal_in_0_1;
      end else if (10'h1fe == _T_15[9:0]) begin
        image_0_510 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_511 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h1ff == _T_37[9:0]) begin
        image_0_511 <= io_pixelVal_in_0_7;
      end else if (10'h1ff == _T_34[9:0]) begin
        image_0_511 <= io_pixelVal_in_0_6;
      end else if (10'h1ff == _T_31[9:0]) begin
        image_0_511 <= io_pixelVal_in_0_5;
      end else if (10'h1ff == _T_28[9:0]) begin
        image_0_511 <= io_pixelVal_in_0_4;
      end else if (10'h1ff == _T_25[9:0]) begin
        image_0_511 <= io_pixelVal_in_0_3;
      end else if (10'h1ff == _T_22[9:0]) begin
        image_0_511 <= io_pixelVal_in_0_2;
      end else if (10'h1ff == _T_19[9:0]) begin
        image_0_511 <= io_pixelVal_in_0_1;
      end else if (10'h1ff == _T_15[9:0]) begin
        image_0_511 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_512 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h200 == _T_37[9:0]) begin
        image_0_512 <= io_pixelVal_in_0_7;
      end else if (10'h200 == _T_34[9:0]) begin
        image_0_512 <= io_pixelVal_in_0_6;
      end else if (10'h200 == _T_31[9:0]) begin
        image_0_512 <= io_pixelVal_in_0_5;
      end else if (10'h200 == _T_28[9:0]) begin
        image_0_512 <= io_pixelVal_in_0_4;
      end else if (10'h200 == _T_25[9:0]) begin
        image_0_512 <= io_pixelVal_in_0_3;
      end else if (10'h200 == _T_22[9:0]) begin
        image_0_512 <= io_pixelVal_in_0_2;
      end else if (10'h200 == _T_19[9:0]) begin
        image_0_512 <= io_pixelVal_in_0_1;
      end else if (10'h200 == _T_15[9:0]) begin
        image_0_512 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_513 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h201 == _T_37[9:0]) begin
        image_0_513 <= io_pixelVal_in_0_7;
      end else if (10'h201 == _T_34[9:0]) begin
        image_0_513 <= io_pixelVal_in_0_6;
      end else if (10'h201 == _T_31[9:0]) begin
        image_0_513 <= io_pixelVal_in_0_5;
      end else if (10'h201 == _T_28[9:0]) begin
        image_0_513 <= io_pixelVal_in_0_4;
      end else if (10'h201 == _T_25[9:0]) begin
        image_0_513 <= io_pixelVal_in_0_3;
      end else if (10'h201 == _T_22[9:0]) begin
        image_0_513 <= io_pixelVal_in_0_2;
      end else if (10'h201 == _T_19[9:0]) begin
        image_0_513 <= io_pixelVal_in_0_1;
      end else if (10'h201 == _T_15[9:0]) begin
        image_0_513 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_514 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h202 == _T_37[9:0]) begin
        image_0_514 <= io_pixelVal_in_0_7;
      end else if (10'h202 == _T_34[9:0]) begin
        image_0_514 <= io_pixelVal_in_0_6;
      end else if (10'h202 == _T_31[9:0]) begin
        image_0_514 <= io_pixelVal_in_0_5;
      end else if (10'h202 == _T_28[9:0]) begin
        image_0_514 <= io_pixelVal_in_0_4;
      end else if (10'h202 == _T_25[9:0]) begin
        image_0_514 <= io_pixelVal_in_0_3;
      end else if (10'h202 == _T_22[9:0]) begin
        image_0_514 <= io_pixelVal_in_0_2;
      end else if (10'h202 == _T_19[9:0]) begin
        image_0_514 <= io_pixelVal_in_0_1;
      end else if (10'h202 == _T_15[9:0]) begin
        image_0_514 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_515 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h203 == _T_37[9:0]) begin
        image_0_515 <= io_pixelVal_in_0_7;
      end else if (10'h203 == _T_34[9:0]) begin
        image_0_515 <= io_pixelVal_in_0_6;
      end else if (10'h203 == _T_31[9:0]) begin
        image_0_515 <= io_pixelVal_in_0_5;
      end else if (10'h203 == _T_28[9:0]) begin
        image_0_515 <= io_pixelVal_in_0_4;
      end else if (10'h203 == _T_25[9:0]) begin
        image_0_515 <= io_pixelVal_in_0_3;
      end else if (10'h203 == _T_22[9:0]) begin
        image_0_515 <= io_pixelVal_in_0_2;
      end else if (10'h203 == _T_19[9:0]) begin
        image_0_515 <= io_pixelVal_in_0_1;
      end else if (10'h203 == _T_15[9:0]) begin
        image_0_515 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_516 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h204 == _T_37[9:0]) begin
        image_0_516 <= io_pixelVal_in_0_7;
      end else if (10'h204 == _T_34[9:0]) begin
        image_0_516 <= io_pixelVal_in_0_6;
      end else if (10'h204 == _T_31[9:0]) begin
        image_0_516 <= io_pixelVal_in_0_5;
      end else if (10'h204 == _T_28[9:0]) begin
        image_0_516 <= io_pixelVal_in_0_4;
      end else if (10'h204 == _T_25[9:0]) begin
        image_0_516 <= io_pixelVal_in_0_3;
      end else if (10'h204 == _T_22[9:0]) begin
        image_0_516 <= io_pixelVal_in_0_2;
      end else if (10'h204 == _T_19[9:0]) begin
        image_0_516 <= io_pixelVal_in_0_1;
      end else if (10'h204 == _T_15[9:0]) begin
        image_0_516 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_517 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h205 == _T_37[9:0]) begin
        image_0_517 <= io_pixelVal_in_0_7;
      end else if (10'h205 == _T_34[9:0]) begin
        image_0_517 <= io_pixelVal_in_0_6;
      end else if (10'h205 == _T_31[9:0]) begin
        image_0_517 <= io_pixelVal_in_0_5;
      end else if (10'h205 == _T_28[9:0]) begin
        image_0_517 <= io_pixelVal_in_0_4;
      end else if (10'h205 == _T_25[9:0]) begin
        image_0_517 <= io_pixelVal_in_0_3;
      end else if (10'h205 == _T_22[9:0]) begin
        image_0_517 <= io_pixelVal_in_0_2;
      end else if (10'h205 == _T_19[9:0]) begin
        image_0_517 <= io_pixelVal_in_0_1;
      end else if (10'h205 == _T_15[9:0]) begin
        image_0_517 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_518 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h206 == _T_37[9:0]) begin
        image_0_518 <= io_pixelVal_in_0_7;
      end else if (10'h206 == _T_34[9:0]) begin
        image_0_518 <= io_pixelVal_in_0_6;
      end else if (10'h206 == _T_31[9:0]) begin
        image_0_518 <= io_pixelVal_in_0_5;
      end else if (10'h206 == _T_28[9:0]) begin
        image_0_518 <= io_pixelVal_in_0_4;
      end else if (10'h206 == _T_25[9:0]) begin
        image_0_518 <= io_pixelVal_in_0_3;
      end else if (10'h206 == _T_22[9:0]) begin
        image_0_518 <= io_pixelVal_in_0_2;
      end else if (10'h206 == _T_19[9:0]) begin
        image_0_518 <= io_pixelVal_in_0_1;
      end else if (10'h206 == _T_15[9:0]) begin
        image_0_518 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_519 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h207 == _T_37[9:0]) begin
        image_0_519 <= io_pixelVal_in_0_7;
      end else if (10'h207 == _T_34[9:0]) begin
        image_0_519 <= io_pixelVal_in_0_6;
      end else if (10'h207 == _T_31[9:0]) begin
        image_0_519 <= io_pixelVal_in_0_5;
      end else if (10'h207 == _T_28[9:0]) begin
        image_0_519 <= io_pixelVal_in_0_4;
      end else if (10'h207 == _T_25[9:0]) begin
        image_0_519 <= io_pixelVal_in_0_3;
      end else if (10'h207 == _T_22[9:0]) begin
        image_0_519 <= io_pixelVal_in_0_2;
      end else if (10'h207 == _T_19[9:0]) begin
        image_0_519 <= io_pixelVal_in_0_1;
      end else if (10'h207 == _T_15[9:0]) begin
        image_0_519 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_520 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h208 == _T_37[9:0]) begin
        image_0_520 <= io_pixelVal_in_0_7;
      end else if (10'h208 == _T_34[9:0]) begin
        image_0_520 <= io_pixelVal_in_0_6;
      end else if (10'h208 == _T_31[9:0]) begin
        image_0_520 <= io_pixelVal_in_0_5;
      end else if (10'h208 == _T_28[9:0]) begin
        image_0_520 <= io_pixelVal_in_0_4;
      end else if (10'h208 == _T_25[9:0]) begin
        image_0_520 <= io_pixelVal_in_0_3;
      end else if (10'h208 == _T_22[9:0]) begin
        image_0_520 <= io_pixelVal_in_0_2;
      end else if (10'h208 == _T_19[9:0]) begin
        image_0_520 <= io_pixelVal_in_0_1;
      end else if (10'h208 == _T_15[9:0]) begin
        image_0_520 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_521 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h209 == _T_37[9:0]) begin
        image_0_521 <= io_pixelVal_in_0_7;
      end else if (10'h209 == _T_34[9:0]) begin
        image_0_521 <= io_pixelVal_in_0_6;
      end else if (10'h209 == _T_31[9:0]) begin
        image_0_521 <= io_pixelVal_in_0_5;
      end else if (10'h209 == _T_28[9:0]) begin
        image_0_521 <= io_pixelVal_in_0_4;
      end else if (10'h209 == _T_25[9:0]) begin
        image_0_521 <= io_pixelVal_in_0_3;
      end else if (10'h209 == _T_22[9:0]) begin
        image_0_521 <= io_pixelVal_in_0_2;
      end else if (10'h209 == _T_19[9:0]) begin
        image_0_521 <= io_pixelVal_in_0_1;
      end else if (10'h209 == _T_15[9:0]) begin
        image_0_521 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_522 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h20a == _T_37[9:0]) begin
        image_0_522 <= io_pixelVal_in_0_7;
      end else if (10'h20a == _T_34[9:0]) begin
        image_0_522 <= io_pixelVal_in_0_6;
      end else if (10'h20a == _T_31[9:0]) begin
        image_0_522 <= io_pixelVal_in_0_5;
      end else if (10'h20a == _T_28[9:0]) begin
        image_0_522 <= io_pixelVal_in_0_4;
      end else if (10'h20a == _T_25[9:0]) begin
        image_0_522 <= io_pixelVal_in_0_3;
      end else if (10'h20a == _T_22[9:0]) begin
        image_0_522 <= io_pixelVal_in_0_2;
      end else if (10'h20a == _T_19[9:0]) begin
        image_0_522 <= io_pixelVal_in_0_1;
      end else if (10'h20a == _T_15[9:0]) begin
        image_0_522 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_523 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h20b == _T_37[9:0]) begin
        image_0_523 <= io_pixelVal_in_0_7;
      end else if (10'h20b == _T_34[9:0]) begin
        image_0_523 <= io_pixelVal_in_0_6;
      end else if (10'h20b == _T_31[9:0]) begin
        image_0_523 <= io_pixelVal_in_0_5;
      end else if (10'h20b == _T_28[9:0]) begin
        image_0_523 <= io_pixelVal_in_0_4;
      end else if (10'h20b == _T_25[9:0]) begin
        image_0_523 <= io_pixelVal_in_0_3;
      end else if (10'h20b == _T_22[9:0]) begin
        image_0_523 <= io_pixelVal_in_0_2;
      end else if (10'h20b == _T_19[9:0]) begin
        image_0_523 <= io_pixelVal_in_0_1;
      end else if (10'h20b == _T_15[9:0]) begin
        image_0_523 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_524 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h20c == _T_37[9:0]) begin
        image_0_524 <= io_pixelVal_in_0_7;
      end else if (10'h20c == _T_34[9:0]) begin
        image_0_524 <= io_pixelVal_in_0_6;
      end else if (10'h20c == _T_31[9:0]) begin
        image_0_524 <= io_pixelVal_in_0_5;
      end else if (10'h20c == _T_28[9:0]) begin
        image_0_524 <= io_pixelVal_in_0_4;
      end else if (10'h20c == _T_25[9:0]) begin
        image_0_524 <= io_pixelVal_in_0_3;
      end else if (10'h20c == _T_22[9:0]) begin
        image_0_524 <= io_pixelVal_in_0_2;
      end else if (10'h20c == _T_19[9:0]) begin
        image_0_524 <= io_pixelVal_in_0_1;
      end else if (10'h20c == _T_15[9:0]) begin
        image_0_524 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_525 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h20d == _T_37[9:0]) begin
        image_0_525 <= io_pixelVal_in_0_7;
      end else if (10'h20d == _T_34[9:0]) begin
        image_0_525 <= io_pixelVal_in_0_6;
      end else if (10'h20d == _T_31[9:0]) begin
        image_0_525 <= io_pixelVal_in_0_5;
      end else if (10'h20d == _T_28[9:0]) begin
        image_0_525 <= io_pixelVal_in_0_4;
      end else if (10'h20d == _T_25[9:0]) begin
        image_0_525 <= io_pixelVal_in_0_3;
      end else if (10'h20d == _T_22[9:0]) begin
        image_0_525 <= io_pixelVal_in_0_2;
      end else if (10'h20d == _T_19[9:0]) begin
        image_0_525 <= io_pixelVal_in_0_1;
      end else if (10'h20d == _T_15[9:0]) begin
        image_0_525 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_526 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h20e == _T_37[9:0]) begin
        image_0_526 <= io_pixelVal_in_0_7;
      end else if (10'h20e == _T_34[9:0]) begin
        image_0_526 <= io_pixelVal_in_0_6;
      end else if (10'h20e == _T_31[9:0]) begin
        image_0_526 <= io_pixelVal_in_0_5;
      end else if (10'h20e == _T_28[9:0]) begin
        image_0_526 <= io_pixelVal_in_0_4;
      end else if (10'h20e == _T_25[9:0]) begin
        image_0_526 <= io_pixelVal_in_0_3;
      end else if (10'h20e == _T_22[9:0]) begin
        image_0_526 <= io_pixelVal_in_0_2;
      end else if (10'h20e == _T_19[9:0]) begin
        image_0_526 <= io_pixelVal_in_0_1;
      end else if (10'h20e == _T_15[9:0]) begin
        image_0_526 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_527 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h20f == _T_37[9:0]) begin
        image_0_527 <= io_pixelVal_in_0_7;
      end else if (10'h20f == _T_34[9:0]) begin
        image_0_527 <= io_pixelVal_in_0_6;
      end else if (10'h20f == _T_31[9:0]) begin
        image_0_527 <= io_pixelVal_in_0_5;
      end else if (10'h20f == _T_28[9:0]) begin
        image_0_527 <= io_pixelVal_in_0_4;
      end else if (10'h20f == _T_25[9:0]) begin
        image_0_527 <= io_pixelVal_in_0_3;
      end else if (10'h20f == _T_22[9:0]) begin
        image_0_527 <= io_pixelVal_in_0_2;
      end else if (10'h20f == _T_19[9:0]) begin
        image_0_527 <= io_pixelVal_in_0_1;
      end else if (10'h20f == _T_15[9:0]) begin
        image_0_527 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_528 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h210 == _T_37[9:0]) begin
        image_0_528 <= io_pixelVal_in_0_7;
      end else if (10'h210 == _T_34[9:0]) begin
        image_0_528 <= io_pixelVal_in_0_6;
      end else if (10'h210 == _T_31[9:0]) begin
        image_0_528 <= io_pixelVal_in_0_5;
      end else if (10'h210 == _T_28[9:0]) begin
        image_0_528 <= io_pixelVal_in_0_4;
      end else if (10'h210 == _T_25[9:0]) begin
        image_0_528 <= io_pixelVal_in_0_3;
      end else if (10'h210 == _T_22[9:0]) begin
        image_0_528 <= io_pixelVal_in_0_2;
      end else if (10'h210 == _T_19[9:0]) begin
        image_0_528 <= io_pixelVal_in_0_1;
      end else if (10'h210 == _T_15[9:0]) begin
        image_0_528 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_529 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h211 == _T_37[9:0]) begin
        image_0_529 <= io_pixelVal_in_0_7;
      end else if (10'h211 == _T_34[9:0]) begin
        image_0_529 <= io_pixelVal_in_0_6;
      end else if (10'h211 == _T_31[9:0]) begin
        image_0_529 <= io_pixelVal_in_0_5;
      end else if (10'h211 == _T_28[9:0]) begin
        image_0_529 <= io_pixelVal_in_0_4;
      end else if (10'h211 == _T_25[9:0]) begin
        image_0_529 <= io_pixelVal_in_0_3;
      end else if (10'h211 == _T_22[9:0]) begin
        image_0_529 <= io_pixelVal_in_0_2;
      end else if (10'h211 == _T_19[9:0]) begin
        image_0_529 <= io_pixelVal_in_0_1;
      end else if (10'h211 == _T_15[9:0]) begin
        image_0_529 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_530 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h212 == _T_37[9:0]) begin
        image_0_530 <= io_pixelVal_in_0_7;
      end else if (10'h212 == _T_34[9:0]) begin
        image_0_530 <= io_pixelVal_in_0_6;
      end else if (10'h212 == _T_31[9:0]) begin
        image_0_530 <= io_pixelVal_in_0_5;
      end else if (10'h212 == _T_28[9:0]) begin
        image_0_530 <= io_pixelVal_in_0_4;
      end else if (10'h212 == _T_25[9:0]) begin
        image_0_530 <= io_pixelVal_in_0_3;
      end else if (10'h212 == _T_22[9:0]) begin
        image_0_530 <= io_pixelVal_in_0_2;
      end else if (10'h212 == _T_19[9:0]) begin
        image_0_530 <= io_pixelVal_in_0_1;
      end else if (10'h212 == _T_15[9:0]) begin
        image_0_530 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_531 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h213 == _T_37[9:0]) begin
        image_0_531 <= io_pixelVal_in_0_7;
      end else if (10'h213 == _T_34[9:0]) begin
        image_0_531 <= io_pixelVal_in_0_6;
      end else if (10'h213 == _T_31[9:0]) begin
        image_0_531 <= io_pixelVal_in_0_5;
      end else if (10'h213 == _T_28[9:0]) begin
        image_0_531 <= io_pixelVal_in_0_4;
      end else if (10'h213 == _T_25[9:0]) begin
        image_0_531 <= io_pixelVal_in_0_3;
      end else if (10'h213 == _T_22[9:0]) begin
        image_0_531 <= io_pixelVal_in_0_2;
      end else if (10'h213 == _T_19[9:0]) begin
        image_0_531 <= io_pixelVal_in_0_1;
      end else if (10'h213 == _T_15[9:0]) begin
        image_0_531 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_532 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h214 == _T_37[9:0]) begin
        image_0_532 <= io_pixelVal_in_0_7;
      end else if (10'h214 == _T_34[9:0]) begin
        image_0_532 <= io_pixelVal_in_0_6;
      end else if (10'h214 == _T_31[9:0]) begin
        image_0_532 <= io_pixelVal_in_0_5;
      end else if (10'h214 == _T_28[9:0]) begin
        image_0_532 <= io_pixelVal_in_0_4;
      end else if (10'h214 == _T_25[9:0]) begin
        image_0_532 <= io_pixelVal_in_0_3;
      end else if (10'h214 == _T_22[9:0]) begin
        image_0_532 <= io_pixelVal_in_0_2;
      end else if (10'h214 == _T_19[9:0]) begin
        image_0_532 <= io_pixelVal_in_0_1;
      end else if (10'h214 == _T_15[9:0]) begin
        image_0_532 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_533 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h215 == _T_37[9:0]) begin
        image_0_533 <= io_pixelVal_in_0_7;
      end else if (10'h215 == _T_34[9:0]) begin
        image_0_533 <= io_pixelVal_in_0_6;
      end else if (10'h215 == _T_31[9:0]) begin
        image_0_533 <= io_pixelVal_in_0_5;
      end else if (10'h215 == _T_28[9:0]) begin
        image_0_533 <= io_pixelVal_in_0_4;
      end else if (10'h215 == _T_25[9:0]) begin
        image_0_533 <= io_pixelVal_in_0_3;
      end else if (10'h215 == _T_22[9:0]) begin
        image_0_533 <= io_pixelVal_in_0_2;
      end else if (10'h215 == _T_19[9:0]) begin
        image_0_533 <= io_pixelVal_in_0_1;
      end else if (10'h215 == _T_15[9:0]) begin
        image_0_533 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_534 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h216 == _T_37[9:0]) begin
        image_0_534 <= io_pixelVal_in_0_7;
      end else if (10'h216 == _T_34[9:0]) begin
        image_0_534 <= io_pixelVal_in_0_6;
      end else if (10'h216 == _T_31[9:0]) begin
        image_0_534 <= io_pixelVal_in_0_5;
      end else if (10'h216 == _T_28[9:0]) begin
        image_0_534 <= io_pixelVal_in_0_4;
      end else if (10'h216 == _T_25[9:0]) begin
        image_0_534 <= io_pixelVal_in_0_3;
      end else if (10'h216 == _T_22[9:0]) begin
        image_0_534 <= io_pixelVal_in_0_2;
      end else if (10'h216 == _T_19[9:0]) begin
        image_0_534 <= io_pixelVal_in_0_1;
      end else if (10'h216 == _T_15[9:0]) begin
        image_0_534 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_535 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h217 == _T_37[9:0]) begin
        image_0_535 <= io_pixelVal_in_0_7;
      end else if (10'h217 == _T_34[9:0]) begin
        image_0_535 <= io_pixelVal_in_0_6;
      end else if (10'h217 == _T_31[9:0]) begin
        image_0_535 <= io_pixelVal_in_0_5;
      end else if (10'h217 == _T_28[9:0]) begin
        image_0_535 <= io_pixelVal_in_0_4;
      end else if (10'h217 == _T_25[9:0]) begin
        image_0_535 <= io_pixelVal_in_0_3;
      end else if (10'h217 == _T_22[9:0]) begin
        image_0_535 <= io_pixelVal_in_0_2;
      end else if (10'h217 == _T_19[9:0]) begin
        image_0_535 <= io_pixelVal_in_0_1;
      end else if (10'h217 == _T_15[9:0]) begin
        image_0_535 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_536 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h218 == _T_37[9:0]) begin
        image_0_536 <= io_pixelVal_in_0_7;
      end else if (10'h218 == _T_34[9:0]) begin
        image_0_536 <= io_pixelVal_in_0_6;
      end else if (10'h218 == _T_31[9:0]) begin
        image_0_536 <= io_pixelVal_in_0_5;
      end else if (10'h218 == _T_28[9:0]) begin
        image_0_536 <= io_pixelVal_in_0_4;
      end else if (10'h218 == _T_25[9:0]) begin
        image_0_536 <= io_pixelVal_in_0_3;
      end else if (10'h218 == _T_22[9:0]) begin
        image_0_536 <= io_pixelVal_in_0_2;
      end else if (10'h218 == _T_19[9:0]) begin
        image_0_536 <= io_pixelVal_in_0_1;
      end else if (10'h218 == _T_15[9:0]) begin
        image_0_536 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_537 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h219 == _T_37[9:0]) begin
        image_0_537 <= io_pixelVal_in_0_7;
      end else if (10'h219 == _T_34[9:0]) begin
        image_0_537 <= io_pixelVal_in_0_6;
      end else if (10'h219 == _T_31[9:0]) begin
        image_0_537 <= io_pixelVal_in_0_5;
      end else if (10'h219 == _T_28[9:0]) begin
        image_0_537 <= io_pixelVal_in_0_4;
      end else if (10'h219 == _T_25[9:0]) begin
        image_0_537 <= io_pixelVal_in_0_3;
      end else if (10'h219 == _T_22[9:0]) begin
        image_0_537 <= io_pixelVal_in_0_2;
      end else if (10'h219 == _T_19[9:0]) begin
        image_0_537 <= io_pixelVal_in_0_1;
      end else if (10'h219 == _T_15[9:0]) begin
        image_0_537 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_538 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h21a == _T_37[9:0]) begin
        image_0_538 <= io_pixelVal_in_0_7;
      end else if (10'h21a == _T_34[9:0]) begin
        image_0_538 <= io_pixelVal_in_0_6;
      end else if (10'h21a == _T_31[9:0]) begin
        image_0_538 <= io_pixelVal_in_0_5;
      end else if (10'h21a == _T_28[9:0]) begin
        image_0_538 <= io_pixelVal_in_0_4;
      end else if (10'h21a == _T_25[9:0]) begin
        image_0_538 <= io_pixelVal_in_0_3;
      end else if (10'h21a == _T_22[9:0]) begin
        image_0_538 <= io_pixelVal_in_0_2;
      end else if (10'h21a == _T_19[9:0]) begin
        image_0_538 <= io_pixelVal_in_0_1;
      end else if (10'h21a == _T_15[9:0]) begin
        image_0_538 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_539 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h21b == _T_37[9:0]) begin
        image_0_539 <= io_pixelVal_in_0_7;
      end else if (10'h21b == _T_34[9:0]) begin
        image_0_539 <= io_pixelVal_in_0_6;
      end else if (10'h21b == _T_31[9:0]) begin
        image_0_539 <= io_pixelVal_in_0_5;
      end else if (10'h21b == _T_28[9:0]) begin
        image_0_539 <= io_pixelVal_in_0_4;
      end else if (10'h21b == _T_25[9:0]) begin
        image_0_539 <= io_pixelVal_in_0_3;
      end else if (10'h21b == _T_22[9:0]) begin
        image_0_539 <= io_pixelVal_in_0_2;
      end else if (10'h21b == _T_19[9:0]) begin
        image_0_539 <= io_pixelVal_in_0_1;
      end else if (10'h21b == _T_15[9:0]) begin
        image_0_539 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_540 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h21c == _T_37[9:0]) begin
        image_0_540 <= io_pixelVal_in_0_7;
      end else if (10'h21c == _T_34[9:0]) begin
        image_0_540 <= io_pixelVal_in_0_6;
      end else if (10'h21c == _T_31[9:0]) begin
        image_0_540 <= io_pixelVal_in_0_5;
      end else if (10'h21c == _T_28[9:0]) begin
        image_0_540 <= io_pixelVal_in_0_4;
      end else if (10'h21c == _T_25[9:0]) begin
        image_0_540 <= io_pixelVal_in_0_3;
      end else if (10'h21c == _T_22[9:0]) begin
        image_0_540 <= io_pixelVal_in_0_2;
      end else if (10'h21c == _T_19[9:0]) begin
        image_0_540 <= io_pixelVal_in_0_1;
      end else if (10'h21c == _T_15[9:0]) begin
        image_0_540 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_541 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h21d == _T_37[9:0]) begin
        image_0_541 <= io_pixelVal_in_0_7;
      end else if (10'h21d == _T_34[9:0]) begin
        image_0_541 <= io_pixelVal_in_0_6;
      end else if (10'h21d == _T_31[9:0]) begin
        image_0_541 <= io_pixelVal_in_0_5;
      end else if (10'h21d == _T_28[9:0]) begin
        image_0_541 <= io_pixelVal_in_0_4;
      end else if (10'h21d == _T_25[9:0]) begin
        image_0_541 <= io_pixelVal_in_0_3;
      end else if (10'h21d == _T_22[9:0]) begin
        image_0_541 <= io_pixelVal_in_0_2;
      end else if (10'h21d == _T_19[9:0]) begin
        image_0_541 <= io_pixelVal_in_0_1;
      end else if (10'h21d == _T_15[9:0]) begin
        image_0_541 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_542 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h21e == _T_37[9:0]) begin
        image_0_542 <= io_pixelVal_in_0_7;
      end else if (10'h21e == _T_34[9:0]) begin
        image_0_542 <= io_pixelVal_in_0_6;
      end else if (10'h21e == _T_31[9:0]) begin
        image_0_542 <= io_pixelVal_in_0_5;
      end else if (10'h21e == _T_28[9:0]) begin
        image_0_542 <= io_pixelVal_in_0_4;
      end else if (10'h21e == _T_25[9:0]) begin
        image_0_542 <= io_pixelVal_in_0_3;
      end else if (10'h21e == _T_22[9:0]) begin
        image_0_542 <= io_pixelVal_in_0_2;
      end else if (10'h21e == _T_19[9:0]) begin
        image_0_542 <= io_pixelVal_in_0_1;
      end else if (10'h21e == _T_15[9:0]) begin
        image_0_542 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_543 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h21f == _T_37[9:0]) begin
        image_0_543 <= io_pixelVal_in_0_7;
      end else if (10'h21f == _T_34[9:0]) begin
        image_0_543 <= io_pixelVal_in_0_6;
      end else if (10'h21f == _T_31[9:0]) begin
        image_0_543 <= io_pixelVal_in_0_5;
      end else if (10'h21f == _T_28[9:0]) begin
        image_0_543 <= io_pixelVal_in_0_4;
      end else if (10'h21f == _T_25[9:0]) begin
        image_0_543 <= io_pixelVal_in_0_3;
      end else if (10'h21f == _T_22[9:0]) begin
        image_0_543 <= io_pixelVal_in_0_2;
      end else if (10'h21f == _T_19[9:0]) begin
        image_0_543 <= io_pixelVal_in_0_1;
      end else if (10'h21f == _T_15[9:0]) begin
        image_0_543 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_544 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h220 == _T_37[9:0]) begin
        image_0_544 <= io_pixelVal_in_0_7;
      end else if (10'h220 == _T_34[9:0]) begin
        image_0_544 <= io_pixelVal_in_0_6;
      end else if (10'h220 == _T_31[9:0]) begin
        image_0_544 <= io_pixelVal_in_0_5;
      end else if (10'h220 == _T_28[9:0]) begin
        image_0_544 <= io_pixelVal_in_0_4;
      end else if (10'h220 == _T_25[9:0]) begin
        image_0_544 <= io_pixelVal_in_0_3;
      end else if (10'h220 == _T_22[9:0]) begin
        image_0_544 <= io_pixelVal_in_0_2;
      end else if (10'h220 == _T_19[9:0]) begin
        image_0_544 <= io_pixelVal_in_0_1;
      end else if (10'h220 == _T_15[9:0]) begin
        image_0_544 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_545 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h221 == _T_37[9:0]) begin
        image_0_545 <= io_pixelVal_in_0_7;
      end else if (10'h221 == _T_34[9:0]) begin
        image_0_545 <= io_pixelVal_in_0_6;
      end else if (10'h221 == _T_31[9:0]) begin
        image_0_545 <= io_pixelVal_in_0_5;
      end else if (10'h221 == _T_28[9:0]) begin
        image_0_545 <= io_pixelVal_in_0_4;
      end else if (10'h221 == _T_25[9:0]) begin
        image_0_545 <= io_pixelVal_in_0_3;
      end else if (10'h221 == _T_22[9:0]) begin
        image_0_545 <= io_pixelVal_in_0_2;
      end else if (10'h221 == _T_19[9:0]) begin
        image_0_545 <= io_pixelVal_in_0_1;
      end else if (10'h221 == _T_15[9:0]) begin
        image_0_545 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_546 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h222 == _T_37[9:0]) begin
        image_0_546 <= io_pixelVal_in_0_7;
      end else if (10'h222 == _T_34[9:0]) begin
        image_0_546 <= io_pixelVal_in_0_6;
      end else if (10'h222 == _T_31[9:0]) begin
        image_0_546 <= io_pixelVal_in_0_5;
      end else if (10'h222 == _T_28[9:0]) begin
        image_0_546 <= io_pixelVal_in_0_4;
      end else if (10'h222 == _T_25[9:0]) begin
        image_0_546 <= io_pixelVal_in_0_3;
      end else if (10'h222 == _T_22[9:0]) begin
        image_0_546 <= io_pixelVal_in_0_2;
      end else if (10'h222 == _T_19[9:0]) begin
        image_0_546 <= io_pixelVal_in_0_1;
      end else if (10'h222 == _T_15[9:0]) begin
        image_0_546 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_547 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h223 == _T_37[9:0]) begin
        image_0_547 <= io_pixelVal_in_0_7;
      end else if (10'h223 == _T_34[9:0]) begin
        image_0_547 <= io_pixelVal_in_0_6;
      end else if (10'h223 == _T_31[9:0]) begin
        image_0_547 <= io_pixelVal_in_0_5;
      end else if (10'h223 == _T_28[9:0]) begin
        image_0_547 <= io_pixelVal_in_0_4;
      end else if (10'h223 == _T_25[9:0]) begin
        image_0_547 <= io_pixelVal_in_0_3;
      end else if (10'h223 == _T_22[9:0]) begin
        image_0_547 <= io_pixelVal_in_0_2;
      end else if (10'h223 == _T_19[9:0]) begin
        image_0_547 <= io_pixelVal_in_0_1;
      end else if (10'h223 == _T_15[9:0]) begin
        image_0_547 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_548 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h224 == _T_37[9:0]) begin
        image_0_548 <= io_pixelVal_in_0_7;
      end else if (10'h224 == _T_34[9:0]) begin
        image_0_548 <= io_pixelVal_in_0_6;
      end else if (10'h224 == _T_31[9:0]) begin
        image_0_548 <= io_pixelVal_in_0_5;
      end else if (10'h224 == _T_28[9:0]) begin
        image_0_548 <= io_pixelVal_in_0_4;
      end else if (10'h224 == _T_25[9:0]) begin
        image_0_548 <= io_pixelVal_in_0_3;
      end else if (10'h224 == _T_22[9:0]) begin
        image_0_548 <= io_pixelVal_in_0_2;
      end else if (10'h224 == _T_19[9:0]) begin
        image_0_548 <= io_pixelVal_in_0_1;
      end else if (10'h224 == _T_15[9:0]) begin
        image_0_548 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_549 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h225 == _T_37[9:0]) begin
        image_0_549 <= io_pixelVal_in_0_7;
      end else if (10'h225 == _T_34[9:0]) begin
        image_0_549 <= io_pixelVal_in_0_6;
      end else if (10'h225 == _T_31[9:0]) begin
        image_0_549 <= io_pixelVal_in_0_5;
      end else if (10'h225 == _T_28[9:0]) begin
        image_0_549 <= io_pixelVal_in_0_4;
      end else if (10'h225 == _T_25[9:0]) begin
        image_0_549 <= io_pixelVal_in_0_3;
      end else if (10'h225 == _T_22[9:0]) begin
        image_0_549 <= io_pixelVal_in_0_2;
      end else if (10'h225 == _T_19[9:0]) begin
        image_0_549 <= io_pixelVal_in_0_1;
      end else if (10'h225 == _T_15[9:0]) begin
        image_0_549 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_550 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h226 == _T_37[9:0]) begin
        image_0_550 <= io_pixelVal_in_0_7;
      end else if (10'h226 == _T_34[9:0]) begin
        image_0_550 <= io_pixelVal_in_0_6;
      end else if (10'h226 == _T_31[9:0]) begin
        image_0_550 <= io_pixelVal_in_0_5;
      end else if (10'h226 == _T_28[9:0]) begin
        image_0_550 <= io_pixelVal_in_0_4;
      end else if (10'h226 == _T_25[9:0]) begin
        image_0_550 <= io_pixelVal_in_0_3;
      end else if (10'h226 == _T_22[9:0]) begin
        image_0_550 <= io_pixelVal_in_0_2;
      end else if (10'h226 == _T_19[9:0]) begin
        image_0_550 <= io_pixelVal_in_0_1;
      end else if (10'h226 == _T_15[9:0]) begin
        image_0_550 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_551 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h227 == _T_37[9:0]) begin
        image_0_551 <= io_pixelVal_in_0_7;
      end else if (10'h227 == _T_34[9:0]) begin
        image_0_551 <= io_pixelVal_in_0_6;
      end else if (10'h227 == _T_31[9:0]) begin
        image_0_551 <= io_pixelVal_in_0_5;
      end else if (10'h227 == _T_28[9:0]) begin
        image_0_551 <= io_pixelVal_in_0_4;
      end else if (10'h227 == _T_25[9:0]) begin
        image_0_551 <= io_pixelVal_in_0_3;
      end else if (10'h227 == _T_22[9:0]) begin
        image_0_551 <= io_pixelVal_in_0_2;
      end else if (10'h227 == _T_19[9:0]) begin
        image_0_551 <= io_pixelVal_in_0_1;
      end else if (10'h227 == _T_15[9:0]) begin
        image_0_551 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_552 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h228 == _T_37[9:0]) begin
        image_0_552 <= io_pixelVal_in_0_7;
      end else if (10'h228 == _T_34[9:0]) begin
        image_0_552 <= io_pixelVal_in_0_6;
      end else if (10'h228 == _T_31[9:0]) begin
        image_0_552 <= io_pixelVal_in_0_5;
      end else if (10'h228 == _T_28[9:0]) begin
        image_0_552 <= io_pixelVal_in_0_4;
      end else if (10'h228 == _T_25[9:0]) begin
        image_0_552 <= io_pixelVal_in_0_3;
      end else if (10'h228 == _T_22[9:0]) begin
        image_0_552 <= io_pixelVal_in_0_2;
      end else if (10'h228 == _T_19[9:0]) begin
        image_0_552 <= io_pixelVal_in_0_1;
      end else if (10'h228 == _T_15[9:0]) begin
        image_0_552 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_553 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h229 == _T_37[9:0]) begin
        image_0_553 <= io_pixelVal_in_0_7;
      end else if (10'h229 == _T_34[9:0]) begin
        image_0_553 <= io_pixelVal_in_0_6;
      end else if (10'h229 == _T_31[9:0]) begin
        image_0_553 <= io_pixelVal_in_0_5;
      end else if (10'h229 == _T_28[9:0]) begin
        image_0_553 <= io_pixelVal_in_0_4;
      end else if (10'h229 == _T_25[9:0]) begin
        image_0_553 <= io_pixelVal_in_0_3;
      end else if (10'h229 == _T_22[9:0]) begin
        image_0_553 <= io_pixelVal_in_0_2;
      end else if (10'h229 == _T_19[9:0]) begin
        image_0_553 <= io_pixelVal_in_0_1;
      end else if (10'h229 == _T_15[9:0]) begin
        image_0_553 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_554 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h22a == _T_37[9:0]) begin
        image_0_554 <= io_pixelVal_in_0_7;
      end else if (10'h22a == _T_34[9:0]) begin
        image_0_554 <= io_pixelVal_in_0_6;
      end else if (10'h22a == _T_31[9:0]) begin
        image_0_554 <= io_pixelVal_in_0_5;
      end else if (10'h22a == _T_28[9:0]) begin
        image_0_554 <= io_pixelVal_in_0_4;
      end else if (10'h22a == _T_25[9:0]) begin
        image_0_554 <= io_pixelVal_in_0_3;
      end else if (10'h22a == _T_22[9:0]) begin
        image_0_554 <= io_pixelVal_in_0_2;
      end else if (10'h22a == _T_19[9:0]) begin
        image_0_554 <= io_pixelVal_in_0_1;
      end else if (10'h22a == _T_15[9:0]) begin
        image_0_554 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_555 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h22b == _T_37[9:0]) begin
        image_0_555 <= io_pixelVal_in_0_7;
      end else if (10'h22b == _T_34[9:0]) begin
        image_0_555 <= io_pixelVal_in_0_6;
      end else if (10'h22b == _T_31[9:0]) begin
        image_0_555 <= io_pixelVal_in_0_5;
      end else if (10'h22b == _T_28[9:0]) begin
        image_0_555 <= io_pixelVal_in_0_4;
      end else if (10'h22b == _T_25[9:0]) begin
        image_0_555 <= io_pixelVal_in_0_3;
      end else if (10'h22b == _T_22[9:0]) begin
        image_0_555 <= io_pixelVal_in_0_2;
      end else if (10'h22b == _T_19[9:0]) begin
        image_0_555 <= io_pixelVal_in_0_1;
      end else if (10'h22b == _T_15[9:0]) begin
        image_0_555 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_556 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h22c == _T_37[9:0]) begin
        image_0_556 <= io_pixelVal_in_0_7;
      end else if (10'h22c == _T_34[9:0]) begin
        image_0_556 <= io_pixelVal_in_0_6;
      end else if (10'h22c == _T_31[9:0]) begin
        image_0_556 <= io_pixelVal_in_0_5;
      end else if (10'h22c == _T_28[9:0]) begin
        image_0_556 <= io_pixelVal_in_0_4;
      end else if (10'h22c == _T_25[9:0]) begin
        image_0_556 <= io_pixelVal_in_0_3;
      end else if (10'h22c == _T_22[9:0]) begin
        image_0_556 <= io_pixelVal_in_0_2;
      end else if (10'h22c == _T_19[9:0]) begin
        image_0_556 <= io_pixelVal_in_0_1;
      end else if (10'h22c == _T_15[9:0]) begin
        image_0_556 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_557 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h22d == _T_37[9:0]) begin
        image_0_557 <= io_pixelVal_in_0_7;
      end else if (10'h22d == _T_34[9:0]) begin
        image_0_557 <= io_pixelVal_in_0_6;
      end else if (10'h22d == _T_31[9:0]) begin
        image_0_557 <= io_pixelVal_in_0_5;
      end else if (10'h22d == _T_28[9:0]) begin
        image_0_557 <= io_pixelVal_in_0_4;
      end else if (10'h22d == _T_25[9:0]) begin
        image_0_557 <= io_pixelVal_in_0_3;
      end else if (10'h22d == _T_22[9:0]) begin
        image_0_557 <= io_pixelVal_in_0_2;
      end else if (10'h22d == _T_19[9:0]) begin
        image_0_557 <= io_pixelVal_in_0_1;
      end else if (10'h22d == _T_15[9:0]) begin
        image_0_557 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_558 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h22e == _T_37[9:0]) begin
        image_0_558 <= io_pixelVal_in_0_7;
      end else if (10'h22e == _T_34[9:0]) begin
        image_0_558 <= io_pixelVal_in_0_6;
      end else if (10'h22e == _T_31[9:0]) begin
        image_0_558 <= io_pixelVal_in_0_5;
      end else if (10'h22e == _T_28[9:0]) begin
        image_0_558 <= io_pixelVal_in_0_4;
      end else if (10'h22e == _T_25[9:0]) begin
        image_0_558 <= io_pixelVal_in_0_3;
      end else if (10'h22e == _T_22[9:0]) begin
        image_0_558 <= io_pixelVal_in_0_2;
      end else if (10'h22e == _T_19[9:0]) begin
        image_0_558 <= io_pixelVal_in_0_1;
      end else if (10'h22e == _T_15[9:0]) begin
        image_0_558 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_559 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h22f == _T_37[9:0]) begin
        image_0_559 <= io_pixelVal_in_0_7;
      end else if (10'h22f == _T_34[9:0]) begin
        image_0_559 <= io_pixelVal_in_0_6;
      end else if (10'h22f == _T_31[9:0]) begin
        image_0_559 <= io_pixelVal_in_0_5;
      end else if (10'h22f == _T_28[9:0]) begin
        image_0_559 <= io_pixelVal_in_0_4;
      end else if (10'h22f == _T_25[9:0]) begin
        image_0_559 <= io_pixelVal_in_0_3;
      end else if (10'h22f == _T_22[9:0]) begin
        image_0_559 <= io_pixelVal_in_0_2;
      end else if (10'h22f == _T_19[9:0]) begin
        image_0_559 <= io_pixelVal_in_0_1;
      end else if (10'h22f == _T_15[9:0]) begin
        image_0_559 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_560 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h230 == _T_37[9:0]) begin
        image_0_560 <= io_pixelVal_in_0_7;
      end else if (10'h230 == _T_34[9:0]) begin
        image_0_560 <= io_pixelVal_in_0_6;
      end else if (10'h230 == _T_31[9:0]) begin
        image_0_560 <= io_pixelVal_in_0_5;
      end else if (10'h230 == _T_28[9:0]) begin
        image_0_560 <= io_pixelVal_in_0_4;
      end else if (10'h230 == _T_25[9:0]) begin
        image_0_560 <= io_pixelVal_in_0_3;
      end else if (10'h230 == _T_22[9:0]) begin
        image_0_560 <= io_pixelVal_in_0_2;
      end else if (10'h230 == _T_19[9:0]) begin
        image_0_560 <= io_pixelVal_in_0_1;
      end else if (10'h230 == _T_15[9:0]) begin
        image_0_560 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_561 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h231 == _T_37[9:0]) begin
        image_0_561 <= io_pixelVal_in_0_7;
      end else if (10'h231 == _T_34[9:0]) begin
        image_0_561 <= io_pixelVal_in_0_6;
      end else if (10'h231 == _T_31[9:0]) begin
        image_0_561 <= io_pixelVal_in_0_5;
      end else if (10'h231 == _T_28[9:0]) begin
        image_0_561 <= io_pixelVal_in_0_4;
      end else if (10'h231 == _T_25[9:0]) begin
        image_0_561 <= io_pixelVal_in_0_3;
      end else if (10'h231 == _T_22[9:0]) begin
        image_0_561 <= io_pixelVal_in_0_2;
      end else if (10'h231 == _T_19[9:0]) begin
        image_0_561 <= io_pixelVal_in_0_1;
      end else if (10'h231 == _T_15[9:0]) begin
        image_0_561 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_562 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h232 == _T_37[9:0]) begin
        image_0_562 <= io_pixelVal_in_0_7;
      end else if (10'h232 == _T_34[9:0]) begin
        image_0_562 <= io_pixelVal_in_0_6;
      end else if (10'h232 == _T_31[9:0]) begin
        image_0_562 <= io_pixelVal_in_0_5;
      end else if (10'h232 == _T_28[9:0]) begin
        image_0_562 <= io_pixelVal_in_0_4;
      end else if (10'h232 == _T_25[9:0]) begin
        image_0_562 <= io_pixelVal_in_0_3;
      end else if (10'h232 == _T_22[9:0]) begin
        image_0_562 <= io_pixelVal_in_0_2;
      end else if (10'h232 == _T_19[9:0]) begin
        image_0_562 <= io_pixelVal_in_0_1;
      end else if (10'h232 == _T_15[9:0]) begin
        image_0_562 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_563 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h233 == _T_37[9:0]) begin
        image_0_563 <= io_pixelVal_in_0_7;
      end else if (10'h233 == _T_34[9:0]) begin
        image_0_563 <= io_pixelVal_in_0_6;
      end else if (10'h233 == _T_31[9:0]) begin
        image_0_563 <= io_pixelVal_in_0_5;
      end else if (10'h233 == _T_28[9:0]) begin
        image_0_563 <= io_pixelVal_in_0_4;
      end else if (10'h233 == _T_25[9:0]) begin
        image_0_563 <= io_pixelVal_in_0_3;
      end else if (10'h233 == _T_22[9:0]) begin
        image_0_563 <= io_pixelVal_in_0_2;
      end else if (10'h233 == _T_19[9:0]) begin
        image_0_563 <= io_pixelVal_in_0_1;
      end else if (10'h233 == _T_15[9:0]) begin
        image_0_563 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_564 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h234 == _T_37[9:0]) begin
        image_0_564 <= io_pixelVal_in_0_7;
      end else if (10'h234 == _T_34[9:0]) begin
        image_0_564 <= io_pixelVal_in_0_6;
      end else if (10'h234 == _T_31[9:0]) begin
        image_0_564 <= io_pixelVal_in_0_5;
      end else if (10'h234 == _T_28[9:0]) begin
        image_0_564 <= io_pixelVal_in_0_4;
      end else if (10'h234 == _T_25[9:0]) begin
        image_0_564 <= io_pixelVal_in_0_3;
      end else if (10'h234 == _T_22[9:0]) begin
        image_0_564 <= io_pixelVal_in_0_2;
      end else if (10'h234 == _T_19[9:0]) begin
        image_0_564 <= io_pixelVal_in_0_1;
      end else if (10'h234 == _T_15[9:0]) begin
        image_0_564 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_565 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h235 == _T_37[9:0]) begin
        image_0_565 <= io_pixelVal_in_0_7;
      end else if (10'h235 == _T_34[9:0]) begin
        image_0_565 <= io_pixelVal_in_0_6;
      end else if (10'h235 == _T_31[9:0]) begin
        image_0_565 <= io_pixelVal_in_0_5;
      end else if (10'h235 == _T_28[9:0]) begin
        image_0_565 <= io_pixelVal_in_0_4;
      end else if (10'h235 == _T_25[9:0]) begin
        image_0_565 <= io_pixelVal_in_0_3;
      end else if (10'h235 == _T_22[9:0]) begin
        image_0_565 <= io_pixelVal_in_0_2;
      end else if (10'h235 == _T_19[9:0]) begin
        image_0_565 <= io_pixelVal_in_0_1;
      end else if (10'h235 == _T_15[9:0]) begin
        image_0_565 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_566 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h236 == _T_37[9:0]) begin
        image_0_566 <= io_pixelVal_in_0_7;
      end else if (10'h236 == _T_34[9:0]) begin
        image_0_566 <= io_pixelVal_in_0_6;
      end else if (10'h236 == _T_31[9:0]) begin
        image_0_566 <= io_pixelVal_in_0_5;
      end else if (10'h236 == _T_28[9:0]) begin
        image_0_566 <= io_pixelVal_in_0_4;
      end else if (10'h236 == _T_25[9:0]) begin
        image_0_566 <= io_pixelVal_in_0_3;
      end else if (10'h236 == _T_22[9:0]) begin
        image_0_566 <= io_pixelVal_in_0_2;
      end else if (10'h236 == _T_19[9:0]) begin
        image_0_566 <= io_pixelVal_in_0_1;
      end else if (10'h236 == _T_15[9:0]) begin
        image_0_566 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_567 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h237 == _T_37[9:0]) begin
        image_0_567 <= io_pixelVal_in_0_7;
      end else if (10'h237 == _T_34[9:0]) begin
        image_0_567 <= io_pixelVal_in_0_6;
      end else if (10'h237 == _T_31[9:0]) begin
        image_0_567 <= io_pixelVal_in_0_5;
      end else if (10'h237 == _T_28[9:0]) begin
        image_0_567 <= io_pixelVal_in_0_4;
      end else if (10'h237 == _T_25[9:0]) begin
        image_0_567 <= io_pixelVal_in_0_3;
      end else if (10'h237 == _T_22[9:0]) begin
        image_0_567 <= io_pixelVal_in_0_2;
      end else if (10'h237 == _T_19[9:0]) begin
        image_0_567 <= io_pixelVal_in_0_1;
      end else if (10'h237 == _T_15[9:0]) begin
        image_0_567 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_568 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h238 == _T_37[9:0]) begin
        image_0_568 <= io_pixelVal_in_0_7;
      end else if (10'h238 == _T_34[9:0]) begin
        image_0_568 <= io_pixelVal_in_0_6;
      end else if (10'h238 == _T_31[9:0]) begin
        image_0_568 <= io_pixelVal_in_0_5;
      end else if (10'h238 == _T_28[9:0]) begin
        image_0_568 <= io_pixelVal_in_0_4;
      end else if (10'h238 == _T_25[9:0]) begin
        image_0_568 <= io_pixelVal_in_0_3;
      end else if (10'h238 == _T_22[9:0]) begin
        image_0_568 <= io_pixelVal_in_0_2;
      end else if (10'h238 == _T_19[9:0]) begin
        image_0_568 <= io_pixelVal_in_0_1;
      end else if (10'h238 == _T_15[9:0]) begin
        image_0_568 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_569 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h239 == _T_37[9:0]) begin
        image_0_569 <= io_pixelVal_in_0_7;
      end else if (10'h239 == _T_34[9:0]) begin
        image_0_569 <= io_pixelVal_in_0_6;
      end else if (10'h239 == _T_31[9:0]) begin
        image_0_569 <= io_pixelVal_in_0_5;
      end else if (10'h239 == _T_28[9:0]) begin
        image_0_569 <= io_pixelVal_in_0_4;
      end else if (10'h239 == _T_25[9:0]) begin
        image_0_569 <= io_pixelVal_in_0_3;
      end else if (10'h239 == _T_22[9:0]) begin
        image_0_569 <= io_pixelVal_in_0_2;
      end else if (10'h239 == _T_19[9:0]) begin
        image_0_569 <= io_pixelVal_in_0_1;
      end else if (10'h239 == _T_15[9:0]) begin
        image_0_569 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_570 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h23a == _T_37[9:0]) begin
        image_0_570 <= io_pixelVal_in_0_7;
      end else if (10'h23a == _T_34[9:0]) begin
        image_0_570 <= io_pixelVal_in_0_6;
      end else if (10'h23a == _T_31[9:0]) begin
        image_0_570 <= io_pixelVal_in_0_5;
      end else if (10'h23a == _T_28[9:0]) begin
        image_0_570 <= io_pixelVal_in_0_4;
      end else if (10'h23a == _T_25[9:0]) begin
        image_0_570 <= io_pixelVal_in_0_3;
      end else if (10'h23a == _T_22[9:0]) begin
        image_0_570 <= io_pixelVal_in_0_2;
      end else if (10'h23a == _T_19[9:0]) begin
        image_0_570 <= io_pixelVal_in_0_1;
      end else if (10'h23a == _T_15[9:0]) begin
        image_0_570 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_571 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h23b == _T_37[9:0]) begin
        image_0_571 <= io_pixelVal_in_0_7;
      end else if (10'h23b == _T_34[9:0]) begin
        image_0_571 <= io_pixelVal_in_0_6;
      end else if (10'h23b == _T_31[9:0]) begin
        image_0_571 <= io_pixelVal_in_0_5;
      end else if (10'h23b == _T_28[9:0]) begin
        image_0_571 <= io_pixelVal_in_0_4;
      end else if (10'h23b == _T_25[9:0]) begin
        image_0_571 <= io_pixelVal_in_0_3;
      end else if (10'h23b == _T_22[9:0]) begin
        image_0_571 <= io_pixelVal_in_0_2;
      end else if (10'h23b == _T_19[9:0]) begin
        image_0_571 <= io_pixelVal_in_0_1;
      end else if (10'h23b == _T_15[9:0]) begin
        image_0_571 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_572 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h23c == _T_37[9:0]) begin
        image_0_572 <= io_pixelVal_in_0_7;
      end else if (10'h23c == _T_34[9:0]) begin
        image_0_572 <= io_pixelVal_in_0_6;
      end else if (10'h23c == _T_31[9:0]) begin
        image_0_572 <= io_pixelVal_in_0_5;
      end else if (10'h23c == _T_28[9:0]) begin
        image_0_572 <= io_pixelVal_in_0_4;
      end else if (10'h23c == _T_25[9:0]) begin
        image_0_572 <= io_pixelVal_in_0_3;
      end else if (10'h23c == _T_22[9:0]) begin
        image_0_572 <= io_pixelVal_in_0_2;
      end else if (10'h23c == _T_19[9:0]) begin
        image_0_572 <= io_pixelVal_in_0_1;
      end else if (10'h23c == _T_15[9:0]) begin
        image_0_572 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_573 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h23d == _T_37[9:0]) begin
        image_0_573 <= io_pixelVal_in_0_7;
      end else if (10'h23d == _T_34[9:0]) begin
        image_0_573 <= io_pixelVal_in_0_6;
      end else if (10'h23d == _T_31[9:0]) begin
        image_0_573 <= io_pixelVal_in_0_5;
      end else if (10'h23d == _T_28[9:0]) begin
        image_0_573 <= io_pixelVal_in_0_4;
      end else if (10'h23d == _T_25[9:0]) begin
        image_0_573 <= io_pixelVal_in_0_3;
      end else if (10'h23d == _T_22[9:0]) begin
        image_0_573 <= io_pixelVal_in_0_2;
      end else if (10'h23d == _T_19[9:0]) begin
        image_0_573 <= io_pixelVal_in_0_1;
      end else if (10'h23d == _T_15[9:0]) begin
        image_0_573 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_574 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h23e == _T_37[9:0]) begin
        image_0_574 <= io_pixelVal_in_0_7;
      end else if (10'h23e == _T_34[9:0]) begin
        image_0_574 <= io_pixelVal_in_0_6;
      end else if (10'h23e == _T_31[9:0]) begin
        image_0_574 <= io_pixelVal_in_0_5;
      end else if (10'h23e == _T_28[9:0]) begin
        image_0_574 <= io_pixelVal_in_0_4;
      end else if (10'h23e == _T_25[9:0]) begin
        image_0_574 <= io_pixelVal_in_0_3;
      end else if (10'h23e == _T_22[9:0]) begin
        image_0_574 <= io_pixelVal_in_0_2;
      end else if (10'h23e == _T_19[9:0]) begin
        image_0_574 <= io_pixelVal_in_0_1;
      end else if (10'h23e == _T_15[9:0]) begin
        image_0_574 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_0_575 <= 4'hf;
    end else if (io_valid_in) begin
      if (10'h23f == _T_37[9:0]) begin
        image_0_575 <= io_pixelVal_in_0_7;
      end else if (10'h23f == _T_34[9:0]) begin
        image_0_575 <= io_pixelVal_in_0_6;
      end else if (10'h23f == _T_31[9:0]) begin
        image_0_575 <= io_pixelVal_in_0_5;
      end else if (10'h23f == _T_28[9:0]) begin
        image_0_575 <= io_pixelVal_in_0_4;
      end else if (10'h23f == _T_25[9:0]) begin
        image_0_575 <= io_pixelVal_in_0_3;
      end else if (10'h23f == _T_22[9:0]) begin
        image_0_575 <= io_pixelVal_in_0_2;
      end else if (10'h23f == _T_19[9:0]) begin
        image_0_575 <= io_pixelVal_in_0_1;
      end else if (10'h23f == _T_15[9:0]) begin
        image_0_575 <= io_pixelVal_in_0_0;
      end
    end
    if (reset) begin
      image_1_0 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h0 == _T_37[9:0]) begin
        image_1_0 <= io_pixelVal_in_1_7;
      end else if (10'h0 == _T_34[9:0]) begin
        image_1_0 <= io_pixelVal_in_1_6;
      end else if (10'h0 == _T_31[9:0]) begin
        image_1_0 <= io_pixelVal_in_1_5;
      end else if (10'h0 == _T_28[9:0]) begin
        image_1_0 <= io_pixelVal_in_1_4;
      end else if (10'h0 == _T_25[9:0]) begin
        image_1_0 <= io_pixelVal_in_1_3;
      end else if (10'h0 == _T_22[9:0]) begin
        image_1_0 <= io_pixelVal_in_1_2;
      end else if (10'h0 == _T_19[9:0]) begin
        image_1_0 <= io_pixelVal_in_1_1;
      end else if (10'h0 == _T_15[9:0]) begin
        image_1_0 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_1 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1 == _T_37[9:0]) begin
        image_1_1 <= io_pixelVal_in_1_7;
      end else if (10'h1 == _T_34[9:0]) begin
        image_1_1 <= io_pixelVal_in_1_6;
      end else if (10'h1 == _T_31[9:0]) begin
        image_1_1 <= io_pixelVal_in_1_5;
      end else if (10'h1 == _T_28[9:0]) begin
        image_1_1 <= io_pixelVal_in_1_4;
      end else if (10'h1 == _T_25[9:0]) begin
        image_1_1 <= io_pixelVal_in_1_3;
      end else if (10'h1 == _T_22[9:0]) begin
        image_1_1 <= io_pixelVal_in_1_2;
      end else if (10'h1 == _T_19[9:0]) begin
        image_1_1 <= io_pixelVal_in_1_1;
      end else if (10'h1 == _T_15[9:0]) begin
        image_1_1 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_2 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h2 == _T_37[9:0]) begin
        image_1_2 <= io_pixelVal_in_1_7;
      end else if (10'h2 == _T_34[9:0]) begin
        image_1_2 <= io_pixelVal_in_1_6;
      end else if (10'h2 == _T_31[9:0]) begin
        image_1_2 <= io_pixelVal_in_1_5;
      end else if (10'h2 == _T_28[9:0]) begin
        image_1_2 <= io_pixelVal_in_1_4;
      end else if (10'h2 == _T_25[9:0]) begin
        image_1_2 <= io_pixelVal_in_1_3;
      end else if (10'h2 == _T_22[9:0]) begin
        image_1_2 <= io_pixelVal_in_1_2;
      end else if (10'h2 == _T_19[9:0]) begin
        image_1_2 <= io_pixelVal_in_1_1;
      end else if (10'h2 == _T_15[9:0]) begin
        image_1_2 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_3 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h3 == _T_37[9:0]) begin
        image_1_3 <= io_pixelVal_in_1_7;
      end else if (10'h3 == _T_34[9:0]) begin
        image_1_3 <= io_pixelVal_in_1_6;
      end else if (10'h3 == _T_31[9:0]) begin
        image_1_3 <= io_pixelVal_in_1_5;
      end else if (10'h3 == _T_28[9:0]) begin
        image_1_3 <= io_pixelVal_in_1_4;
      end else if (10'h3 == _T_25[9:0]) begin
        image_1_3 <= io_pixelVal_in_1_3;
      end else if (10'h3 == _T_22[9:0]) begin
        image_1_3 <= io_pixelVal_in_1_2;
      end else if (10'h3 == _T_19[9:0]) begin
        image_1_3 <= io_pixelVal_in_1_1;
      end else if (10'h3 == _T_15[9:0]) begin
        image_1_3 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_4 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h4 == _T_37[9:0]) begin
        image_1_4 <= io_pixelVal_in_1_7;
      end else if (10'h4 == _T_34[9:0]) begin
        image_1_4 <= io_pixelVal_in_1_6;
      end else if (10'h4 == _T_31[9:0]) begin
        image_1_4 <= io_pixelVal_in_1_5;
      end else if (10'h4 == _T_28[9:0]) begin
        image_1_4 <= io_pixelVal_in_1_4;
      end else if (10'h4 == _T_25[9:0]) begin
        image_1_4 <= io_pixelVal_in_1_3;
      end else if (10'h4 == _T_22[9:0]) begin
        image_1_4 <= io_pixelVal_in_1_2;
      end else if (10'h4 == _T_19[9:0]) begin
        image_1_4 <= io_pixelVal_in_1_1;
      end else if (10'h4 == _T_15[9:0]) begin
        image_1_4 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_5 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h5 == _T_37[9:0]) begin
        image_1_5 <= io_pixelVal_in_1_7;
      end else if (10'h5 == _T_34[9:0]) begin
        image_1_5 <= io_pixelVal_in_1_6;
      end else if (10'h5 == _T_31[9:0]) begin
        image_1_5 <= io_pixelVal_in_1_5;
      end else if (10'h5 == _T_28[9:0]) begin
        image_1_5 <= io_pixelVal_in_1_4;
      end else if (10'h5 == _T_25[9:0]) begin
        image_1_5 <= io_pixelVal_in_1_3;
      end else if (10'h5 == _T_22[9:0]) begin
        image_1_5 <= io_pixelVal_in_1_2;
      end else if (10'h5 == _T_19[9:0]) begin
        image_1_5 <= io_pixelVal_in_1_1;
      end else if (10'h5 == _T_15[9:0]) begin
        image_1_5 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_6 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h6 == _T_37[9:0]) begin
        image_1_6 <= io_pixelVal_in_1_7;
      end else if (10'h6 == _T_34[9:0]) begin
        image_1_6 <= io_pixelVal_in_1_6;
      end else if (10'h6 == _T_31[9:0]) begin
        image_1_6 <= io_pixelVal_in_1_5;
      end else if (10'h6 == _T_28[9:0]) begin
        image_1_6 <= io_pixelVal_in_1_4;
      end else if (10'h6 == _T_25[9:0]) begin
        image_1_6 <= io_pixelVal_in_1_3;
      end else if (10'h6 == _T_22[9:0]) begin
        image_1_6 <= io_pixelVal_in_1_2;
      end else if (10'h6 == _T_19[9:0]) begin
        image_1_6 <= io_pixelVal_in_1_1;
      end else if (10'h6 == _T_15[9:0]) begin
        image_1_6 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_7 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h7 == _T_37[9:0]) begin
        image_1_7 <= io_pixelVal_in_1_7;
      end else if (10'h7 == _T_34[9:0]) begin
        image_1_7 <= io_pixelVal_in_1_6;
      end else if (10'h7 == _T_31[9:0]) begin
        image_1_7 <= io_pixelVal_in_1_5;
      end else if (10'h7 == _T_28[9:0]) begin
        image_1_7 <= io_pixelVal_in_1_4;
      end else if (10'h7 == _T_25[9:0]) begin
        image_1_7 <= io_pixelVal_in_1_3;
      end else if (10'h7 == _T_22[9:0]) begin
        image_1_7 <= io_pixelVal_in_1_2;
      end else if (10'h7 == _T_19[9:0]) begin
        image_1_7 <= io_pixelVal_in_1_1;
      end else if (10'h7 == _T_15[9:0]) begin
        image_1_7 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_8 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h8 == _T_37[9:0]) begin
        image_1_8 <= io_pixelVal_in_1_7;
      end else if (10'h8 == _T_34[9:0]) begin
        image_1_8 <= io_pixelVal_in_1_6;
      end else if (10'h8 == _T_31[9:0]) begin
        image_1_8 <= io_pixelVal_in_1_5;
      end else if (10'h8 == _T_28[9:0]) begin
        image_1_8 <= io_pixelVal_in_1_4;
      end else if (10'h8 == _T_25[9:0]) begin
        image_1_8 <= io_pixelVal_in_1_3;
      end else if (10'h8 == _T_22[9:0]) begin
        image_1_8 <= io_pixelVal_in_1_2;
      end else if (10'h8 == _T_19[9:0]) begin
        image_1_8 <= io_pixelVal_in_1_1;
      end else if (10'h8 == _T_15[9:0]) begin
        image_1_8 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_9 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h9 == _T_37[9:0]) begin
        image_1_9 <= io_pixelVal_in_1_7;
      end else if (10'h9 == _T_34[9:0]) begin
        image_1_9 <= io_pixelVal_in_1_6;
      end else if (10'h9 == _T_31[9:0]) begin
        image_1_9 <= io_pixelVal_in_1_5;
      end else if (10'h9 == _T_28[9:0]) begin
        image_1_9 <= io_pixelVal_in_1_4;
      end else if (10'h9 == _T_25[9:0]) begin
        image_1_9 <= io_pixelVal_in_1_3;
      end else if (10'h9 == _T_22[9:0]) begin
        image_1_9 <= io_pixelVal_in_1_2;
      end else if (10'h9 == _T_19[9:0]) begin
        image_1_9 <= io_pixelVal_in_1_1;
      end else if (10'h9 == _T_15[9:0]) begin
        image_1_9 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_10 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha == _T_37[9:0]) begin
        image_1_10 <= io_pixelVal_in_1_7;
      end else if (10'ha == _T_34[9:0]) begin
        image_1_10 <= io_pixelVal_in_1_6;
      end else if (10'ha == _T_31[9:0]) begin
        image_1_10 <= io_pixelVal_in_1_5;
      end else if (10'ha == _T_28[9:0]) begin
        image_1_10 <= io_pixelVal_in_1_4;
      end else if (10'ha == _T_25[9:0]) begin
        image_1_10 <= io_pixelVal_in_1_3;
      end else if (10'ha == _T_22[9:0]) begin
        image_1_10 <= io_pixelVal_in_1_2;
      end else if (10'ha == _T_19[9:0]) begin
        image_1_10 <= io_pixelVal_in_1_1;
      end else if (10'ha == _T_15[9:0]) begin
        image_1_10 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_11 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb == _T_37[9:0]) begin
        image_1_11 <= io_pixelVal_in_1_7;
      end else if (10'hb == _T_34[9:0]) begin
        image_1_11 <= io_pixelVal_in_1_6;
      end else if (10'hb == _T_31[9:0]) begin
        image_1_11 <= io_pixelVal_in_1_5;
      end else if (10'hb == _T_28[9:0]) begin
        image_1_11 <= io_pixelVal_in_1_4;
      end else if (10'hb == _T_25[9:0]) begin
        image_1_11 <= io_pixelVal_in_1_3;
      end else if (10'hb == _T_22[9:0]) begin
        image_1_11 <= io_pixelVal_in_1_2;
      end else if (10'hb == _T_19[9:0]) begin
        image_1_11 <= io_pixelVal_in_1_1;
      end else if (10'hb == _T_15[9:0]) begin
        image_1_11 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_12 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc == _T_37[9:0]) begin
        image_1_12 <= io_pixelVal_in_1_7;
      end else if (10'hc == _T_34[9:0]) begin
        image_1_12 <= io_pixelVal_in_1_6;
      end else if (10'hc == _T_31[9:0]) begin
        image_1_12 <= io_pixelVal_in_1_5;
      end else if (10'hc == _T_28[9:0]) begin
        image_1_12 <= io_pixelVal_in_1_4;
      end else if (10'hc == _T_25[9:0]) begin
        image_1_12 <= io_pixelVal_in_1_3;
      end else if (10'hc == _T_22[9:0]) begin
        image_1_12 <= io_pixelVal_in_1_2;
      end else if (10'hc == _T_19[9:0]) begin
        image_1_12 <= io_pixelVal_in_1_1;
      end else if (10'hc == _T_15[9:0]) begin
        image_1_12 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_13 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd == _T_37[9:0]) begin
        image_1_13 <= io_pixelVal_in_1_7;
      end else if (10'hd == _T_34[9:0]) begin
        image_1_13 <= io_pixelVal_in_1_6;
      end else if (10'hd == _T_31[9:0]) begin
        image_1_13 <= io_pixelVal_in_1_5;
      end else if (10'hd == _T_28[9:0]) begin
        image_1_13 <= io_pixelVal_in_1_4;
      end else if (10'hd == _T_25[9:0]) begin
        image_1_13 <= io_pixelVal_in_1_3;
      end else if (10'hd == _T_22[9:0]) begin
        image_1_13 <= io_pixelVal_in_1_2;
      end else if (10'hd == _T_19[9:0]) begin
        image_1_13 <= io_pixelVal_in_1_1;
      end else if (10'hd == _T_15[9:0]) begin
        image_1_13 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_14 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he == _T_37[9:0]) begin
        image_1_14 <= io_pixelVal_in_1_7;
      end else if (10'he == _T_34[9:0]) begin
        image_1_14 <= io_pixelVal_in_1_6;
      end else if (10'he == _T_31[9:0]) begin
        image_1_14 <= io_pixelVal_in_1_5;
      end else if (10'he == _T_28[9:0]) begin
        image_1_14 <= io_pixelVal_in_1_4;
      end else if (10'he == _T_25[9:0]) begin
        image_1_14 <= io_pixelVal_in_1_3;
      end else if (10'he == _T_22[9:0]) begin
        image_1_14 <= io_pixelVal_in_1_2;
      end else if (10'he == _T_19[9:0]) begin
        image_1_14 <= io_pixelVal_in_1_1;
      end else if (10'he == _T_15[9:0]) begin
        image_1_14 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_15 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf == _T_37[9:0]) begin
        image_1_15 <= io_pixelVal_in_1_7;
      end else if (10'hf == _T_34[9:0]) begin
        image_1_15 <= io_pixelVal_in_1_6;
      end else if (10'hf == _T_31[9:0]) begin
        image_1_15 <= io_pixelVal_in_1_5;
      end else if (10'hf == _T_28[9:0]) begin
        image_1_15 <= io_pixelVal_in_1_4;
      end else if (10'hf == _T_25[9:0]) begin
        image_1_15 <= io_pixelVal_in_1_3;
      end else if (10'hf == _T_22[9:0]) begin
        image_1_15 <= io_pixelVal_in_1_2;
      end else if (10'hf == _T_19[9:0]) begin
        image_1_15 <= io_pixelVal_in_1_1;
      end else if (10'hf == _T_15[9:0]) begin
        image_1_15 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_16 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h10 == _T_37[9:0]) begin
        image_1_16 <= io_pixelVal_in_1_7;
      end else if (10'h10 == _T_34[9:0]) begin
        image_1_16 <= io_pixelVal_in_1_6;
      end else if (10'h10 == _T_31[9:0]) begin
        image_1_16 <= io_pixelVal_in_1_5;
      end else if (10'h10 == _T_28[9:0]) begin
        image_1_16 <= io_pixelVal_in_1_4;
      end else if (10'h10 == _T_25[9:0]) begin
        image_1_16 <= io_pixelVal_in_1_3;
      end else if (10'h10 == _T_22[9:0]) begin
        image_1_16 <= io_pixelVal_in_1_2;
      end else if (10'h10 == _T_19[9:0]) begin
        image_1_16 <= io_pixelVal_in_1_1;
      end else if (10'h10 == _T_15[9:0]) begin
        image_1_16 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_17 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h11 == _T_37[9:0]) begin
        image_1_17 <= io_pixelVal_in_1_7;
      end else if (10'h11 == _T_34[9:0]) begin
        image_1_17 <= io_pixelVal_in_1_6;
      end else if (10'h11 == _T_31[9:0]) begin
        image_1_17 <= io_pixelVal_in_1_5;
      end else if (10'h11 == _T_28[9:0]) begin
        image_1_17 <= io_pixelVal_in_1_4;
      end else if (10'h11 == _T_25[9:0]) begin
        image_1_17 <= io_pixelVal_in_1_3;
      end else if (10'h11 == _T_22[9:0]) begin
        image_1_17 <= io_pixelVal_in_1_2;
      end else if (10'h11 == _T_19[9:0]) begin
        image_1_17 <= io_pixelVal_in_1_1;
      end else if (10'h11 == _T_15[9:0]) begin
        image_1_17 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_18 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h12 == _T_37[9:0]) begin
        image_1_18 <= io_pixelVal_in_1_7;
      end else if (10'h12 == _T_34[9:0]) begin
        image_1_18 <= io_pixelVal_in_1_6;
      end else if (10'h12 == _T_31[9:0]) begin
        image_1_18 <= io_pixelVal_in_1_5;
      end else if (10'h12 == _T_28[9:0]) begin
        image_1_18 <= io_pixelVal_in_1_4;
      end else if (10'h12 == _T_25[9:0]) begin
        image_1_18 <= io_pixelVal_in_1_3;
      end else if (10'h12 == _T_22[9:0]) begin
        image_1_18 <= io_pixelVal_in_1_2;
      end else if (10'h12 == _T_19[9:0]) begin
        image_1_18 <= io_pixelVal_in_1_1;
      end else if (10'h12 == _T_15[9:0]) begin
        image_1_18 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_19 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h13 == _T_37[9:0]) begin
        image_1_19 <= io_pixelVal_in_1_7;
      end else if (10'h13 == _T_34[9:0]) begin
        image_1_19 <= io_pixelVal_in_1_6;
      end else if (10'h13 == _T_31[9:0]) begin
        image_1_19 <= io_pixelVal_in_1_5;
      end else if (10'h13 == _T_28[9:0]) begin
        image_1_19 <= io_pixelVal_in_1_4;
      end else if (10'h13 == _T_25[9:0]) begin
        image_1_19 <= io_pixelVal_in_1_3;
      end else if (10'h13 == _T_22[9:0]) begin
        image_1_19 <= io_pixelVal_in_1_2;
      end else if (10'h13 == _T_19[9:0]) begin
        image_1_19 <= io_pixelVal_in_1_1;
      end else if (10'h13 == _T_15[9:0]) begin
        image_1_19 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_20 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h14 == _T_37[9:0]) begin
        image_1_20 <= io_pixelVal_in_1_7;
      end else if (10'h14 == _T_34[9:0]) begin
        image_1_20 <= io_pixelVal_in_1_6;
      end else if (10'h14 == _T_31[9:0]) begin
        image_1_20 <= io_pixelVal_in_1_5;
      end else if (10'h14 == _T_28[9:0]) begin
        image_1_20 <= io_pixelVal_in_1_4;
      end else if (10'h14 == _T_25[9:0]) begin
        image_1_20 <= io_pixelVal_in_1_3;
      end else if (10'h14 == _T_22[9:0]) begin
        image_1_20 <= io_pixelVal_in_1_2;
      end else if (10'h14 == _T_19[9:0]) begin
        image_1_20 <= io_pixelVal_in_1_1;
      end else if (10'h14 == _T_15[9:0]) begin
        image_1_20 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_21 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h15 == _T_37[9:0]) begin
        image_1_21 <= io_pixelVal_in_1_7;
      end else if (10'h15 == _T_34[9:0]) begin
        image_1_21 <= io_pixelVal_in_1_6;
      end else if (10'h15 == _T_31[9:0]) begin
        image_1_21 <= io_pixelVal_in_1_5;
      end else if (10'h15 == _T_28[9:0]) begin
        image_1_21 <= io_pixelVal_in_1_4;
      end else if (10'h15 == _T_25[9:0]) begin
        image_1_21 <= io_pixelVal_in_1_3;
      end else if (10'h15 == _T_22[9:0]) begin
        image_1_21 <= io_pixelVal_in_1_2;
      end else if (10'h15 == _T_19[9:0]) begin
        image_1_21 <= io_pixelVal_in_1_1;
      end else if (10'h15 == _T_15[9:0]) begin
        image_1_21 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_22 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h16 == _T_37[9:0]) begin
        image_1_22 <= io_pixelVal_in_1_7;
      end else if (10'h16 == _T_34[9:0]) begin
        image_1_22 <= io_pixelVal_in_1_6;
      end else if (10'h16 == _T_31[9:0]) begin
        image_1_22 <= io_pixelVal_in_1_5;
      end else if (10'h16 == _T_28[9:0]) begin
        image_1_22 <= io_pixelVal_in_1_4;
      end else if (10'h16 == _T_25[9:0]) begin
        image_1_22 <= io_pixelVal_in_1_3;
      end else if (10'h16 == _T_22[9:0]) begin
        image_1_22 <= io_pixelVal_in_1_2;
      end else if (10'h16 == _T_19[9:0]) begin
        image_1_22 <= io_pixelVal_in_1_1;
      end else if (10'h16 == _T_15[9:0]) begin
        image_1_22 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_23 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h17 == _T_37[9:0]) begin
        image_1_23 <= io_pixelVal_in_1_7;
      end else if (10'h17 == _T_34[9:0]) begin
        image_1_23 <= io_pixelVal_in_1_6;
      end else if (10'h17 == _T_31[9:0]) begin
        image_1_23 <= io_pixelVal_in_1_5;
      end else if (10'h17 == _T_28[9:0]) begin
        image_1_23 <= io_pixelVal_in_1_4;
      end else if (10'h17 == _T_25[9:0]) begin
        image_1_23 <= io_pixelVal_in_1_3;
      end else if (10'h17 == _T_22[9:0]) begin
        image_1_23 <= io_pixelVal_in_1_2;
      end else if (10'h17 == _T_19[9:0]) begin
        image_1_23 <= io_pixelVal_in_1_1;
      end else if (10'h17 == _T_15[9:0]) begin
        image_1_23 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_24 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h18 == _T_37[9:0]) begin
        image_1_24 <= io_pixelVal_in_1_7;
      end else if (10'h18 == _T_34[9:0]) begin
        image_1_24 <= io_pixelVal_in_1_6;
      end else if (10'h18 == _T_31[9:0]) begin
        image_1_24 <= io_pixelVal_in_1_5;
      end else if (10'h18 == _T_28[9:0]) begin
        image_1_24 <= io_pixelVal_in_1_4;
      end else if (10'h18 == _T_25[9:0]) begin
        image_1_24 <= io_pixelVal_in_1_3;
      end else if (10'h18 == _T_22[9:0]) begin
        image_1_24 <= io_pixelVal_in_1_2;
      end else if (10'h18 == _T_19[9:0]) begin
        image_1_24 <= io_pixelVal_in_1_1;
      end else if (10'h18 == _T_15[9:0]) begin
        image_1_24 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_25 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h19 == _T_37[9:0]) begin
        image_1_25 <= io_pixelVal_in_1_7;
      end else if (10'h19 == _T_34[9:0]) begin
        image_1_25 <= io_pixelVal_in_1_6;
      end else if (10'h19 == _T_31[9:0]) begin
        image_1_25 <= io_pixelVal_in_1_5;
      end else if (10'h19 == _T_28[9:0]) begin
        image_1_25 <= io_pixelVal_in_1_4;
      end else if (10'h19 == _T_25[9:0]) begin
        image_1_25 <= io_pixelVal_in_1_3;
      end else if (10'h19 == _T_22[9:0]) begin
        image_1_25 <= io_pixelVal_in_1_2;
      end else if (10'h19 == _T_19[9:0]) begin
        image_1_25 <= io_pixelVal_in_1_1;
      end else if (10'h19 == _T_15[9:0]) begin
        image_1_25 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_26 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a == _T_37[9:0]) begin
        image_1_26 <= io_pixelVal_in_1_7;
      end else if (10'h1a == _T_34[9:0]) begin
        image_1_26 <= io_pixelVal_in_1_6;
      end else if (10'h1a == _T_31[9:0]) begin
        image_1_26 <= io_pixelVal_in_1_5;
      end else if (10'h1a == _T_28[9:0]) begin
        image_1_26 <= io_pixelVal_in_1_4;
      end else if (10'h1a == _T_25[9:0]) begin
        image_1_26 <= io_pixelVal_in_1_3;
      end else if (10'h1a == _T_22[9:0]) begin
        image_1_26 <= io_pixelVal_in_1_2;
      end else if (10'h1a == _T_19[9:0]) begin
        image_1_26 <= io_pixelVal_in_1_1;
      end else if (10'h1a == _T_15[9:0]) begin
        image_1_26 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_27 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b == _T_37[9:0]) begin
        image_1_27 <= io_pixelVal_in_1_7;
      end else if (10'h1b == _T_34[9:0]) begin
        image_1_27 <= io_pixelVal_in_1_6;
      end else if (10'h1b == _T_31[9:0]) begin
        image_1_27 <= io_pixelVal_in_1_5;
      end else if (10'h1b == _T_28[9:0]) begin
        image_1_27 <= io_pixelVal_in_1_4;
      end else if (10'h1b == _T_25[9:0]) begin
        image_1_27 <= io_pixelVal_in_1_3;
      end else if (10'h1b == _T_22[9:0]) begin
        image_1_27 <= io_pixelVal_in_1_2;
      end else if (10'h1b == _T_19[9:0]) begin
        image_1_27 <= io_pixelVal_in_1_1;
      end else if (10'h1b == _T_15[9:0]) begin
        image_1_27 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_28 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c == _T_37[9:0]) begin
        image_1_28 <= io_pixelVal_in_1_7;
      end else if (10'h1c == _T_34[9:0]) begin
        image_1_28 <= io_pixelVal_in_1_6;
      end else if (10'h1c == _T_31[9:0]) begin
        image_1_28 <= io_pixelVal_in_1_5;
      end else if (10'h1c == _T_28[9:0]) begin
        image_1_28 <= io_pixelVal_in_1_4;
      end else if (10'h1c == _T_25[9:0]) begin
        image_1_28 <= io_pixelVal_in_1_3;
      end else if (10'h1c == _T_22[9:0]) begin
        image_1_28 <= io_pixelVal_in_1_2;
      end else if (10'h1c == _T_19[9:0]) begin
        image_1_28 <= io_pixelVal_in_1_1;
      end else if (10'h1c == _T_15[9:0]) begin
        image_1_28 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_29 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d == _T_37[9:0]) begin
        image_1_29 <= io_pixelVal_in_1_7;
      end else if (10'h1d == _T_34[9:0]) begin
        image_1_29 <= io_pixelVal_in_1_6;
      end else if (10'h1d == _T_31[9:0]) begin
        image_1_29 <= io_pixelVal_in_1_5;
      end else if (10'h1d == _T_28[9:0]) begin
        image_1_29 <= io_pixelVal_in_1_4;
      end else if (10'h1d == _T_25[9:0]) begin
        image_1_29 <= io_pixelVal_in_1_3;
      end else if (10'h1d == _T_22[9:0]) begin
        image_1_29 <= io_pixelVal_in_1_2;
      end else if (10'h1d == _T_19[9:0]) begin
        image_1_29 <= io_pixelVal_in_1_1;
      end else if (10'h1d == _T_15[9:0]) begin
        image_1_29 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_30 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e == _T_37[9:0]) begin
        image_1_30 <= io_pixelVal_in_1_7;
      end else if (10'h1e == _T_34[9:0]) begin
        image_1_30 <= io_pixelVal_in_1_6;
      end else if (10'h1e == _T_31[9:0]) begin
        image_1_30 <= io_pixelVal_in_1_5;
      end else if (10'h1e == _T_28[9:0]) begin
        image_1_30 <= io_pixelVal_in_1_4;
      end else if (10'h1e == _T_25[9:0]) begin
        image_1_30 <= io_pixelVal_in_1_3;
      end else if (10'h1e == _T_22[9:0]) begin
        image_1_30 <= io_pixelVal_in_1_2;
      end else if (10'h1e == _T_19[9:0]) begin
        image_1_30 <= io_pixelVal_in_1_1;
      end else if (10'h1e == _T_15[9:0]) begin
        image_1_30 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_31 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f == _T_37[9:0]) begin
        image_1_31 <= io_pixelVal_in_1_7;
      end else if (10'h1f == _T_34[9:0]) begin
        image_1_31 <= io_pixelVal_in_1_6;
      end else if (10'h1f == _T_31[9:0]) begin
        image_1_31 <= io_pixelVal_in_1_5;
      end else if (10'h1f == _T_28[9:0]) begin
        image_1_31 <= io_pixelVal_in_1_4;
      end else if (10'h1f == _T_25[9:0]) begin
        image_1_31 <= io_pixelVal_in_1_3;
      end else if (10'h1f == _T_22[9:0]) begin
        image_1_31 <= io_pixelVal_in_1_2;
      end else if (10'h1f == _T_19[9:0]) begin
        image_1_31 <= io_pixelVal_in_1_1;
      end else if (10'h1f == _T_15[9:0]) begin
        image_1_31 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_32 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h20 == _T_37[9:0]) begin
        image_1_32 <= io_pixelVal_in_1_7;
      end else if (10'h20 == _T_34[9:0]) begin
        image_1_32 <= io_pixelVal_in_1_6;
      end else if (10'h20 == _T_31[9:0]) begin
        image_1_32 <= io_pixelVal_in_1_5;
      end else if (10'h20 == _T_28[9:0]) begin
        image_1_32 <= io_pixelVal_in_1_4;
      end else if (10'h20 == _T_25[9:0]) begin
        image_1_32 <= io_pixelVal_in_1_3;
      end else if (10'h20 == _T_22[9:0]) begin
        image_1_32 <= io_pixelVal_in_1_2;
      end else if (10'h20 == _T_19[9:0]) begin
        image_1_32 <= io_pixelVal_in_1_1;
      end else if (10'h20 == _T_15[9:0]) begin
        image_1_32 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_33 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h21 == _T_37[9:0]) begin
        image_1_33 <= io_pixelVal_in_1_7;
      end else if (10'h21 == _T_34[9:0]) begin
        image_1_33 <= io_pixelVal_in_1_6;
      end else if (10'h21 == _T_31[9:0]) begin
        image_1_33 <= io_pixelVal_in_1_5;
      end else if (10'h21 == _T_28[9:0]) begin
        image_1_33 <= io_pixelVal_in_1_4;
      end else if (10'h21 == _T_25[9:0]) begin
        image_1_33 <= io_pixelVal_in_1_3;
      end else if (10'h21 == _T_22[9:0]) begin
        image_1_33 <= io_pixelVal_in_1_2;
      end else if (10'h21 == _T_19[9:0]) begin
        image_1_33 <= io_pixelVal_in_1_1;
      end else if (10'h21 == _T_15[9:0]) begin
        image_1_33 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_34 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h22 == _T_37[9:0]) begin
        image_1_34 <= io_pixelVal_in_1_7;
      end else if (10'h22 == _T_34[9:0]) begin
        image_1_34 <= io_pixelVal_in_1_6;
      end else if (10'h22 == _T_31[9:0]) begin
        image_1_34 <= io_pixelVal_in_1_5;
      end else if (10'h22 == _T_28[9:0]) begin
        image_1_34 <= io_pixelVal_in_1_4;
      end else if (10'h22 == _T_25[9:0]) begin
        image_1_34 <= io_pixelVal_in_1_3;
      end else if (10'h22 == _T_22[9:0]) begin
        image_1_34 <= io_pixelVal_in_1_2;
      end else if (10'h22 == _T_19[9:0]) begin
        image_1_34 <= io_pixelVal_in_1_1;
      end else if (10'h22 == _T_15[9:0]) begin
        image_1_34 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_35 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h23 == _T_37[9:0]) begin
        image_1_35 <= io_pixelVal_in_1_7;
      end else if (10'h23 == _T_34[9:0]) begin
        image_1_35 <= io_pixelVal_in_1_6;
      end else if (10'h23 == _T_31[9:0]) begin
        image_1_35 <= io_pixelVal_in_1_5;
      end else if (10'h23 == _T_28[9:0]) begin
        image_1_35 <= io_pixelVal_in_1_4;
      end else if (10'h23 == _T_25[9:0]) begin
        image_1_35 <= io_pixelVal_in_1_3;
      end else if (10'h23 == _T_22[9:0]) begin
        image_1_35 <= io_pixelVal_in_1_2;
      end else if (10'h23 == _T_19[9:0]) begin
        image_1_35 <= io_pixelVal_in_1_1;
      end else if (10'h23 == _T_15[9:0]) begin
        image_1_35 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_36 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h24 == _T_37[9:0]) begin
        image_1_36 <= io_pixelVal_in_1_7;
      end else if (10'h24 == _T_34[9:0]) begin
        image_1_36 <= io_pixelVal_in_1_6;
      end else if (10'h24 == _T_31[9:0]) begin
        image_1_36 <= io_pixelVal_in_1_5;
      end else if (10'h24 == _T_28[9:0]) begin
        image_1_36 <= io_pixelVal_in_1_4;
      end else if (10'h24 == _T_25[9:0]) begin
        image_1_36 <= io_pixelVal_in_1_3;
      end else if (10'h24 == _T_22[9:0]) begin
        image_1_36 <= io_pixelVal_in_1_2;
      end else if (10'h24 == _T_19[9:0]) begin
        image_1_36 <= io_pixelVal_in_1_1;
      end else if (10'h24 == _T_15[9:0]) begin
        image_1_36 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_37 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h25 == _T_37[9:0]) begin
        image_1_37 <= io_pixelVal_in_1_7;
      end else if (10'h25 == _T_34[9:0]) begin
        image_1_37 <= io_pixelVal_in_1_6;
      end else if (10'h25 == _T_31[9:0]) begin
        image_1_37 <= io_pixelVal_in_1_5;
      end else if (10'h25 == _T_28[9:0]) begin
        image_1_37 <= io_pixelVal_in_1_4;
      end else if (10'h25 == _T_25[9:0]) begin
        image_1_37 <= io_pixelVal_in_1_3;
      end else if (10'h25 == _T_22[9:0]) begin
        image_1_37 <= io_pixelVal_in_1_2;
      end else if (10'h25 == _T_19[9:0]) begin
        image_1_37 <= io_pixelVal_in_1_1;
      end else if (10'h25 == _T_15[9:0]) begin
        image_1_37 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_38 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h26 == _T_37[9:0]) begin
        image_1_38 <= io_pixelVal_in_1_7;
      end else if (10'h26 == _T_34[9:0]) begin
        image_1_38 <= io_pixelVal_in_1_6;
      end else if (10'h26 == _T_31[9:0]) begin
        image_1_38 <= io_pixelVal_in_1_5;
      end else if (10'h26 == _T_28[9:0]) begin
        image_1_38 <= io_pixelVal_in_1_4;
      end else if (10'h26 == _T_25[9:0]) begin
        image_1_38 <= io_pixelVal_in_1_3;
      end else if (10'h26 == _T_22[9:0]) begin
        image_1_38 <= io_pixelVal_in_1_2;
      end else if (10'h26 == _T_19[9:0]) begin
        image_1_38 <= io_pixelVal_in_1_1;
      end else if (10'h26 == _T_15[9:0]) begin
        image_1_38 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_39 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h27 == _T_37[9:0]) begin
        image_1_39 <= io_pixelVal_in_1_7;
      end else if (10'h27 == _T_34[9:0]) begin
        image_1_39 <= io_pixelVal_in_1_6;
      end else if (10'h27 == _T_31[9:0]) begin
        image_1_39 <= io_pixelVal_in_1_5;
      end else if (10'h27 == _T_28[9:0]) begin
        image_1_39 <= io_pixelVal_in_1_4;
      end else if (10'h27 == _T_25[9:0]) begin
        image_1_39 <= io_pixelVal_in_1_3;
      end else if (10'h27 == _T_22[9:0]) begin
        image_1_39 <= io_pixelVal_in_1_2;
      end else if (10'h27 == _T_19[9:0]) begin
        image_1_39 <= io_pixelVal_in_1_1;
      end else if (10'h27 == _T_15[9:0]) begin
        image_1_39 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_40 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h28 == _T_37[9:0]) begin
        image_1_40 <= io_pixelVal_in_1_7;
      end else if (10'h28 == _T_34[9:0]) begin
        image_1_40 <= io_pixelVal_in_1_6;
      end else if (10'h28 == _T_31[9:0]) begin
        image_1_40 <= io_pixelVal_in_1_5;
      end else if (10'h28 == _T_28[9:0]) begin
        image_1_40 <= io_pixelVal_in_1_4;
      end else if (10'h28 == _T_25[9:0]) begin
        image_1_40 <= io_pixelVal_in_1_3;
      end else if (10'h28 == _T_22[9:0]) begin
        image_1_40 <= io_pixelVal_in_1_2;
      end else if (10'h28 == _T_19[9:0]) begin
        image_1_40 <= io_pixelVal_in_1_1;
      end else if (10'h28 == _T_15[9:0]) begin
        image_1_40 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_41 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h29 == _T_37[9:0]) begin
        image_1_41 <= io_pixelVal_in_1_7;
      end else if (10'h29 == _T_34[9:0]) begin
        image_1_41 <= io_pixelVal_in_1_6;
      end else if (10'h29 == _T_31[9:0]) begin
        image_1_41 <= io_pixelVal_in_1_5;
      end else if (10'h29 == _T_28[9:0]) begin
        image_1_41 <= io_pixelVal_in_1_4;
      end else if (10'h29 == _T_25[9:0]) begin
        image_1_41 <= io_pixelVal_in_1_3;
      end else if (10'h29 == _T_22[9:0]) begin
        image_1_41 <= io_pixelVal_in_1_2;
      end else if (10'h29 == _T_19[9:0]) begin
        image_1_41 <= io_pixelVal_in_1_1;
      end else if (10'h29 == _T_15[9:0]) begin
        image_1_41 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_42 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h2a == _T_37[9:0]) begin
        image_1_42 <= io_pixelVal_in_1_7;
      end else if (10'h2a == _T_34[9:0]) begin
        image_1_42 <= io_pixelVal_in_1_6;
      end else if (10'h2a == _T_31[9:0]) begin
        image_1_42 <= io_pixelVal_in_1_5;
      end else if (10'h2a == _T_28[9:0]) begin
        image_1_42 <= io_pixelVal_in_1_4;
      end else if (10'h2a == _T_25[9:0]) begin
        image_1_42 <= io_pixelVal_in_1_3;
      end else if (10'h2a == _T_22[9:0]) begin
        image_1_42 <= io_pixelVal_in_1_2;
      end else if (10'h2a == _T_19[9:0]) begin
        image_1_42 <= io_pixelVal_in_1_1;
      end else if (10'h2a == _T_15[9:0]) begin
        image_1_42 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_43 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h2b == _T_37[9:0]) begin
        image_1_43 <= io_pixelVal_in_1_7;
      end else if (10'h2b == _T_34[9:0]) begin
        image_1_43 <= io_pixelVal_in_1_6;
      end else if (10'h2b == _T_31[9:0]) begin
        image_1_43 <= io_pixelVal_in_1_5;
      end else if (10'h2b == _T_28[9:0]) begin
        image_1_43 <= io_pixelVal_in_1_4;
      end else if (10'h2b == _T_25[9:0]) begin
        image_1_43 <= io_pixelVal_in_1_3;
      end else if (10'h2b == _T_22[9:0]) begin
        image_1_43 <= io_pixelVal_in_1_2;
      end else if (10'h2b == _T_19[9:0]) begin
        image_1_43 <= io_pixelVal_in_1_1;
      end else if (10'h2b == _T_15[9:0]) begin
        image_1_43 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_44 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h2c == _T_37[9:0]) begin
        image_1_44 <= io_pixelVal_in_1_7;
      end else if (10'h2c == _T_34[9:0]) begin
        image_1_44 <= io_pixelVal_in_1_6;
      end else if (10'h2c == _T_31[9:0]) begin
        image_1_44 <= io_pixelVal_in_1_5;
      end else if (10'h2c == _T_28[9:0]) begin
        image_1_44 <= io_pixelVal_in_1_4;
      end else if (10'h2c == _T_25[9:0]) begin
        image_1_44 <= io_pixelVal_in_1_3;
      end else if (10'h2c == _T_22[9:0]) begin
        image_1_44 <= io_pixelVal_in_1_2;
      end else if (10'h2c == _T_19[9:0]) begin
        image_1_44 <= io_pixelVal_in_1_1;
      end else if (10'h2c == _T_15[9:0]) begin
        image_1_44 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_45 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h2d == _T_37[9:0]) begin
        image_1_45 <= io_pixelVal_in_1_7;
      end else if (10'h2d == _T_34[9:0]) begin
        image_1_45 <= io_pixelVal_in_1_6;
      end else if (10'h2d == _T_31[9:0]) begin
        image_1_45 <= io_pixelVal_in_1_5;
      end else if (10'h2d == _T_28[9:0]) begin
        image_1_45 <= io_pixelVal_in_1_4;
      end else if (10'h2d == _T_25[9:0]) begin
        image_1_45 <= io_pixelVal_in_1_3;
      end else if (10'h2d == _T_22[9:0]) begin
        image_1_45 <= io_pixelVal_in_1_2;
      end else if (10'h2d == _T_19[9:0]) begin
        image_1_45 <= io_pixelVal_in_1_1;
      end else if (10'h2d == _T_15[9:0]) begin
        image_1_45 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_46 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h2e == _T_37[9:0]) begin
        image_1_46 <= io_pixelVal_in_1_7;
      end else if (10'h2e == _T_34[9:0]) begin
        image_1_46 <= io_pixelVal_in_1_6;
      end else if (10'h2e == _T_31[9:0]) begin
        image_1_46 <= io_pixelVal_in_1_5;
      end else if (10'h2e == _T_28[9:0]) begin
        image_1_46 <= io_pixelVal_in_1_4;
      end else if (10'h2e == _T_25[9:0]) begin
        image_1_46 <= io_pixelVal_in_1_3;
      end else if (10'h2e == _T_22[9:0]) begin
        image_1_46 <= io_pixelVal_in_1_2;
      end else if (10'h2e == _T_19[9:0]) begin
        image_1_46 <= io_pixelVal_in_1_1;
      end else if (10'h2e == _T_15[9:0]) begin
        image_1_46 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_47 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h2f == _T_37[9:0]) begin
        image_1_47 <= io_pixelVal_in_1_7;
      end else if (10'h2f == _T_34[9:0]) begin
        image_1_47 <= io_pixelVal_in_1_6;
      end else if (10'h2f == _T_31[9:0]) begin
        image_1_47 <= io_pixelVal_in_1_5;
      end else if (10'h2f == _T_28[9:0]) begin
        image_1_47 <= io_pixelVal_in_1_4;
      end else if (10'h2f == _T_25[9:0]) begin
        image_1_47 <= io_pixelVal_in_1_3;
      end else if (10'h2f == _T_22[9:0]) begin
        image_1_47 <= io_pixelVal_in_1_2;
      end else if (10'h2f == _T_19[9:0]) begin
        image_1_47 <= io_pixelVal_in_1_1;
      end else if (10'h2f == _T_15[9:0]) begin
        image_1_47 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_48 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h30 == _T_37[9:0]) begin
        image_1_48 <= io_pixelVal_in_1_7;
      end else if (10'h30 == _T_34[9:0]) begin
        image_1_48 <= io_pixelVal_in_1_6;
      end else if (10'h30 == _T_31[9:0]) begin
        image_1_48 <= io_pixelVal_in_1_5;
      end else if (10'h30 == _T_28[9:0]) begin
        image_1_48 <= io_pixelVal_in_1_4;
      end else if (10'h30 == _T_25[9:0]) begin
        image_1_48 <= io_pixelVal_in_1_3;
      end else if (10'h30 == _T_22[9:0]) begin
        image_1_48 <= io_pixelVal_in_1_2;
      end else if (10'h30 == _T_19[9:0]) begin
        image_1_48 <= io_pixelVal_in_1_1;
      end else if (10'h30 == _T_15[9:0]) begin
        image_1_48 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_49 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h31 == _T_37[9:0]) begin
        image_1_49 <= io_pixelVal_in_1_7;
      end else if (10'h31 == _T_34[9:0]) begin
        image_1_49 <= io_pixelVal_in_1_6;
      end else if (10'h31 == _T_31[9:0]) begin
        image_1_49 <= io_pixelVal_in_1_5;
      end else if (10'h31 == _T_28[9:0]) begin
        image_1_49 <= io_pixelVal_in_1_4;
      end else if (10'h31 == _T_25[9:0]) begin
        image_1_49 <= io_pixelVal_in_1_3;
      end else if (10'h31 == _T_22[9:0]) begin
        image_1_49 <= io_pixelVal_in_1_2;
      end else if (10'h31 == _T_19[9:0]) begin
        image_1_49 <= io_pixelVal_in_1_1;
      end else if (10'h31 == _T_15[9:0]) begin
        image_1_49 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_50 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h32 == _T_37[9:0]) begin
        image_1_50 <= io_pixelVal_in_1_7;
      end else if (10'h32 == _T_34[9:0]) begin
        image_1_50 <= io_pixelVal_in_1_6;
      end else if (10'h32 == _T_31[9:0]) begin
        image_1_50 <= io_pixelVal_in_1_5;
      end else if (10'h32 == _T_28[9:0]) begin
        image_1_50 <= io_pixelVal_in_1_4;
      end else if (10'h32 == _T_25[9:0]) begin
        image_1_50 <= io_pixelVal_in_1_3;
      end else if (10'h32 == _T_22[9:0]) begin
        image_1_50 <= io_pixelVal_in_1_2;
      end else if (10'h32 == _T_19[9:0]) begin
        image_1_50 <= io_pixelVal_in_1_1;
      end else if (10'h32 == _T_15[9:0]) begin
        image_1_50 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_51 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h33 == _T_37[9:0]) begin
        image_1_51 <= io_pixelVal_in_1_7;
      end else if (10'h33 == _T_34[9:0]) begin
        image_1_51 <= io_pixelVal_in_1_6;
      end else if (10'h33 == _T_31[9:0]) begin
        image_1_51 <= io_pixelVal_in_1_5;
      end else if (10'h33 == _T_28[9:0]) begin
        image_1_51 <= io_pixelVal_in_1_4;
      end else if (10'h33 == _T_25[9:0]) begin
        image_1_51 <= io_pixelVal_in_1_3;
      end else if (10'h33 == _T_22[9:0]) begin
        image_1_51 <= io_pixelVal_in_1_2;
      end else if (10'h33 == _T_19[9:0]) begin
        image_1_51 <= io_pixelVal_in_1_1;
      end else if (10'h33 == _T_15[9:0]) begin
        image_1_51 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_52 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h34 == _T_37[9:0]) begin
        image_1_52 <= io_pixelVal_in_1_7;
      end else if (10'h34 == _T_34[9:0]) begin
        image_1_52 <= io_pixelVal_in_1_6;
      end else if (10'h34 == _T_31[9:0]) begin
        image_1_52 <= io_pixelVal_in_1_5;
      end else if (10'h34 == _T_28[9:0]) begin
        image_1_52 <= io_pixelVal_in_1_4;
      end else if (10'h34 == _T_25[9:0]) begin
        image_1_52 <= io_pixelVal_in_1_3;
      end else if (10'h34 == _T_22[9:0]) begin
        image_1_52 <= io_pixelVal_in_1_2;
      end else if (10'h34 == _T_19[9:0]) begin
        image_1_52 <= io_pixelVal_in_1_1;
      end else if (10'h34 == _T_15[9:0]) begin
        image_1_52 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_53 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h35 == _T_37[9:0]) begin
        image_1_53 <= io_pixelVal_in_1_7;
      end else if (10'h35 == _T_34[9:0]) begin
        image_1_53 <= io_pixelVal_in_1_6;
      end else if (10'h35 == _T_31[9:0]) begin
        image_1_53 <= io_pixelVal_in_1_5;
      end else if (10'h35 == _T_28[9:0]) begin
        image_1_53 <= io_pixelVal_in_1_4;
      end else if (10'h35 == _T_25[9:0]) begin
        image_1_53 <= io_pixelVal_in_1_3;
      end else if (10'h35 == _T_22[9:0]) begin
        image_1_53 <= io_pixelVal_in_1_2;
      end else if (10'h35 == _T_19[9:0]) begin
        image_1_53 <= io_pixelVal_in_1_1;
      end else if (10'h35 == _T_15[9:0]) begin
        image_1_53 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_54 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h36 == _T_37[9:0]) begin
        image_1_54 <= io_pixelVal_in_1_7;
      end else if (10'h36 == _T_34[9:0]) begin
        image_1_54 <= io_pixelVal_in_1_6;
      end else if (10'h36 == _T_31[9:0]) begin
        image_1_54 <= io_pixelVal_in_1_5;
      end else if (10'h36 == _T_28[9:0]) begin
        image_1_54 <= io_pixelVal_in_1_4;
      end else if (10'h36 == _T_25[9:0]) begin
        image_1_54 <= io_pixelVal_in_1_3;
      end else if (10'h36 == _T_22[9:0]) begin
        image_1_54 <= io_pixelVal_in_1_2;
      end else if (10'h36 == _T_19[9:0]) begin
        image_1_54 <= io_pixelVal_in_1_1;
      end else if (10'h36 == _T_15[9:0]) begin
        image_1_54 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_55 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h37 == _T_37[9:0]) begin
        image_1_55 <= io_pixelVal_in_1_7;
      end else if (10'h37 == _T_34[9:0]) begin
        image_1_55 <= io_pixelVal_in_1_6;
      end else if (10'h37 == _T_31[9:0]) begin
        image_1_55 <= io_pixelVal_in_1_5;
      end else if (10'h37 == _T_28[9:0]) begin
        image_1_55 <= io_pixelVal_in_1_4;
      end else if (10'h37 == _T_25[9:0]) begin
        image_1_55 <= io_pixelVal_in_1_3;
      end else if (10'h37 == _T_22[9:0]) begin
        image_1_55 <= io_pixelVal_in_1_2;
      end else if (10'h37 == _T_19[9:0]) begin
        image_1_55 <= io_pixelVal_in_1_1;
      end else if (10'h37 == _T_15[9:0]) begin
        image_1_55 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_56 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h38 == _T_37[9:0]) begin
        image_1_56 <= io_pixelVal_in_1_7;
      end else if (10'h38 == _T_34[9:0]) begin
        image_1_56 <= io_pixelVal_in_1_6;
      end else if (10'h38 == _T_31[9:0]) begin
        image_1_56 <= io_pixelVal_in_1_5;
      end else if (10'h38 == _T_28[9:0]) begin
        image_1_56 <= io_pixelVal_in_1_4;
      end else if (10'h38 == _T_25[9:0]) begin
        image_1_56 <= io_pixelVal_in_1_3;
      end else if (10'h38 == _T_22[9:0]) begin
        image_1_56 <= io_pixelVal_in_1_2;
      end else if (10'h38 == _T_19[9:0]) begin
        image_1_56 <= io_pixelVal_in_1_1;
      end else if (10'h38 == _T_15[9:0]) begin
        image_1_56 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_57 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h39 == _T_37[9:0]) begin
        image_1_57 <= io_pixelVal_in_1_7;
      end else if (10'h39 == _T_34[9:0]) begin
        image_1_57 <= io_pixelVal_in_1_6;
      end else if (10'h39 == _T_31[9:0]) begin
        image_1_57 <= io_pixelVal_in_1_5;
      end else if (10'h39 == _T_28[9:0]) begin
        image_1_57 <= io_pixelVal_in_1_4;
      end else if (10'h39 == _T_25[9:0]) begin
        image_1_57 <= io_pixelVal_in_1_3;
      end else if (10'h39 == _T_22[9:0]) begin
        image_1_57 <= io_pixelVal_in_1_2;
      end else if (10'h39 == _T_19[9:0]) begin
        image_1_57 <= io_pixelVal_in_1_1;
      end else if (10'h39 == _T_15[9:0]) begin
        image_1_57 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_58 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h3a == _T_37[9:0]) begin
        image_1_58 <= io_pixelVal_in_1_7;
      end else if (10'h3a == _T_34[9:0]) begin
        image_1_58 <= io_pixelVal_in_1_6;
      end else if (10'h3a == _T_31[9:0]) begin
        image_1_58 <= io_pixelVal_in_1_5;
      end else if (10'h3a == _T_28[9:0]) begin
        image_1_58 <= io_pixelVal_in_1_4;
      end else if (10'h3a == _T_25[9:0]) begin
        image_1_58 <= io_pixelVal_in_1_3;
      end else if (10'h3a == _T_22[9:0]) begin
        image_1_58 <= io_pixelVal_in_1_2;
      end else if (10'h3a == _T_19[9:0]) begin
        image_1_58 <= io_pixelVal_in_1_1;
      end else if (10'h3a == _T_15[9:0]) begin
        image_1_58 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_59 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h3b == _T_37[9:0]) begin
        image_1_59 <= io_pixelVal_in_1_7;
      end else if (10'h3b == _T_34[9:0]) begin
        image_1_59 <= io_pixelVal_in_1_6;
      end else if (10'h3b == _T_31[9:0]) begin
        image_1_59 <= io_pixelVal_in_1_5;
      end else if (10'h3b == _T_28[9:0]) begin
        image_1_59 <= io_pixelVal_in_1_4;
      end else if (10'h3b == _T_25[9:0]) begin
        image_1_59 <= io_pixelVal_in_1_3;
      end else if (10'h3b == _T_22[9:0]) begin
        image_1_59 <= io_pixelVal_in_1_2;
      end else if (10'h3b == _T_19[9:0]) begin
        image_1_59 <= io_pixelVal_in_1_1;
      end else if (10'h3b == _T_15[9:0]) begin
        image_1_59 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_60 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h3c == _T_37[9:0]) begin
        image_1_60 <= io_pixelVal_in_1_7;
      end else if (10'h3c == _T_34[9:0]) begin
        image_1_60 <= io_pixelVal_in_1_6;
      end else if (10'h3c == _T_31[9:0]) begin
        image_1_60 <= io_pixelVal_in_1_5;
      end else if (10'h3c == _T_28[9:0]) begin
        image_1_60 <= io_pixelVal_in_1_4;
      end else if (10'h3c == _T_25[9:0]) begin
        image_1_60 <= io_pixelVal_in_1_3;
      end else if (10'h3c == _T_22[9:0]) begin
        image_1_60 <= io_pixelVal_in_1_2;
      end else if (10'h3c == _T_19[9:0]) begin
        image_1_60 <= io_pixelVal_in_1_1;
      end else if (10'h3c == _T_15[9:0]) begin
        image_1_60 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_61 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h3d == _T_37[9:0]) begin
        image_1_61 <= io_pixelVal_in_1_7;
      end else if (10'h3d == _T_34[9:0]) begin
        image_1_61 <= io_pixelVal_in_1_6;
      end else if (10'h3d == _T_31[9:0]) begin
        image_1_61 <= io_pixelVal_in_1_5;
      end else if (10'h3d == _T_28[9:0]) begin
        image_1_61 <= io_pixelVal_in_1_4;
      end else if (10'h3d == _T_25[9:0]) begin
        image_1_61 <= io_pixelVal_in_1_3;
      end else if (10'h3d == _T_22[9:0]) begin
        image_1_61 <= io_pixelVal_in_1_2;
      end else if (10'h3d == _T_19[9:0]) begin
        image_1_61 <= io_pixelVal_in_1_1;
      end else if (10'h3d == _T_15[9:0]) begin
        image_1_61 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_62 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h3e == _T_37[9:0]) begin
        image_1_62 <= io_pixelVal_in_1_7;
      end else if (10'h3e == _T_34[9:0]) begin
        image_1_62 <= io_pixelVal_in_1_6;
      end else if (10'h3e == _T_31[9:0]) begin
        image_1_62 <= io_pixelVal_in_1_5;
      end else if (10'h3e == _T_28[9:0]) begin
        image_1_62 <= io_pixelVal_in_1_4;
      end else if (10'h3e == _T_25[9:0]) begin
        image_1_62 <= io_pixelVal_in_1_3;
      end else if (10'h3e == _T_22[9:0]) begin
        image_1_62 <= io_pixelVal_in_1_2;
      end else if (10'h3e == _T_19[9:0]) begin
        image_1_62 <= io_pixelVal_in_1_1;
      end else if (10'h3e == _T_15[9:0]) begin
        image_1_62 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_63 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h3f == _T_37[9:0]) begin
        image_1_63 <= io_pixelVal_in_1_7;
      end else if (10'h3f == _T_34[9:0]) begin
        image_1_63 <= io_pixelVal_in_1_6;
      end else if (10'h3f == _T_31[9:0]) begin
        image_1_63 <= io_pixelVal_in_1_5;
      end else if (10'h3f == _T_28[9:0]) begin
        image_1_63 <= io_pixelVal_in_1_4;
      end else if (10'h3f == _T_25[9:0]) begin
        image_1_63 <= io_pixelVal_in_1_3;
      end else if (10'h3f == _T_22[9:0]) begin
        image_1_63 <= io_pixelVal_in_1_2;
      end else if (10'h3f == _T_19[9:0]) begin
        image_1_63 <= io_pixelVal_in_1_1;
      end else if (10'h3f == _T_15[9:0]) begin
        image_1_63 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_64 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h40 == _T_37[9:0]) begin
        image_1_64 <= io_pixelVal_in_1_7;
      end else if (10'h40 == _T_34[9:0]) begin
        image_1_64 <= io_pixelVal_in_1_6;
      end else if (10'h40 == _T_31[9:0]) begin
        image_1_64 <= io_pixelVal_in_1_5;
      end else if (10'h40 == _T_28[9:0]) begin
        image_1_64 <= io_pixelVal_in_1_4;
      end else if (10'h40 == _T_25[9:0]) begin
        image_1_64 <= io_pixelVal_in_1_3;
      end else if (10'h40 == _T_22[9:0]) begin
        image_1_64 <= io_pixelVal_in_1_2;
      end else if (10'h40 == _T_19[9:0]) begin
        image_1_64 <= io_pixelVal_in_1_1;
      end else if (10'h40 == _T_15[9:0]) begin
        image_1_64 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_65 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h41 == _T_37[9:0]) begin
        image_1_65 <= io_pixelVal_in_1_7;
      end else if (10'h41 == _T_34[9:0]) begin
        image_1_65 <= io_pixelVal_in_1_6;
      end else if (10'h41 == _T_31[9:0]) begin
        image_1_65 <= io_pixelVal_in_1_5;
      end else if (10'h41 == _T_28[9:0]) begin
        image_1_65 <= io_pixelVal_in_1_4;
      end else if (10'h41 == _T_25[9:0]) begin
        image_1_65 <= io_pixelVal_in_1_3;
      end else if (10'h41 == _T_22[9:0]) begin
        image_1_65 <= io_pixelVal_in_1_2;
      end else if (10'h41 == _T_19[9:0]) begin
        image_1_65 <= io_pixelVal_in_1_1;
      end else if (10'h41 == _T_15[9:0]) begin
        image_1_65 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_66 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h42 == _T_37[9:0]) begin
        image_1_66 <= io_pixelVal_in_1_7;
      end else if (10'h42 == _T_34[9:0]) begin
        image_1_66 <= io_pixelVal_in_1_6;
      end else if (10'h42 == _T_31[9:0]) begin
        image_1_66 <= io_pixelVal_in_1_5;
      end else if (10'h42 == _T_28[9:0]) begin
        image_1_66 <= io_pixelVal_in_1_4;
      end else if (10'h42 == _T_25[9:0]) begin
        image_1_66 <= io_pixelVal_in_1_3;
      end else if (10'h42 == _T_22[9:0]) begin
        image_1_66 <= io_pixelVal_in_1_2;
      end else if (10'h42 == _T_19[9:0]) begin
        image_1_66 <= io_pixelVal_in_1_1;
      end else if (10'h42 == _T_15[9:0]) begin
        image_1_66 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_67 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h43 == _T_37[9:0]) begin
        image_1_67 <= io_pixelVal_in_1_7;
      end else if (10'h43 == _T_34[9:0]) begin
        image_1_67 <= io_pixelVal_in_1_6;
      end else if (10'h43 == _T_31[9:0]) begin
        image_1_67 <= io_pixelVal_in_1_5;
      end else if (10'h43 == _T_28[9:0]) begin
        image_1_67 <= io_pixelVal_in_1_4;
      end else if (10'h43 == _T_25[9:0]) begin
        image_1_67 <= io_pixelVal_in_1_3;
      end else if (10'h43 == _T_22[9:0]) begin
        image_1_67 <= io_pixelVal_in_1_2;
      end else if (10'h43 == _T_19[9:0]) begin
        image_1_67 <= io_pixelVal_in_1_1;
      end else if (10'h43 == _T_15[9:0]) begin
        image_1_67 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_68 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h44 == _T_37[9:0]) begin
        image_1_68 <= io_pixelVal_in_1_7;
      end else if (10'h44 == _T_34[9:0]) begin
        image_1_68 <= io_pixelVal_in_1_6;
      end else if (10'h44 == _T_31[9:0]) begin
        image_1_68 <= io_pixelVal_in_1_5;
      end else if (10'h44 == _T_28[9:0]) begin
        image_1_68 <= io_pixelVal_in_1_4;
      end else if (10'h44 == _T_25[9:0]) begin
        image_1_68 <= io_pixelVal_in_1_3;
      end else if (10'h44 == _T_22[9:0]) begin
        image_1_68 <= io_pixelVal_in_1_2;
      end else if (10'h44 == _T_19[9:0]) begin
        image_1_68 <= io_pixelVal_in_1_1;
      end else if (10'h44 == _T_15[9:0]) begin
        image_1_68 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_69 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h45 == _T_37[9:0]) begin
        image_1_69 <= io_pixelVal_in_1_7;
      end else if (10'h45 == _T_34[9:0]) begin
        image_1_69 <= io_pixelVal_in_1_6;
      end else if (10'h45 == _T_31[9:0]) begin
        image_1_69 <= io_pixelVal_in_1_5;
      end else if (10'h45 == _T_28[9:0]) begin
        image_1_69 <= io_pixelVal_in_1_4;
      end else if (10'h45 == _T_25[9:0]) begin
        image_1_69 <= io_pixelVal_in_1_3;
      end else if (10'h45 == _T_22[9:0]) begin
        image_1_69 <= io_pixelVal_in_1_2;
      end else if (10'h45 == _T_19[9:0]) begin
        image_1_69 <= io_pixelVal_in_1_1;
      end else if (10'h45 == _T_15[9:0]) begin
        image_1_69 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_70 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h46 == _T_37[9:0]) begin
        image_1_70 <= io_pixelVal_in_1_7;
      end else if (10'h46 == _T_34[9:0]) begin
        image_1_70 <= io_pixelVal_in_1_6;
      end else if (10'h46 == _T_31[9:0]) begin
        image_1_70 <= io_pixelVal_in_1_5;
      end else if (10'h46 == _T_28[9:0]) begin
        image_1_70 <= io_pixelVal_in_1_4;
      end else if (10'h46 == _T_25[9:0]) begin
        image_1_70 <= io_pixelVal_in_1_3;
      end else if (10'h46 == _T_22[9:0]) begin
        image_1_70 <= io_pixelVal_in_1_2;
      end else if (10'h46 == _T_19[9:0]) begin
        image_1_70 <= io_pixelVal_in_1_1;
      end else if (10'h46 == _T_15[9:0]) begin
        image_1_70 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_71 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h47 == _T_37[9:0]) begin
        image_1_71 <= io_pixelVal_in_1_7;
      end else if (10'h47 == _T_34[9:0]) begin
        image_1_71 <= io_pixelVal_in_1_6;
      end else if (10'h47 == _T_31[9:0]) begin
        image_1_71 <= io_pixelVal_in_1_5;
      end else if (10'h47 == _T_28[9:0]) begin
        image_1_71 <= io_pixelVal_in_1_4;
      end else if (10'h47 == _T_25[9:0]) begin
        image_1_71 <= io_pixelVal_in_1_3;
      end else if (10'h47 == _T_22[9:0]) begin
        image_1_71 <= io_pixelVal_in_1_2;
      end else if (10'h47 == _T_19[9:0]) begin
        image_1_71 <= io_pixelVal_in_1_1;
      end else if (10'h47 == _T_15[9:0]) begin
        image_1_71 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_72 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h48 == _T_37[9:0]) begin
        image_1_72 <= io_pixelVal_in_1_7;
      end else if (10'h48 == _T_34[9:0]) begin
        image_1_72 <= io_pixelVal_in_1_6;
      end else if (10'h48 == _T_31[9:0]) begin
        image_1_72 <= io_pixelVal_in_1_5;
      end else if (10'h48 == _T_28[9:0]) begin
        image_1_72 <= io_pixelVal_in_1_4;
      end else if (10'h48 == _T_25[9:0]) begin
        image_1_72 <= io_pixelVal_in_1_3;
      end else if (10'h48 == _T_22[9:0]) begin
        image_1_72 <= io_pixelVal_in_1_2;
      end else if (10'h48 == _T_19[9:0]) begin
        image_1_72 <= io_pixelVal_in_1_1;
      end else if (10'h48 == _T_15[9:0]) begin
        image_1_72 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_73 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h49 == _T_37[9:0]) begin
        image_1_73 <= io_pixelVal_in_1_7;
      end else if (10'h49 == _T_34[9:0]) begin
        image_1_73 <= io_pixelVal_in_1_6;
      end else if (10'h49 == _T_31[9:0]) begin
        image_1_73 <= io_pixelVal_in_1_5;
      end else if (10'h49 == _T_28[9:0]) begin
        image_1_73 <= io_pixelVal_in_1_4;
      end else if (10'h49 == _T_25[9:0]) begin
        image_1_73 <= io_pixelVal_in_1_3;
      end else if (10'h49 == _T_22[9:0]) begin
        image_1_73 <= io_pixelVal_in_1_2;
      end else if (10'h49 == _T_19[9:0]) begin
        image_1_73 <= io_pixelVal_in_1_1;
      end else if (10'h49 == _T_15[9:0]) begin
        image_1_73 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_74 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h4a == _T_37[9:0]) begin
        image_1_74 <= io_pixelVal_in_1_7;
      end else if (10'h4a == _T_34[9:0]) begin
        image_1_74 <= io_pixelVal_in_1_6;
      end else if (10'h4a == _T_31[9:0]) begin
        image_1_74 <= io_pixelVal_in_1_5;
      end else if (10'h4a == _T_28[9:0]) begin
        image_1_74 <= io_pixelVal_in_1_4;
      end else if (10'h4a == _T_25[9:0]) begin
        image_1_74 <= io_pixelVal_in_1_3;
      end else if (10'h4a == _T_22[9:0]) begin
        image_1_74 <= io_pixelVal_in_1_2;
      end else if (10'h4a == _T_19[9:0]) begin
        image_1_74 <= io_pixelVal_in_1_1;
      end else if (10'h4a == _T_15[9:0]) begin
        image_1_74 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_75 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h4b == _T_37[9:0]) begin
        image_1_75 <= io_pixelVal_in_1_7;
      end else if (10'h4b == _T_34[9:0]) begin
        image_1_75 <= io_pixelVal_in_1_6;
      end else if (10'h4b == _T_31[9:0]) begin
        image_1_75 <= io_pixelVal_in_1_5;
      end else if (10'h4b == _T_28[9:0]) begin
        image_1_75 <= io_pixelVal_in_1_4;
      end else if (10'h4b == _T_25[9:0]) begin
        image_1_75 <= io_pixelVal_in_1_3;
      end else if (10'h4b == _T_22[9:0]) begin
        image_1_75 <= io_pixelVal_in_1_2;
      end else if (10'h4b == _T_19[9:0]) begin
        image_1_75 <= io_pixelVal_in_1_1;
      end else if (10'h4b == _T_15[9:0]) begin
        image_1_75 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_76 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h4c == _T_37[9:0]) begin
        image_1_76 <= io_pixelVal_in_1_7;
      end else if (10'h4c == _T_34[9:0]) begin
        image_1_76 <= io_pixelVal_in_1_6;
      end else if (10'h4c == _T_31[9:0]) begin
        image_1_76 <= io_pixelVal_in_1_5;
      end else if (10'h4c == _T_28[9:0]) begin
        image_1_76 <= io_pixelVal_in_1_4;
      end else if (10'h4c == _T_25[9:0]) begin
        image_1_76 <= io_pixelVal_in_1_3;
      end else if (10'h4c == _T_22[9:0]) begin
        image_1_76 <= io_pixelVal_in_1_2;
      end else if (10'h4c == _T_19[9:0]) begin
        image_1_76 <= io_pixelVal_in_1_1;
      end else if (10'h4c == _T_15[9:0]) begin
        image_1_76 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_77 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h4d == _T_37[9:0]) begin
        image_1_77 <= io_pixelVal_in_1_7;
      end else if (10'h4d == _T_34[9:0]) begin
        image_1_77 <= io_pixelVal_in_1_6;
      end else if (10'h4d == _T_31[9:0]) begin
        image_1_77 <= io_pixelVal_in_1_5;
      end else if (10'h4d == _T_28[9:0]) begin
        image_1_77 <= io_pixelVal_in_1_4;
      end else if (10'h4d == _T_25[9:0]) begin
        image_1_77 <= io_pixelVal_in_1_3;
      end else if (10'h4d == _T_22[9:0]) begin
        image_1_77 <= io_pixelVal_in_1_2;
      end else if (10'h4d == _T_19[9:0]) begin
        image_1_77 <= io_pixelVal_in_1_1;
      end else if (10'h4d == _T_15[9:0]) begin
        image_1_77 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_78 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h4e == _T_37[9:0]) begin
        image_1_78 <= io_pixelVal_in_1_7;
      end else if (10'h4e == _T_34[9:0]) begin
        image_1_78 <= io_pixelVal_in_1_6;
      end else if (10'h4e == _T_31[9:0]) begin
        image_1_78 <= io_pixelVal_in_1_5;
      end else if (10'h4e == _T_28[9:0]) begin
        image_1_78 <= io_pixelVal_in_1_4;
      end else if (10'h4e == _T_25[9:0]) begin
        image_1_78 <= io_pixelVal_in_1_3;
      end else if (10'h4e == _T_22[9:0]) begin
        image_1_78 <= io_pixelVal_in_1_2;
      end else if (10'h4e == _T_19[9:0]) begin
        image_1_78 <= io_pixelVal_in_1_1;
      end else if (10'h4e == _T_15[9:0]) begin
        image_1_78 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_79 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h4f == _T_37[9:0]) begin
        image_1_79 <= io_pixelVal_in_1_7;
      end else if (10'h4f == _T_34[9:0]) begin
        image_1_79 <= io_pixelVal_in_1_6;
      end else if (10'h4f == _T_31[9:0]) begin
        image_1_79 <= io_pixelVal_in_1_5;
      end else if (10'h4f == _T_28[9:0]) begin
        image_1_79 <= io_pixelVal_in_1_4;
      end else if (10'h4f == _T_25[9:0]) begin
        image_1_79 <= io_pixelVal_in_1_3;
      end else if (10'h4f == _T_22[9:0]) begin
        image_1_79 <= io_pixelVal_in_1_2;
      end else if (10'h4f == _T_19[9:0]) begin
        image_1_79 <= io_pixelVal_in_1_1;
      end else if (10'h4f == _T_15[9:0]) begin
        image_1_79 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_80 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h50 == _T_37[9:0]) begin
        image_1_80 <= io_pixelVal_in_1_7;
      end else if (10'h50 == _T_34[9:0]) begin
        image_1_80 <= io_pixelVal_in_1_6;
      end else if (10'h50 == _T_31[9:0]) begin
        image_1_80 <= io_pixelVal_in_1_5;
      end else if (10'h50 == _T_28[9:0]) begin
        image_1_80 <= io_pixelVal_in_1_4;
      end else if (10'h50 == _T_25[9:0]) begin
        image_1_80 <= io_pixelVal_in_1_3;
      end else if (10'h50 == _T_22[9:0]) begin
        image_1_80 <= io_pixelVal_in_1_2;
      end else if (10'h50 == _T_19[9:0]) begin
        image_1_80 <= io_pixelVal_in_1_1;
      end else if (10'h50 == _T_15[9:0]) begin
        image_1_80 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_81 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h51 == _T_37[9:0]) begin
        image_1_81 <= io_pixelVal_in_1_7;
      end else if (10'h51 == _T_34[9:0]) begin
        image_1_81 <= io_pixelVal_in_1_6;
      end else if (10'h51 == _T_31[9:0]) begin
        image_1_81 <= io_pixelVal_in_1_5;
      end else if (10'h51 == _T_28[9:0]) begin
        image_1_81 <= io_pixelVal_in_1_4;
      end else if (10'h51 == _T_25[9:0]) begin
        image_1_81 <= io_pixelVal_in_1_3;
      end else if (10'h51 == _T_22[9:0]) begin
        image_1_81 <= io_pixelVal_in_1_2;
      end else if (10'h51 == _T_19[9:0]) begin
        image_1_81 <= io_pixelVal_in_1_1;
      end else if (10'h51 == _T_15[9:0]) begin
        image_1_81 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_82 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h52 == _T_37[9:0]) begin
        image_1_82 <= io_pixelVal_in_1_7;
      end else if (10'h52 == _T_34[9:0]) begin
        image_1_82 <= io_pixelVal_in_1_6;
      end else if (10'h52 == _T_31[9:0]) begin
        image_1_82 <= io_pixelVal_in_1_5;
      end else if (10'h52 == _T_28[9:0]) begin
        image_1_82 <= io_pixelVal_in_1_4;
      end else if (10'h52 == _T_25[9:0]) begin
        image_1_82 <= io_pixelVal_in_1_3;
      end else if (10'h52 == _T_22[9:0]) begin
        image_1_82 <= io_pixelVal_in_1_2;
      end else if (10'h52 == _T_19[9:0]) begin
        image_1_82 <= io_pixelVal_in_1_1;
      end else if (10'h52 == _T_15[9:0]) begin
        image_1_82 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_83 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h53 == _T_37[9:0]) begin
        image_1_83 <= io_pixelVal_in_1_7;
      end else if (10'h53 == _T_34[9:0]) begin
        image_1_83 <= io_pixelVal_in_1_6;
      end else if (10'h53 == _T_31[9:0]) begin
        image_1_83 <= io_pixelVal_in_1_5;
      end else if (10'h53 == _T_28[9:0]) begin
        image_1_83 <= io_pixelVal_in_1_4;
      end else if (10'h53 == _T_25[9:0]) begin
        image_1_83 <= io_pixelVal_in_1_3;
      end else if (10'h53 == _T_22[9:0]) begin
        image_1_83 <= io_pixelVal_in_1_2;
      end else if (10'h53 == _T_19[9:0]) begin
        image_1_83 <= io_pixelVal_in_1_1;
      end else if (10'h53 == _T_15[9:0]) begin
        image_1_83 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_84 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h54 == _T_37[9:0]) begin
        image_1_84 <= io_pixelVal_in_1_7;
      end else if (10'h54 == _T_34[9:0]) begin
        image_1_84 <= io_pixelVal_in_1_6;
      end else if (10'h54 == _T_31[9:0]) begin
        image_1_84 <= io_pixelVal_in_1_5;
      end else if (10'h54 == _T_28[9:0]) begin
        image_1_84 <= io_pixelVal_in_1_4;
      end else if (10'h54 == _T_25[9:0]) begin
        image_1_84 <= io_pixelVal_in_1_3;
      end else if (10'h54 == _T_22[9:0]) begin
        image_1_84 <= io_pixelVal_in_1_2;
      end else if (10'h54 == _T_19[9:0]) begin
        image_1_84 <= io_pixelVal_in_1_1;
      end else if (10'h54 == _T_15[9:0]) begin
        image_1_84 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_85 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h55 == _T_37[9:0]) begin
        image_1_85 <= io_pixelVal_in_1_7;
      end else if (10'h55 == _T_34[9:0]) begin
        image_1_85 <= io_pixelVal_in_1_6;
      end else if (10'h55 == _T_31[9:0]) begin
        image_1_85 <= io_pixelVal_in_1_5;
      end else if (10'h55 == _T_28[9:0]) begin
        image_1_85 <= io_pixelVal_in_1_4;
      end else if (10'h55 == _T_25[9:0]) begin
        image_1_85 <= io_pixelVal_in_1_3;
      end else if (10'h55 == _T_22[9:0]) begin
        image_1_85 <= io_pixelVal_in_1_2;
      end else if (10'h55 == _T_19[9:0]) begin
        image_1_85 <= io_pixelVal_in_1_1;
      end else if (10'h55 == _T_15[9:0]) begin
        image_1_85 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_86 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h56 == _T_37[9:0]) begin
        image_1_86 <= io_pixelVal_in_1_7;
      end else if (10'h56 == _T_34[9:0]) begin
        image_1_86 <= io_pixelVal_in_1_6;
      end else if (10'h56 == _T_31[9:0]) begin
        image_1_86 <= io_pixelVal_in_1_5;
      end else if (10'h56 == _T_28[9:0]) begin
        image_1_86 <= io_pixelVal_in_1_4;
      end else if (10'h56 == _T_25[9:0]) begin
        image_1_86 <= io_pixelVal_in_1_3;
      end else if (10'h56 == _T_22[9:0]) begin
        image_1_86 <= io_pixelVal_in_1_2;
      end else if (10'h56 == _T_19[9:0]) begin
        image_1_86 <= io_pixelVal_in_1_1;
      end else if (10'h56 == _T_15[9:0]) begin
        image_1_86 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_87 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h57 == _T_37[9:0]) begin
        image_1_87 <= io_pixelVal_in_1_7;
      end else if (10'h57 == _T_34[9:0]) begin
        image_1_87 <= io_pixelVal_in_1_6;
      end else if (10'h57 == _T_31[9:0]) begin
        image_1_87 <= io_pixelVal_in_1_5;
      end else if (10'h57 == _T_28[9:0]) begin
        image_1_87 <= io_pixelVal_in_1_4;
      end else if (10'h57 == _T_25[9:0]) begin
        image_1_87 <= io_pixelVal_in_1_3;
      end else if (10'h57 == _T_22[9:0]) begin
        image_1_87 <= io_pixelVal_in_1_2;
      end else if (10'h57 == _T_19[9:0]) begin
        image_1_87 <= io_pixelVal_in_1_1;
      end else if (10'h57 == _T_15[9:0]) begin
        image_1_87 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_88 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h58 == _T_37[9:0]) begin
        image_1_88 <= io_pixelVal_in_1_7;
      end else if (10'h58 == _T_34[9:0]) begin
        image_1_88 <= io_pixelVal_in_1_6;
      end else if (10'h58 == _T_31[9:0]) begin
        image_1_88 <= io_pixelVal_in_1_5;
      end else if (10'h58 == _T_28[9:0]) begin
        image_1_88 <= io_pixelVal_in_1_4;
      end else if (10'h58 == _T_25[9:0]) begin
        image_1_88 <= io_pixelVal_in_1_3;
      end else if (10'h58 == _T_22[9:0]) begin
        image_1_88 <= io_pixelVal_in_1_2;
      end else if (10'h58 == _T_19[9:0]) begin
        image_1_88 <= io_pixelVal_in_1_1;
      end else if (10'h58 == _T_15[9:0]) begin
        image_1_88 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_89 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h59 == _T_37[9:0]) begin
        image_1_89 <= io_pixelVal_in_1_7;
      end else if (10'h59 == _T_34[9:0]) begin
        image_1_89 <= io_pixelVal_in_1_6;
      end else if (10'h59 == _T_31[9:0]) begin
        image_1_89 <= io_pixelVal_in_1_5;
      end else if (10'h59 == _T_28[9:0]) begin
        image_1_89 <= io_pixelVal_in_1_4;
      end else if (10'h59 == _T_25[9:0]) begin
        image_1_89 <= io_pixelVal_in_1_3;
      end else if (10'h59 == _T_22[9:0]) begin
        image_1_89 <= io_pixelVal_in_1_2;
      end else if (10'h59 == _T_19[9:0]) begin
        image_1_89 <= io_pixelVal_in_1_1;
      end else if (10'h59 == _T_15[9:0]) begin
        image_1_89 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_90 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h5a == _T_37[9:0]) begin
        image_1_90 <= io_pixelVal_in_1_7;
      end else if (10'h5a == _T_34[9:0]) begin
        image_1_90 <= io_pixelVal_in_1_6;
      end else if (10'h5a == _T_31[9:0]) begin
        image_1_90 <= io_pixelVal_in_1_5;
      end else if (10'h5a == _T_28[9:0]) begin
        image_1_90 <= io_pixelVal_in_1_4;
      end else if (10'h5a == _T_25[9:0]) begin
        image_1_90 <= io_pixelVal_in_1_3;
      end else if (10'h5a == _T_22[9:0]) begin
        image_1_90 <= io_pixelVal_in_1_2;
      end else if (10'h5a == _T_19[9:0]) begin
        image_1_90 <= io_pixelVal_in_1_1;
      end else if (10'h5a == _T_15[9:0]) begin
        image_1_90 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_91 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h5b == _T_37[9:0]) begin
        image_1_91 <= io_pixelVal_in_1_7;
      end else if (10'h5b == _T_34[9:0]) begin
        image_1_91 <= io_pixelVal_in_1_6;
      end else if (10'h5b == _T_31[9:0]) begin
        image_1_91 <= io_pixelVal_in_1_5;
      end else if (10'h5b == _T_28[9:0]) begin
        image_1_91 <= io_pixelVal_in_1_4;
      end else if (10'h5b == _T_25[9:0]) begin
        image_1_91 <= io_pixelVal_in_1_3;
      end else if (10'h5b == _T_22[9:0]) begin
        image_1_91 <= io_pixelVal_in_1_2;
      end else if (10'h5b == _T_19[9:0]) begin
        image_1_91 <= io_pixelVal_in_1_1;
      end else if (10'h5b == _T_15[9:0]) begin
        image_1_91 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_92 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h5c == _T_37[9:0]) begin
        image_1_92 <= io_pixelVal_in_1_7;
      end else if (10'h5c == _T_34[9:0]) begin
        image_1_92 <= io_pixelVal_in_1_6;
      end else if (10'h5c == _T_31[9:0]) begin
        image_1_92 <= io_pixelVal_in_1_5;
      end else if (10'h5c == _T_28[9:0]) begin
        image_1_92 <= io_pixelVal_in_1_4;
      end else if (10'h5c == _T_25[9:0]) begin
        image_1_92 <= io_pixelVal_in_1_3;
      end else if (10'h5c == _T_22[9:0]) begin
        image_1_92 <= io_pixelVal_in_1_2;
      end else if (10'h5c == _T_19[9:0]) begin
        image_1_92 <= io_pixelVal_in_1_1;
      end else if (10'h5c == _T_15[9:0]) begin
        image_1_92 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_93 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h5d == _T_37[9:0]) begin
        image_1_93 <= io_pixelVal_in_1_7;
      end else if (10'h5d == _T_34[9:0]) begin
        image_1_93 <= io_pixelVal_in_1_6;
      end else if (10'h5d == _T_31[9:0]) begin
        image_1_93 <= io_pixelVal_in_1_5;
      end else if (10'h5d == _T_28[9:0]) begin
        image_1_93 <= io_pixelVal_in_1_4;
      end else if (10'h5d == _T_25[9:0]) begin
        image_1_93 <= io_pixelVal_in_1_3;
      end else if (10'h5d == _T_22[9:0]) begin
        image_1_93 <= io_pixelVal_in_1_2;
      end else if (10'h5d == _T_19[9:0]) begin
        image_1_93 <= io_pixelVal_in_1_1;
      end else if (10'h5d == _T_15[9:0]) begin
        image_1_93 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_94 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h5e == _T_37[9:0]) begin
        image_1_94 <= io_pixelVal_in_1_7;
      end else if (10'h5e == _T_34[9:0]) begin
        image_1_94 <= io_pixelVal_in_1_6;
      end else if (10'h5e == _T_31[9:0]) begin
        image_1_94 <= io_pixelVal_in_1_5;
      end else if (10'h5e == _T_28[9:0]) begin
        image_1_94 <= io_pixelVal_in_1_4;
      end else if (10'h5e == _T_25[9:0]) begin
        image_1_94 <= io_pixelVal_in_1_3;
      end else if (10'h5e == _T_22[9:0]) begin
        image_1_94 <= io_pixelVal_in_1_2;
      end else if (10'h5e == _T_19[9:0]) begin
        image_1_94 <= io_pixelVal_in_1_1;
      end else if (10'h5e == _T_15[9:0]) begin
        image_1_94 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_95 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h5f == _T_37[9:0]) begin
        image_1_95 <= io_pixelVal_in_1_7;
      end else if (10'h5f == _T_34[9:0]) begin
        image_1_95 <= io_pixelVal_in_1_6;
      end else if (10'h5f == _T_31[9:0]) begin
        image_1_95 <= io_pixelVal_in_1_5;
      end else if (10'h5f == _T_28[9:0]) begin
        image_1_95 <= io_pixelVal_in_1_4;
      end else if (10'h5f == _T_25[9:0]) begin
        image_1_95 <= io_pixelVal_in_1_3;
      end else if (10'h5f == _T_22[9:0]) begin
        image_1_95 <= io_pixelVal_in_1_2;
      end else if (10'h5f == _T_19[9:0]) begin
        image_1_95 <= io_pixelVal_in_1_1;
      end else if (10'h5f == _T_15[9:0]) begin
        image_1_95 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_96 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h60 == _T_37[9:0]) begin
        image_1_96 <= io_pixelVal_in_1_7;
      end else if (10'h60 == _T_34[9:0]) begin
        image_1_96 <= io_pixelVal_in_1_6;
      end else if (10'h60 == _T_31[9:0]) begin
        image_1_96 <= io_pixelVal_in_1_5;
      end else if (10'h60 == _T_28[9:0]) begin
        image_1_96 <= io_pixelVal_in_1_4;
      end else if (10'h60 == _T_25[9:0]) begin
        image_1_96 <= io_pixelVal_in_1_3;
      end else if (10'h60 == _T_22[9:0]) begin
        image_1_96 <= io_pixelVal_in_1_2;
      end else if (10'h60 == _T_19[9:0]) begin
        image_1_96 <= io_pixelVal_in_1_1;
      end else if (10'h60 == _T_15[9:0]) begin
        image_1_96 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_97 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h61 == _T_37[9:0]) begin
        image_1_97 <= io_pixelVal_in_1_7;
      end else if (10'h61 == _T_34[9:0]) begin
        image_1_97 <= io_pixelVal_in_1_6;
      end else if (10'h61 == _T_31[9:0]) begin
        image_1_97 <= io_pixelVal_in_1_5;
      end else if (10'h61 == _T_28[9:0]) begin
        image_1_97 <= io_pixelVal_in_1_4;
      end else if (10'h61 == _T_25[9:0]) begin
        image_1_97 <= io_pixelVal_in_1_3;
      end else if (10'h61 == _T_22[9:0]) begin
        image_1_97 <= io_pixelVal_in_1_2;
      end else if (10'h61 == _T_19[9:0]) begin
        image_1_97 <= io_pixelVal_in_1_1;
      end else if (10'h61 == _T_15[9:0]) begin
        image_1_97 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_98 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h62 == _T_37[9:0]) begin
        image_1_98 <= io_pixelVal_in_1_7;
      end else if (10'h62 == _T_34[9:0]) begin
        image_1_98 <= io_pixelVal_in_1_6;
      end else if (10'h62 == _T_31[9:0]) begin
        image_1_98 <= io_pixelVal_in_1_5;
      end else if (10'h62 == _T_28[9:0]) begin
        image_1_98 <= io_pixelVal_in_1_4;
      end else if (10'h62 == _T_25[9:0]) begin
        image_1_98 <= io_pixelVal_in_1_3;
      end else if (10'h62 == _T_22[9:0]) begin
        image_1_98 <= io_pixelVal_in_1_2;
      end else if (10'h62 == _T_19[9:0]) begin
        image_1_98 <= io_pixelVal_in_1_1;
      end else if (10'h62 == _T_15[9:0]) begin
        image_1_98 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_99 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h63 == _T_37[9:0]) begin
        image_1_99 <= io_pixelVal_in_1_7;
      end else if (10'h63 == _T_34[9:0]) begin
        image_1_99 <= io_pixelVal_in_1_6;
      end else if (10'h63 == _T_31[9:0]) begin
        image_1_99 <= io_pixelVal_in_1_5;
      end else if (10'h63 == _T_28[9:0]) begin
        image_1_99 <= io_pixelVal_in_1_4;
      end else if (10'h63 == _T_25[9:0]) begin
        image_1_99 <= io_pixelVal_in_1_3;
      end else if (10'h63 == _T_22[9:0]) begin
        image_1_99 <= io_pixelVal_in_1_2;
      end else if (10'h63 == _T_19[9:0]) begin
        image_1_99 <= io_pixelVal_in_1_1;
      end else if (10'h63 == _T_15[9:0]) begin
        image_1_99 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_100 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h64 == _T_37[9:0]) begin
        image_1_100 <= io_pixelVal_in_1_7;
      end else if (10'h64 == _T_34[9:0]) begin
        image_1_100 <= io_pixelVal_in_1_6;
      end else if (10'h64 == _T_31[9:0]) begin
        image_1_100 <= io_pixelVal_in_1_5;
      end else if (10'h64 == _T_28[9:0]) begin
        image_1_100 <= io_pixelVal_in_1_4;
      end else if (10'h64 == _T_25[9:0]) begin
        image_1_100 <= io_pixelVal_in_1_3;
      end else if (10'h64 == _T_22[9:0]) begin
        image_1_100 <= io_pixelVal_in_1_2;
      end else if (10'h64 == _T_19[9:0]) begin
        image_1_100 <= io_pixelVal_in_1_1;
      end else if (10'h64 == _T_15[9:0]) begin
        image_1_100 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_101 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h65 == _T_37[9:0]) begin
        image_1_101 <= io_pixelVal_in_1_7;
      end else if (10'h65 == _T_34[9:0]) begin
        image_1_101 <= io_pixelVal_in_1_6;
      end else if (10'h65 == _T_31[9:0]) begin
        image_1_101 <= io_pixelVal_in_1_5;
      end else if (10'h65 == _T_28[9:0]) begin
        image_1_101 <= io_pixelVal_in_1_4;
      end else if (10'h65 == _T_25[9:0]) begin
        image_1_101 <= io_pixelVal_in_1_3;
      end else if (10'h65 == _T_22[9:0]) begin
        image_1_101 <= io_pixelVal_in_1_2;
      end else if (10'h65 == _T_19[9:0]) begin
        image_1_101 <= io_pixelVal_in_1_1;
      end else if (10'h65 == _T_15[9:0]) begin
        image_1_101 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_102 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h66 == _T_37[9:0]) begin
        image_1_102 <= io_pixelVal_in_1_7;
      end else if (10'h66 == _T_34[9:0]) begin
        image_1_102 <= io_pixelVal_in_1_6;
      end else if (10'h66 == _T_31[9:0]) begin
        image_1_102 <= io_pixelVal_in_1_5;
      end else if (10'h66 == _T_28[9:0]) begin
        image_1_102 <= io_pixelVal_in_1_4;
      end else if (10'h66 == _T_25[9:0]) begin
        image_1_102 <= io_pixelVal_in_1_3;
      end else if (10'h66 == _T_22[9:0]) begin
        image_1_102 <= io_pixelVal_in_1_2;
      end else if (10'h66 == _T_19[9:0]) begin
        image_1_102 <= io_pixelVal_in_1_1;
      end else if (10'h66 == _T_15[9:0]) begin
        image_1_102 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_103 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h67 == _T_37[9:0]) begin
        image_1_103 <= io_pixelVal_in_1_7;
      end else if (10'h67 == _T_34[9:0]) begin
        image_1_103 <= io_pixelVal_in_1_6;
      end else if (10'h67 == _T_31[9:0]) begin
        image_1_103 <= io_pixelVal_in_1_5;
      end else if (10'h67 == _T_28[9:0]) begin
        image_1_103 <= io_pixelVal_in_1_4;
      end else if (10'h67 == _T_25[9:0]) begin
        image_1_103 <= io_pixelVal_in_1_3;
      end else if (10'h67 == _T_22[9:0]) begin
        image_1_103 <= io_pixelVal_in_1_2;
      end else if (10'h67 == _T_19[9:0]) begin
        image_1_103 <= io_pixelVal_in_1_1;
      end else if (10'h67 == _T_15[9:0]) begin
        image_1_103 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_104 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h68 == _T_37[9:0]) begin
        image_1_104 <= io_pixelVal_in_1_7;
      end else if (10'h68 == _T_34[9:0]) begin
        image_1_104 <= io_pixelVal_in_1_6;
      end else if (10'h68 == _T_31[9:0]) begin
        image_1_104 <= io_pixelVal_in_1_5;
      end else if (10'h68 == _T_28[9:0]) begin
        image_1_104 <= io_pixelVal_in_1_4;
      end else if (10'h68 == _T_25[9:0]) begin
        image_1_104 <= io_pixelVal_in_1_3;
      end else if (10'h68 == _T_22[9:0]) begin
        image_1_104 <= io_pixelVal_in_1_2;
      end else if (10'h68 == _T_19[9:0]) begin
        image_1_104 <= io_pixelVal_in_1_1;
      end else if (10'h68 == _T_15[9:0]) begin
        image_1_104 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_105 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h69 == _T_37[9:0]) begin
        image_1_105 <= io_pixelVal_in_1_7;
      end else if (10'h69 == _T_34[9:0]) begin
        image_1_105 <= io_pixelVal_in_1_6;
      end else if (10'h69 == _T_31[9:0]) begin
        image_1_105 <= io_pixelVal_in_1_5;
      end else if (10'h69 == _T_28[9:0]) begin
        image_1_105 <= io_pixelVal_in_1_4;
      end else if (10'h69 == _T_25[9:0]) begin
        image_1_105 <= io_pixelVal_in_1_3;
      end else if (10'h69 == _T_22[9:0]) begin
        image_1_105 <= io_pixelVal_in_1_2;
      end else if (10'h69 == _T_19[9:0]) begin
        image_1_105 <= io_pixelVal_in_1_1;
      end else if (10'h69 == _T_15[9:0]) begin
        image_1_105 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_106 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h6a == _T_37[9:0]) begin
        image_1_106 <= io_pixelVal_in_1_7;
      end else if (10'h6a == _T_34[9:0]) begin
        image_1_106 <= io_pixelVal_in_1_6;
      end else if (10'h6a == _T_31[9:0]) begin
        image_1_106 <= io_pixelVal_in_1_5;
      end else if (10'h6a == _T_28[9:0]) begin
        image_1_106 <= io_pixelVal_in_1_4;
      end else if (10'h6a == _T_25[9:0]) begin
        image_1_106 <= io_pixelVal_in_1_3;
      end else if (10'h6a == _T_22[9:0]) begin
        image_1_106 <= io_pixelVal_in_1_2;
      end else if (10'h6a == _T_19[9:0]) begin
        image_1_106 <= io_pixelVal_in_1_1;
      end else if (10'h6a == _T_15[9:0]) begin
        image_1_106 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_107 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h6b == _T_37[9:0]) begin
        image_1_107 <= io_pixelVal_in_1_7;
      end else if (10'h6b == _T_34[9:0]) begin
        image_1_107 <= io_pixelVal_in_1_6;
      end else if (10'h6b == _T_31[9:0]) begin
        image_1_107 <= io_pixelVal_in_1_5;
      end else if (10'h6b == _T_28[9:0]) begin
        image_1_107 <= io_pixelVal_in_1_4;
      end else if (10'h6b == _T_25[9:0]) begin
        image_1_107 <= io_pixelVal_in_1_3;
      end else if (10'h6b == _T_22[9:0]) begin
        image_1_107 <= io_pixelVal_in_1_2;
      end else if (10'h6b == _T_19[9:0]) begin
        image_1_107 <= io_pixelVal_in_1_1;
      end else if (10'h6b == _T_15[9:0]) begin
        image_1_107 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_108 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h6c == _T_37[9:0]) begin
        image_1_108 <= io_pixelVal_in_1_7;
      end else if (10'h6c == _T_34[9:0]) begin
        image_1_108 <= io_pixelVal_in_1_6;
      end else if (10'h6c == _T_31[9:0]) begin
        image_1_108 <= io_pixelVal_in_1_5;
      end else if (10'h6c == _T_28[9:0]) begin
        image_1_108 <= io_pixelVal_in_1_4;
      end else if (10'h6c == _T_25[9:0]) begin
        image_1_108 <= io_pixelVal_in_1_3;
      end else if (10'h6c == _T_22[9:0]) begin
        image_1_108 <= io_pixelVal_in_1_2;
      end else if (10'h6c == _T_19[9:0]) begin
        image_1_108 <= io_pixelVal_in_1_1;
      end else if (10'h6c == _T_15[9:0]) begin
        image_1_108 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_109 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h6d == _T_37[9:0]) begin
        image_1_109 <= io_pixelVal_in_1_7;
      end else if (10'h6d == _T_34[9:0]) begin
        image_1_109 <= io_pixelVal_in_1_6;
      end else if (10'h6d == _T_31[9:0]) begin
        image_1_109 <= io_pixelVal_in_1_5;
      end else if (10'h6d == _T_28[9:0]) begin
        image_1_109 <= io_pixelVal_in_1_4;
      end else if (10'h6d == _T_25[9:0]) begin
        image_1_109 <= io_pixelVal_in_1_3;
      end else if (10'h6d == _T_22[9:0]) begin
        image_1_109 <= io_pixelVal_in_1_2;
      end else if (10'h6d == _T_19[9:0]) begin
        image_1_109 <= io_pixelVal_in_1_1;
      end else if (10'h6d == _T_15[9:0]) begin
        image_1_109 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_110 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h6e == _T_37[9:0]) begin
        image_1_110 <= io_pixelVal_in_1_7;
      end else if (10'h6e == _T_34[9:0]) begin
        image_1_110 <= io_pixelVal_in_1_6;
      end else if (10'h6e == _T_31[9:0]) begin
        image_1_110 <= io_pixelVal_in_1_5;
      end else if (10'h6e == _T_28[9:0]) begin
        image_1_110 <= io_pixelVal_in_1_4;
      end else if (10'h6e == _T_25[9:0]) begin
        image_1_110 <= io_pixelVal_in_1_3;
      end else if (10'h6e == _T_22[9:0]) begin
        image_1_110 <= io_pixelVal_in_1_2;
      end else if (10'h6e == _T_19[9:0]) begin
        image_1_110 <= io_pixelVal_in_1_1;
      end else if (10'h6e == _T_15[9:0]) begin
        image_1_110 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_111 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h6f == _T_37[9:0]) begin
        image_1_111 <= io_pixelVal_in_1_7;
      end else if (10'h6f == _T_34[9:0]) begin
        image_1_111 <= io_pixelVal_in_1_6;
      end else if (10'h6f == _T_31[9:0]) begin
        image_1_111 <= io_pixelVal_in_1_5;
      end else if (10'h6f == _T_28[9:0]) begin
        image_1_111 <= io_pixelVal_in_1_4;
      end else if (10'h6f == _T_25[9:0]) begin
        image_1_111 <= io_pixelVal_in_1_3;
      end else if (10'h6f == _T_22[9:0]) begin
        image_1_111 <= io_pixelVal_in_1_2;
      end else if (10'h6f == _T_19[9:0]) begin
        image_1_111 <= io_pixelVal_in_1_1;
      end else if (10'h6f == _T_15[9:0]) begin
        image_1_111 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_112 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h70 == _T_37[9:0]) begin
        image_1_112 <= io_pixelVal_in_1_7;
      end else if (10'h70 == _T_34[9:0]) begin
        image_1_112 <= io_pixelVal_in_1_6;
      end else if (10'h70 == _T_31[9:0]) begin
        image_1_112 <= io_pixelVal_in_1_5;
      end else if (10'h70 == _T_28[9:0]) begin
        image_1_112 <= io_pixelVal_in_1_4;
      end else if (10'h70 == _T_25[9:0]) begin
        image_1_112 <= io_pixelVal_in_1_3;
      end else if (10'h70 == _T_22[9:0]) begin
        image_1_112 <= io_pixelVal_in_1_2;
      end else if (10'h70 == _T_19[9:0]) begin
        image_1_112 <= io_pixelVal_in_1_1;
      end else if (10'h70 == _T_15[9:0]) begin
        image_1_112 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_113 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h71 == _T_37[9:0]) begin
        image_1_113 <= io_pixelVal_in_1_7;
      end else if (10'h71 == _T_34[9:0]) begin
        image_1_113 <= io_pixelVal_in_1_6;
      end else if (10'h71 == _T_31[9:0]) begin
        image_1_113 <= io_pixelVal_in_1_5;
      end else if (10'h71 == _T_28[9:0]) begin
        image_1_113 <= io_pixelVal_in_1_4;
      end else if (10'h71 == _T_25[9:0]) begin
        image_1_113 <= io_pixelVal_in_1_3;
      end else if (10'h71 == _T_22[9:0]) begin
        image_1_113 <= io_pixelVal_in_1_2;
      end else if (10'h71 == _T_19[9:0]) begin
        image_1_113 <= io_pixelVal_in_1_1;
      end else if (10'h71 == _T_15[9:0]) begin
        image_1_113 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_114 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h72 == _T_37[9:0]) begin
        image_1_114 <= io_pixelVal_in_1_7;
      end else if (10'h72 == _T_34[9:0]) begin
        image_1_114 <= io_pixelVal_in_1_6;
      end else if (10'h72 == _T_31[9:0]) begin
        image_1_114 <= io_pixelVal_in_1_5;
      end else if (10'h72 == _T_28[9:0]) begin
        image_1_114 <= io_pixelVal_in_1_4;
      end else if (10'h72 == _T_25[9:0]) begin
        image_1_114 <= io_pixelVal_in_1_3;
      end else if (10'h72 == _T_22[9:0]) begin
        image_1_114 <= io_pixelVal_in_1_2;
      end else if (10'h72 == _T_19[9:0]) begin
        image_1_114 <= io_pixelVal_in_1_1;
      end else if (10'h72 == _T_15[9:0]) begin
        image_1_114 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_115 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h73 == _T_37[9:0]) begin
        image_1_115 <= io_pixelVal_in_1_7;
      end else if (10'h73 == _T_34[9:0]) begin
        image_1_115 <= io_pixelVal_in_1_6;
      end else if (10'h73 == _T_31[9:0]) begin
        image_1_115 <= io_pixelVal_in_1_5;
      end else if (10'h73 == _T_28[9:0]) begin
        image_1_115 <= io_pixelVal_in_1_4;
      end else if (10'h73 == _T_25[9:0]) begin
        image_1_115 <= io_pixelVal_in_1_3;
      end else if (10'h73 == _T_22[9:0]) begin
        image_1_115 <= io_pixelVal_in_1_2;
      end else if (10'h73 == _T_19[9:0]) begin
        image_1_115 <= io_pixelVal_in_1_1;
      end else if (10'h73 == _T_15[9:0]) begin
        image_1_115 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_116 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h74 == _T_37[9:0]) begin
        image_1_116 <= io_pixelVal_in_1_7;
      end else if (10'h74 == _T_34[9:0]) begin
        image_1_116 <= io_pixelVal_in_1_6;
      end else if (10'h74 == _T_31[9:0]) begin
        image_1_116 <= io_pixelVal_in_1_5;
      end else if (10'h74 == _T_28[9:0]) begin
        image_1_116 <= io_pixelVal_in_1_4;
      end else if (10'h74 == _T_25[9:0]) begin
        image_1_116 <= io_pixelVal_in_1_3;
      end else if (10'h74 == _T_22[9:0]) begin
        image_1_116 <= io_pixelVal_in_1_2;
      end else if (10'h74 == _T_19[9:0]) begin
        image_1_116 <= io_pixelVal_in_1_1;
      end else if (10'h74 == _T_15[9:0]) begin
        image_1_116 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_117 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h75 == _T_37[9:0]) begin
        image_1_117 <= io_pixelVal_in_1_7;
      end else if (10'h75 == _T_34[9:0]) begin
        image_1_117 <= io_pixelVal_in_1_6;
      end else if (10'h75 == _T_31[9:0]) begin
        image_1_117 <= io_pixelVal_in_1_5;
      end else if (10'h75 == _T_28[9:0]) begin
        image_1_117 <= io_pixelVal_in_1_4;
      end else if (10'h75 == _T_25[9:0]) begin
        image_1_117 <= io_pixelVal_in_1_3;
      end else if (10'h75 == _T_22[9:0]) begin
        image_1_117 <= io_pixelVal_in_1_2;
      end else if (10'h75 == _T_19[9:0]) begin
        image_1_117 <= io_pixelVal_in_1_1;
      end else if (10'h75 == _T_15[9:0]) begin
        image_1_117 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_118 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h76 == _T_37[9:0]) begin
        image_1_118 <= io_pixelVal_in_1_7;
      end else if (10'h76 == _T_34[9:0]) begin
        image_1_118 <= io_pixelVal_in_1_6;
      end else if (10'h76 == _T_31[9:0]) begin
        image_1_118 <= io_pixelVal_in_1_5;
      end else if (10'h76 == _T_28[9:0]) begin
        image_1_118 <= io_pixelVal_in_1_4;
      end else if (10'h76 == _T_25[9:0]) begin
        image_1_118 <= io_pixelVal_in_1_3;
      end else if (10'h76 == _T_22[9:0]) begin
        image_1_118 <= io_pixelVal_in_1_2;
      end else if (10'h76 == _T_19[9:0]) begin
        image_1_118 <= io_pixelVal_in_1_1;
      end else if (10'h76 == _T_15[9:0]) begin
        image_1_118 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_119 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h77 == _T_37[9:0]) begin
        image_1_119 <= io_pixelVal_in_1_7;
      end else if (10'h77 == _T_34[9:0]) begin
        image_1_119 <= io_pixelVal_in_1_6;
      end else if (10'h77 == _T_31[9:0]) begin
        image_1_119 <= io_pixelVal_in_1_5;
      end else if (10'h77 == _T_28[9:0]) begin
        image_1_119 <= io_pixelVal_in_1_4;
      end else if (10'h77 == _T_25[9:0]) begin
        image_1_119 <= io_pixelVal_in_1_3;
      end else if (10'h77 == _T_22[9:0]) begin
        image_1_119 <= io_pixelVal_in_1_2;
      end else if (10'h77 == _T_19[9:0]) begin
        image_1_119 <= io_pixelVal_in_1_1;
      end else if (10'h77 == _T_15[9:0]) begin
        image_1_119 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_120 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h78 == _T_37[9:0]) begin
        image_1_120 <= io_pixelVal_in_1_7;
      end else if (10'h78 == _T_34[9:0]) begin
        image_1_120 <= io_pixelVal_in_1_6;
      end else if (10'h78 == _T_31[9:0]) begin
        image_1_120 <= io_pixelVal_in_1_5;
      end else if (10'h78 == _T_28[9:0]) begin
        image_1_120 <= io_pixelVal_in_1_4;
      end else if (10'h78 == _T_25[9:0]) begin
        image_1_120 <= io_pixelVal_in_1_3;
      end else if (10'h78 == _T_22[9:0]) begin
        image_1_120 <= io_pixelVal_in_1_2;
      end else if (10'h78 == _T_19[9:0]) begin
        image_1_120 <= io_pixelVal_in_1_1;
      end else if (10'h78 == _T_15[9:0]) begin
        image_1_120 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_121 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h79 == _T_37[9:0]) begin
        image_1_121 <= io_pixelVal_in_1_7;
      end else if (10'h79 == _T_34[9:0]) begin
        image_1_121 <= io_pixelVal_in_1_6;
      end else if (10'h79 == _T_31[9:0]) begin
        image_1_121 <= io_pixelVal_in_1_5;
      end else if (10'h79 == _T_28[9:0]) begin
        image_1_121 <= io_pixelVal_in_1_4;
      end else if (10'h79 == _T_25[9:0]) begin
        image_1_121 <= io_pixelVal_in_1_3;
      end else if (10'h79 == _T_22[9:0]) begin
        image_1_121 <= io_pixelVal_in_1_2;
      end else if (10'h79 == _T_19[9:0]) begin
        image_1_121 <= io_pixelVal_in_1_1;
      end else if (10'h79 == _T_15[9:0]) begin
        image_1_121 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_122 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h7a == _T_37[9:0]) begin
        image_1_122 <= io_pixelVal_in_1_7;
      end else if (10'h7a == _T_34[9:0]) begin
        image_1_122 <= io_pixelVal_in_1_6;
      end else if (10'h7a == _T_31[9:0]) begin
        image_1_122 <= io_pixelVal_in_1_5;
      end else if (10'h7a == _T_28[9:0]) begin
        image_1_122 <= io_pixelVal_in_1_4;
      end else if (10'h7a == _T_25[9:0]) begin
        image_1_122 <= io_pixelVal_in_1_3;
      end else if (10'h7a == _T_22[9:0]) begin
        image_1_122 <= io_pixelVal_in_1_2;
      end else if (10'h7a == _T_19[9:0]) begin
        image_1_122 <= io_pixelVal_in_1_1;
      end else if (10'h7a == _T_15[9:0]) begin
        image_1_122 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_123 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h7b == _T_37[9:0]) begin
        image_1_123 <= io_pixelVal_in_1_7;
      end else if (10'h7b == _T_34[9:0]) begin
        image_1_123 <= io_pixelVal_in_1_6;
      end else if (10'h7b == _T_31[9:0]) begin
        image_1_123 <= io_pixelVal_in_1_5;
      end else if (10'h7b == _T_28[9:0]) begin
        image_1_123 <= io_pixelVal_in_1_4;
      end else if (10'h7b == _T_25[9:0]) begin
        image_1_123 <= io_pixelVal_in_1_3;
      end else if (10'h7b == _T_22[9:0]) begin
        image_1_123 <= io_pixelVal_in_1_2;
      end else if (10'h7b == _T_19[9:0]) begin
        image_1_123 <= io_pixelVal_in_1_1;
      end else if (10'h7b == _T_15[9:0]) begin
        image_1_123 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_124 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h7c == _T_37[9:0]) begin
        image_1_124 <= io_pixelVal_in_1_7;
      end else if (10'h7c == _T_34[9:0]) begin
        image_1_124 <= io_pixelVal_in_1_6;
      end else if (10'h7c == _T_31[9:0]) begin
        image_1_124 <= io_pixelVal_in_1_5;
      end else if (10'h7c == _T_28[9:0]) begin
        image_1_124 <= io_pixelVal_in_1_4;
      end else if (10'h7c == _T_25[9:0]) begin
        image_1_124 <= io_pixelVal_in_1_3;
      end else if (10'h7c == _T_22[9:0]) begin
        image_1_124 <= io_pixelVal_in_1_2;
      end else if (10'h7c == _T_19[9:0]) begin
        image_1_124 <= io_pixelVal_in_1_1;
      end else if (10'h7c == _T_15[9:0]) begin
        image_1_124 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_125 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h7d == _T_37[9:0]) begin
        image_1_125 <= io_pixelVal_in_1_7;
      end else if (10'h7d == _T_34[9:0]) begin
        image_1_125 <= io_pixelVal_in_1_6;
      end else if (10'h7d == _T_31[9:0]) begin
        image_1_125 <= io_pixelVal_in_1_5;
      end else if (10'h7d == _T_28[9:0]) begin
        image_1_125 <= io_pixelVal_in_1_4;
      end else if (10'h7d == _T_25[9:0]) begin
        image_1_125 <= io_pixelVal_in_1_3;
      end else if (10'h7d == _T_22[9:0]) begin
        image_1_125 <= io_pixelVal_in_1_2;
      end else if (10'h7d == _T_19[9:0]) begin
        image_1_125 <= io_pixelVal_in_1_1;
      end else if (10'h7d == _T_15[9:0]) begin
        image_1_125 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_126 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h7e == _T_37[9:0]) begin
        image_1_126 <= io_pixelVal_in_1_7;
      end else if (10'h7e == _T_34[9:0]) begin
        image_1_126 <= io_pixelVal_in_1_6;
      end else if (10'h7e == _T_31[9:0]) begin
        image_1_126 <= io_pixelVal_in_1_5;
      end else if (10'h7e == _T_28[9:0]) begin
        image_1_126 <= io_pixelVal_in_1_4;
      end else if (10'h7e == _T_25[9:0]) begin
        image_1_126 <= io_pixelVal_in_1_3;
      end else if (10'h7e == _T_22[9:0]) begin
        image_1_126 <= io_pixelVal_in_1_2;
      end else if (10'h7e == _T_19[9:0]) begin
        image_1_126 <= io_pixelVal_in_1_1;
      end else if (10'h7e == _T_15[9:0]) begin
        image_1_126 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_127 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h7f == _T_37[9:0]) begin
        image_1_127 <= io_pixelVal_in_1_7;
      end else if (10'h7f == _T_34[9:0]) begin
        image_1_127 <= io_pixelVal_in_1_6;
      end else if (10'h7f == _T_31[9:0]) begin
        image_1_127 <= io_pixelVal_in_1_5;
      end else if (10'h7f == _T_28[9:0]) begin
        image_1_127 <= io_pixelVal_in_1_4;
      end else if (10'h7f == _T_25[9:0]) begin
        image_1_127 <= io_pixelVal_in_1_3;
      end else if (10'h7f == _T_22[9:0]) begin
        image_1_127 <= io_pixelVal_in_1_2;
      end else if (10'h7f == _T_19[9:0]) begin
        image_1_127 <= io_pixelVal_in_1_1;
      end else if (10'h7f == _T_15[9:0]) begin
        image_1_127 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_128 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h80 == _T_37[9:0]) begin
        image_1_128 <= io_pixelVal_in_1_7;
      end else if (10'h80 == _T_34[9:0]) begin
        image_1_128 <= io_pixelVal_in_1_6;
      end else if (10'h80 == _T_31[9:0]) begin
        image_1_128 <= io_pixelVal_in_1_5;
      end else if (10'h80 == _T_28[9:0]) begin
        image_1_128 <= io_pixelVal_in_1_4;
      end else if (10'h80 == _T_25[9:0]) begin
        image_1_128 <= io_pixelVal_in_1_3;
      end else if (10'h80 == _T_22[9:0]) begin
        image_1_128 <= io_pixelVal_in_1_2;
      end else if (10'h80 == _T_19[9:0]) begin
        image_1_128 <= io_pixelVal_in_1_1;
      end else if (10'h80 == _T_15[9:0]) begin
        image_1_128 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_129 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h81 == _T_37[9:0]) begin
        image_1_129 <= io_pixelVal_in_1_7;
      end else if (10'h81 == _T_34[9:0]) begin
        image_1_129 <= io_pixelVal_in_1_6;
      end else if (10'h81 == _T_31[9:0]) begin
        image_1_129 <= io_pixelVal_in_1_5;
      end else if (10'h81 == _T_28[9:0]) begin
        image_1_129 <= io_pixelVal_in_1_4;
      end else if (10'h81 == _T_25[9:0]) begin
        image_1_129 <= io_pixelVal_in_1_3;
      end else if (10'h81 == _T_22[9:0]) begin
        image_1_129 <= io_pixelVal_in_1_2;
      end else if (10'h81 == _T_19[9:0]) begin
        image_1_129 <= io_pixelVal_in_1_1;
      end else if (10'h81 == _T_15[9:0]) begin
        image_1_129 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_130 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h82 == _T_37[9:0]) begin
        image_1_130 <= io_pixelVal_in_1_7;
      end else if (10'h82 == _T_34[9:0]) begin
        image_1_130 <= io_pixelVal_in_1_6;
      end else if (10'h82 == _T_31[9:0]) begin
        image_1_130 <= io_pixelVal_in_1_5;
      end else if (10'h82 == _T_28[9:0]) begin
        image_1_130 <= io_pixelVal_in_1_4;
      end else if (10'h82 == _T_25[9:0]) begin
        image_1_130 <= io_pixelVal_in_1_3;
      end else if (10'h82 == _T_22[9:0]) begin
        image_1_130 <= io_pixelVal_in_1_2;
      end else if (10'h82 == _T_19[9:0]) begin
        image_1_130 <= io_pixelVal_in_1_1;
      end else if (10'h82 == _T_15[9:0]) begin
        image_1_130 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_131 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h83 == _T_37[9:0]) begin
        image_1_131 <= io_pixelVal_in_1_7;
      end else if (10'h83 == _T_34[9:0]) begin
        image_1_131 <= io_pixelVal_in_1_6;
      end else if (10'h83 == _T_31[9:0]) begin
        image_1_131 <= io_pixelVal_in_1_5;
      end else if (10'h83 == _T_28[9:0]) begin
        image_1_131 <= io_pixelVal_in_1_4;
      end else if (10'h83 == _T_25[9:0]) begin
        image_1_131 <= io_pixelVal_in_1_3;
      end else if (10'h83 == _T_22[9:0]) begin
        image_1_131 <= io_pixelVal_in_1_2;
      end else if (10'h83 == _T_19[9:0]) begin
        image_1_131 <= io_pixelVal_in_1_1;
      end else if (10'h83 == _T_15[9:0]) begin
        image_1_131 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_132 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h84 == _T_37[9:0]) begin
        image_1_132 <= io_pixelVal_in_1_7;
      end else if (10'h84 == _T_34[9:0]) begin
        image_1_132 <= io_pixelVal_in_1_6;
      end else if (10'h84 == _T_31[9:0]) begin
        image_1_132 <= io_pixelVal_in_1_5;
      end else if (10'h84 == _T_28[9:0]) begin
        image_1_132 <= io_pixelVal_in_1_4;
      end else if (10'h84 == _T_25[9:0]) begin
        image_1_132 <= io_pixelVal_in_1_3;
      end else if (10'h84 == _T_22[9:0]) begin
        image_1_132 <= io_pixelVal_in_1_2;
      end else if (10'h84 == _T_19[9:0]) begin
        image_1_132 <= io_pixelVal_in_1_1;
      end else if (10'h84 == _T_15[9:0]) begin
        image_1_132 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_133 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h85 == _T_37[9:0]) begin
        image_1_133 <= io_pixelVal_in_1_7;
      end else if (10'h85 == _T_34[9:0]) begin
        image_1_133 <= io_pixelVal_in_1_6;
      end else if (10'h85 == _T_31[9:0]) begin
        image_1_133 <= io_pixelVal_in_1_5;
      end else if (10'h85 == _T_28[9:0]) begin
        image_1_133 <= io_pixelVal_in_1_4;
      end else if (10'h85 == _T_25[9:0]) begin
        image_1_133 <= io_pixelVal_in_1_3;
      end else if (10'h85 == _T_22[9:0]) begin
        image_1_133 <= io_pixelVal_in_1_2;
      end else if (10'h85 == _T_19[9:0]) begin
        image_1_133 <= io_pixelVal_in_1_1;
      end else if (10'h85 == _T_15[9:0]) begin
        image_1_133 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_134 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h86 == _T_37[9:0]) begin
        image_1_134 <= io_pixelVal_in_1_7;
      end else if (10'h86 == _T_34[9:0]) begin
        image_1_134 <= io_pixelVal_in_1_6;
      end else if (10'h86 == _T_31[9:0]) begin
        image_1_134 <= io_pixelVal_in_1_5;
      end else if (10'h86 == _T_28[9:0]) begin
        image_1_134 <= io_pixelVal_in_1_4;
      end else if (10'h86 == _T_25[9:0]) begin
        image_1_134 <= io_pixelVal_in_1_3;
      end else if (10'h86 == _T_22[9:0]) begin
        image_1_134 <= io_pixelVal_in_1_2;
      end else if (10'h86 == _T_19[9:0]) begin
        image_1_134 <= io_pixelVal_in_1_1;
      end else if (10'h86 == _T_15[9:0]) begin
        image_1_134 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_135 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h87 == _T_37[9:0]) begin
        image_1_135 <= io_pixelVal_in_1_7;
      end else if (10'h87 == _T_34[9:0]) begin
        image_1_135 <= io_pixelVal_in_1_6;
      end else if (10'h87 == _T_31[9:0]) begin
        image_1_135 <= io_pixelVal_in_1_5;
      end else if (10'h87 == _T_28[9:0]) begin
        image_1_135 <= io_pixelVal_in_1_4;
      end else if (10'h87 == _T_25[9:0]) begin
        image_1_135 <= io_pixelVal_in_1_3;
      end else if (10'h87 == _T_22[9:0]) begin
        image_1_135 <= io_pixelVal_in_1_2;
      end else if (10'h87 == _T_19[9:0]) begin
        image_1_135 <= io_pixelVal_in_1_1;
      end else if (10'h87 == _T_15[9:0]) begin
        image_1_135 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_136 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h88 == _T_37[9:0]) begin
        image_1_136 <= io_pixelVal_in_1_7;
      end else if (10'h88 == _T_34[9:0]) begin
        image_1_136 <= io_pixelVal_in_1_6;
      end else if (10'h88 == _T_31[9:0]) begin
        image_1_136 <= io_pixelVal_in_1_5;
      end else if (10'h88 == _T_28[9:0]) begin
        image_1_136 <= io_pixelVal_in_1_4;
      end else if (10'h88 == _T_25[9:0]) begin
        image_1_136 <= io_pixelVal_in_1_3;
      end else if (10'h88 == _T_22[9:0]) begin
        image_1_136 <= io_pixelVal_in_1_2;
      end else if (10'h88 == _T_19[9:0]) begin
        image_1_136 <= io_pixelVal_in_1_1;
      end else if (10'h88 == _T_15[9:0]) begin
        image_1_136 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_137 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h89 == _T_37[9:0]) begin
        image_1_137 <= io_pixelVal_in_1_7;
      end else if (10'h89 == _T_34[9:0]) begin
        image_1_137 <= io_pixelVal_in_1_6;
      end else if (10'h89 == _T_31[9:0]) begin
        image_1_137 <= io_pixelVal_in_1_5;
      end else if (10'h89 == _T_28[9:0]) begin
        image_1_137 <= io_pixelVal_in_1_4;
      end else if (10'h89 == _T_25[9:0]) begin
        image_1_137 <= io_pixelVal_in_1_3;
      end else if (10'h89 == _T_22[9:0]) begin
        image_1_137 <= io_pixelVal_in_1_2;
      end else if (10'h89 == _T_19[9:0]) begin
        image_1_137 <= io_pixelVal_in_1_1;
      end else if (10'h89 == _T_15[9:0]) begin
        image_1_137 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_138 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h8a == _T_37[9:0]) begin
        image_1_138 <= io_pixelVal_in_1_7;
      end else if (10'h8a == _T_34[9:0]) begin
        image_1_138 <= io_pixelVal_in_1_6;
      end else if (10'h8a == _T_31[9:0]) begin
        image_1_138 <= io_pixelVal_in_1_5;
      end else if (10'h8a == _T_28[9:0]) begin
        image_1_138 <= io_pixelVal_in_1_4;
      end else if (10'h8a == _T_25[9:0]) begin
        image_1_138 <= io_pixelVal_in_1_3;
      end else if (10'h8a == _T_22[9:0]) begin
        image_1_138 <= io_pixelVal_in_1_2;
      end else if (10'h8a == _T_19[9:0]) begin
        image_1_138 <= io_pixelVal_in_1_1;
      end else if (10'h8a == _T_15[9:0]) begin
        image_1_138 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_139 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h8b == _T_37[9:0]) begin
        image_1_139 <= io_pixelVal_in_1_7;
      end else if (10'h8b == _T_34[9:0]) begin
        image_1_139 <= io_pixelVal_in_1_6;
      end else if (10'h8b == _T_31[9:0]) begin
        image_1_139 <= io_pixelVal_in_1_5;
      end else if (10'h8b == _T_28[9:0]) begin
        image_1_139 <= io_pixelVal_in_1_4;
      end else if (10'h8b == _T_25[9:0]) begin
        image_1_139 <= io_pixelVal_in_1_3;
      end else if (10'h8b == _T_22[9:0]) begin
        image_1_139 <= io_pixelVal_in_1_2;
      end else if (10'h8b == _T_19[9:0]) begin
        image_1_139 <= io_pixelVal_in_1_1;
      end else if (10'h8b == _T_15[9:0]) begin
        image_1_139 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_140 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h8c == _T_37[9:0]) begin
        image_1_140 <= io_pixelVal_in_1_7;
      end else if (10'h8c == _T_34[9:0]) begin
        image_1_140 <= io_pixelVal_in_1_6;
      end else if (10'h8c == _T_31[9:0]) begin
        image_1_140 <= io_pixelVal_in_1_5;
      end else if (10'h8c == _T_28[9:0]) begin
        image_1_140 <= io_pixelVal_in_1_4;
      end else if (10'h8c == _T_25[9:0]) begin
        image_1_140 <= io_pixelVal_in_1_3;
      end else if (10'h8c == _T_22[9:0]) begin
        image_1_140 <= io_pixelVal_in_1_2;
      end else if (10'h8c == _T_19[9:0]) begin
        image_1_140 <= io_pixelVal_in_1_1;
      end else if (10'h8c == _T_15[9:0]) begin
        image_1_140 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_141 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h8d == _T_37[9:0]) begin
        image_1_141 <= io_pixelVal_in_1_7;
      end else if (10'h8d == _T_34[9:0]) begin
        image_1_141 <= io_pixelVal_in_1_6;
      end else if (10'h8d == _T_31[9:0]) begin
        image_1_141 <= io_pixelVal_in_1_5;
      end else if (10'h8d == _T_28[9:0]) begin
        image_1_141 <= io_pixelVal_in_1_4;
      end else if (10'h8d == _T_25[9:0]) begin
        image_1_141 <= io_pixelVal_in_1_3;
      end else if (10'h8d == _T_22[9:0]) begin
        image_1_141 <= io_pixelVal_in_1_2;
      end else if (10'h8d == _T_19[9:0]) begin
        image_1_141 <= io_pixelVal_in_1_1;
      end else if (10'h8d == _T_15[9:0]) begin
        image_1_141 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_142 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h8e == _T_37[9:0]) begin
        image_1_142 <= io_pixelVal_in_1_7;
      end else if (10'h8e == _T_34[9:0]) begin
        image_1_142 <= io_pixelVal_in_1_6;
      end else if (10'h8e == _T_31[9:0]) begin
        image_1_142 <= io_pixelVal_in_1_5;
      end else if (10'h8e == _T_28[9:0]) begin
        image_1_142 <= io_pixelVal_in_1_4;
      end else if (10'h8e == _T_25[9:0]) begin
        image_1_142 <= io_pixelVal_in_1_3;
      end else if (10'h8e == _T_22[9:0]) begin
        image_1_142 <= io_pixelVal_in_1_2;
      end else if (10'h8e == _T_19[9:0]) begin
        image_1_142 <= io_pixelVal_in_1_1;
      end else if (10'h8e == _T_15[9:0]) begin
        image_1_142 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_143 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h8f == _T_37[9:0]) begin
        image_1_143 <= io_pixelVal_in_1_7;
      end else if (10'h8f == _T_34[9:0]) begin
        image_1_143 <= io_pixelVal_in_1_6;
      end else if (10'h8f == _T_31[9:0]) begin
        image_1_143 <= io_pixelVal_in_1_5;
      end else if (10'h8f == _T_28[9:0]) begin
        image_1_143 <= io_pixelVal_in_1_4;
      end else if (10'h8f == _T_25[9:0]) begin
        image_1_143 <= io_pixelVal_in_1_3;
      end else if (10'h8f == _T_22[9:0]) begin
        image_1_143 <= io_pixelVal_in_1_2;
      end else if (10'h8f == _T_19[9:0]) begin
        image_1_143 <= io_pixelVal_in_1_1;
      end else if (10'h8f == _T_15[9:0]) begin
        image_1_143 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_144 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h90 == _T_37[9:0]) begin
        image_1_144 <= io_pixelVal_in_1_7;
      end else if (10'h90 == _T_34[9:0]) begin
        image_1_144 <= io_pixelVal_in_1_6;
      end else if (10'h90 == _T_31[9:0]) begin
        image_1_144 <= io_pixelVal_in_1_5;
      end else if (10'h90 == _T_28[9:0]) begin
        image_1_144 <= io_pixelVal_in_1_4;
      end else if (10'h90 == _T_25[9:0]) begin
        image_1_144 <= io_pixelVal_in_1_3;
      end else if (10'h90 == _T_22[9:0]) begin
        image_1_144 <= io_pixelVal_in_1_2;
      end else if (10'h90 == _T_19[9:0]) begin
        image_1_144 <= io_pixelVal_in_1_1;
      end else if (10'h90 == _T_15[9:0]) begin
        image_1_144 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_145 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h91 == _T_37[9:0]) begin
        image_1_145 <= io_pixelVal_in_1_7;
      end else if (10'h91 == _T_34[9:0]) begin
        image_1_145 <= io_pixelVal_in_1_6;
      end else if (10'h91 == _T_31[9:0]) begin
        image_1_145 <= io_pixelVal_in_1_5;
      end else if (10'h91 == _T_28[9:0]) begin
        image_1_145 <= io_pixelVal_in_1_4;
      end else if (10'h91 == _T_25[9:0]) begin
        image_1_145 <= io_pixelVal_in_1_3;
      end else if (10'h91 == _T_22[9:0]) begin
        image_1_145 <= io_pixelVal_in_1_2;
      end else if (10'h91 == _T_19[9:0]) begin
        image_1_145 <= io_pixelVal_in_1_1;
      end else if (10'h91 == _T_15[9:0]) begin
        image_1_145 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_146 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h92 == _T_37[9:0]) begin
        image_1_146 <= io_pixelVal_in_1_7;
      end else if (10'h92 == _T_34[9:0]) begin
        image_1_146 <= io_pixelVal_in_1_6;
      end else if (10'h92 == _T_31[9:0]) begin
        image_1_146 <= io_pixelVal_in_1_5;
      end else if (10'h92 == _T_28[9:0]) begin
        image_1_146 <= io_pixelVal_in_1_4;
      end else if (10'h92 == _T_25[9:0]) begin
        image_1_146 <= io_pixelVal_in_1_3;
      end else if (10'h92 == _T_22[9:0]) begin
        image_1_146 <= io_pixelVal_in_1_2;
      end else if (10'h92 == _T_19[9:0]) begin
        image_1_146 <= io_pixelVal_in_1_1;
      end else if (10'h92 == _T_15[9:0]) begin
        image_1_146 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_147 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h93 == _T_37[9:0]) begin
        image_1_147 <= io_pixelVal_in_1_7;
      end else if (10'h93 == _T_34[9:0]) begin
        image_1_147 <= io_pixelVal_in_1_6;
      end else if (10'h93 == _T_31[9:0]) begin
        image_1_147 <= io_pixelVal_in_1_5;
      end else if (10'h93 == _T_28[9:0]) begin
        image_1_147 <= io_pixelVal_in_1_4;
      end else if (10'h93 == _T_25[9:0]) begin
        image_1_147 <= io_pixelVal_in_1_3;
      end else if (10'h93 == _T_22[9:0]) begin
        image_1_147 <= io_pixelVal_in_1_2;
      end else if (10'h93 == _T_19[9:0]) begin
        image_1_147 <= io_pixelVal_in_1_1;
      end else if (10'h93 == _T_15[9:0]) begin
        image_1_147 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_148 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h94 == _T_37[9:0]) begin
        image_1_148 <= io_pixelVal_in_1_7;
      end else if (10'h94 == _T_34[9:0]) begin
        image_1_148 <= io_pixelVal_in_1_6;
      end else if (10'h94 == _T_31[9:0]) begin
        image_1_148 <= io_pixelVal_in_1_5;
      end else if (10'h94 == _T_28[9:0]) begin
        image_1_148 <= io_pixelVal_in_1_4;
      end else if (10'h94 == _T_25[9:0]) begin
        image_1_148 <= io_pixelVal_in_1_3;
      end else if (10'h94 == _T_22[9:0]) begin
        image_1_148 <= io_pixelVal_in_1_2;
      end else if (10'h94 == _T_19[9:0]) begin
        image_1_148 <= io_pixelVal_in_1_1;
      end else if (10'h94 == _T_15[9:0]) begin
        image_1_148 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_149 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h95 == _T_37[9:0]) begin
        image_1_149 <= io_pixelVal_in_1_7;
      end else if (10'h95 == _T_34[9:0]) begin
        image_1_149 <= io_pixelVal_in_1_6;
      end else if (10'h95 == _T_31[9:0]) begin
        image_1_149 <= io_pixelVal_in_1_5;
      end else if (10'h95 == _T_28[9:0]) begin
        image_1_149 <= io_pixelVal_in_1_4;
      end else if (10'h95 == _T_25[9:0]) begin
        image_1_149 <= io_pixelVal_in_1_3;
      end else if (10'h95 == _T_22[9:0]) begin
        image_1_149 <= io_pixelVal_in_1_2;
      end else if (10'h95 == _T_19[9:0]) begin
        image_1_149 <= io_pixelVal_in_1_1;
      end else if (10'h95 == _T_15[9:0]) begin
        image_1_149 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_150 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h96 == _T_37[9:0]) begin
        image_1_150 <= io_pixelVal_in_1_7;
      end else if (10'h96 == _T_34[9:0]) begin
        image_1_150 <= io_pixelVal_in_1_6;
      end else if (10'h96 == _T_31[9:0]) begin
        image_1_150 <= io_pixelVal_in_1_5;
      end else if (10'h96 == _T_28[9:0]) begin
        image_1_150 <= io_pixelVal_in_1_4;
      end else if (10'h96 == _T_25[9:0]) begin
        image_1_150 <= io_pixelVal_in_1_3;
      end else if (10'h96 == _T_22[9:0]) begin
        image_1_150 <= io_pixelVal_in_1_2;
      end else if (10'h96 == _T_19[9:0]) begin
        image_1_150 <= io_pixelVal_in_1_1;
      end else if (10'h96 == _T_15[9:0]) begin
        image_1_150 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_151 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h97 == _T_37[9:0]) begin
        image_1_151 <= io_pixelVal_in_1_7;
      end else if (10'h97 == _T_34[9:0]) begin
        image_1_151 <= io_pixelVal_in_1_6;
      end else if (10'h97 == _T_31[9:0]) begin
        image_1_151 <= io_pixelVal_in_1_5;
      end else if (10'h97 == _T_28[9:0]) begin
        image_1_151 <= io_pixelVal_in_1_4;
      end else if (10'h97 == _T_25[9:0]) begin
        image_1_151 <= io_pixelVal_in_1_3;
      end else if (10'h97 == _T_22[9:0]) begin
        image_1_151 <= io_pixelVal_in_1_2;
      end else if (10'h97 == _T_19[9:0]) begin
        image_1_151 <= io_pixelVal_in_1_1;
      end else if (10'h97 == _T_15[9:0]) begin
        image_1_151 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_152 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h98 == _T_37[9:0]) begin
        image_1_152 <= io_pixelVal_in_1_7;
      end else if (10'h98 == _T_34[9:0]) begin
        image_1_152 <= io_pixelVal_in_1_6;
      end else if (10'h98 == _T_31[9:0]) begin
        image_1_152 <= io_pixelVal_in_1_5;
      end else if (10'h98 == _T_28[9:0]) begin
        image_1_152 <= io_pixelVal_in_1_4;
      end else if (10'h98 == _T_25[9:0]) begin
        image_1_152 <= io_pixelVal_in_1_3;
      end else if (10'h98 == _T_22[9:0]) begin
        image_1_152 <= io_pixelVal_in_1_2;
      end else if (10'h98 == _T_19[9:0]) begin
        image_1_152 <= io_pixelVal_in_1_1;
      end else if (10'h98 == _T_15[9:0]) begin
        image_1_152 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_153 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h99 == _T_37[9:0]) begin
        image_1_153 <= io_pixelVal_in_1_7;
      end else if (10'h99 == _T_34[9:0]) begin
        image_1_153 <= io_pixelVal_in_1_6;
      end else if (10'h99 == _T_31[9:0]) begin
        image_1_153 <= io_pixelVal_in_1_5;
      end else if (10'h99 == _T_28[9:0]) begin
        image_1_153 <= io_pixelVal_in_1_4;
      end else if (10'h99 == _T_25[9:0]) begin
        image_1_153 <= io_pixelVal_in_1_3;
      end else if (10'h99 == _T_22[9:0]) begin
        image_1_153 <= io_pixelVal_in_1_2;
      end else if (10'h99 == _T_19[9:0]) begin
        image_1_153 <= io_pixelVal_in_1_1;
      end else if (10'h99 == _T_15[9:0]) begin
        image_1_153 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_154 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h9a == _T_37[9:0]) begin
        image_1_154 <= io_pixelVal_in_1_7;
      end else if (10'h9a == _T_34[9:0]) begin
        image_1_154 <= io_pixelVal_in_1_6;
      end else if (10'h9a == _T_31[9:0]) begin
        image_1_154 <= io_pixelVal_in_1_5;
      end else if (10'h9a == _T_28[9:0]) begin
        image_1_154 <= io_pixelVal_in_1_4;
      end else if (10'h9a == _T_25[9:0]) begin
        image_1_154 <= io_pixelVal_in_1_3;
      end else if (10'h9a == _T_22[9:0]) begin
        image_1_154 <= io_pixelVal_in_1_2;
      end else if (10'h9a == _T_19[9:0]) begin
        image_1_154 <= io_pixelVal_in_1_1;
      end else if (10'h9a == _T_15[9:0]) begin
        image_1_154 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_155 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h9b == _T_37[9:0]) begin
        image_1_155 <= io_pixelVal_in_1_7;
      end else if (10'h9b == _T_34[9:0]) begin
        image_1_155 <= io_pixelVal_in_1_6;
      end else if (10'h9b == _T_31[9:0]) begin
        image_1_155 <= io_pixelVal_in_1_5;
      end else if (10'h9b == _T_28[9:0]) begin
        image_1_155 <= io_pixelVal_in_1_4;
      end else if (10'h9b == _T_25[9:0]) begin
        image_1_155 <= io_pixelVal_in_1_3;
      end else if (10'h9b == _T_22[9:0]) begin
        image_1_155 <= io_pixelVal_in_1_2;
      end else if (10'h9b == _T_19[9:0]) begin
        image_1_155 <= io_pixelVal_in_1_1;
      end else if (10'h9b == _T_15[9:0]) begin
        image_1_155 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_156 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h9c == _T_37[9:0]) begin
        image_1_156 <= io_pixelVal_in_1_7;
      end else if (10'h9c == _T_34[9:0]) begin
        image_1_156 <= io_pixelVal_in_1_6;
      end else if (10'h9c == _T_31[9:0]) begin
        image_1_156 <= io_pixelVal_in_1_5;
      end else if (10'h9c == _T_28[9:0]) begin
        image_1_156 <= io_pixelVal_in_1_4;
      end else if (10'h9c == _T_25[9:0]) begin
        image_1_156 <= io_pixelVal_in_1_3;
      end else if (10'h9c == _T_22[9:0]) begin
        image_1_156 <= io_pixelVal_in_1_2;
      end else if (10'h9c == _T_19[9:0]) begin
        image_1_156 <= io_pixelVal_in_1_1;
      end else if (10'h9c == _T_15[9:0]) begin
        image_1_156 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_157 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h9d == _T_37[9:0]) begin
        image_1_157 <= io_pixelVal_in_1_7;
      end else if (10'h9d == _T_34[9:0]) begin
        image_1_157 <= io_pixelVal_in_1_6;
      end else if (10'h9d == _T_31[9:0]) begin
        image_1_157 <= io_pixelVal_in_1_5;
      end else if (10'h9d == _T_28[9:0]) begin
        image_1_157 <= io_pixelVal_in_1_4;
      end else if (10'h9d == _T_25[9:0]) begin
        image_1_157 <= io_pixelVal_in_1_3;
      end else if (10'h9d == _T_22[9:0]) begin
        image_1_157 <= io_pixelVal_in_1_2;
      end else if (10'h9d == _T_19[9:0]) begin
        image_1_157 <= io_pixelVal_in_1_1;
      end else if (10'h9d == _T_15[9:0]) begin
        image_1_157 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_158 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h9e == _T_37[9:0]) begin
        image_1_158 <= io_pixelVal_in_1_7;
      end else if (10'h9e == _T_34[9:0]) begin
        image_1_158 <= io_pixelVal_in_1_6;
      end else if (10'h9e == _T_31[9:0]) begin
        image_1_158 <= io_pixelVal_in_1_5;
      end else if (10'h9e == _T_28[9:0]) begin
        image_1_158 <= io_pixelVal_in_1_4;
      end else if (10'h9e == _T_25[9:0]) begin
        image_1_158 <= io_pixelVal_in_1_3;
      end else if (10'h9e == _T_22[9:0]) begin
        image_1_158 <= io_pixelVal_in_1_2;
      end else if (10'h9e == _T_19[9:0]) begin
        image_1_158 <= io_pixelVal_in_1_1;
      end else if (10'h9e == _T_15[9:0]) begin
        image_1_158 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_159 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h9f == _T_37[9:0]) begin
        image_1_159 <= io_pixelVal_in_1_7;
      end else if (10'h9f == _T_34[9:0]) begin
        image_1_159 <= io_pixelVal_in_1_6;
      end else if (10'h9f == _T_31[9:0]) begin
        image_1_159 <= io_pixelVal_in_1_5;
      end else if (10'h9f == _T_28[9:0]) begin
        image_1_159 <= io_pixelVal_in_1_4;
      end else if (10'h9f == _T_25[9:0]) begin
        image_1_159 <= io_pixelVal_in_1_3;
      end else if (10'h9f == _T_22[9:0]) begin
        image_1_159 <= io_pixelVal_in_1_2;
      end else if (10'h9f == _T_19[9:0]) begin
        image_1_159 <= io_pixelVal_in_1_1;
      end else if (10'h9f == _T_15[9:0]) begin
        image_1_159 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_160 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha0 == _T_37[9:0]) begin
        image_1_160 <= io_pixelVal_in_1_7;
      end else if (10'ha0 == _T_34[9:0]) begin
        image_1_160 <= io_pixelVal_in_1_6;
      end else if (10'ha0 == _T_31[9:0]) begin
        image_1_160 <= io_pixelVal_in_1_5;
      end else if (10'ha0 == _T_28[9:0]) begin
        image_1_160 <= io_pixelVal_in_1_4;
      end else if (10'ha0 == _T_25[9:0]) begin
        image_1_160 <= io_pixelVal_in_1_3;
      end else if (10'ha0 == _T_22[9:0]) begin
        image_1_160 <= io_pixelVal_in_1_2;
      end else if (10'ha0 == _T_19[9:0]) begin
        image_1_160 <= io_pixelVal_in_1_1;
      end else if (10'ha0 == _T_15[9:0]) begin
        image_1_160 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_161 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha1 == _T_37[9:0]) begin
        image_1_161 <= io_pixelVal_in_1_7;
      end else if (10'ha1 == _T_34[9:0]) begin
        image_1_161 <= io_pixelVal_in_1_6;
      end else if (10'ha1 == _T_31[9:0]) begin
        image_1_161 <= io_pixelVal_in_1_5;
      end else if (10'ha1 == _T_28[9:0]) begin
        image_1_161 <= io_pixelVal_in_1_4;
      end else if (10'ha1 == _T_25[9:0]) begin
        image_1_161 <= io_pixelVal_in_1_3;
      end else if (10'ha1 == _T_22[9:0]) begin
        image_1_161 <= io_pixelVal_in_1_2;
      end else if (10'ha1 == _T_19[9:0]) begin
        image_1_161 <= io_pixelVal_in_1_1;
      end else if (10'ha1 == _T_15[9:0]) begin
        image_1_161 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_162 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha2 == _T_37[9:0]) begin
        image_1_162 <= io_pixelVal_in_1_7;
      end else if (10'ha2 == _T_34[9:0]) begin
        image_1_162 <= io_pixelVal_in_1_6;
      end else if (10'ha2 == _T_31[9:0]) begin
        image_1_162 <= io_pixelVal_in_1_5;
      end else if (10'ha2 == _T_28[9:0]) begin
        image_1_162 <= io_pixelVal_in_1_4;
      end else if (10'ha2 == _T_25[9:0]) begin
        image_1_162 <= io_pixelVal_in_1_3;
      end else if (10'ha2 == _T_22[9:0]) begin
        image_1_162 <= io_pixelVal_in_1_2;
      end else if (10'ha2 == _T_19[9:0]) begin
        image_1_162 <= io_pixelVal_in_1_1;
      end else if (10'ha2 == _T_15[9:0]) begin
        image_1_162 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_163 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha3 == _T_37[9:0]) begin
        image_1_163 <= io_pixelVal_in_1_7;
      end else if (10'ha3 == _T_34[9:0]) begin
        image_1_163 <= io_pixelVal_in_1_6;
      end else if (10'ha3 == _T_31[9:0]) begin
        image_1_163 <= io_pixelVal_in_1_5;
      end else if (10'ha3 == _T_28[9:0]) begin
        image_1_163 <= io_pixelVal_in_1_4;
      end else if (10'ha3 == _T_25[9:0]) begin
        image_1_163 <= io_pixelVal_in_1_3;
      end else if (10'ha3 == _T_22[9:0]) begin
        image_1_163 <= io_pixelVal_in_1_2;
      end else if (10'ha3 == _T_19[9:0]) begin
        image_1_163 <= io_pixelVal_in_1_1;
      end else if (10'ha3 == _T_15[9:0]) begin
        image_1_163 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_164 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha4 == _T_37[9:0]) begin
        image_1_164 <= io_pixelVal_in_1_7;
      end else if (10'ha4 == _T_34[9:0]) begin
        image_1_164 <= io_pixelVal_in_1_6;
      end else if (10'ha4 == _T_31[9:0]) begin
        image_1_164 <= io_pixelVal_in_1_5;
      end else if (10'ha4 == _T_28[9:0]) begin
        image_1_164 <= io_pixelVal_in_1_4;
      end else if (10'ha4 == _T_25[9:0]) begin
        image_1_164 <= io_pixelVal_in_1_3;
      end else if (10'ha4 == _T_22[9:0]) begin
        image_1_164 <= io_pixelVal_in_1_2;
      end else if (10'ha4 == _T_19[9:0]) begin
        image_1_164 <= io_pixelVal_in_1_1;
      end else if (10'ha4 == _T_15[9:0]) begin
        image_1_164 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_165 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha5 == _T_37[9:0]) begin
        image_1_165 <= io_pixelVal_in_1_7;
      end else if (10'ha5 == _T_34[9:0]) begin
        image_1_165 <= io_pixelVal_in_1_6;
      end else if (10'ha5 == _T_31[9:0]) begin
        image_1_165 <= io_pixelVal_in_1_5;
      end else if (10'ha5 == _T_28[9:0]) begin
        image_1_165 <= io_pixelVal_in_1_4;
      end else if (10'ha5 == _T_25[9:0]) begin
        image_1_165 <= io_pixelVal_in_1_3;
      end else if (10'ha5 == _T_22[9:0]) begin
        image_1_165 <= io_pixelVal_in_1_2;
      end else if (10'ha5 == _T_19[9:0]) begin
        image_1_165 <= io_pixelVal_in_1_1;
      end else if (10'ha5 == _T_15[9:0]) begin
        image_1_165 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_166 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha6 == _T_37[9:0]) begin
        image_1_166 <= io_pixelVal_in_1_7;
      end else if (10'ha6 == _T_34[9:0]) begin
        image_1_166 <= io_pixelVal_in_1_6;
      end else if (10'ha6 == _T_31[9:0]) begin
        image_1_166 <= io_pixelVal_in_1_5;
      end else if (10'ha6 == _T_28[9:0]) begin
        image_1_166 <= io_pixelVal_in_1_4;
      end else if (10'ha6 == _T_25[9:0]) begin
        image_1_166 <= io_pixelVal_in_1_3;
      end else if (10'ha6 == _T_22[9:0]) begin
        image_1_166 <= io_pixelVal_in_1_2;
      end else if (10'ha6 == _T_19[9:0]) begin
        image_1_166 <= io_pixelVal_in_1_1;
      end else if (10'ha6 == _T_15[9:0]) begin
        image_1_166 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_167 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha7 == _T_37[9:0]) begin
        image_1_167 <= io_pixelVal_in_1_7;
      end else if (10'ha7 == _T_34[9:0]) begin
        image_1_167 <= io_pixelVal_in_1_6;
      end else if (10'ha7 == _T_31[9:0]) begin
        image_1_167 <= io_pixelVal_in_1_5;
      end else if (10'ha7 == _T_28[9:0]) begin
        image_1_167 <= io_pixelVal_in_1_4;
      end else if (10'ha7 == _T_25[9:0]) begin
        image_1_167 <= io_pixelVal_in_1_3;
      end else if (10'ha7 == _T_22[9:0]) begin
        image_1_167 <= io_pixelVal_in_1_2;
      end else if (10'ha7 == _T_19[9:0]) begin
        image_1_167 <= io_pixelVal_in_1_1;
      end else if (10'ha7 == _T_15[9:0]) begin
        image_1_167 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_168 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha8 == _T_37[9:0]) begin
        image_1_168 <= io_pixelVal_in_1_7;
      end else if (10'ha8 == _T_34[9:0]) begin
        image_1_168 <= io_pixelVal_in_1_6;
      end else if (10'ha8 == _T_31[9:0]) begin
        image_1_168 <= io_pixelVal_in_1_5;
      end else if (10'ha8 == _T_28[9:0]) begin
        image_1_168 <= io_pixelVal_in_1_4;
      end else if (10'ha8 == _T_25[9:0]) begin
        image_1_168 <= io_pixelVal_in_1_3;
      end else if (10'ha8 == _T_22[9:0]) begin
        image_1_168 <= io_pixelVal_in_1_2;
      end else if (10'ha8 == _T_19[9:0]) begin
        image_1_168 <= io_pixelVal_in_1_1;
      end else if (10'ha8 == _T_15[9:0]) begin
        image_1_168 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_169 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha9 == _T_37[9:0]) begin
        image_1_169 <= io_pixelVal_in_1_7;
      end else if (10'ha9 == _T_34[9:0]) begin
        image_1_169 <= io_pixelVal_in_1_6;
      end else if (10'ha9 == _T_31[9:0]) begin
        image_1_169 <= io_pixelVal_in_1_5;
      end else if (10'ha9 == _T_28[9:0]) begin
        image_1_169 <= io_pixelVal_in_1_4;
      end else if (10'ha9 == _T_25[9:0]) begin
        image_1_169 <= io_pixelVal_in_1_3;
      end else if (10'ha9 == _T_22[9:0]) begin
        image_1_169 <= io_pixelVal_in_1_2;
      end else if (10'ha9 == _T_19[9:0]) begin
        image_1_169 <= io_pixelVal_in_1_1;
      end else if (10'ha9 == _T_15[9:0]) begin
        image_1_169 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_170 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'haa == _T_37[9:0]) begin
        image_1_170 <= io_pixelVal_in_1_7;
      end else if (10'haa == _T_34[9:0]) begin
        image_1_170 <= io_pixelVal_in_1_6;
      end else if (10'haa == _T_31[9:0]) begin
        image_1_170 <= io_pixelVal_in_1_5;
      end else if (10'haa == _T_28[9:0]) begin
        image_1_170 <= io_pixelVal_in_1_4;
      end else if (10'haa == _T_25[9:0]) begin
        image_1_170 <= io_pixelVal_in_1_3;
      end else if (10'haa == _T_22[9:0]) begin
        image_1_170 <= io_pixelVal_in_1_2;
      end else if (10'haa == _T_19[9:0]) begin
        image_1_170 <= io_pixelVal_in_1_1;
      end else if (10'haa == _T_15[9:0]) begin
        image_1_170 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_171 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hab == _T_37[9:0]) begin
        image_1_171 <= io_pixelVal_in_1_7;
      end else if (10'hab == _T_34[9:0]) begin
        image_1_171 <= io_pixelVal_in_1_6;
      end else if (10'hab == _T_31[9:0]) begin
        image_1_171 <= io_pixelVal_in_1_5;
      end else if (10'hab == _T_28[9:0]) begin
        image_1_171 <= io_pixelVal_in_1_4;
      end else if (10'hab == _T_25[9:0]) begin
        image_1_171 <= io_pixelVal_in_1_3;
      end else if (10'hab == _T_22[9:0]) begin
        image_1_171 <= io_pixelVal_in_1_2;
      end else if (10'hab == _T_19[9:0]) begin
        image_1_171 <= io_pixelVal_in_1_1;
      end else if (10'hab == _T_15[9:0]) begin
        image_1_171 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_172 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hac == _T_37[9:0]) begin
        image_1_172 <= io_pixelVal_in_1_7;
      end else if (10'hac == _T_34[9:0]) begin
        image_1_172 <= io_pixelVal_in_1_6;
      end else if (10'hac == _T_31[9:0]) begin
        image_1_172 <= io_pixelVal_in_1_5;
      end else if (10'hac == _T_28[9:0]) begin
        image_1_172 <= io_pixelVal_in_1_4;
      end else if (10'hac == _T_25[9:0]) begin
        image_1_172 <= io_pixelVal_in_1_3;
      end else if (10'hac == _T_22[9:0]) begin
        image_1_172 <= io_pixelVal_in_1_2;
      end else if (10'hac == _T_19[9:0]) begin
        image_1_172 <= io_pixelVal_in_1_1;
      end else if (10'hac == _T_15[9:0]) begin
        image_1_172 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_173 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'had == _T_37[9:0]) begin
        image_1_173 <= io_pixelVal_in_1_7;
      end else if (10'had == _T_34[9:0]) begin
        image_1_173 <= io_pixelVal_in_1_6;
      end else if (10'had == _T_31[9:0]) begin
        image_1_173 <= io_pixelVal_in_1_5;
      end else if (10'had == _T_28[9:0]) begin
        image_1_173 <= io_pixelVal_in_1_4;
      end else if (10'had == _T_25[9:0]) begin
        image_1_173 <= io_pixelVal_in_1_3;
      end else if (10'had == _T_22[9:0]) begin
        image_1_173 <= io_pixelVal_in_1_2;
      end else if (10'had == _T_19[9:0]) begin
        image_1_173 <= io_pixelVal_in_1_1;
      end else if (10'had == _T_15[9:0]) begin
        image_1_173 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_174 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hae == _T_37[9:0]) begin
        image_1_174 <= io_pixelVal_in_1_7;
      end else if (10'hae == _T_34[9:0]) begin
        image_1_174 <= io_pixelVal_in_1_6;
      end else if (10'hae == _T_31[9:0]) begin
        image_1_174 <= io_pixelVal_in_1_5;
      end else if (10'hae == _T_28[9:0]) begin
        image_1_174 <= io_pixelVal_in_1_4;
      end else if (10'hae == _T_25[9:0]) begin
        image_1_174 <= io_pixelVal_in_1_3;
      end else if (10'hae == _T_22[9:0]) begin
        image_1_174 <= io_pixelVal_in_1_2;
      end else if (10'hae == _T_19[9:0]) begin
        image_1_174 <= io_pixelVal_in_1_1;
      end else if (10'hae == _T_15[9:0]) begin
        image_1_174 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_175 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'haf == _T_37[9:0]) begin
        image_1_175 <= io_pixelVal_in_1_7;
      end else if (10'haf == _T_34[9:0]) begin
        image_1_175 <= io_pixelVal_in_1_6;
      end else if (10'haf == _T_31[9:0]) begin
        image_1_175 <= io_pixelVal_in_1_5;
      end else if (10'haf == _T_28[9:0]) begin
        image_1_175 <= io_pixelVal_in_1_4;
      end else if (10'haf == _T_25[9:0]) begin
        image_1_175 <= io_pixelVal_in_1_3;
      end else if (10'haf == _T_22[9:0]) begin
        image_1_175 <= io_pixelVal_in_1_2;
      end else if (10'haf == _T_19[9:0]) begin
        image_1_175 <= io_pixelVal_in_1_1;
      end else if (10'haf == _T_15[9:0]) begin
        image_1_175 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_176 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb0 == _T_37[9:0]) begin
        image_1_176 <= io_pixelVal_in_1_7;
      end else if (10'hb0 == _T_34[9:0]) begin
        image_1_176 <= io_pixelVal_in_1_6;
      end else if (10'hb0 == _T_31[9:0]) begin
        image_1_176 <= io_pixelVal_in_1_5;
      end else if (10'hb0 == _T_28[9:0]) begin
        image_1_176 <= io_pixelVal_in_1_4;
      end else if (10'hb0 == _T_25[9:0]) begin
        image_1_176 <= io_pixelVal_in_1_3;
      end else if (10'hb0 == _T_22[9:0]) begin
        image_1_176 <= io_pixelVal_in_1_2;
      end else if (10'hb0 == _T_19[9:0]) begin
        image_1_176 <= io_pixelVal_in_1_1;
      end else if (10'hb0 == _T_15[9:0]) begin
        image_1_176 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_177 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb1 == _T_37[9:0]) begin
        image_1_177 <= io_pixelVal_in_1_7;
      end else if (10'hb1 == _T_34[9:0]) begin
        image_1_177 <= io_pixelVal_in_1_6;
      end else if (10'hb1 == _T_31[9:0]) begin
        image_1_177 <= io_pixelVal_in_1_5;
      end else if (10'hb1 == _T_28[9:0]) begin
        image_1_177 <= io_pixelVal_in_1_4;
      end else if (10'hb1 == _T_25[9:0]) begin
        image_1_177 <= io_pixelVal_in_1_3;
      end else if (10'hb1 == _T_22[9:0]) begin
        image_1_177 <= io_pixelVal_in_1_2;
      end else if (10'hb1 == _T_19[9:0]) begin
        image_1_177 <= io_pixelVal_in_1_1;
      end else if (10'hb1 == _T_15[9:0]) begin
        image_1_177 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_178 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb2 == _T_37[9:0]) begin
        image_1_178 <= io_pixelVal_in_1_7;
      end else if (10'hb2 == _T_34[9:0]) begin
        image_1_178 <= io_pixelVal_in_1_6;
      end else if (10'hb2 == _T_31[9:0]) begin
        image_1_178 <= io_pixelVal_in_1_5;
      end else if (10'hb2 == _T_28[9:0]) begin
        image_1_178 <= io_pixelVal_in_1_4;
      end else if (10'hb2 == _T_25[9:0]) begin
        image_1_178 <= io_pixelVal_in_1_3;
      end else if (10'hb2 == _T_22[9:0]) begin
        image_1_178 <= io_pixelVal_in_1_2;
      end else if (10'hb2 == _T_19[9:0]) begin
        image_1_178 <= io_pixelVal_in_1_1;
      end else if (10'hb2 == _T_15[9:0]) begin
        image_1_178 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_179 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb3 == _T_37[9:0]) begin
        image_1_179 <= io_pixelVal_in_1_7;
      end else if (10'hb3 == _T_34[9:0]) begin
        image_1_179 <= io_pixelVal_in_1_6;
      end else if (10'hb3 == _T_31[9:0]) begin
        image_1_179 <= io_pixelVal_in_1_5;
      end else if (10'hb3 == _T_28[9:0]) begin
        image_1_179 <= io_pixelVal_in_1_4;
      end else if (10'hb3 == _T_25[9:0]) begin
        image_1_179 <= io_pixelVal_in_1_3;
      end else if (10'hb3 == _T_22[9:0]) begin
        image_1_179 <= io_pixelVal_in_1_2;
      end else if (10'hb3 == _T_19[9:0]) begin
        image_1_179 <= io_pixelVal_in_1_1;
      end else if (10'hb3 == _T_15[9:0]) begin
        image_1_179 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_180 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb4 == _T_37[9:0]) begin
        image_1_180 <= io_pixelVal_in_1_7;
      end else if (10'hb4 == _T_34[9:0]) begin
        image_1_180 <= io_pixelVal_in_1_6;
      end else if (10'hb4 == _T_31[9:0]) begin
        image_1_180 <= io_pixelVal_in_1_5;
      end else if (10'hb4 == _T_28[9:0]) begin
        image_1_180 <= io_pixelVal_in_1_4;
      end else if (10'hb4 == _T_25[9:0]) begin
        image_1_180 <= io_pixelVal_in_1_3;
      end else if (10'hb4 == _T_22[9:0]) begin
        image_1_180 <= io_pixelVal_in_1_2;
      end else if (10'hb4 == _T_19[9:0]) begin
        image_1_180 <= io_pixelVal_in_1_1;
      end else if (10'hb4 == _T_15[9:0]) begin
        image_1_180 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_181 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb5 == _T_37[9:0]) begin
        image_1_181 <= io_pixelVal_in_1_7;
      end else if (10'hb5 == _T_34[9:0]) begin
        image_1_181 <= io_pixelVal_in_1_6;
      end else if (10'hb5 == _T_31[9:0]) begin
        image_1_181 <= io_pixelVal_in_1_5;
      end else if (10'hb5 == _T_28[9:0]) begin
        image_1_181 <= io_pixelVal_in_1_4;
      end else if (10'hb5 == _T_25[9:0]) begin
        image_1_181 <= io_pixelVal_in_1_3;
      end else if (10'hb5 == _T_22[9:0]) begin
        image_1_181 <= io_pixelVal_in_1_2;
      end else if (10'hb5 == _T_19[9:0]) begin
        image_1_181 <= io_pixelVal_in_1_1;
      end else if (10'hb5 == _T_15[9:0]) begin
        image_1_181 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_182 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb6 == _T_37[9:0]) begin
        image_1_182 <= io_pixelVal_in_1_7;
      end else if (10'hb6 == _T_34[9:0]) begin
        image_1_182 <= io_pixelVal_in_1_6;
      end else if (10'hb6 == _T_31[9:0]) begin
        image_1_182 <= io_pixelVal_in_1_5;
      end else if (10'hb6 == _T_28[9:0]) begin
        image_1_182 <= io_pixelVal_in_1_4;
      end else if (10'hb6 == _T_25[9:0]) begin
        image_1_182 <= io_pixelVal_in_1_3;
      end else if (10'hb6 == _T_22[9:0]) begin
        image_1_182 <= io_pixelVal_in_1_2;
      end else if (10'hb6 == _T_19[9:0]) begin
        image_1_182 <= io_pixelVal_in_1_1;
      end else if (10'hb6 == _T_15[9:0]) begin
        image_1_182 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_183 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb7 == _T_37[9:0]) begin
        image_1_183 <= io_pixelVal_in_1_7;
      end else if (10'hb7 == _T_34[9:0]) begin
        image_1_183 <= io_pixelVal_in_1_6;
      end else if (10'hb7 == _T_31[9:0]) begin
        image_1_183 <= io_pixelVal_in_1_5;
      end else if (10'hb7 == _T_28[9:0]) begin
        image_1_183 <= io_pixelVal_in_1_4;
      end else if (10'hb7 == _T_25[9:0]) begin
        image_1_183 <= io_pixelVal_in_1_3;
      end else if (10'hb7 == _T_22[9:0]) begin
        image_1_183 <= io_pixelVal_in_1_2;
      end else if (10'hb7 == _T_19[9:0]) begin
        image_1_183 <= io_pixelVal_in_1_1;
      end else if (10'hb7 == _T_15[9:0]) begin
        image_1_183 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_184 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb8 == _T_37[9:0]) begin
        image_1_184 <= io_pixelVal_in_1_7;
      end else if (10'hb8 == _T_34[9:0]) begin
        image_1_184 <= io_pixelVal_in_1_6;
      end else if (10'hb8 == _T_31[9:0]) begin
        image_1_184 <= io_pixelVal_in_1_5;
      end else if (10'hb8 == _T_28[9:0]) begin
        image_1_184 <= io_pixelVal_in_1_4;
      end else if (10'hb8 == _T_25[9:0]) begin
        image_1_184 <= io_pixelVal_in_1_3;
      end else if (10'hb8 == _T_22[9:0]) begin
        image_1_184 <= io_pixelVal_in_1_2;
      end else if (10'hb8 == _T_19[9:0]) begin
        image_1_184 <= io_pixelVal_in_1_1;
      end else if (10'hb8 == _T_15[9:0]) begin
        image_1_184 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_185 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb9 == _T_37[9:0]) begin
        image_1_185 <= io_pixelVal_in_1_7;
      end else if (10'hb9 == _T_34[9:0]) begin
        image_1_185 <= io_pixelVal_in_1_6;
      end else if (10'hb9 == _T_31[9:0]) begin
        image_1_185 <= io_pixelVal_in_1_5;
      end else if (10'hb9 == _T_28[9:0]) begin
        image_1_185 <= io_pixelVal_in_1_4;
      end else if (10'hb9 == _T_25[9:0]) begin
        image_1_185 <= io_pixelVal_in_1_3;
      end else if (10'hb9 == _T_22[9:0]) begin
        image_1_185 <= io_pixelVal_in_1_2;
      end else if (10'hb9 == _T_19[9:0]) begin
        image_1_185 <= io_pixelVal_in_1_1;
      end else if (10'hb9 == _T_15[9:0]) begin
        image_1_185 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_186 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hba == _T_37[9:0]) begin
        image_1_186 <= io_pixelVal_in_1_7;
      end else if (10'hba == _T_34[9:0]) begin
        image_1_186 <= io_pixelVal_in_1_6;
      end else if (10'hba == _T_31[9:0]) begin
        image_1_186 <= io_pixelVal_in_1_5;
      end else if (10'hba == _T_28[9:0]) begin
        image_1_186 <= io_pixelVal_in_1_4;
      end else if (10'hba == _T_25[9:0]) begin
        image_1_186 <= io_pixelVal_in_1_3;
      end else if (10'hba == _T_22[9:0]) begin
        image_1_186 <= io_pixelVal_in_1_2;
      end else if (10'hba == _T_19[9:0]) begin
        image_1_186 <= io_pixelVal_in_1_1;
      end else if (10'hba == _T_15[9:0]) begin
        image_1_186 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_187 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hbb == _T_37[9:0]) begin
        image_1_187 <= io_pixelVal_in_1_7;
      end else if (10'hbb == _T_34[9:0]) begin
        image_1_187 <= io_pixelVal_in_1_6;
      end else if (10'hbb == _T_31[9:0]) begin
        image_1_187 <= io_pixelVal_in_1_5;
      end else if (10'hbb == _T_28[9:0]) begin
        image_1_187 <= io_pixelVal_in_1_4;
      end else if (10'hbb == _T_25[9:0]) begin
        image_1_187 <= io_pixelVal_in_1_3;
      end else if (10'hbb == _T_22[9:0]) begin
        image_1_187 <= io_pixelVal_in_1_2;
      end else if (10'hbb == _T_19[9:0]) begin
        image_1_187 <= io_pixelVal_in_1_1;
      end else if (10'hbb == _T_15[9:0]) begin
        image_1_187 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_188 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hbc == _T_37[9:0]) begin
        image_1_188 <= io_pixelVal_in_1_7;
      end else if (10'hbc == _T_34[9:0]) begin
        image_1_188 <= io_pixelVal_in_1_6;
      end else if (10'hbc == _T_31[9:0]) begin
        image_1_188 <= io_pixelVal_in_1_5;
      end else if (10'hbc == _T_28[9:0]) begin
        image_1_188 <= io_pixelVal_in_1_4;
      end else if (10'hbc == _T_25[9:0]) begin
        image_1_188 <= io_pixelVal_in_1_3;
      end else if (10'hbc == _T_22[9:0]) begin
        image_1_188 <= io_pixelVal_in_1_2;
      end else if (10'hbc == _T_19[9:0]) begin
        image_1_188 <= io_pixelVal_in_1_1;
      end else if (10'hbc == _T_15[9:0]) begin
        image_1_188 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_189 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hbd == _T_37[9:0]) begin
        image_1_189 <= io_pixelVal_in_1_7;
      end else if (10'hbd == _T_34[9:0]) begin
        image_1_189 <= io_pixelVal_in_1_6;
      end else if (10'hbd == _T_31[9:0]) begin
        image_1_189 <= io_pixelVal_in_1_5;
      end else if (10'hbd == _T_28[9:0]) begin
        image_1_189 <= io_pixelVal_in_1_4;
      end else if (10'hbd == _T_25[9:0]) begin
        image_1_189 <= io_pixelVal_in_1_3;
      end else if (10'hbd == _T_22[9:0]) begin
        image_1_189 <= io_pixelVal_in_1_2;
      end else if (10'hbd == _T_19[9:0]) begin
        image_1_189 <= io_pixelVal_in_1_1;
      end else if (10'hbd == _T_15[9:0]) begin
        image_1_189 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_190 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hbe == _T_37[9:0]) begin
        image_1_190 <= io_pixelVal_in_1_7;
      end else if (10'hbe == _T_34[9:0]) begin
        image_1_190 <= io_pixelVal_in_1_6;
      end else if (10'hbe == _T_31[9:0]) begin
        image_1_190 <= io_pixelVal_in_1_5;
      end else if (10'hbe == _T_28[9:0]) begin
        image_1_190 <= io_pixelVal_in_1_4;
      end else if (10'hbe == _T_25[9:0]) begin
        image_1_190 <= io_pixelVal_in_1_3;
      end else if (10'hbe == _T_22[9:0]) begin
        image_1_190 <= io_pixelVal_in_1_2;
      end else if (10'hbe == _T_19[9:0]) begin
        image_1_190 <= io_pixelVal_in_1_1;
      end else if (10'hbe == _T_15[9:0]) begin
        image_1_190 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_191 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hbf == _T_37[9:0]) begin
        image_1_191 <= io_pixelVal_in_1_7;
      end else if (10'hbf == _T_34[9:0]) begin
        image_1_191 <= io_pixelVal_in_1_6;
      end else if (10'hbf == _T_31[9:0]) begin
        image_1_191 <= io_pixelVal_in_1_5;
      end else if (10'hbf == _T_28[9:0]) begin
        image_1_191 <= io_pixelVal_in_1_4;
      end else if (10'hbf == _T_25[9:0]) begin
        image_1_191 <= io_pixelVal_in_1_3;
      end else if (10'hbf == _T_22[9:0]) begin
        image_1_191 <= io_pixelVal_in_1_2;
      end else if (10'hbf == _T_19[9:0]) begin
        image_1_191 <= io_pixelVal_in_1_1;
      end else if (10'hbf == _T_15[9:0]) begin
        image_1_191 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_192 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc0 == _T_37[9:0]) begin
        image_1_192 <= io_pixelVal_in_1_7;
      end else if (10'hc0 == _T_34[9:0]) begin
        image_1_192 <= io_pixelVal_in_1_6;
      end else if (10'hc0 == _T_31[9:0]) begin
        image_1_192 <= io_pixelVal_in_1_5;
      end else if (10'hc0 == _T_28[9:0]) begin
        image_1_192 <= io_pixelVal_in_1_4;
      end else if (10'hc0 == _T_25[9:0]) begin
        image_1_192 <= io_pixelVal_in_1_3;
      end else if (10'hc0 == _T_22[9:0]) begin
        image_1_192 <= io_pixelVal_in_1_2;
      end else if (10'hc0 == _T_19[9:0]) begin
        image_1_192 <= io_pixelVal_in_1_1;
      end else if (10'hc0 == _T_15[9:0]) begin
        image_1_192 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_193 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc1 == _T_37[9:0]) begin
        image_1_193 <= io_pixelVal_in_1_7;
      end else if (10'hc1 == _T_34[9:0]) begin
        image_1_193 <= io_pixelVal_in_1_6;
      end else if (10'hc1 == _T_31[9:0]) begin
        image_1_193 <= io_pixelVal_in_1_5;
      end else if (10'hc1 == _T_28[9:0]) begin
        image_1_193 <= io_pixelVal_in_1_4;
      end else if (10'hc1 == _T_25[9:0]) begin
        image_1_193 <= io_pixelVal_in_1_3;
      end else if (10'hc1 == _T_22[9:0]) begin
        image_1_193 <= io_pixelVal_in_1_2;
      end else if (10'hc1 == _T_19[9:0]) begin
        image_1_193 <= io_pixelVal_in_1_1;
      end else if (10'hc1 == _T_15[9:0]) begin
        image_1_193 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_194 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc2 == _T_37[9:0]) begin
        image_1_194 <= io_pixelVal_in_1_7;
      end else if (10'hc2 == _T_34[9:0]) begin
        image_1_194 <= io_pixelVal_in_1_6;
      end else if (10'hc2 == _T_31[9:0]) begin
        image_1_194 <= io_pixelVal_in_1_5;
      end else if (10'hc2 == _T_28[9:0]) begin
        image_1_194 <= io_pixelVal_in_1_4;
      end else if (10'hc2 == _T_25[9:0]) begin
        image_1_194 <= io_pixelVal_in_1_3;
      end else if (10'hc2 == _T_22[9:0]) begin
        image_1_194 <= io_pixelVal_in_1_2;
      end else if (10'hc2 == _T_19[9:0]) begin
        image_1_194 <= io_pixelVal_in_1_1;
      end else if (10'hc2 == _T_15[9:0]) begin
        image_1_194 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_195 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc3 == _T_37[9:0]) begin
        image_1_195 <= io_pixelVal_in_1_7;
      end else if (10'hc3 == _T_34[9:0]) begin
        image_1_195 <= io_pixelVal_in_1_6;
      end else if (10'hc3 == _T_31[9:0]) begin
        image_1_195 <= io_pixelVal_in_1_5;
      end else if (10'hc3 == _T_28[9:0]) begin
        image_1_195 <= io_pixelVal_in_1_4;
      end else if (10'hc3 == _T_25[9:0]) begin
        image_1_195 <= io_pixelVal_in_1_3;
      end else if (10'hc3 == _T_22[9:0]) begin
        image_1_195 <= io_pixelVal_in_1_2;
      end else if (10'hc3 == _T_19[9:0]) begin
        image_1_195 <= io_pixelVal_in_1_1;
      end else if (10'hc3 == _T_15[9:0]) begin
        image_1_195 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_196 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc4 == _T_37[9:0]) begin
        image_1_196 <= io_pixelVal_in_1_7;
      end else if (10'hc4 == _T_34[9:0]) begin
        image_1_196 <= io_pixelVal_in_1_6;
      end else if (10'hc4 == _T_31[9:0]) begin
        image_1_196 <= io_pixelVal_in_1_5;
      end else if (10'hc4 == _T_28[9:0]) begin
        image_1_196 <= io_pixelVal_in_1_4;
      end else if (10'hc4 == _T_25[9:0]) begin
        image_1_196 <= io_pixelVal_in_1_3;
      end else if (10'hc4 == _T_22[9:0]) begin
        image_1_196 <= io_pixelVal_in_1_2;
      end else if (10'hc4 == _T_19[9:0]) begin
        image_1_196 <= io_pixelVal_in_1_1;
      end else if (10'hc4 == _T_15[9:0]) begin
        image_1_196 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_197 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc5 == _T_37[9:0]) begin
        image_1_197 <= io_pixelVal_in_1_7;
      end else if (10'hc5 == _T_34[9:0]) begin
        image_1_197 <= io_pixelVal_in_1_6;
      end else if (10'hc5 == _T_31[9:0]) begin
        image_1_197 <= io_pixelVal_in_1_5;
      end else if (10'hc5 == _T_28[9:0]) begin
        image_1_197 <= io_pixelVal_in_1_4;
      end else if (10'hc5 == _T_25[9:0]) begin
        image_1_197 <= io_pixelVal_in_1_3;
      end else if (10'hc5 == _T_22[9:0]) begin
        image_1_197 <= io_pixelVal_in_1_2;
      end else if (10'hc5 == _T_19[9:0]) begin
        image_1_197 <= io_pixelVal_in_1_1;
      end else if (10'hc5 == _T_15[9:0]) begin
        image_1_197 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_198 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc6 == _T_37[9:0]) begin
        image_1_198 <= io_pixelVal_in_1_7;
      end else if (10'hc6 == _T_34[9:0]) begin
        image_1_198 <= io_pixelVal_in_1_6;
      end else if (10'hc6 == _T_31[9:0]) begin
        image_1_198 <= io_pixelVal_in_1_5;
      end else if (10'hc6 == _T_28[9:0]) begin
        image_1_198 <= io_pixelVal_in_1_4;
      end else if (10'hc6 == _T_25[9:0]) begin
        image_1_198 <= io_pixelVal_in_1_3;
      end else if (10'hc6 == _T_22[9:0]) begin
        image_1_198 <= io_pixelVal_in_1_2;
      end else if (10'hc6 == _T_19[9:0]) begin
        image_1_198 <= io_pixelVal_in_1_1;
      end else if (10'hc6 == _T_15[9:0]) begin
        image_1_198 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_199 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc7 == _T_37[9:0]) begin
        image_1_199 <= io_pixelVal_in_1_7;
      end else if (10'hc7 == _T_34[9:0]) begin
        image_1_199 <= io_pixelVal_in_1_6;
      end else if (10'hc7 == _T_31[9:0]) begin
        image_1_199 <= io_pixelVal_in_1_5;
      end else if (10'hc7 == _T_28[9:0]) begin
        image_1_199 <= io_pixelVal_in_1_4;
      end else if (10'hc7 == _T_25[9:0]) begin
        image_1_199 <= io_pixelVal_in_1_3;
      end else if (10'hc7 == _T_22[9:0]) begin
        image_1_199 <= io_pixelVal_in_1_2;
      end else if (10'hc7 == _T_19[9:0]) begin
        image_1_199 <= io_pixelVal_in_1_1;
      end else if (10'hc7 == _T_15[9:0]) begin
        image_1_199 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_200 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc8 == _T_37[9:0]) begin
        image_1_200 <= io_pixelVal_in_1_7;
      end else if (10'hc8 == _T_34[9:0]) begin
        image_1_200 <= io_pixelVal_in_1_6;
      end else if (10'hc8 == _T_31[9:0]) begin
        image_1_200 <= io_pixelVal_in_1_5;
      end else if (10'hc8 == _T_28[9:0]) begin
        image_1_200 <= io_pixelVal_in_1_4;
      end else if (10'hc8 == _T_25[9:0]) begin
        image_1_200 <= io_pixelVal_in_1_3;
      end else if (10'hc8 == _T_22[9:0]) begin
        image_1_200 <= io_pixelVal_in_1_2;
      end else if (10'hc8 == _T_19[9:0]) begin
        image_1_200 <= io_pixelVal_in_1_1;
      end else if (10'hc8 == _T_15[9:0]) begin
        image_1_200 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_201 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc9 == _T_37[9:0]) begin
        image_1_201 <= io_pixelVal_in_1_7;
      end else if (10'hc9 == _T_34[9:0]) begin
        image_1_201 <= io_pixelVal_in_1_6;
      end else if (10'hc9 == _T_31[9:0]) begin
        image_1_201 <= io_pixelVal_in_1_5;
      end else if (10'hc9 == _T_28[9:0]) begin
        image_1_201 <= io_pixelVal_in_1_4;
      end else if (10'hc9 == _T_25[9:0]) begin
        image_1_201 <= io_pixelVal_in_1_3;
      end else if (10'hc9 == _T_22[9:0]) begin
        image_1_201 <= io_pixelVal_in_1_2;
      end else if (10'hc9 == _T_19[9:0]) begin
        image_1_201 <= io_pixelVal_in_1_1;
      end else if (10'hc9 == _T_15[9:0]) begin
        image_1_201 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_202 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hca == _T_37[9:0]) begin
        image_1_202 <= io_pixelVal_in_1_7;
      end else if (10'hca == _T_34[9:0]) begin
        image_1_202 <= io_pixelVal_in_1_6;
      end else if (10'hca == _T_31[9:0]) begin
        image_1_202 <= io_pixelVal_in_1_5;
      end else if (10'hca == _T_28[9:0]) begin
        image_1_202 <= io_pixelVal_in_1_4;
      end else if (10'hca == _T_25[9:0]) begin
        image_1_202 <= io_pixelVal_in_1_3;
      end else if (10'hca == _T_22[9:0]) begin
        image_1_202 <= io_pixelVal_in_1_2;
      end else if (10'hca == _T_19[9:0]) begin
        image_1_202 <= io_pixelVal_in_1_1;
      end else if (10'hca == _T_15[9:0]) begin
        image_1_202 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_203 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hcb == _T_37[9:0]) begin
        image_1_203 <= io_pixelVal_in_1_7;
      end else if (10'hcb == _T_34[9:0]) begin
        image_1_203 <= io_pixelVal_in_1_6;
      end else if (10'hcb == _T_31[9:0]) begin
        image_1_203 <= io_pixelVal_in_1_5;
      end else if (10'hcb == _T_28[9:0]) begin
        image_1_203 <= io_pixelVal_in_1_4;
      end else if (10'hcb == _T_25[9:0]) begin
        image_1_203 <= io_pixelVal_in_1_3;
      end else if (10'hcb == _T_22[9:0]) begin
        image_1_203 <= io_pixelVal_in_1_2;
      end else if (10'hcb == _T_19[9:0]) begin
        image_1_203 <= io_pixelVal_in_1_1;
      end else if (10'hcb == _T_15[9:0]) begin
        image_1_203 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_204 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hcc == _T_37[9:0]) begin
        image_1_204 <= io_pixelVal_in_1_7;
      end else if (10'hcc == _T_34[9:0]) begin
        image_1_204 <= io_pixelVal_in_1_6;
      end else if (10'hcc == _T_31[9:0]) begin
        image_1_204 <= io_pixelVal_in_1_5;
      end else if (10'hcc == _T_28[9:0]) begin
        image_1_204 <= io_pixelVal_in_1_4;
      end else if (10'hcc == _T_25[9:0]) begin
        image_1_204 <= io_pixelVal_in_1_3;
      end else if (10'hcc == _T_22[9:0]) begin
        image_1_204 <= io_pixelVal_in_1_2;
      end else if (10'hcc == _T_19[9:0]) begin
        image_1_204 <= io_pixelVal_in_1_1;
      end else if (10'hcc == _T_15[9:0]) begin
        image_1_204 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_205 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hcd == _T_37[9:0]) begin
        image_1_205 <= io_pixelVal_in_1_7;
      end else if (10'hcd == _T_34[9:0]) begin
        image_1_205 <= io_pixelVal_in_1_6;
      end else if (10'hcd == _T_31[9:0]) begin
        image_1_205 <= io_pixelVal_in_1_5;
      end else if (10'hcd == _T_28[9:0]) begin
        image_1_205 <= io_pixelVal_in_1_4;
      end else if (10'hcd == _T_25[9:0]) begin
        image_1_205 <= io_pixelVal_in_1_3;
      end else if (10'hcd == _T_22[9:0]) begin
        image_1_205 <= io_pixelVal_in_1_2;
      end else if (10'hcd == _T_19[9:0]) begin
        image_1_205 <= io_pixelVal_in_1_1;
      end else if (10'hcd == _T_15[9:0]) begin
        image_1_205 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_206 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hce == _T_37[9:0]) begin
        image_1_206 <= io_pixelVal_in_1_7;
      end else if (10'hce == _T_34[9:0]) begin
        image_1_206 <= io_pixelVal_in_1_6;
      end else if (10'hce == _T_31[9:0]) begin
        image_1_206 <= io_pixelVal_in_1_5;
      end else if (10'hce == _T_28[9:0]) begin
        image_1_206 <= io_pixelVal_in_1_4;
      end else if (10'hce == _T_25[9:0]) begin
        image_1_206 <= io_pixelVal_in_1_3;
      end else if (10'hce == _T_22[9:0]) begin
        image_1_206 <= io_pixelVal_in_1_2;
      end else if (10'hce == _T_19[9:0]) begin
        image_1_206 <= io_pixelVal_in_1_1;
      end else if (10'hce == _T_15[9:0]) begin
        image_1_206 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_207 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hcf == _T_37[9:0]) begin
        image_1_207 <= io_pixelVal_in_1_7;
      end else if (10'hcf == _T_34[9:0]) begin
        image_1_207 <= io_pixelVal_in_1_6;
      end else if (10'hcf == _T_31[9:0]) begin
        image_1_207 <= io_pixelVal_in_1_5;
      end else if (10'hcf == _T_28[9:0]) begin
        image_1_207 <= io_pixelVal_in_1_4;
      end else if (10'hcf == _T_25[9:0]) begin
        image_1_207 <= io_pixelVal_in_1_3;
      end else if (10'hcf == _T_22[9:0]) begin
        image_1_207 <= io_pixelVal_in_1_2;
      end else if (10'hcf == _T_19[9:0]) begin
        image_1_207 <= io_pixelVal_in_1_1;
      end else if (10'hcf == _T_15[9:0]) begin
        image_1_207 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_208 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd0 == _T_37[9:0]) begin
        image_1_208 <= io_pixelVal_in_1_7;
      end else if (10'hd0 == _T_34[9:0]) begin
        image_1_208 <= io_pixelVal_in_1_6;
      end else if (10'hd0 == _T_31[9:0]) begin
        image_1_208 <= io_pixelVal_in_1_5;
      end else if (10'hd0 == _T_28[9:0]) begin
        image_1_208 <= io_pixelVal_in_1_4;
      end else if (10'hd0 == _T_25[9:0]) begin
        image_1_208 <= io_pixelVal_in_1_3;
      end else if (10'hd0 == _T_22[9:0]) begin
        image_1_208 <= io_pixelVal_in_1_2;
      end else if (10'hd0 == _T_19[9:0]) begin
        image_1_208 <= io_pixelVal_in_1_1;
      end else if (10'hd0 == _T_15[9:0]) begin
        image_1_208 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_209 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd1 == _T_37[9:0]) begin
        image_1_209 <= io_pixelVal_in_1_7;
      end else if (10'hd1 == _T_34[9:0]) begin
        image_1_209 <= io_pixelVal_in_1_6;
      end else if (10'hd1 == _T_31[9:0]) begin
        image_1_209 <= io_pixelVal_in_1_5;
      end else if (10'hd1 == _T_28[9:0]) begin
        image_1_209 <= io_pixelVal_in_1_4;
      end else if (10'hd1 == _T_25[9:0]) begin
        image_1_209 <= io_pixelVal_in_1_3;
      end else if (10'hd1 == _T_22[9:0]) begin
        image_1_209 <= io_pixelVal_in_1_2;
      end else if (10'hd1 == _T_19[9:0]) begin
        image_1_209 <= io_pixelVal_in_1_1;
      end else if (10'hd1 == _T_15[9:0]) begin
        image_1_209 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_210 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd2 == _T_37[9:0]) begin
        image_1_210 <= io_pixelVal_in_1_7;
      end else if (10'hd2 == _T_34[9:0]) begin
        image_1_210 <= io_pixelVal_in_1_6;
      end else if (10'hd2 == _T_31[9:0]) begin
        image_1_210 <= io_pixelVal_in_1_5;
      end else if (10'hd2 == _T_28[9:0]) begin
        image_1_210 <= io_pixelVal_in_1_4;
      end else if (10'hd2 == _T_25[9:0]) begin
        image_1_210 <= io_pixelVal_in_1_3;
      end else if (10'hd2 == _T_22[9:0]) begin
        image_1_210 <= io_pixelVal_in_1_2;
      end else if (10'hd2 == _T_19[9:0]) begin
        image_1_210 <= io_pixelVal_in_1_1;
      end else if (10'hd2 == _T_15[9:0]) begin
        image_1_210 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_211 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd3 == _T_37[9:0]) begin
        image_1_211 <= io_pixelVal_in_1_7;
      end else if (10'hd3 == _T_34[9:0]) begin
        image_1_211 <= io_pixelVal_in_1_6;
      end else if (10'hd3 == _T_31[9:0]) begin
        image_1_211 <= io_pixelVal_in_1_5;
      end else if (10'hd3 == _T_28[9:0]) begin
        image_1_211 <= io_pixelVal_in_1_4;
      end else if (10'hd3 == _T_25[9:0]) begin
        image_1_211 <= io_pixelVal_in_1_3;
      end else if (10'hd3 == _T_22[9:0]) begin
        image_1_211 <= io_pixelVal_in_1_2;
      end else if (10'hd3 == _T_19[9:0]) begin
        image_1_211 <= io_pixelVal_in_1_1;
      end else if (10'hd3 == _T_15[9:0]) begin
        image_1_211 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_212 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd4 == _T_37[9:0]) begin
        image_1_212 <= io_pixelVal_in_1_7;
      end else if (10'hd4 == _T_34[9:0]) begin
        image_1_212 <= io_pixelVal_in_1_6;
      end else if (10'hd4 == _T_31[9:0]) begin
        image_1_212 <= io_pixelVal_in_1_5;
      end else if (10'hd4 == _T_28[9:0]) begin
        image_1_212 <= io_pixelVal_in_1_4;
      end else if (10'hd4 == _T_25[9:0]) begin
        image_1_212 <= io_pixelVal_in_1_3;
      end else if (10'hd4 == _T_22[9:0]) begin
        image_1_212 <= io_pixelVal_in_1_2;
      end else if (10'hd4 == _T_19[9:0]) begin
        image_1_212 <= io_pixelVal_in_1_1;
      end else if (10'hd4 == _T_15[9:0]) begin
        image_1_212 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_213 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd5 == _T_37[9:0]) begin
        image_1_213 <= io_pixelVal_in_1_7;
      end else if (10'hd5 == _T_34[9:0]) begin
        image_1_213 <= io_pixelVal_in_1_6;
      end else if (10'hd5 == _T_31[9:0]) begin
        image_1_213 <= io_pixelVal_in_1_5;
      end else if (10'hd5 == _T_28[9:0]) begin
        image_1_213 <= io_pixelVal_in_1_4;
      end else if (10'hd5 == _T_25[9:0]) begin
        image_1_213 <= io_pixelVal_in_1_3;
      end else if (10'hd5 == _T_22[9:0]) begin
        image_1_213 <= io_pixelVal_in_1_2;
      end else if (10'hd5 == _T_19[9:0]) begin
        image_1_213 <= io_pixelVal_in_1_1;
      end else if (10'hd5 == _T_15[9:0]) begin
        image_1_213 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_214 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd6 == _T_37[9:0]) begin
        image_1_214 <= io_pixelVal_in_1_7;
      end else if (10'hd6 == _T_34[9:0]) begin
        image_1_214 <= io_pixelVal_in_1_6;
      end else if (10'hd6 == _T_31[9:0]) begin
        image_1_214 <= io_pixelVal_in_1_5;
      end else if (10'hd6 == _T_28[9:0]) begin
        image_1_214 <= io_pixelVal_in_1_4;
      end else if (10'hd6 == _T_25[9:0]) begin
        image_1_214 <= io_pixelVal_in_1_3;
      end else if (10'hd6 == _T_22[9:0]) begin
        image_1_214 <= io_pixelVal_in_1_2;
      end else if (10'hd6 == _T_19[9:0]) begin
        image_1_214 <= io_pixelVal_in_1_1;
      end else if (10'hd6 == _T_15[9:0]) begin
        image_1_214 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_215 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd7 == _T_37[9:0]) begin
        image_1_215 <= io_pixelVal_in_1_7;
      end else if (10'hd7 == _T_34[9:0]) begin
        image_1_215 <= io_pixelVal_in_1_6;
      end else if (10'hd7 == _T_31[9:0]) begin
        image_1_215 <= io_pixelVal_in_1_5;
      end else if (10'hd7 == _T_28[9:0]) begin
        image_1_215 <= io_pixelVal_in_1_4;
      end else if (10'hd7 == _T_25[9:0]) begin
        image_1_215 <= io_pixelVal_in_1_3;
      end else if (10'hd7 == _T_22[9:0]) begin
        image_1_215 <= io_pixelVal_in_1_2;
      end else if (10'hd7 == _T_19[9:0]) begin
        image_1_215 <= io_pixelVal_in_1_1;
      end else if (10'hd7 == _T_15[9:0]) begin
        image_1_215 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_216 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd8 == _T_37[9:0]) begin
        image_1_216 <= io_pixelVal_in_1_7;
      end else if (10'hd8 == _T_34[9:0]) begin
        image_1_216 <= io_pixelVal_in_1_6;
      end else if (10'hd8 == _T_31[9:0]) begin
        image_1_216 <= io_pixelVal_in_1_5;
      end else if (10'hd8 == _T_28[9:0]) begin
        image_1_216 <= io_pixelVal_in_1_4;
      end else if (10'hd8 == _T_25[9:0]) begin
        image_1_216 <= io_pixelVal_in_1_3;
      end else if (10'hd8 == _T_22[9:0]) begin
        image_1_216 <= io_pixelVal_in_1_2;
      end else if (10'hd8 == _T_19[9:0]) begin
        image_1_216 <= io_pixelVal_in_1_1;
      end else if (10'hd8 == _T_15[9:0]) begin
        image_1_216 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_217 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd9 == _T_37[9:0]) begin
        image_1_217 <= io_pixelVal_in_1_7;
      end else if (10'hd9 == _T_34[9:0]) begin
        image_1_217 <= io_pixelVal_in_1_6;
      end else if (10'hd9 == _T_31[9:0]) begin
        image_1_217 <= io_pixelVal_in_1_5;
      end else if (10'hd9 == _T_28[9:0]) begin
        image_1_217 <= io_pixelVal_in_1_4;
      end else if (10'hd9 == _T_25[9:0]) begin
        image_1_217 <= io_pixelVal_in_1_3;
      end else if (10'hd9 == _T_22[9:0]) begin
        image_1_217 <= io_pixelVal_in_1_2;
      end else if (10'hd9 == _T_19[9:0]) begin
        image_1_217 <= io_pixelVal_in_1_1;
      end else if (10'hd9 == _T_15[9:0]) begin
        image_1_217 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_218 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hda == _T_37[9:0]) begin
        image_1_218 <= io_pixelVal_in_1_7;
      end else if (10'hda == _T_34[9:0]) begin
        image_1_218 <= io_pixelVal_in_1_6;
      end else if (10'hda == _T_31[9:0]) begin
        image_1_218 <= io_pixelVal_in_1_5;
      end else if (10'hda == _T_28[9:0]) begin
        image_1_218 <= io_pixelVal_in_1_4;
      end else if (10'hda == _T_25[9:0]) begin
        image_1_218 <= io_pixelVal_in_1_3;
      end else if (10'hda == _T_22[9:0]) begin
        image_1_218 <= io_pixelVal_in_1_2;
      end else if (10'hda == _T_19[9:0]) begin
        image_1_218 <= io_pixelVal_in_1_1;
      end else if (10'hda == _T_15[9:0]) begin
        image_1_218 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_219 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hdb == _T_37[9:0]) begin
        image_1_219 <= io_pixelVal_in_1_7;
      end else if (10'hdb == _T_34[9:0]) begin
        image_1_219 <= io_pixelVal_in_1_6;
      end else if (10'hdb == _T_31[9:0]) begin
        image_1_219 <= io_pixelVal_in_1_5;
      end else if (10'hdb == _T_28[9:0]) begin
        image_1_219 <= io_pixelVal_in_1_4;
      end else if (10'hdb == _T_25[9:0]) begin
        image_1_219 <= io_pixelVal_in_1_3;
      end else if (10'hdb == _T_22[9:0]) begin
        image_1_219 <= io_pixelVal_in_1_2;
      end else if (10'hdb == _T_19[9:0]) begin
        image_1_219 <= io_pixelVal_in_1_1;
      end else if (10'hdb == _T_15[9:0]) begin
        image_1_219 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_220 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hdc == _T_37[9:0]) begin
        image_1_220 <= io_pixelVal_in_1_7;
      end else if (10'hdc == _T_34[9:0]) begin
        image_1_220 <= io_pixelVal_in_1_6;
      end else if (10'hdc == _T_31[9:0]) begin
        image_1_220 <= io_pixelVal_in_1_5;
      end else if (10'hdc == _T_28[9:0]) begin
        image_1_220 <= io_pixelVal_in_1_4;
      end else if (10'hdc == _T_25[9:0]) begin
        image_1_220 <= io_pixelVal_in_1_3;
      end else if (10'hdc == _T_22[9:0]) begin
        image_1_220 <= io_pixelVal_in_1_2;
      end else if (10'hdc == _T_19[9:0]) begin
        image_1_220 <= io_pixelVal_in_1_1;
      end else if (10'hdc == _T_15[9:0]) begin
        image_1_220 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_221 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hdd == _T_37[9:0]) begin
        image_1_221 <= io_pixelVal_in_1_7;
      end else if (10'hdd == _T_34[9:0]) begin
        image_1_221 <= io_pixelVal_in_1_6;
      end else if (10'hdd == _T_31[9:0]) begin
        image_1_221 <= io_pixelVal_in_1_5;
      end else if (10'hdd == _T_28[9:0]) begin
        image_1_221 <= io_pixelVal_in_1_4;
      end else if (10'hdd == _T_25[9:0]) begin
        image_1_221 <= io_pixelVal_in_1_3;
      end else if (10'hdd == _T_22[9:0]) begin
        image_1_221 <= io_pixelVal_in_1_2;
      end else if (10'hdd == _T_19[9:0]) begin
        image_1_221 <= io_pixelVal_in_1_1;
      end else if (10'hdd == _T_15[9:0]) begin
        image_1_221 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_222 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hde == _T_37[9:0]) begin
        image_1_222 <= io_pixelVal_in_1_7;
      end else if (10'hde == _T_34[9:0]) begin
        image_1_222 <= io_pixelVal_in_1_6;
      end else if (10'hde == _T_31[9:0]) begin
        image_1_222 <= io_pixelVal_in_1_5;
      end else if (10'hde == _T_28[9:0]) begin
        image_1_222 <= io_pixelVal_in_1_4;
      end else if (10'hde == _T_25[9:0]) begin
        image_1_222 <= io_pixelVal_in_1_3;
      end else if (10'hde == _T_22[9:0]) begin
        image_1_222 <= io_pixelVal_in_1_2;
      end else if (10'hde == _T_19[9:0]) begin
        image_1_222 <= io_pixelVal_in_1_1;
      end else if (10'hde == _T_15[9:0]) begin
        image_1_222 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_223 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hdf == _T_37[9:0]) begin
        image_1_223 <= io_pixelVal_in_1_7;
      end else if (10'hdf == _T_34[9:0]) begin
        image_1_223 <= io_pixelVal_in_1_6;
      end else if (10'hdf == _T_31[9:0]) begin
        image_1_223 <= io_pixelVal_in_1_5;
      end else if (10'hdf == _T_28[9:0]) begin
        image_1_223 <= io_pixelVal_in_1_4;
      end else if (10'hdf == _T_25[9:0]) begin
        image_1_223 <= io_pixelVal_in_1_3;
      end else if (10'hdf == _T_22[9:0]) begin
        image_1_223 <= io_pixelVal_in_1_2;
      end else if (10'hdf == _T_19[9:0]) begin
        image_1_223 <= io_pixelVal_in_1_1;
      end else if (10'hdf == _T_15[9:0]) begin
        image_1_223 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_224 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he0 == _T_37[9:0]) begin
        image_1_224 <= io_pixelVal_in_1_7;
      end else if (10'he0 == _T_34[9:0]) begin
        image_1_224 <= io_pixelVal_in_1_6;
      end else if (10'he0 == _T_31[9:0]) begin
        image_1_224 <= io_pixelVal_in_1_5;
      end else if (10'he0 == _T_28[9:0]) begin
        image_1_224 <= io_pixelVal_in_1_4;
      end else if (10'he0 == _T_25[9:0]) begin
        image_1_224 <= io_pixelVal_in_1_3;
      end else if (10'he0 == _T_22[9:0]) begin
        image_1_224 <= io_pixelVal_in_1_2;
      end else if (10'he0 == _T_19[9:0]) begin
        image_1_224 <= io_pixelVal_in_1_1;
      end else if (10'he0 == _T_15[9:0]) begin
        image_1_224 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_225 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he1 == _T_37[9:0]) begin
        image_1_225 <= io_pixelVal_in_1_7;
      end else if (10'he1 == _T_34[9:0]) begin
        image_1_225 <= io_pixelVal_in_1_6;
      end else if (10'he1 == _T_31[9:0]) begin
        image_1_225 <= io_pixelVal_in_1_5;
      end else if (10'he1 == _T_28[9:0]) begin
        image_1_225 <= io_pixelVal_in_1_4;
      end else if (10'he1 == _T_25[9:0]) begin
        image_1_225 <= io_pixelVal_in_1_3;
      end else if (10'he1 == _T_22[9:0]) begin
        image_1_225 <= io_pixelVal_in_1_2;
      end else if (10'he1 == _T_19[9:0]) begin
        image_1_225 <= io_pixelVal_in_1_1;
      end else if (10'he1 == _T_15[9:0]) begin
        image_1_225 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_226 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he2 == _T_37[9:0]) begin
        image_1_226 <= io_pixelVal_in_1_7;
      end else if (10'he2 == _T_34[9:0]) begin
        image_1_226 <= io_pixelVal_in_1_6;
      end else if (10'he2 == _T_31[9:0]) begin
        image_1_226 <= io_pixelVal_in_1_5;
      end else if (10'he2 == _T_28[9:0]) begin
        image_1_226 <= io_pixelVal_in_1_4;
      end else if (10'he2 == _T_25[9:0]) begin
        image_1_226 <= io_pixelVal_in_1_3;
      end else if (10'he2 == _T_22[9:0]) begin
        image_1_226 <= io_pixelVal_in_1_2;
      end else if (10'he2 == _T_19[9:0]) begin
        image_1_226 <= io_pixelVal_in_1_1;
      end else if (10'he2 == _T_15[9:0]) begin
        image_1_226 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_227 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he3 == _T_37[9:0]) begin
        image_1_227 <= io_pixelVal_in_1_7;
      end else if (10'he3 == _T_34[9:0]) begin
        image_1_227 <= io_pixelVal_in_1_6;
      end else if (10'he3 == _T_31[9:0]) begin
        image_1_227 <= io_pixelVal_in_1_5;
      end else if (10'he3 == _T_28[9:0]) begin
        image_1_227 <= io_pixelVal_in_1_4;
      end else if (10'he3 == _T_25[9:0]) begin
        image_1_227 <= io_pixelVal_in_1_3;
      end else if (10'he3 == _T_22[9:0]) begin
        image_1_227 <= io_pixelVal_in_1_2;
      end else if (10'he3 == _T_19[9:0]) begin
        image_1_227 <= io_pixelVal_in_1_1;
      end else if (10'he3 == _T_15[9:0]) begin
        image_1_227 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_228 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he4 == _T_37[9:0]) begin
        image_1_228 <= io_pixelVal_in_1_7;
      end else if (10'he4 == _T_34[9:0]) begin
        image_1_228 <= io_pixelVal_in_1_6;
      end else if (10'he4 == _T_31[9:0]) begin
        image_1_228 <= io_pixelVal_in_1_5;
      end else if (10'he4 == _T_28[9:0]) begin
        image_1_228 <= io_pixelVal_in_1_4;
      end else if (10'he4 == _T_25[9:0]) begin
        image_1_228 <= io_pixelVal_in_1_3;
      end else if (10'he4 == _T_22[9:0]) begin
        image_1_228 <= io_pixelVal_in_1_2;
      end else if (10'he4 == _T_19[9:0]) begin
        image_1_228 <= io_pixelVal_in_1_1;
      end else if (10'he4 == _T_15[9:0]) begin
        image_1_228 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_229 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he5 == _T_37[9:0]) begin
        image_1_229 <= io_pixelVal_in_1_7;
      end else if (10'he5 == _T_34[9:0]) begin
        image_1_229 <= io_pixelVal_in_1_6;
      end else if (10'he5 == _T_31[9:0]) begin
        image_1_229 <= io_pixelVal_in_1_5;
      end else if (10'he5 == _T_28[9:0]) begin
        image_1_229 <= io_pixelVal_in_1_4;
      end else if (10'he5 == _T_25[9:0]) begin
        image_1_229 <= io_pixelVal_in_1_3;
      end else if (10'he5 == _T_22[9:0]) begin
        image_1_229 <= io_pixelVal_in_1_2;
      end else if (10'he5 == _T_19[9:0]) begin
        image_1_229 <= io_pixelVal_in_1_1;
      end else if (10'he5 == _T_15[9:0]) begin
        image_1_229 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_230 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he6 == _T_37[9:0]) begin
        image_1_230 <= io_pixelVal_in_1_7;
      end else if (10'he6 == _T_34[9:0]) begin
        image_1_230 <= io_pixelVal_in_1_6;
      end else if (10'he6 == _T_31[9:0]) begin
        image_1_230 <= io_pixelVal_in_1_5;
      end else if (10'he6 == _T_28[9:0]) begin
        image_1_230 <= io_pixelVal_in_1_4;
      end else if (10'he6 == _T_25[9:0]) begin
        image_1_230 <= io_pixelVal_in_1_3;
      end else if (10'he6 == _T_22[9:0]) begin
        image_1_230 <= io_pixelVal_in_1_2;
      end else if (10'he6 == _T_19[9:0]) begin
        image_1_230 <= io_pixelVal_in_1_1;
      end else if (10'he6 == _T_15[9:0]) begin
        image_1_230 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_231 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he7 == _T_37[9:0]) begin
        image_1_231 <= io_pixelVal_in_1_7;
      end else if (10'he7 == _T_34[9:0]) begin
        image_1_231 <= io_pixelVal_in_1_6;
      end else if (10'he7 == _T_31[9:0]) begin
        image_1_231 <= io_pixelVal_in_1_5;
      end else if (10'he7 == _T_28[9:0]) begin
        image_1_231 <= io_pixelVal_in_1_4;
      end else if (10'he7 == _T_25[9:0]) begin
        image_1_231 <= io_pixelVal_in_1_3;
      end else if (10'he7 == _T_22[9:0]) begin
        image_1_231 <= io_pixelVal_in_1_2;
      end else if (10'he7 == _T_19[9:0]) begin
        image_1_231 <= io_pixelVal_in_1_1;
      end else if (10'he7 == _T_15[9:0]) begin
        image_1_231 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_232 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he8 == _T_37[9:0]) begin
        image_1_232 <= io_pixelVal_in_1_7;
      end else if (10'he8 == _T_34[9:0]) begin
        image_1_232 <= io_pixelVal_in_1_6;
      end else if (10'he8 == _T_31[9:0]) begin
        image_1_232 <= io_pixelVal_in_1_5;
      end else if (10'he8 == _T_28[9:0]) begin
        image_1_232 <= io_pixelVal_in_1_4;
      end else if (10'he8 == _T_25[9:0]) begin
        image_1_232 <= io_pixelVal_in_1_3;
      end else if (10'he8 == _T_22[9:0]) begin
        image_1_232 <= io_pixelVal_in_1_2;
      end else if (10'he8 == _T_19[9:0]) begin
        image_1_232 <= io_pixelVal_in_1_1;
      end else if (10'he8 == _T_15[9:0]) begin
        image_1_232 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_233 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he9 == _T_37[9:0]) begin
        image_1_233 <= io_pixelVal_in_1_7;
      end else if (10'he9 == _T_34[9:0]) begin
        image_1_233 <= io_pixelVal_in_1_6;
      end else if (10'he9 == _T_31[9:0]) begin
        image_1_233 <= io_pixelVal_in_1_5;
      end else if (10'he9 == _T_28[9:0]) begin
        image_1_233 <= io_pixelVal_in_1_4;
      end else if (10'he9 == _T_25[9:0]) begin
        image_1_233 <= io_pixelVal_in_1_3;
      end else if (10'he9 == _T_22[9:0]) begin
        image_1_233 <= io_pixelVal_in_1_2;
      end else if (10'he9 == _T_19[9:0]) begin
        image_1_233 <= io_pixelVal_in_1_1;
      end else if (10'he9 == _T_15[9:0]) begin
        image_1_233 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_234 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hea == _T_37[9:0]) begin
        image_1_234 <= io_pixelVal_in_1_7;
      end else if (10'hea == _T_34[9:0]) begin
        image_1_234 <= io_pixelVal_in_1_6;
      end else if (10'hea == _T_31[9:0]) begin
        image_1_234 <= io_pixelVal_in_1_5;
      end else if (10'hea == _T_28[9:0]) begin
        image_1_234 <= io_pixelVal_in_1_4;
      end else if (10'hea == _T_25[9:0]) begin
        image_1_234 <= io_pixelVal_in_1_3;
      end else if (10'hea == _T_22[9:0]) begin
        image_1_234 <= io_pixelVal_in_1_2;
      end else if (10'hea == _T_19[9:0]) begin
        image_1_234 <= io_pixelVal_in_1_1;
      end else if (10'hea == _T_15[9:0]) begin
        image_1_234 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_235 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'heb == _T_37[9:0]) begin
        image_1_235 <= io_pixelVal_in_1_7;
      end else if (10'heb == _T_34[9:0]) begin
        image_1_235 <= io_pixelVal_in_1_6;
      end else if (10'heb == _T_31[9:0]) begin
        image_1_235 <= io_pixelVal_in_1_5;
      end else if (10'heb == _T_28[9:0]) begin
        image_1_235 <= io_pixelVal_in_1_4;
      end else if (10'heb == _T_25[9:0]) begin
        image_1_235 <= io_pixelVal_in_1_3;
      end else if (10'heb == _T_22[9:0]) begin
        image_1_235 <= io_pixelVal_in_1_2;
      end else if (10'heb == _T_19[9:0]) begin
        image_1_235 <= io_pixelVal_in_1_1;
      end else if (10'heb == _T_15[9:0]) begin
        image_1_235 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_236 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hec == _T_37[9:0]) begin
        image_1_236 <= io_pixelVal_in_1_7;
      end else if (10'hec == _T_34[9:0]) begin
        image_1_236 <= io_pixelVal_in_1_6;
      end else if (10'hec == _T_31[9:0]) begin
        image_1_236 <= io_pixelVal_in_1_5;
      end else if (10'hec == _T_28[9:0]) begin
        image_1_236 <= io_pixelVal_in_1_4;
      end else if (10'hec == _T_25[9:0]) begin
        image_1_236 <= io_pixelVal_in_1_3;
      end else if (10'hec == _T_22[9:0]) begin
        image_1_236 <= io_pixelVal_in_1_2;
      end else if (10'hec == _T_19[9:0]) begin
        image_1_236 <= io_pixelVal_in_1_1;
      end else if (10'hec == _T_15[9:0]) begin
        image_1_236 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_237 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hed == _T_37[9:0]) begin
        image_1_237 <= io_pixelVal_in_1_7;
      end else if (10'hed == _T_34[9:0]) begin
        image_1_237 <= io_pixelVal_in_1_6;
      end else if (10'hed == _T_31[9:0]) begin
        image_1_237 <= io_pixelVal_in_1_5;
      end else if (10'hed == _T_28[9:0]) begin
        image_1_237 <= io_pixelVal_in_1_4;
      end else if (10'hed == _T_25[9:0]) begin
        image_1_237 <= io_pixelVal_in_1_3;
      end else if (10'hed == _T_22[9:0]) begin
        image_1_237 <= io_pixelVal_in_1_2;
      end else if (10'hed == _T_19[9:0]) begin
        image_1_237 <= io_pixelVal_in_1_1;
      end else if (10'hed == _T_15[9:0]) begin
        image_1_237 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_238 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hee == _T_37[9:0]) begin
        image_1_238 <= io_pixelVal_in_1_7;
      end else if (10'hee == _T_34[9:0]) begin
        image_1_238 <= io_pixelVal_in_1_6;
      end else if (10'hee == _T_31[9:0]) begin
        image_1_238 <= io_pixelVal_in_1_5;
      end else if (10'hee == _T_28[9:0]) begin
        image_1_238 <= io_pixelVal_in_1_4;
      end else if (10'hee == _T_25[9:0]) begin
        image_1_238 <= io_pixelVal_in_1_3;
      end else if (10'hee == _T_22[9:0]) begin
        image_1_238 <= io_pixelVal_in_1_2;
      end else if (10'hee == _T_19[9:0]) begin
        image_1_238 <= io_pixelVal_in_1_1;
      end else if (10'hee == _T_15[9:0]) begin
        image_1_238 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_239 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hef == _T_37[9:0]) begin
        image_1_239 <= io_pixelVal_in_1_7;
      end else if (10'hef == _T_34[9:0]) begin
        image_1_239 <= io_pixelVal_in_1_6;
      end else if (10'hef == _T_31[9:0]) begin
        image_1_239 <= io_pixelVal_in_1_5;
      end else if (10'hef == _T_28[9:0]) begin
        image_1_239 <= io_pixelVal_in_1_4;
      end else if (10'hef == _T_25[9:0]) begin
        image_1_239 <= io_pixelVal_in_1_3;
      end else if (10'hef == _T_22[9:0]) begin
        image_1_239 <= io_pixelVal_in_1_2;
      end else if (10'hef == _T_19[9:0]) begin
        image_1_239 <= io_pixelVal_in_1_1;
      end else if (10'hef == _T_15[9:0]) begin
        image_1_239 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_240 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf0 == _T_37[9:0]) begin
        image_1_240 <= io_pixelVal_in_1_7;
      end else if (10'hf0 == _T_34[9:0]) begin
        image_1_240 <= io_pixelVal_in_1_6;
      end else if (10'hf0 == _T_31[9:0]) begin
        image_1_240 <= io_pixelVal_in_1_5;
      end else if (10'hf0 == _T_28[9:0]) begin
        image_1_240 <= io_pixelVal_in_1_4;
      end else if (10'hf0 == _T_25[9:0]) begin
        image_1_240 <= io_pixelVal_in_1_3;
      end else if (10'hf0 == _T_22[9:0]) begin
        image_1_240 <= io_pixelVal_in_1_2;
      end else if (10'hf0 == _T_19[9:0]) begin
        image_1_240 <= io_pixelVal_in_1_1;
      end else if (10'hf0 == _T_15[9:0]) begin
        image_1_240 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_241 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf1 == _T_37[9:0]) begin
        image_1_241 <= io_pixelVal_in_1_7;
      end else if (10'hf1 == _T_34[9:0]) begin
        image_1_241 <= io_pixelVal_in_1_6;
      end else if (10'hf1 == _T_31[9:0]) begin
        image_1_241 <= io_pixelVal_in_1_5;
      end else if (10'hf1 == _T_28[9:0]) begin
        image_1_241 <= io_pixelVal_in_1_4;
      end else if (10'hf1 == _T_25[9:0]) begin
        image_1_241 <= io_pixelVal_in_1_3;
      end else if (10'hf1 == _T_22[9:0]) begin
        image_1_241 <= io_pixelVal_in_1_2;
      end else if (10'hf1 == _T_19[9:0]) begin
        image_1_241 <= io_pixelVal_in_1_1;
      end else if (10'hf1 == _T_15[9:0]) begin
        image_1_241 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_242 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf2 == _T_37[9:0]) begin
        image_1_242 <= io_pixelVal_in_1_7;
      end else if (10'hf2 == _T_34[9:0]) begin
        image_1_242 <= io_pixelVal_in_1_6;
      end else if (10'hf2 == _T_31[9:0]) begin
        image_1_242 <= io_pixelVal_in_1_5;
      end else if (10'hf2 == _T_28[9:0]) begin
        image_1_242 <= io_pixelVal_in_1_4;
      end else if (10'hf2 == _T_25[9:0]) begin
        image_1_242 <= io_pixelVal_in_1_3;
      end else if (10'hf2 == _T_22[9:0]) begin
        image_1_242 <= io_pixelVal_in_1_2;
      end else if (10'hf2 == _T_19[9:0]) begin
        image_1_242 <= io_pixelVal_in_1_1;
      end else if (10'hf2 == _T_15[9:0]) begin
        image_1_242 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_243 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf3 == _T_37[9:0]) begin
        image_1_243 <= io_pixelVal_in_1_7;
      end else if (10'hf3 == _T_34[9:0]) begin
        image_1_243 <= io_pixelVal_in_1_6;
      end else if (10'hf3 == _T_31[9:0]) begin
        image_1_243 <= io_pixelVal_in_1_5;
      end else if (10'hf3 == _T_28[9:0]) begin
        image_1_243 <= io_pixelVal_in_1_4;
      end else if (10'hf3 == _T_25[9:0]) begin
        image_1_243 <= io_pixelVal_in_1_3;
      end else if (10'hf3 == _T_22[9:0]) begin
        image_1_243 <= io_pixelVal_in_1_2;
      end else if (10'hf3 == _T_19[9:0]) begin
        image_1_243 <= io_pixelVal_in_1_1;
      end else if (10'hf3 == _T_15[9:0]) begin
        image_1_243 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_244 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf4 == _T_37[9:0]) begin
        image_1_244 <= io_pixelVal_in_1_7;
      end else if (10'hf4 == _T_34[9:0]) begin
        image_1_244 <= io_pixelVal_in_1_6;
      end else if (10'hf4 == _T_31[9:0]) begin
        image_1_244 <= io_pixelVal_in_1_5;
      end else if (10'hf4 == _T_28[9:0]) begin
        image_1_244 <= io_pixelVal_in_1_4;
      end else if (10'hf4 == _T_25[9:0]) begin
        image_1_244 <= io_pixelVal_in_1_3;
      end else if (10'hf4 == _T_22[9:0]) begin
        image_1_244 <= io_pixelVal_in_1_2;
      end else if (10'hf4 == _T_19[9:0]) begin
        image_1_244 <= io_pixelVal_in_1_1;
      end else if (10'hf4 == _T_15[9:0]) begin
        image_1_244 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_245 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf5 == _T_37[9:0]) begin
        image_1_245 <= io_pixelVal_in_1_7;
      end else if (10'hf5 == _T_34[9:0]) begin
        image_1_245 <= io_pixelVal_in_1_6;
      end else if (10'hf5 == _T_31[9:0]) begin
        image_1_245 <= io_pixelVal_in_1_5;
      end else if (10'hf5 == _T_28[9:0]) begin
        image_1_245 <= io_pixelVal_in_1_4;
      end else if (10'hf5 == _T_25[9:0]) begin
        image_1_245 <= io_pixelVal_in_1_3;
      end else if (10'hf5 == _T_22[9:0]) begin
        image_1_245 <= io_pixelVal_in_1_2;
      end else if (10'hf5 == _T_19[9:0]) begin
        image_1_245 <= io_pixelVal_in_1_1;
      end else if (10'hf5 == _T_15[9:0]) begin
        image_1_245 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_246 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf6 == _T_37[9:0]) begin
        image_1_246 <= io_pixelVal_in_1_7;
      end else if (10'hf6 == _T_34[9:0]) begin
        image_1_246 <= io_pixelVal_in_1_6;
      end else if (10'hf6 == _T_31[9:0]) begin
        image_1_246 <= io_pixelVal_in_1_5;
      end else if (10'hf6 == _T_28[9:0]) begin
        image_1_246 <= io_pixelVal_in_1_4;
      end else if (10'hf6 == _T_25[9:0]) begin
        image_1_246 <= io_pixelVal_in_1_3;
      end else if (10'hf6 == _T_22[9:0]) begin
        image_1_246 <= io_pixelVal_in_1_2;
      end else if (10'hf6 == _T_19[9:0]) begin
        image_1_246 <= io_pixelVal_in_1_1;
      end else if (10'hf6 == _T_15[9:0]) begin
        image_1_246 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_247 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf7 == _T_37[9:0]) begin
        image_1_247 <= io_pixelVal_in_1_7;
      end else if (10'hf7 == _T_34[9:0]) begin
        image_1_247 <= io_pixelVal_in_1_6;
      end else if (10'hf7 == _T_31[9:0]) begin
        image_1_247 <= io_pixelVal_in_1_5;
      end else if (10'hf7 == _T_28[9:0]) begin
        image_1_247 <= io_pixelVal_in_1_4;
      end else if (10'hf7 == _T_25[9:0]) begin
        image_1_247 <= io_pixelVal_in_1_3;
      end else if (10'hf7 == _T_22[9:0]) begin
        image_1_247 <= io_pixelVal_in_1_2;
      end else if (10'hf7 == _T_19[9:0]) begin
        image_1_247 <= io_pixelVal_in_1_1;
      end else if (10'hf7 == _T_15[9:0]) begin
        image_1_247 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_248 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf8 == _T_37[9:0]) begin
        image_1_248 <= io_pixelVal_in_1_7;
      end else if (10'hf8 == _T_34[9:0]) begin
        image_1_248 <= io_pixelVal_in_1_6;
      end else if (10'hf8 == _T_31[9:0]) begin
        image_1_248 <= io_pixelVal_in_1_5;
      end else if (10'hf8 == _T_28[9:0]) begin
        image_1_248 <= io_pixelVal_in_1_4;
      end else if (10'hf8 == _T_25[9:0]) begin
        image_1_248 <= io_pixelVal_in_1_3;
      end else if (10'hf8 == _T_22[9:0]) begin
        image_1_248 <= io_pixelVal_in_1_2;
      end else if (10'hf8 == _T_19[9:0]) begin
        image_1_248 <= io_pixelVal_in_1_1;
      end else if (10'hf8 == _T_15[9:0]) begin
        image_1_248 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_249 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf9 == _T_37[9:0]) begin
        image_1_249 <= io_pixelVal_in_1_7;
      end else if (10'hf9 == _T_34[9:0]) begin
        image_1_249 <= io_pixelVal_in_1_6;
      end else if (10'hf9 == _T_31[9:0]) begin
        image_1_249 <= io_pixelVal_in_1_5;
      end else if (10'hf9 == _T_28[9:0]) begin
        image_1_249 <= io_pixelVal_in_1_4;
      end else if (10'hf9 == _T_25[9:0]) begin
        image_1_249 <= io_pixelVal_in_1_3;
      end else if (10'hf9 == _T_22[9:0]) begin
        image_1_249 <= io_pixelVal_in_1_2;
      end else if (10'hf9 == _T_19[9:0]) begin
        image_1_249 <= io_pixelVal_in_1_1;
      end else if (10'hf9 == _T_15[9:0]) begin
        image_1_249 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_250 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hfa == _T_37[9:0]) begin
        image_1_250 <= io_pixelVal_in_1_7;
      end else if (10'hfa == _T_34[9:0]) begin
        image_1_250 <= io_pixelVal_in_1_6;
      end else if (10'hfa == _T_31[9:0]) begin
        image_1_250 <= io_pixelVal_in_1_5;
      end else if (10'hfa == _T_28[9:0]) begin
        image_1_250 <= io_pixelVal_in_1_4;
      end else if (10'hfa == _T_25[9:0]) begin
        image_1_250 <= io_pixelVal_in_1_3;
      end else if (10'hfa == _T_22[9:0]) begin
        image_1_250 <= io_pixelVal_in_1_2;
      end else if (10'hfa == _T_19[9:0]) begin
        image_1_250 <= io_pixelVal_in_1_1;
      end else if (10'hfa == _T_15[9:0]) begin
        image_1_250 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_251 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hfb == _T_37[9:0]) begin
        image_1_251 <= io_pixelVal_in_1_7;
      end else if (10'hfb == _T_34[9:0]) begin
        image_1_251 <= io_pixelVal_in_1_6;
      end else if (10'hfb == _T_31[9:0]) begin
        image_1_251 <= io_pixelVal_in_1_5;
      end else if (10'hfb == _T_28[9:0]) begin
        image_1_251 <= io_pixelVal_in_1_4;
      end else if (10'hfb == _T_25[9:0]) begin
        image_1_251 <= io_pixelVal_in_1_3;
      end else if (10'hfb == _T_22[9:0]) begin
        image_1_251 <= io_pixelVal_in_1_2;
      end else if (10'hfb == _T_19[9:0]) begin
        image_1_251 <= io_pixelVal_in_1_1;
      end else if (10'hfb == _T_15[9:0]) begin
        image_1_251 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_252 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hfc == _T_37[9:0]) begin
        image_1_252 <= io_pixelVal_in_1_7;
      end else if (10'hfc == _T_34[9:0]) begin
        image_1_252 <= io_pixelVal_in_1_6;
      end else if (10'hfc == _T_31[9:0]) begin
        image_1_252 <= io_pixelVal_in_1_5;
      end else if (10'hfc == _T_28[9:0]) begin
        image_1_252 <= io_pixelVal_in_1_4;
      end else if (10'hfc == _T_25[9:0]) begin
        image_1_252 <= io_pixelVal_in_1_3;
      end else if (10'hfc == _T_22[9:0]) begin
        image_1_252 <= io_pixelVal_in_1_2;
      end else if (10'hfc == _T_19[9:0]) begin
        image_1_252 <= io_pixelVal_in_1_1;
      end else if (10'hfc == _T_15[9:0]) begin
        image_1_252 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_253 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hfd == _T_37[9:0]) begin
        image_1_253 <= io_pixelVal_in_1_7;
      end else if (10'hfd == _T_34[9:0]) begin
        image_1_253 <= io_pixelVal_in_1_6;
      end else if (10'hfd == _T_31[9:0]) begin
        image_1_253 <= io_pixelVal_in_1_5;
      end else if (10'hfd == _T_28[9:0]) begin
        image_1_253 <= io_pixelVal_in_1_4;
      end else if (10'hfd == _T_25[9:0]) begin
        image_1_253 <= io_pixelVal_in_1_3;
      end else if (10'hfd == _T_22[9:0]) begin
        image_1_253 <= io_pixelVal_in_1_2;
      end else if (10'hfd == _T_19[9:0]) begin
        image_1_253 <= io_pixelVal_in_1_1;
      end else if (10'hfd == _T_15[9:0]) begin
        image_1_253 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_254 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hfe == _T_37[9:0]) begin
        image_1_254 <= io_pixelVal_in_1_7;
      end else if (10'hfe == _T_34[9:0]) begin
        image_1_254 <= io_pixelVal_in_1_6;
      end else if (10'hfe == _T_31[9:0]) begin
        image_1_254 <= io_pixelVal_in_1_5;
      end else if (10'hfe == _T_28[9:0]) begin
        image_1_254 <= io_pixelVal_in_1_4;
      end else if (10'hfe == _T_25[9:0]) begin
        image_1_254 <= io_pixelVal_in_1_3;
      end else if (10'hfe == _T_22[9:0]) begin
        image_1_254 <= io_pixelVal_in_1_2;
      end else if (10'hfe == _T_19[9:0]) begin
        image_1_254 <= io_pixelVal_in_1_1;
      end else if (10'hfe == _T_15[9:0]) begin
        image_1_254 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_255 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hff == _T_37[9:0]) begin
        image_1_255 <= io_pixelVal_in_1_7;
      end else if (10'hff == _T_34[9:0]) begin
        image_1_255 <= io_pixelVal_in_1_6;
      end else if (10'hff == _T_31[9:0]) begin
        image_1_255 <= io_pixelVal_in_1_5;
      end else if (10'hff == _T_28[9:0]) begin
        image_1_255 <= io_pixelVal_in_1_4;
      end else if (10'hff == _T_25[9:0]) begin
        image_1_255 <= io_pixelVal_in_1_3;
      end else if (10'hff == _T_22[9:0]) begin
        image_1_255 <= io_pixelVal_in_1_2;
      end else if (10'hff == _T_19[9:0]) begin
        image_1_255 <= io_pixelVal_in_1_1;
      end else if (10'hff == _T_15[9:0]) begin
        image_1_255 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_256 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h100 == _T_37[9:0]) begin
        image_1_256 <= io_pixelVal_in_1_7;
      end else if (10'h100 == _T_34[9:0]) begin
        image_1_256 <= io_pixelVal_in_1_6;
      end else if (10'h100 == _T_31[9:0]) begin
        image_1_256 <= io_pixelVal_in_1_5;
      end else if (10'h100 == _T_28[9:0]) begin
        image_1_256 <= io_pixelVal_in_1_4;
      end else if (10'h100 == _T_25[9:0]) begin
        image_1_256 <= io_pixelVal_in_1_3;
      end else if (10'h100 == _T_22[9:0]) begin
        image_1_256 <= io_pixelVal_in_1_2;
      end else if (10'h100 == _T_19[9:0]) begin
        image_1_256 <= io_pixelVal_in_1_1;
      end else if (10'h100 == _T_15[9:0]) begin
        image_1_256 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_257 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h101 == _T_37[9:0]) begin
        image_1_257 <= io_pixelVal_in_1_7;
      end else if (10'h101 == _T_34[9:0]) begin
        image_1_257 <= io_pixelVal_in_1_6;
      end else if (10'h101 == _T_31[9:0]) begin
        image_1_257 <= io_pixelVal_in_1_5;
      end else if (10'h101 == _T_28[9:0]) begin
        image_1_257 <= io_pixelVal_in_1_4;
      end else if (10'h101 == _T_25[9:0]) begin
        image_1_257 <= io_pixelVal_in_1_3;
      end else if (10'h101 == _T_22[9:0]) begin
        image_1_257 <= io_pixelVal_in_1_2;
      end else if (10'h101 == _T_19[9:0]) begin
        image_1_257 <= io_pixelVal_in_1_1;
      end else if (10'h101 == _T_15[9:0]) begin
        image_1_257 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_258 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h102 == _T_37[9:0]) begin
        image_1_258 <= io_pixelVal_in_1_7;
      end else if (10'h102 == _T_34[9:0]) begin
        image_1_258 <= io_pixelVal_in_1_6;
      end else if (10'h102 == _T_31[9:0]) begin
        image_1_258 <= io_pixelVal_in_1_5;
      end else if (10'h102 == _T_28[9:0]) begin
        image_1_258 <= io_pixelVal_in_1_4;
      end else if (10'h102 == _T_25[9:0]) begin
        image_1_258 <= io_pixelVal_in_1_3;
      end else if (10'h102 == _T_22[9:0]) begin
        image_1_258 <= io_pixelVal_in_1_2;
      end else if (10'h102 == _T_19[9:0]) begin
        image_1_258 <= io_pixelVal_in_1_1;
      end else if (10'h102 == _T_15[9:0]) begin
        image_1_258 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_259 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h103 == _T_37[9:0]) begin
        image_1_259 <= io_pixelVal_in_1_7;
      end else if (10'h103 == _T_34[9:0]) begin
        image_1_259 <= io_pixelVal_in_1_6;
      end else if (10'h103 == _T_31[9:0]) begin
        image_1_259 <= io_pixelVal_in_1_5;
      end else if (10'h103 == _T_28[9:0]) begin
        image_1_259 <= io_pixelVal_in_1_4;
      end else if (10'h103 == _T_25[9:0]) begin
        image_1_259 <= io_pixelVal_in_1_3;
      end else if (10'h103 == _T_22[9:0]) begin
        image_1_259 <= io_pixelVal_in_1_2;
      end else if (10'h103 == _T_19[9:0]) begin
        image_1_259 <= io_pixelVal_in_1_1;
      end else if (10'h103 == _T_15[9:0]) begin
        image_1_259 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_260 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h104 == _T_37[9:0]) begin
        image_1_260 <= io_pixelVal_in_1_7;
      end else if (10'h104 == _T_34[9:0]) begin
        image_1_260 <= io_pixelVal_in_1_6;
      end else if (10'h104 == _T_31[9:0]) begin
        image_1_260 <= io_pixelVal_in_1_5;
      end else if (10'h104 == _T_28[9:0]) begin
        image_1_260 <= io_pixelVal_in_1_4;
      end else if (10'h104 == _T_25[9:0]) begin
        image_1_260 <= io_pixelVal_in_1_3;
      end else if (10'h104 == _T_22[9:0]) begin
        image_1_260 <= io_pixelVal_in_1_2;
      end else if (10'h104 == _T_19[9:0]) begin
        image_1_260 <= io_pixelVal_in_1_1;
      end else if (10'h104 == _T_15[9:0]) begin
        image_1_260 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_261 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h105 == _T_37[9:0]) begin
        image_1_261 <= io_pixelVal_in_1_7;
      end else if (10'h105 == _T_34[9:0]) begin
        image_1_261 <= io_pixelVal_in_1_6;
      end else if (10'h105 == _T_31[9:0]) begin
        image_1_261 <= io_pixelVal_in_1_5;
      end else if (10'h105 == _T_28[9:0]) begin
        image_1_261 <= io_pixelVal_in_1_4;
      end else if (10'h105 == _T_25[9:0]) begin
        image_1_261 <= io_pixelVal_in_1_3;
      end else if (10'h105 == _T_22[9:0]) begin
        image_1_261 <= io_pixelVal_in_1_2;
      end else if (10'h105 == _T_19[9:0]) begin
        image_1_261 <= io_pixelVal_in_1_1;
      end else if (10'h105 == _T_15[9:0]) begin
        image_1_261 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_262 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h106 == _T_37[9:0]) begin
        image_1_262 <= io_pixelVal_in_1_7;
      end else if (10'h106 == _T_34[9:0]) begin
        image_1_262 <= io_pixelVal_in_1_6;
      end else if (10'h106 == _T_31[9:0]) begin
        image_1_262 <= io_pixelVal_in_1_5;
      end else if (10'h106 == _T_28[9:0]) begin
        image_1_262 <= io_pixelVal_in_1_4;
      end else if (10'h106 == _T_25[9:0]) begin
        image_1_262 <= io_pixelVal_in_1_3;
      end else if (10'h106 == _T_22[9:0]) begin
        image_1_262 <= io_pixelVal_in_1_2;
      end else if (10'h106 == _T_19[9:0]) begin
        image_1_262 <= io_pixelVal_in_1_1;
      end else if (10'h106 == _T_15[9:0]) begin
        image_1_262 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_263 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h107 == _T_37[9:0]) begin
        image_1_263 <= io_pixelVal_in_1_7;
      end else if (10'h107 == _T_34[9:0]) begin
        image_1_263 <= io_pixelVal_in_1_6;
      end else if (10'h107 == _T_31[9:0]) begin
        image_1_263 <= io_pixelVal_in_1_5;
      end else if (10'h107 == _T_28[9:0]) begin
        image_1_263 <= io_pixelVal_in_1_4;
      end else if (10'h107 == _T_25[9:0]) begin
        image_1_263 <= io_pixelVal_in_1_3;
      end else if (10'h107 == _T_22[9:0]) begin
        image_1_263 <= io_pixelVal_in_1_2;
      end else if (10'h107 == _T_19[9:0]) begin
        image_1_263 <= io_pixelVal_in_1_1;
      end else if (10'h107 == _T_15[9:0]) begin
        image_1_263 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_264 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h108 == _T_37[9:0]) begin
        image_1_264 <= io_pixelVal_in_1_7;
      end else if (10'h108 == _T_34[9:0]) begin
        image_1_264 <= io_pixelVal_in_1_6;
      end else if (10'h108 == _T_31[9:0]) begin
        image_1_264 <= io_pixelVal_in_1_5;
      end else if (10'h108 == _T_28[9:0]) begin
        image_1_264 <= io_pixelVal_in_1_4;
      end else if (10'h108 == _T_25[9:0]) begin
        image_1_264 <= io_pixelVal_in_1_3;
      end else if (10'h108 == _T_22[9:0]) begin
        image_1_264 <= io_pixelVal_in_1_2;
      end else if (10'h108 == _T_19[9:0]) begin
        image_1_264 <= io_pixelVal_in_1_1;
      end else if (10'h108 == _T_15[9:0]) begin
        image_1_264 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_265 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h109 == _T_37[9:0]) begin
        image_1_265 <= io_pixelVal_in_1_7;
      end else if (10'h109 == _T_34[9:0]) begin
        image_1_265 <= io_pixelVal_in_1_6;
      end else if (10'h109 == _T_31[9:0]) begin
        image_1_265 <= io_pixelVal_in_1_5;
      end else if (10'h109 == _T_28[9:0]) begin
        image_1_265 <= io_pixelVal_in_1_4;
      end else if (10'h109 == _T_25[9:0]) begin
        image_1_265 <= io_pixelVal_in_1_3;
      end else if (10'h109 == _T_22[9:0]) begin
        image_1_265 <= io_pixelVal_in_1_2;
      end else if (10'h109 == _T_19[9:0]) begin
        image_1_265 <= io_pixelVal_in_1_1;
      end else if (10'h109 == _T_15[9:0]) begin
        image_1_265 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_266 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h10a == _T_37[9:0]) begin
        image_1_266 <= io_pixelVal_in_1_7;
      end else if (10'h10a == _T_34[9:0]) begin
        image_1_266 <= io_pixelVal_in_1_6;
      end else if (10'h10a == _T_31[9:0]) begin
        image_1_266 <= io_pixelVal_in_1_5;
      end else if (10'h10a == _T_28[9:0]) begin
        image_1_266 <= io_pixelVal_in_1_4;
      end else if (10'h10a == _T_25[9:0]) begin
        image_1_266 <= io_pixelVal_in_1_3;
      end else if (10'h10a == _T_22[9:0]) begin
        image_1_266 <= io_pixelVal_in_1_2;
      end else if (10'h10a == _T_19[9:0]) begin
        image_1_266 <= io_pixelVal_in_1_1;
      end else if (10'h10a == _T_15[9:0]) begin
        image_1_266 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_267 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h10b == _T_37[9:0]) begin
        image_1_267 <= io_pixelVal_in_1_7;
      end else if (10'h10b == _T_34[9:0]) begin
        image_1_267 <= io_pixelVal_in_1_6;
      end else if (10'h10b == _T_31[9:0]) begin
        image_1_267 <= io_pixelVal_in_1_5;
      end else if (10'h10b == _T_28[9:0]) begin
        image_1_267 <= io_pixelVal_in_1_4;
      end else if (10'h10b == _T_25[9:0]) begin
        image_1_267 <= io_pixelVal_in_1_3;
      end else if (10'h10b == _T_22[9:0]) begin
        image_1_267 <= io_pixelVal_in_1_2;
      end else if (10'h10b == _T_19[9:0]) begin
        image_1_267 <= io_pixelVal_in_1_1;
      end else if (10'h10b == _T_15[9:0]) begin
        image_1_267 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_268 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h10c == _T_37[9:0]) begin
        image_1_268 <= io_pixelVal_in_1_7;
      end else if (10'h10c == _T_34[9:0]) begin
        image_1_268 <= io_pixelVal_in_1_6;
      end else if (10'h10c == _T_31[9:0]) begin
        image_1_268 <= io_pixelVal_in_1_5;
      end else if (10'h10c == _T_28[9:0]) begin
        image_1_268 <= io_pixelVal_in_1_4;
      end else if (10'h10c == _T_25[9:0]) begin
        image_1_268 <= io_pixelVal_in_1_3;
      end else if (10'h10c == _T_22[9:0]) begin
        image_1_268 <= io_pixelVal_in_1_2;
      end else if (10'h10c == _T_19[9:0]) begin
        image_1_268 <= io_pixelVal_in_1_1;
      end else if (10'h10c == _T_15[9:0]) begin
        image_1_268 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_269 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h10d == _T_37[9:0]) begin
        image_1_269 <= io_pixelVal_in_1_7;
      end else if (10'h10d == _T_34[9:0]) begin
        image_1_269 <= io_pixelVal_in_1_6;
      end else if (10'h10d == _T_31[9:0]) begin
        image_1_269 <= io_pixelVal_in_1_5;
      end else if (10'h10d == _T_28[9:0]) begin
        image_1_269 <= io_pixelVal_in_1_4;
      end else if (10'h10d == _T_25[9:0]) begin
        image_1_269 <= io_pixelVal_in_1_3;
      end else if (10'h10d == _T_22[9:0]) begin
        image_1_269 <= io_pixelVal_in_1_2;
      end else if (10'h10d == _T_19[9:0]) begin
        image_1_269 <= io_pixelVal_in_1_1;
      end else if (10'h10d == _T_15[9:0]) begin
        image_1_269 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_270 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h10e == _T_37[9:0]) begin
        image_1_270 <= io_pixelVal_in_1_7;
      end else if (10'h10e == _T_34[9:0]) begin
        image_1_270 <= io_pixelVal_in_1_6;
      end else if (10'h10e == _T_31[9:0]) begin
        image_1_270 <= io_pixelVal_in_1_5;
      end else if (10'h10e == _T_28[9:0]) begin
        image_1_270 <= io_pixelVal_in_1_4;
      end else if (10'h10e == _T_25[9:0]) begin
        image_1_270 <= io_pixelVal_in_1_3;
      end else if (10'h10e == _T_22[9:0]) begin
        image_1_270 <= io_pixelVal_in_1_2;
      end else if (10'h10e == _T_19[9:0]) begin
        image_1_270 <= io_pixelVal_in_1_1;
      end else if (10'h10e == _T_15[9:0]) begin
        image_1_270 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_271 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h10f == _T_37[9:0]) begin
        image_1_271 <= io_pixelVal_in_1_7;
      end else if (10'h10f == _T_34[9:0]) begin
        image_1_271 <= io_pixelVal_in_1_6;
      end else if (10'h10f == _T_31[9:0]) begin
        image_1_271 <= io_pixelVal_in_1_5;
      end else if (10'h10f == _T_28[9:0]) begin
        image_1_271 <= io_pixelVal_in_1_4;
      end else if (10'h10f == _T_25[9:0]) begin
        image_1_271 <= io_pixelVal_in_1_3;
      end else if (10'h10f == _T_22[9:0]) begin
        image_1_271 <= io_pixelVal_in_1_2;
      end else if (10'h10f == _T_19[9:0]) begin
        image_1_271 <= io_pixelVal_in_1_1;
      end else if (10'h10f == _T_15[9:0]) begin
        image_1_271 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_272 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h110 == _T_37[9:0]) begin
        image_1_272 <= io_pixelVal_in_1_7;
      end else if (10'h110 == _T_34[9:0]) begin
        image_1_272 <= io_pixelVal_in_1_6;
      end else if (10'h110 == _T_31[9:0]) begin
        image_1_272 <= io_pixelVal_in_1_5;
      end else if (10'h110 == _T_28[9:0]) begin
        image_1_272 <= io_pixelVal_in_1_4;
      end else if (10'h110 == _T_25[9:0]) begin
        image_1_272 <= io_pixelVal_in_1_3;
      end else if (10'h110 == _T_22[9:0]) begin
        image_1_272 <= io_pixelVal_in_1_2;
      end else if (10'h110 == _T_19[9:0]) begin
        image_1_272 <= io_pixelVal_in_1_1;
      end else if (10'h110 == _T_15[9:0]) begin
        image_1_272 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_273 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h111 == _T_37[9:0]) begin
        image_1_273 <= io_pixelVal_in_1_7;
      end else if (10'h111 == _T_34[9:0]) begin
        image_1_273 <= io_pixelVal_in_1_6;
      end else if (10'h111 == _T_31[9:0]) begin
        image_1_273 <= io_pixelVal_in_1_5;
      end else if (10'h111 == _T_28[9:0]) begin
        image_1_273 <= io_pixelVal_in_1_4;
      end else if (10'h111 == _T_25[9:0]) begin
        image_1_273 <= io_pixelVal_in_1_3;
      end else if (10'h111 == _T_22[9:0]) begin
        image_1_273 <= io_pixelVal_in_1_2;
      end else if (10'h111 == _T_19[9:0]) begin
        image_1_273 <= io_pixelVal_in_1_1;
      end else if (10'h111 == _T_15[9:0]) begin
        image_1_273 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_274 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h112 == _T_37[9:0]) begin
        image_1_274 <= io_pixelVal_in_1_7;
      end else if (10'h112 == _T_34[9:0]) begin
        image_1_274 <= io_pixelVal_in_1_6;
      end else if (10'h112 == _T_31[9:0]) begin
        image_1_274 <= io_pixelVal_in_1_5;
      end else if (10'h112 == _T_28[9:0]) begin
        image_1_274 <= io_pixelVal_in_1_4;
      end else if (10'h112 == _T_25[9:0]) begin
        image_1_274 <= io_pixelVal_in_1_3;
      end else if (10'h112 == _T_22[9:0]) begin
        image_1_274 <= io_pixelVal_in_1_2;
      end else if (10'h112 == _T_19[9:0]) begin
        image_1_274 <= io_pixelVal_in_1_1;
      end else if (10'h112 == _T_15[9:0]) begin
        image_1_274 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_275 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h113 == _T_37[9:0]) begin
        image_1_275 <= io_pixelVal_in_1_7;
      end else if (10'h113 == _T_34[9:0]) begin
        image_1_275 <= io_pixelVal_in_1_6;
      end else if (10'h113 == _T_31[9:0]) begin
        image_1_275 <= io_pixelVal_in_1_5;
      end else if (10'h113 == _T_28[9:0]) begin
        image_1_275 <= io_pixelVal_in_1_4;
      end else if (10'h113 == _T_25[9:0]) begin
        image_1_275 <= io_pixelVal_in_1_3;
      end else if (10'h113 == _T_22[9:0]) begin
        image_1_275 <= io_pixelVal_in_1_2;
      end else if (10'h113 == _T_19[9:0]) begin
        image_1_275 <= io_pixelVal_in_1_1;
      end else if (10'h113 == _T_15[9:0]) begin
        image_1_275 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_276 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h114 == _T_37[9:0]) begin
        image_1_276 <= io_pixelVal_in_1_7;
      end else if (10'h114 == _T_34[9:0]) begin
        image_1_276 <= io_pixelVal_in_1_6;
      end else if (10'h114 == _T_31[9:0]) begin
        image_1_276 <= io_pixelVal_in_1_5;
      end else if (10'h114 == _T_28[9:0]) begin
        image_1_276 <= io_pixelVal_in_1_4;
      end else if (10'h114 == _T_25[9:0]) begin
        image_1_276 <= io_pixelVal_in_1_3;
      end else if (10'h114 == _T_22[9:0]) begin
        image_1_276 <= io_pixelVal_in_1_2;
      end else if (10'h114 == _T_19[9:0]) begin
        image_1_276 <= io_pixelVal_in_1_1;
      end else if (10'h114 == _T_15[9:0]) begin
        image_1_276 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_277 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h115 == _T_37[9:0]) begin
        image_1_277 <= io_pixelVal_in_1_7;
      end else if (10'h115 == _T_34[9:0]) begin
        image_1_277 <= io_pixelVal_in_1_6;
      end else if (10'h115 == _T_31[9:0]) begin
        image_1_277 <= io_pixelVal_in_1_5;
      end else if (10'h115 == _T_28[9:0]) begin
        image_1_277 <= io_pixelVal_in_1_4;
      end else if (10'h115 == _T_25[9:0]) begin
        image_1_277 <= io_pixelVal_in_1_3;
      end else if (10'h115 == _T_22[9:0]) begin
        image_1_277 <= io_pixelVal_in_1_2;
      end else if (10'h115 == _T_19[9:0]) begin
        image_1_277 <= io_pixelVal_in_1_1;
      end else if (10'h115 == _T_15[9:0]) begin
        image_1_277 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_278 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h116 == _T_37[9:0]) begin
        image_1_278 <= io_pixelVal_in_1_7;
      end else if (10'h116 == _T_34[9:0]) begin
        image_1_278 <= io_pixelVal_in_1_6;
      end else if (10'h116 == _T_31[9:0]) begin
        image_1_278 <= io_pixelVal_in_1_5;
      end else if (10'h116 == _T_28[9:0]) begin
        image_1_278 <= io_pixelVal_in_1_4;
      end else if (10'h116 == _T_25[9:0]) begin
        image_1_278 <= io_pixelVal_in_1_3;
      end else if (10'h116 == _T_22[9:0]) begin
        image_1_278 <= io_pixelVal_in_1_2;
      end else if (10'h116 == _T_19[9:0]) begin
        image_1_278 <= io_pixelVal_in_1_1;
      end else if (10'h116 == _T_15[9:0]) begin
        image_1_278 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_279 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h117 == _T_37[9:0]) begin
        image_1_279 <= io_pixelVal_in_1_7;
      end else if (10'h117 == _T_34[9:0]) begin
        image_1_279 <= io_pixelVal_in_1_6;
      end else if (10'h117 == _T_31[9:0]) begin
        image_1_279 <= io_pixelVal_in_1_5;
      end else if (10'h117 == _T_28[9:0]) begin
        image_1_279 <= io_pixelVal_in_1_4;
      end else if (10'h117 == _T_25[9:0]) begin
        image_1_279 <= io_pixelVal_in_1_3;
      end else if (10'h117 == _T_22[9:0]) begin
        image_1_279 <= io_pixelVal_in_1_2;
      end else if (10'h117 == _T_19[9:0]) begin
        image_1_279 <= io_pixelVal_in_1_1;
      end else if (10'h117 == _T_15[9:0]) begin
        image_1_279 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_280 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h118 == _T_37[9:0]) begin
        image_1_280 <= io_pixelVal_in_1_7;
      end else if (10'h118 == _T_34[9:0]) begin
        image_1_280 <= io_pixelVal_in_1_6;
      end else if (10'h118 == _T_31[9:0]) begin
        image_1_280 <= io_pixelVal_in_1_5;
      end else if (10'h118 == _T_28[9:0]) begin
        image_1_280 <= io_pixelVal_in_1_4;
      end else if (10'h118 == _T_25[9:0]) begin
        image_1_280 <= io_pixelVal_in_1_3;
      end else if (10'h118 == _T_22[9:0]) begin
        image_1_280 <= io_pixelVal_in_1_2;
      end else if (10'h118 == _T_19[9:0]) begin
        image_1_280 <= io_pixelVal_in_1_1;
      end else if (10'h118 == _T_15[9:0]) begin
        image_1_280 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_281 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h119 == _T_37[9:0]) begin
        image_1_281 <= io_pixelVal_in_1_7;
      end else if (10'h119 == _T_34[9:0]) begin
        image_1_281 <= io_pixelVal_in_1_6;
      end else if (10'h119 == _T_31[9:0]) begin
        image_1_281 <= io_pixelVal_in_1_5;
      end else if (10'h119 == _T_28[9:0]) begin
        image_1_281 <= io_pixelVal_in_1_4;
      end else if (10'h119 == _T_25[9:0]) begin
        image_1_281 <= io_pixelVal_in_1_3;
      end else if (10'h119 == _T_22[9:0]) begin
        image_1_281 <= io_pixelVal_in_1_2;
      end else if (10'h119 == _T_19[9:0]) begin
        image_1_281 <= io_pixelVal_in_1_1;
      end else if (10'h119 == _T_15[9:0]) begin
        image_1_281 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_282 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h11a == _T_37[9:0]) begin
        image_1_282 <= io_pixelVal_in_1_7;
      end else if (10'h11a == _T_34[9:0]) begin
        image_1_282 <= io_pixelVal_in_1_6;
      end else if (10'h11a == _T_31[9:0]) begin
        image_1_282 <= io_pixelVal_in_1_5;
      end else if (10'h11a == _T_28[9:0]) begin
        image_1_282 <= io_pixelVal_in_1_4;
      end else if (10'h11a == _T_25[9:0]) begin
        image_1_282 <= io_pixelVal_in_1_3;
      end else if (10'h11a == _T_22[9:0]) begin
        image_1_282 <= io_pixelVal_in_1_2;
      end else if (10'h11a == _T_19[9:0]) begin
        image_1_282 <= io_pixelVal_in_1_1;
      end else if (10'h11a == _T_15[9:0]) begin
        image_1_282 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_283 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h11b == _T_37[9:0]) begin
        image_1_283 <= io_pixelVal_in_1_7;
      end else if (10'h11b == _T_34[9:0]) begin
        image_1_283 <= io_pixelVal_in_1_6;
      end else if (10'h11b == _T_31[9:0]) begin
        image_1_283 <= io_pixelVal_in_1_5;
      end else if (10'h11b == _T_28[9:0]) begin
        image_1_283 <= io_pixelVal_in_1_4;
      end else if (10'h11b == _T_25[9:0]) begin
        image_1_283 <= io_pixelVal_in_1_3;
      end else if (10'h11b == _T_22[9:0]) begin
        image_1_283 <= io_pixelVal_in_1_2;
      end else if (10'h11b == _T_19[9:0]) begin
        image_1_283 <= io_pixelVal_in_1_1;
      end else if (10'h11b == _T_15[9:0]) begin
        image_1_283 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_284 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h11c == _T_37[9:0]) begin
        image_1_284 <= io_pixelVal_in_1_7;
      end else if (10'h11c == _T_34[9:0]) begin
        image_1_284 <= io_pixelVal_in_1_6;
      end else if (10'h11c == _T_31[9:0]) begin
        image_1_284 <= io_pixelVal_in_1_5;
      end else if (10'h11c == _T_28[9:0]) begin
        image_1_284 <= io_pixelVal_in_1_4;
      end else if (10'h11c == _T_25[9:0]) begin
        image_1_284 <= io_pixelVal_in_1_3;
      end else if (10'h11c == _T_22[9:0]) begin
        image_1_284 <= io_pixelVal_in_1_2;
      end else if (10'h11c == _T_19[9:0]) begin
        image_1_284 <= io_pixelVal_in_1_1;
      end else if (10'h11c == _T_15[9:0]) begin
        image_1_284 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_285 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h11d == _T_37[9:0]) begin
        image_1_285 <= io_pixelVal_in_1_7;
      end else if (10'h11d == _T_34[9:0]) begin
        image_1_285 <= io_pixelVal_in_1_6;
      end else if (10'h11d == _T_31[9:0]) begin
        image_1_285 <= io_pixelVal_in_1_5;
      end else if (10'h11d == _T_28[9:0]) begin
        image_1_285 <= io_pixelVal_in_1_4;
      end else if (10'h11d == _T_25[9:0]) begin
        image_1_285 <= io_pixelVal_in_1_3;
      end else if (10'h11d == _T_22[9:0]) begin
        image_1_285 <= io_pixelVal_in_1_2;
      end else if (10'h11d == _T_19[9:0]) begin
        image_1_285 <= io_pixelVal_in_1_1;
      end else if (10'h11d == _T_15[9:0]) begin
        image_1_285 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_286 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h11e == _T_37[9:0]) begin
        image_1_286 <= io_pixelVal_in_1_7;
      end else if (10'h11e == _T_34[9:0]) begin
        image_1_286 <= io_pixelVal_in_1_6;
      end else if (10'h11e == _T_31[9:0]) begin
        image_1_286 <= io_pixelVal_in_1_5;
      end else if (10'h11e == _T_28[9:0]) begin
        image_1_286 <= io_pixelVal_in_1_4;
      end else if (10'h11e == _T_25[9:0]) begin
        image_1_286 <= io_pixelVal_in_1_3;
      end else if (10'h11e == _T_22[9:0]) begin
        image_1_286 <= io_pixelVal_in_1_2;
      end else if (10'h11e == _T_19[9:0]) begin
        image_1_286 <= io_pixelVal_in_1_1;
      end else if (10'h11e == _T_15[9:0]) begin
        image_1_286 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_287 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h11f == _T_37[9:0]) begin
        image_1_287 <= io_pixelVal_in_1_7;
      end else if (10'h11f == _T_34[9:0]) begin
        image_1_287 <= io_pixelVal_in_1_6;
      end else if (10'h11f == _T_31[9:0]) begin
        image_1_287 <= io_pixelVal_in_1_5;
      end else if (10'h11f == _T_28[9:0]) begin
        image_1_287 <= io_pixelVal_in_1_4;
      end else if (10'h11f == _T_25[9:0]) begin
        image_1_287 <= io_pixelVal_in_1_3;
      end else if (10'h11f == _T_22[9:0]) begin
        image_1_287 <= io_pixelVal_in_1_2;
      end else if (10'h11f == _T_19[9:0]) begin
        image_1_287 <= io_pixelVal_in_1_1;
      end else if (10'h11f == _T_15[9:0]) begin
        image_1_287 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_288 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h120 == _T_37[9:0]) begin
        image_1_288 <= io_pixelVal_in_1_7;
      end else if (10'h120 == _T_34[9:0]) begin
        image_1_288 <= io_pixelVal_in_1_6;
      end else if (10'h120 == _T_31[9:0]) begin
        image_1_288 <= io_pixelVal_in_1_5;
      end else if (10'h120 == _T_28[9:0]) begin
        image_1_288 <= io_pixelVal_in_1_4;
      end else if (10'h120 == _T_25[9:0]) begin
        image_1_288 <= io_pixelVal_in_1_3;
      end else if (10'h120 == _T_22[9:0]) begin
        image_1_288 <= io_pixelVal_in_1_2;
      end else if (10'h120 == _T_19[9:0]) begin
        image_1_288 <= io_pixelVal_in_1_1;
      end else if (10'h120 == _T_15[9:0]) begin
        image_1_288 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_289 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h121 == _T_37[9:0]) begin
        image_1_289 <= io_pixelVal_in_1_7;
      end else if (10'h121 == _T_34[9:0]) begin
        image_1_289 <= io_pixelVal_in_1_6;
      end else if (10'h121 == _T_31[9:0]) begin
        image_1_289 <= io_pixelVal_in_1_5;
      end else if (10'h121 == _T_28[9:0]) begin
        image_1_289 <= io_pixelVal_in_1_4;
      end else if (10'h121 == _T_25[9:0]) begin
        image_1_289 <= io_pixelVal_in_1_3;
      end else if (10'h121 == _T_22[9:0]) begin
        image_1_289 <= io_pixelVal_in_1_2;
      end else if (10'h121 == _T_19[9:0]) begin
        image_1_289 <= io_pixelVal_in_1_1;
      end else if (10'h121 == _T_15[9:0]) begin
        image_1_289 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_290 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h122 == _T_37[9:0]) begin
        image_1_290 <= io_pixelVal_in_1_7;
      end else if (10'h122 == _T_34[9:0]) begin
        image_1_290 <= io_pixelVal_in_1_6;
      end else if (10'h122 == _T_31[9:0]) begin
        image_1_290 <= io_pixelVal_in_1_5;
      end else if (10'h122 == _T_28[9:0]) begin
        image_1_290 <= io_pixelVal_in_1_4;
      end else if (10'h122 == _T_25[9:0]) begin
        image_1_290 <= io_pixelVal_in_1_3;
      end else if (10'h122 == _T_22[9:0]) begin
        image_1_290 <= io_pixelVal_in_1_2;
      end else if (10'h122 == _T_19[9:0]) begin
        image_1_290 <= io_pixelVal_in_1_1;
      end else if (10'h122 == _T_15[9:0]) begin
        image_1_290 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_291 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h123 == _T_37[9:0]) begin
        image_1_291 <= io_pixelVal_in_1_7;
      end else if (10'h123 == _T_34[9:0]) begin
        image_1_291 <= io_pixelVal_in_1_6;
      end else if (10'h123 == _T_31[9:0]) begin
        image_1_291 <= io_pixelVal_in_1_5;
      end else if (10'h123 == _T_28[9:0]) begin
        image_1_291 <= io_pixelVal_in_1_4;
      end else if (10'h123 == _T_25[9:0]) begin
        image_1_291 <= io_pixelVal_in_1_3;
      end else if (10'h123 == _T_22[9:0]) begin
        image_1_291 <= io_pixelVal_in_1_2;
      end else if (10'h123 == _T_19[9:0]) begin
        image_1_291 <= io_pixelVal_in_1_1;
      end else if (10'h123 == _T_15[9:0]) begin
        image_1_291 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_292 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h124 == _T_37[9:0]) begin
        image_1_292 <= io_pixelVal_in_1_7;
      end else if (10'h124 == _T_34[9:0]) begin
        image_1_292 <= io_pixelVal_in_1_6;
      end else if (10'h124 == _T_31[9:0]) begin
        image_1_292 <= io_pixelVal_in_1_5;
      end else if (10'h124 == _T_28[9:0]) begin
        image_1_292 <= io_pixelVal_in_1_4;
      end else if (10'h124 == _T_25[9:0]) begin
        image_1_292 <= io_pixelVal_in_1_3;
      end else if (10'h124 == _T_22[9:0]) begin
        image_1_292 <= io_pixelVal_in_1_2;
      end else if (10'h124 == _T_19[9:0]) begin
        image_1_292 <= io_pixelVal_in_1_1;
      end else if (10'h124 == _T_15[9:0]) begin
        image_1_292 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_293 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h125 == _T_37[9:0]) begin
        image_1_293 <= io_pixelVal_in_1_7;
      end else if (10'h125 == _T_34[9:0]) begin
        image_1_293 <= io_pixelVal_in_1_6;
      end else if (10'h125 == _T_31[9:0]) begin
        image_1_293 <= io_pixelVal_in_1_5;
      end else if (10'h125 == _T_28[9:0]) begin
        image_1_293 <= io_pixelVal_in_1_4;
      end else if (10'h125 == _T_25[9:0]) begin
        image_1_293 <= io_pixelVal_in_1_3;
      end else if (10'h125 == _T_22[9:0]) begin
        image_1_293 <= io_pixelVal_in_1_2;
      end else if (10'h125 == _T_19[9:0]) begin
        image_1_293 <= io_pixelVal_in_1_1;
      end else if (10'h125 == _T_15[9:0]) begin
        image_1_293 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_294 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h126 == _T_37[9:0]) begin
        image_1_294 <= io_pixelVal_in_1_7;
      end else if (10'h126 == _T_34[9:0]) begin
        image_1_294 <= io_pixelVal_in_1_6;
      end else if (10'h126 == _T_31[9:0]) begin
        image_1_294 <= io_pixelVal_in_1_5;
      end else if (10'h126 == _T_28[9:0]) begin
        image_1_294 <= io_pixelVal_in_1_4;
      end else if (10'h126 == _T_25[9:0]) begin
        image_1_294 <= io_pixelVal_in_1_3;
      end else if (10'h126 == _T_22[9:0]) begin
        image_1_294 <= io_pixelVal_in_1_2;
      end else if (10'h126 == _T_19[9:0]) begin
        image_1_294 <= io_pixelVal_in_1_1;
      end else if (10'h126 == _T_15[9:0]) begin
        image_1_294 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_295 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h127 == _T_37[9:0]) begin
        image_1_295 <= io_pixelVal_in_1_7;
      end else if (10'h127 == _T_34[9:0]) begin
        image_1_295 <= io_pixelVal_in_1_6;
      end else if (10'h127 == _T_31[9:0]) begin
        image_1_295 <= io_pixelVal_in_1_5;
      end else if (10'h127 == _T_28[9:0]) begin
        image_1_295 <= io_pixelVal_in_1_4;
      end else if (10'h127 == _T_25[9:0]) begin
        image_1_295 <= io_pixelVal_in_1_3;
      end else if (10'h127 == _T_22[9:0]) begin
        image_1_295 <= io_pixelVal_in_1_2;
      end else if (10'h127 == _T_19[9:0]) begin
        image_1_295 <= io_pixelVal_in_1_1;
      end else if (10'h127 == _T_15[9:0]) begin
        image_1_295 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_296 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h128 == _T_37[9:0]) begin
        image_1_296 <= io_pixelVal_in_1_7;
      end else if (10'h128 == _T_34[9:0]) begin
        image_1_296 <= io_pixelVal_in_1_6;
      end else if (10'h128 == _T_31[9:0]) begin
        image_1_296 <= io_pixelVal_in_1_5;
      end else if (10'h128 == _T_28[9:0]) begin
        image_1_296 <= io_pixelVal_in_1_4;
      end else if (10'h128 == _T_25[9:0]) begin
        image_1_296 <= io_pixelVal_in_1_3;
      end else if (10'h128 == _T_22[9:0]) begin
        image_1_296 <= io_pixelVal_in_1_2;
      end else if (10'h128 == _T_19[9:0]) begin
        image_1_296 <= io_pixelVal_in_1_1;
      end else if (10'h128 == _T_15[9:0]) begin
        image_1_296 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_297 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h129 == _T_37[9:0]) begin
        image_1_297 <= io_pixelVal_in_1_7;
      end else if (10'h129 == _T_34[9:0]) begin
        image_1_297 <= io_pixelVal_in_1_6;
      end else if (10'h129 == _T_31[9:0]) begin
        image_1_297 <= io_pixelVal_in_1_5;
      end else if (10'h129 == _T_28[9:0]) begin
        image_1_297 <= io_pixelVal_in_1_4;
      end else if (10'h129 == _T_25[9:0]) begin
        image_1_297 <= io_pixelVal_in_1_3;
      end else if (10'h129 == _T_22[9:0]) begin
        image_1_297 <= io_pixelVal_in_1_2;
      end else if (10'h129 == _T_19[9:0]) begin
        image_1_297 <= io_pixelVal_in_1_1;
      end else if (10'h129 == _T_15[9:0]) begin
        image_1_297 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_298 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h12a == _T_37[9:0]) begin
        image_1_298 <= io_pixelVal_in_1_7;
      end else if (10'h12a == _T_34[9:0]) begin
        image_1_298 <= io_pixelVal_in_1_6;
      end else if (10'h12a == _T_31[9:0]) begin
        image_1_298 <= io_pixelVal_in_1_5;
      end else if (10'h12a == _T_28[9:0]) begin
        image_1_298 <= io_pixelVal_in_1_4;
      end else if (10'h12a == _T_25[9:0]) begin
        image_1_298 <= io_pixelVal_in_1_3;
      end else if (10'h12a == _T_22[9:0]) begin
        image_1_298 <= io_pixelVal_in_1_2;
      end else if (10'h12a == _T_19[9:0]) begin
        image_1_298 <= io_pixelVal_in_1_1;
      end else if (10'h12a == _T_15[9:0]) begin
        image_1_298 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_299 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h12b == _T_37[9:0]) begin
        image_1_299 <= io_pixelVal_in_1_7;
      end else if (10'h12b == _T_34[9:0]) begin
        image_1_299 <= io_pixelVal_in_1_6;
      end else if (10'h12b == _T_31[9:0]) begin
        image_1_299 <= io_pixelVal_in_1_5;
      end else if (10'h12b == _T_28[9:0]) begin
        image_1_299 <= io_pixelVal_in_1_4;
      end else if (10'h12b == _T_25[9:0]) begin
        image_1_299 <= io_pixelVal_in_1_3;
      end else if (10'h12b == _T_22[9:0]) begin
        image_1_299 <= io_pixelVal_in_1_2;
      end else if (10'h12b == _T_19[9:0]) begin
        image_1_299 <= io_pixelVal_in_1_1;
      end else if (10'h12b == _T_15[9:0]) begin
        image_1_299 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_300 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h12c == _T_37[9:0]) begin
        image_1_300 <= io_pixelVal_in_1_7;
      end else if (10'h12c == _T_34[9:0]) begin
        image_1_300 <= io_pixelVal_in_1_6;
      end else if (10'h12c == _T_31[9:0]) begin
        image_1_300 <= io_pixelVal_in_1_5;
      end else if (10'h12c == _T_28[9:0]) begin
        image_1_300 <= io_pixelVal_in_1_4;
      end else if (10'h12c == _T_25[9:0]) begin
        image_1_300 <= io_pixelVal_in_1_3;
      end else if (10'h12c == _T_22[9:0]) begin
        image_1_300 <= io_pixelVal_in_1_2;
      end else if (10'h12c == _T_19[9:0]) begin
        image_1_300 <= io_pixelVal_in_1_1;
      end else if (10'h12c == _T_15[9:0]) begin
        image_1_300 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_301 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h12d == _T_37[9:0]) begin
        image_1_301 <= io_pixelVal_in_1_7;
      end else if (10'h12d == _T_34[9:0]) begin
        image_1_301 <= io_pixelVal_in_1_6;
      end else if (10'h12d == _T_31[9:0]) begin
        image_1_301 <= io_pixelVal_in_1_5;
      end else if (10'h12d == _T_28[9:0]) begin
        image_1_301 <= io_pixelVal_in_1_4;
      end else if (10'h12d == _T_25[9:0]) begin
        image_1_301 <= io_pixelVal_in_1_3;
      end else if (10'h12d == _T_22[9:0]) begin
        image_1_301 <= io_pixelVal_in_1_2;
      end else if (10'h12d == _T_19[9:0]) begin
        image_1_301 <= io_pixelVal_in_1_1;
      end else if (10'h12d == _T_15[9:0]) begin
        image_1_301 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_302 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h12e == _T_37[9:0]) begin
        image_1_302 <= io_pixelVal_in_1_7;
      end else if (10'h12e == _T_34[9:0]) begin
        image_1_302 <= io_pixelVal_in_1_6;
      end else if (10'h12e == _T_31[9:0]) begin
        image_1_302 <= io_pixelVal_in_1_5;
      end else if (10'h12e == _T_28[9:0]) begin
        image_1_302 <= io_pixelVal_in_1_4;
      end else if (10'h12e == _T_25[9:0]) begin
        image_1_302 <= io_pixelVal_in_1_3;
      end else if (10'h12e == _T_22[9:0]) begin
        image_1_302 <= io_pixelVal_in_1_2;
      end else if (10'h12e == _T_19[9:0]) begin
        image_1_302 <= io_pixelVal_in_1_1;
      end else if (10'h12e == _T_15[9:0]) begin
        image_1_302 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_303 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h12f == _T_37[9:0]) begin
        image_1_303 <= io_pixelVal_in_1_7;
      end else if (10'h12f == _T_34[9:0]) begin
        image_1_303 <= io_pixelVal_in_1_6;
      end else if (10'h12f == _T_31[9:0]) begin
        image_1_303 <= io_pixelVal_in_1_5;
      end else if (10'h12f == _T_28[9:0]) begin
        image_1_303 <= io_pixelVal_in_1_4;
      end else if (10'h12f == _T_25[9:0]) begin
        image_1_303 <= io_pixelVal_in_1_3;
      end else if (10'h12f == _T_22[9:0]) begin
        image_1_303 <= io_pixelVal_in_1_2;
      end else if (10'h12f == _T_19[9:0]) begin
        image_1_303 <= io_pixelVal_in_1_1;
      end else if (10'h12f == _T_15[9:0]) begin
        image_1_303 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_304 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h130 == _T_37[9:0]) begin
        image_1_304 <= io_pixelVal_in_1_7;
      end else if (10'h130 == _T_34[9:0]) begin
        image_1_304 <= io_pixelVal_in_1_6;
      end else if (10'h130 == _T_31[9:0]) begin
        image_1_304 <= io_pixelVal_in_1_5;
      end else if (10'h130 == _T_28[9:0]) begin
        image_1_304 <= io_pixelVal_in_1_4;
      end else if (10'h130 == _T_25[9:0]) begin
        image_1_304 <= io_pixelVal_in_1_3;
      end else if (10'h130 == _T_22[9:0]) begin
        image_1_304 <= io_pixelVal_in_1_2;
      end else if (10'h130 == _T_19[9:0]) begin
        image_1_304 <= io_pixelVal_in_1_1;
      end else if (10'h130 == _T_15[9:0]) begin
        image_1_304 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_305 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h131 == _T_37[9:0]) begin
        image_1_305 <= io_pixelVal_in_1_7;
      end else if (10'h131 == _T_34[9:0]) begin
        image_1_305 <= io_pixelVal_in_1_6;
      end else if (10'h131 == _T_31[9:0]) begin
        image_1_305 <= io_pixelVal_in_1_5;
      end else if (10'h131 == _T_28[9:0]) begin
        image_1_305 <= io_pixelVal_in_1_4;
      end else if (10'h131 == _T_25[9:0]) begin
        image_1_305 <= io_pixelVal_in_1_3;
      end else if (10'h131 == _T_22[9:0]) begin
        image_1_305 <= io_pixelVal_in_1_2;
      end else if (10'h131 == _T_19[9:0]) begin
        image_1_305 <= io_pixelVal_in_1_1;
      end else if (10'h131 == _T_15[9:0]) begin
        image_1_305 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_306 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h132 == _T_37[9:0]) begin
        image_1_306 <= io_pixelVal_in_1_7;
      end else if (10'h132 == _T_34[9:0]) begin
        image_1_306 <= io_pixelVal_in_1_6;
      end else if (10'h132 == _T_31[9:0]) begin
        image_1_306 <= io_pixelVal_in_1_5;
      end else if (10'h132 == _T_28[9:0]) begin
        image_1_306 <= io_pixelVal_in_1_4;
      end else if (10'h132 == _T_25[9:0]) begin
        image_1_306 <= io_pixelVal_in_1_3;
      end else if (10'h132 == _T_22[9:0]) begin
        image_1_306 <= io_pixelVal_in_1_2;
      end else if (10'h132 == _T_19[9:0]) begin
        image_1_306 <= io_pixelVal_in_1_1;
      end else if (10'h132 == _T_15[9:0]) begin
        image_1_306 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_307 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h133 == _T_37[9:0]) begin
        image_1_307 <= io_pixelVal_in_1_7;
      end else if (10'h133 == _T_34[9:0]) begin
        image_1_307 <= io_pixelVal_in_1_6;
      end else if (10'h133 == _T_31[9:0]) begin
        image_1_307 <= io_pixelVal_in_1_5;
      end else if (10'h133 == _T_28[9:0]) begin
        image_1_307 <= io_pixelVal_in_1_4;
      end else if (10'h133 == _T_25[9:0]) begin
        image_1_307 <= io_pixelVal_in_1_3;
      end else if (10'h133 == _T_22[9:0]) begin
        image_1_307 <= io_pixelVal_in_1_2;
      end else if (10'h133 == _T_19[9:0]) begin
        image_1_307 <= io_pixelVal_in_1_1;
      end else if (10'h133 == _T_15[9:0]) begin
        image_1_307 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_308 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h134 == _T_37[9:0]) begin
        image_1_308 <= io_pixelVal_in_1_7;
      end else if (10'h134 == _T_34[9:0]) begin
        image_1_308 <= io_pixelVal_in_1_6;
      end else if (10'h134 == _T_31[9:0]) begin
        image_1_308 <= io_pixelVal_in_1_5;
      end else if (10'h134 == _T_28[9:0]) begin
        image_1_308 <= io_pixelVal_in_1_4;
      end else if (10'h134 == _T_25[9:0]) begin
        image_1_308 <= io_pixelVal_in_1_3;
      end else if (10'h134 == _T_22[9:0]) begin
        image_1_308 <= io_pixelVal_in_1_2;
      end else if (10'h134 == _T_19[9:0]) begin
        image_1_308 <= io_pixelVal_in_1_1;
      end else if (10'h134 == _T_15[9:0]) begin
        image_1_308 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_309 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h135 == _T_37[9:0]) begin
        image_1_309 <= io_pixelVal_in_1_7;
      end else if (10'h135 == _T_34[9:0]) begin
        image_1_309 <= io_pixelVal_in_1_6;
      end else if (10'h135 == _T_31[9:0]) begin
        image_1_309 <= io_pixelVal_in_1_5;
      end else if (10'h135 == _T_28[9:0]) begin
        image_1_309 <= io_pixelVal_in_1_4;
      end else if (10'h135 == _T_25[9:0]) begin
        image_1_309 <= io_pixelVal_in_1_3;
      end else if (10'h135 == _T_22[9:0]) begin
        image_1_309 <= io_pixelVal_in_1_2;
      end else if (10'h135 == _T_19[9:0]) begin
        image_1_309 <= io_pixelVal_in_1_1;
      end else if (10'h135 == _T_15[9:0]) begin
        image_1_309 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_310 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h136 == _T_37[9:0]) begin
        image_1_310 <= io_pixelVal_in_1_7;
      end else if (10'h136 == _T_34[9:0]) begin
        image_1_310 <= io_pixelVal_in_1_6;
      end else if (10'h136 == _T_31[9:0]) begin
        image_1_310 <= io_pixelVal_in_1_5;
      end else if (10'h136 == _T_28[9:0]) begin
        image_1_310 <= io_pixelVal_in_1_4;
      end else if (10'h136 == _T_25[9:0]) begin
        image_1_310 <= io_pixelVal_in_1_3;
      end else if (10'h136 == _T_22[9:0]) begin
        image_1_310 <= io_pixelVal_in_1_2;
      end else if (10'h136 == _T_19[9:0]) begin
        image_1_310 <= io_pixelVal_in_1_1;
      end else if (10'h136 == _T_15[9:0]) begin
        image_1_310 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_311 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h137 == _T_37[9:0]) begin
        image_1_311 <= io_pixelVal_in_1_7;
      end else if (10'h137 == _T_34[9:0]) begin
        image_1_311 <= io_pixelVal_in_1_6;
      end else if (10'h137 == _T_31[9:0]) begin
        image_1_311 <= io_pixelVal_in_1_5;
      end else if (10'h137 == _T_28[9:0]) begin
        image_1_311 <= io_pixelVal_in_1_4;
      end else if (10'h137 == _T_25[9:0]) begin
        image_1_311 <= io_pixelVal_in_1_3;
      end else if (10'h137 == _T_22[9:0]) begin
        image_1_311 <= io_pixelVal_in_1_2;
      end else if (10'h137 == _T_19[9:0]) begin
        image_1_311 <= io_pixelVal_in_1_1;
      end else if (10'h137 == _T_15[9:0]) begin
        image_1_311 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_312 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h138 == _T_37[9:0]) begin
        image_1_312 <= io_pixelVal_in_1_7;
      end else if (10'h138 == _T_34[9:0]) begin
        image_1_312 <= io_pixelVal_in_1_6;
      end else if (10'h138 == _T_31[9:0]) begin
        image_1_312 <= io_pixelVal_in_1_5;
      end else if (10'h138 == _T_28[9:0]) begin
        image_1_312 <= io_pixelVal_in_1_4;
      end else if (10'h138 == _T_25[9:0]) begin
        image_1_312 <= io_pixelVal_in_1_3;
      end else if (10'h138 == _T_22[9:0]) begin
        image_1_312 <= io_pixelVal_in_1_2;
      end else if (10'h138 == _T_19[9:0]) begin
        image_1_312 <= io_pixelVal_in_1_1;
      end else if (10'h138 == _T_15[9:0]) begin
        image_1_312 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_313 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h139 == _T_37[9:0]) begin
        image_1_313 <= io_pixelVal_in_1_7;
      end else if (10'h139 == _T_34[9:0]) begin
        image_1_313 <= io_pixelVal_in_1_6;
      end else if (10'h139 == _T_31[9:0]) begin
        image_1_313 <= io_pixelVal_in_1_5;
      end else if (10'h139 == _T_28[9:0]) begin
        image_1_313 <= io_pixelVal_in_1_4;
      end else if (10'h139 == _T_25[9:0]) begin
        image_1_313 <= io_pixelVal_in_1_3;
      end else if (10'h139 == _T_22[9:0]) begin
        image_1_313 <= io_pixelVal_in_1_2;
      end else if (10'h139 == _T_19[9:0]) begin
        image_1_313 <= io_pixelVal_in_1_1;
      end else if (10'h139 == _T_15[9:0]) begin
        image_1_313 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_314 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h13a == _T_37[9:0]) begin
        image_1_314 <= io_pixelVal_in_1_7;
      end else if (10'h13a == _T_34[9:0]) begin
        image_1_314 <= io_pixelVal_in_1_6;
      end else if (10'h13a == _T_31[9:0]) begin
        image_1_314 <= io_pixelVal_in_1_5;
      end else if (10'h13a == _T_28[9:0]) begin
        image_1_314 <= io_pixelVal_in_1_4;
      end else if (10'h13a == _T_25[9:0]) begin
        image_1_314 <= io_pixelVal_in_1_3;
      end else if (10'h13a == _T_22[9:0]) begin
        image_1_314 <= io_pixelVal_in_1_2;
      end else if (10'h13a == _T_19[9:0]) begin
        image_1_314 <= io_pixelVal_in_1_1;
      end else if (10'h13a == _T_15[9:0]) begin
        image_1_314 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_315 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h13b == _T_37[9:0]) begin
        image_1_315 <= io_pixelVal_in_1_7;
      end else if (10'h13b == _T_34[9:0]) begin
        image_1_315 <= io_pixelVal_in_1_6;
      end else if (10'h13b == _T_31[9:0]) begin
        image_1_315 <= io_pixelVal_in_1_5;
      end else if (10'h13b == _T_28[9:0]) begin
        image_1_315 <= io_pixelVal_in_1_4;
      end else if (10'h13b == _T_25[9:0]) begin
        image_1_315 <= io_pixelVal_in_1_3;
      end else if (10'h13b == _T_22[9:0]) begin
        image_1_315 <= io_pixelVal_in_1_2;
      end else if (10'h13b == _T_19[9:0]) begin
        image_1_315 <= io_pixelVal_in_1_1;
      end else if (10'h13b == _T_15[9:0]) begin
        image_1_315 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_316 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h13c == _T_37[9:0]) begin
        image_1_316 <= io_pixelVal_in_1_7;
      end else if (10'h13c == _T_34[9:0]) begin
        image_1_316 <= io_pixelVal_in_1_6;
      end else if (10'h13c == _T_31[9:0]) begin
        image_1_316 <= io_pixelVal_in_1_5;
      end else if (10'h13c == _T_28[9:0]) begin
        image_1_316 <= io_pixelVal_in_1_4;
      end else if (10'h13c == _T_25[9:0]) begin
        image_1_316 <= io_pixelVal_in_1_3;
      end else if (10'h13c == _T_22[9:0]) begin
        image_1_316 <= io_pixelVal_in_1_2;
      end else if (10'h13c == _T_19[9:0]) begin
        image_1_316 <= io_pixelVal_in_1_1;
      end else if (10'h13c == _T_15[9:0]) begin
        image_1_316 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_317 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h13d == _T_37[9:0]) begin
        image_1_317 <= io_pixelVal_in_1_7;
      end else if (10'h13d == _T_34[9:0]) begin
        image_1_317 <= io_pixelVal_in_1_6;
      end else if (10'h13d == _T_31[9:0]) begin
        image_1_317 <= io_pixelVal_in_1_5;
      end else if (10'h13d == _T_28[9:0]) begin
        image_1_317 <= io_pixelVal_in_1_4;
      end else if (10'h13d == _T_25[9:0]) begin
        image_1_317 <= io_pixelVal_in_1_3;
      end else if (10'h13d == _T_22[9:0]) begin
        image_1_317 <= io_pixelVal_in_1_2;
      end else if (10'h13d == _T_19[9:0]) begin
        image_1_317 <= io_pixelVal_in_1_1;
      end else if (10'h13d == _T_15[9:0]) begin
        image_1_317 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_318 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h13e == _T_37[9:0]) begin
        image_1_318 <= io_pixelVal_in_1_7;
      end else if (10'h13e == _T_34[9:0]) begin
        image_1_318 <= io_pixelVal_in_1_6;
      end else if (10'h13e == _T_31[9:0]) begin
        image_1_318 <= io_pixelVal_in_1_5;
      end else if (10'h13e == _T_28[9:0]) begin
        image_1_318 <= io_pixelVal_in_1_4;
      end else if (10'h13e == _T_25[9:0]) begin
        image_1_318 <= io_pixelVal_in_1_3;
      end else if (10'h13e == _T_22[9:0]) begin
        image_1_318 <= io_pixelVal_in_1_2;
      end else if (10'h13e == _T_19[9:0]) begin
        image_1_318 <= io_pixelVal_in_1_1;
      end else if (10'h13e == _T_15[9:0]) begin
        image_1_318 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_319 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h13f == _T_37[9:0]) begin
        image_1_319 <= io_pixelVal_in_1_7;
      end else if (10'h13f == _T_34[9:0]) begin
        image_1_319 <= io_pixelVal_in_1_6;
      end else if (10'h13f == _T_31[9:0]) begin
        image_1_319 <= io_pixelVal_in_1_5;
      end else if (10'h13f == _T_28[9:0]) begin
        image_1_319 <= io_pixelVal_in_1_4;
      end else if (10'h13f == _T_25[9:0]) begin
        image_1_319 <= io_pixelVal_in_1_3;
      end else if (10'h13f == _T_22[9:0]) begin
        image_1_319 <= io_pixelVal_in_1_2;
      end else if (10'h13f == _T_19[9:0]) begin
        image_1_319 <= io_pixelVal_in_1_1;
      end else if (10'h13f == _T_15[9:0]) begin
        image_1_319 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_320 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h140 == _T_37[9:0]) begin
        image_1_320 <= io_pixelVal_in_1_7;
      end else if (10'h140 == _T_34[9:0]) begin
        image_1_320 <= io_pixelVal_in_1_6;
      end else if (10'h140 == _T_31[9:0]) begin
        image_1_320 <= io_pixelVal_in_1_5;
      end else if (10'h140 == _T_28[9:0]) begin
        image_1_320 <= io_pixelVal_in_1_4;
      end else if (10'h140 == _T_25[9:0]) begin
        image_1_320 <= io_pixelVal_in_1_3;
      end else if (10'h140 == _T_22[9:0]) begin
        image_1_320 <= io_pixelVal_in_1_2;
      end else if (10'h140 == _T_19[9:0]) begin
        image_1_320 <= io_pixelVal_in_1_1;
      end else if (10'h140 == _T_15[9:0]) begin
        image_1_320 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_321 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h141 == _T_37[9:0]) begin
        image_1_321 <= io_pixelVal_in_1_7;
      end else if (10'h141 == _T_34[9:0]) begin
        image_1_321 <= io_pixelVal_in_1_6;
      end else if (10'h141 == _T_31[9:0]) begin
        image_1_321 <= io_pixelVal_in_1_5;
      end else if (10'h141 == _T_28[9:0]) begin
        image_1_321 <= io_pixelVal_in_1_4;
      end else if (10'h141 == _T_25[9:0]) begin
        image_1_321 <= io_pixelVal_in_1_3;
      end else if (10'h141 == _T_22[9:0]) begin
        image_1_321 <= io_pixelVal_in_1_2;
      end else if (10'h141 == _T_19[9:0]) begin
        image_1_321 <= io_pixelVal_in_1_1;
      end else if (10'h141 == _T_15[9:0]) begin
        image_1_321 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_322 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h142 == _T_37[9:0]) begin
        image_1_322 <= io_pixelVal_in_1_7;
      end else if (10'h142 == _T_34[9:0]) begin
        image_1_322 <= io_pixelVal_in_1_6;
      end else if (10'h142 == _T_31[9:0]) begin
        image_1_322 <= io_pixelVal_in_1_5;
      end else if (10'h142 == _T_28[9:0]) begin
        image_1_322 <= io_pixelVal_in_1_4;
      end else if (10'h142 == _T_25[9:0]) begin
        image_1_322 <= io_pixelVal_in_1_3;
      end else if (10'h142 == _T_22[9:0]) begin
        image_1_322 <= io_pixelVal_in_1_2;
      end else if (10'h142 == _T_19[9:0]) begin
        image_1_322 <= io_pixelVal_in_1_1;
      end else if (10'h142 == _T_15[9:0]) begin
        image_1_322 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_323 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h143 == _T_37[9:0]) begin
        image_1_323 <= io_pixelVal_in_1_7;
      end else if (10'h143 == _T_34[9:0]) begin
        image_1_323 <= io_pixelVal_in_1_6;
      end else if (10'h143 == _T_31[9:0]) begin
        image_1_323 <= io_pixelVal_in_1_5;
      end else if (10'h143 == _T_28[9:0]) begin
        image_1_323 <= io_pixelVal_in_1_4;
      end else if (10'h143 == _T_25[9:0]) begin
        image_1_323 <= io_pixelVal_in_1_3;
      end else if (10'h143 == _T_22[9:0]) begin
        image_1_323 <= io_pixelVal_in_1_2;
      end else if (10'h143 == _T_19[9:0]) begin
        image_1_323 <= io_pixelVal_in_1_1;
      end else if (10'h143 == _T_15[9:0]) begin
        image_1_323 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_324 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h144 == _T_37[9:0]) begin
        image_1_324 <= io_pixelVal_in_1_7;
      end else if (10'h144 == _T_34[9:0]) begin
        image_1_324 <= io_pixelVal_in_1_6;
      end else if (10'h144 == _T_31[9:0]) begin
        image_1_324 <= io_pixelVal_in_1_5;
      end else if (10'h144 == _T_28[9:0]) begin
        image_1_324 <= io_pixelVal_in_1_4;
      end else if (10'h144 == _T_25[9:0]) begin
        image_1_324 <= io_pixelVal_in_1_3;
      end else if (10'h144 == _T_22[9:0]) begin
        image_1_324 <= io_pixelVal_in_1_2;
      end else if (10'h144 == _T_19[9:0]) begin
        image_1_324 <= io_pixelVal_in_1_1;
      end else if (10'h144 == _T_15[9:0]) begin
        image_1_324 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_325 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h145 == _T_37[9:0]) begin
        image_1_325 <= io_pixelVal_in_1_7;
      end else if (10'h145 == _T_34[9:0]) begin
        image_1_325 <= io_pixelVal_in_1_6;
      end else if (10'h145 == _T_31[9:0]) begin
        image_1_325 <= io_pixelVal_in_1_5;
      end else if (10'h145 == _T_28[9:0]) begin
        image_1_325 <= io_pixelVal_in_1_4;
      end else if (10'h145 == _T_25[9:0]) begin
        image_1_325 <= io_pixelVal_in_1_3;
      end else if (10'h145 == _T_22[9:0]) begin
        image_1_325 <= io_pixelVal_in_1_2;
      end else if (10'h145 == _T_19[9:0]) begin
        image_1_325 <= io_pixelVal_in_1_1;
      end else if (10'h145 == _T_15[9:0]) begin
        image_1_325 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_326 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h146 == _T_37[9:0]) begin
        image_1_326 <= io_pixelVal_in_1_7;
      end else if (10'h146 == _T_34[9:0]) begin
        image_1_326 <= io_pixelVal_in_1_6;
      end else if (10'h146 == _T_31[9:0]) begin
        image_1_326 <= io_pixelVal_in_1_5;
      end else if (10'h146 == _T_28[9:0]) begin
        image_1_326 <= io_pixelVal_in_1_4;
      end else if (10'h146 == _T_25[9:0]) begin
        image_1_326 <= io_pixelVal_in_1_3;
      end else if (10'h146 == _T_22[9:0]) begin
        image_1_326 <= io_pixelVal_in_1_2;
      end else if (10'h146 == _T_19[9:0]) begin
        image_1_326 <= io_pixelVal_in_1_1;
      end else if (10'h146 == _T_15[9:0]) begin
        image_1_326 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_327 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h147 == _T_37[9:0]) begin
        image_1_327 <= io_pixelVal_in_1_7;
      end else if (10'h147 == _T_34[9:0]) begin
        image_1_327 <= io_pixelVal_in_1_6;
      end else if (10'h147 == _T_31[9:0]) begin
        image_1_327 <= io_pixelVal_in_1_5;
      end else if (10'h147 == _T_28[9:0]) begin
        image_1_327 <= io_pixelVal_in_1_4;
      end else if (10'h147 == _T_25[9:0]) begin
        image_1_327 <= io_pixelVal_in_1_3;
      end else if (10'h147 == _T_22[9:0]) begin
        image_1_327 <= io_pixelVal_in_1_2;
      end else if (10'h147 == _T_19[9:0]) begin
        image_1_327 <= io_pixelVal_in_1_1;
      end else if (10'h147 == _T_15[9:0]) begin
        image_1_327 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_328 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h148 == _T_37[9:0]) begin
        image_1_328 <= io_pixelVal_in_1_7;
      end else if (10'h148 == _T_34[9:0]) begin
        image_1_328 <= io_pixelVal_in_1_6;
      end else if (10'h148 == _T_31[9:0]) begin
        image_1_328 <= io_pixelVal_in_1_5;
      end else if (10'h148 == _T_28[9:0]) begin
        image_1_328 <= io_pixelVal_in_1_4;
      end else if (10'h148 == _T_25[9:0]) begin
        image_1_328 <= io_pixelVal_in_1_3;
      end else if (10'h148 == _T_22[9:0]) begin
        image_1_328 <= io_pixelVal_in_1_2;
      end else if (10'h148 == _T_19[9:0]) begin
        image_1_328 <= io_pixelVal_in_1_1;
      end else if (10'h148 == _T_15[9:0]) begin
        image_1_328 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_329 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h149 == _T_37[9:0]) begin
        image_1_329 <= io_pixelVal_in_1_7;
      end else if (10'h149 == _T_34[9:0]) begin
        image_1_329 <= io_pixelVal_in_1_6;
      end else if (10'h149 == _T_31[9:0]) begin
        image_1_329 <= io_pixelVal_in_1_5;
      end else if (10'h149 == _T_28[9:0]) begin
        image_1_329 <= io_pixelVal_in_1_4;
      end else if (10'h149 == _T_25[9:0]) begin
        image_1_329 <= io_pixelVal_in_1_3;
      end else if (10'h149 == _T_22[9:0]) begin
        image_1_329 <= io_pixelVal_in_1_2;
      end else if (10'h149 == _T_19[9:0]) begin
        image_1_329 <= io_pixelVal_in_1_1;
      end else if (10'h149 == _T_15[9:0]) begin
        image_1_329 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_330 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h14a == _T_37[9:0]) begin
        image_1_330 <= io_pixelVal_in_1_7;
      end else if (10'h14a == _T_34[9:0]) begin
        image_1_330 <= io_pixelVal_in_1_6;
      end else if (10'h14a == _T_31[9:0]) begin
        image_1_330 <= io_pixelVal_in_1_5;
      end else if (10'h14a == _T_28[9:0]) begin
        image_1_330 <= io_pixelVal_in_1_4;
      end else if (10'h14a == _T_25[9:0]) begin
        image_1_330 <= io_pixelVal_in_1_3;
      end else if (10'h14a == _T_22[9:0]) begin
        image_1_330 <= io_pixelVal_in_1_2;
      end else if (10'h14a == _T_19[9:0]) begin
        image_1_330 <= io_pixelVal_in_1_1;
      end else if (10'h14a == _T_15[9:0]) begin
        image_1_330 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_331 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h14b == _T_37[9:0]) begin
        image_1_331 <= io_pixelVal_in_1_7;
      end else if (10'h14b == _T_34[9:0]) begin
        image_1_331 <= io_pixelVal_in_1_6;
      end else if (10'h14b == _T_31[9:0]) begin
        image_1_331 <= io_pixelVal_in_1_5;
      end else if (10'h14b == _T_28[9:0]) begin
        image_1_331 <= io_pixelVal_in_1_4;
      end else if (10'h14b == _T_25[9:0]) begin
        image_1_331 <= io_pixelVal_in_1_3;
      end else if (10'h14b == _T_22[9:0]) begin
        image_1_331 <= io_pixelVal_in_1_2;
      end else if (10'h14b == _T_19[9:0]) begin
        image_1_331 <= io_pixelVal_in_1_1;
      end else if (10'h14b == _T_15[9:0]) begin
        image_1_331 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_332 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h14c == _T_37[9:0]) begin
        image_1_332 <= io_pixelVal_in_1_7;
      end else if (10'h14c == _T_34[9:0]) begin
        image_1_332 <= io_pixelVal_in_1_6;
      end else if (10'h14c == _T_31[9:0]) begin
        image_1_332 <= io_pixelVal_in_1_5;
      end else if (10'h14c == _T_28[9:0]) begin
        image_1_332 <= io_pixelVal_in_1_4;
      end else if (10'h14c == _T_25[9:0]) begin
        image_1_332 <= io_pixelVal_in_1_3;
      end else if (10'h14c == _T_22[9:0]) begin
        image_1_332 <= io_pixelVal_in_1_2;
      end else if (10'h14c == _T_19[9:0]) begin
        image_1_332 <= io_pixelVal_in_1_1;
      end else if (10'h14c == _T_15[9:0]) begin
        image_1_332 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_333 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h14d == _T_37[9:0]) begin
        image_1_333 <= io_pixelVal_in_1_7;
      end else if (10'h14d == _T_34[9:0]) begin
        image_1_333 <= io_pixelVal_in_1_6;
      end else if (10'h14d == _T_31[9:0]) begin
        image_1_333 <= io_pixelVal_in_1_5;
      end else if (10'h14d == _T_28[9:0]) begin
        image_1_333 <= io_pixelVal_in_1_4;
      end else if (10'h14d == _T_25[9:0]) begin
        image_1_333 <= io_pixelVal_in_1_3;
      end else if (10'h14d == _T_22[9:0]) begin
        image_1_333 <= io_pixelVal_in_1_2;
      end else if (10'h14d == _T_19[9:0]) begin
        image_1_333 <= io_pixelVal_in_1_1;
      end else if (10'h14d == _T_15[9:0]) begin
        image_1_333 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_334 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h14e == _T_37[9:0]) begin
        image_1_334 <= io_pixelVal_in_1_7;
      end else if (10'h14e == _T_34[9:0]) begin
        image_1_334 <= io_pixelVal_in_1_6;
      end else if (10'h14e == _T_31[9:0]) begin
        image_1_334 <= io_pixelVal_in_1_5;
      end else if (10'h14e == _T_28[9:0]) begin
        image_1_334 <= io_pixelVal_in_1_4;
      end else if (10'h14e == _T_25[9:0]) begin
        image_1_334 <= io_pixelVal_in_1_3;
      end else if (10'h14e == _T_22[9:0]) begin
        image_1_334 <= io_pixelVal_in_1_2;
      end else if (10'h14e == _T_19[9:0]) begin
        image_1_334 <= io_pixelVal_in_1_1;
      end else if (10'h14e == _T_15[9:0]) begin
        image_1_334 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_335 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h14f == _T_37[9:0]) begin
        image_1_335 <= io_pixelVal_in_1_7;
      end else if (10'h14f == _T_34[9:0]) begin
        image_1_335 <= io_pixelVal_in_1_6;
      end else if (10'h14f == _T_31[9:0]) begin
        image_1_335 <= io_pixelVal_in_1_5;
      end else if (10'h14f == _T_28[9:0]) begin
        image_1_335 <= io_pixelVal_in_1_4;
      end else if (10'h14f == _T_25[9:0]) begin
        image_1_335 <= io_pixelVal_in_1_3;
      end else if (10'h14f == _T_22[9:0]) begin
        image_1_335 <= io_pixelVal_in_1_2;
      end else if (10'h14f == _T_19[9:0]) begin
        image_1_335 <= io_pixelVal_in_1_1;
      end else if (10'h14f == _T_15[9:0]) begin
        image_1_335 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_336 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h150 == _T_37[9:0]) begin
        image_1_336 <= io_pixelVal_in_1_7;
      end else if (10'h150 == _T_34[9:0]) begin
        image_1_336 <= io_pixelVal_in_1_6;
      end else if (10'h150 == _T_31[9:0]) begin
        image_1_336 <= io_pixelVal_in_1_5;
      end else if (10'h150 == _T_28[9:0]) begin
        image_1_336 <= io_pixelVal_in_1_4;
      end else if (10'h150 == _T_25[9:0]) begin
        image_1_336 <= io_pixelVal_in_1_3;
      end else if (10'h150 == _T_22[9:0]) begin
        image_1_336 <= io_pixelVal_in_1_2;
      end else if (10'h150 == _T_19[9:0]) begin
        image_1_336 <= io_pixelVal_in_1_1;
      end else if (10'h150 == _T_15[9:0]) begin
        image_1_336 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_337 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h151 == _T_37[9:0]) begin
        image_1_337 <= io_pixelVal_in_1_7;
      end else if (10'h151 == _T_34[9:0]) begin
        image_1_337 <= io_pixelVal_in_1_6;
      end else if (10'h151 == _T_31[9:0]) begin
        image_1_337 <= io_pixelVal_in_1_5;
      end else if (10'h151 == _T_28[9:0]) begin
        image_1_337 <= io_pixelVal_in_1_4;
      end else if (10'h151 == _T_25[9:0]) begin
        image_1_337 <= io_pixelVal_in_1_3;
      end else if (10'h151 == _T_22[9:0]) begin
        image_1_337 <= io_pixelVal_in_1_2;
      end else if (10'h151 == _T_19[9:0]) begin
        image_1_337 <= io_pixelVal_in_1_1;
      end else if (10'h151 == _T_15[9:0]) begin
        image_1_337 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_338 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h152 == _T_37[9:0]) begin
        image_1_338 <= io_pixelVal_in_1_7;
      end else if (10'h152 == _T_34[9:0]) begin
        image_1_338 <= io_pixelVal_in_1_6;
      end else if (10'h152 == _T_31[9:0]) begin
        image_1_338 <= io_pixelVal_in_1_5;
      end else if (10'h152 == _T_28[9:0]) begin
        image_1_338 <= io_pixelVal_in_1_4;
      end else if (10'h152 == _T_25[9:0]) begin
        image_1_338 <= io_pixelVal_in_1_3;
      end else if (10'h152 == _T_22[9:0]) begin
        image_1_338 <= io_pixelVal_in_1_2;
      end else if (10'h152 == _T_19[9:0]) begin
        image_1_338 <= io_pixelVal_in_1_1;
      end else if (10'h152 == _T_15[9:0]) begin
        image_1_338 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_339 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h153 == _T_37[9:0]) begin
        image_1_339 <= io_pixelVal_in_1_7;
      end else if (10'h153 == _T_34[9:0]) begin
        image_1_339 <= io_pixelVal_in_1_6;
      end else if (10'h153 == _T_31[9:0]) begin
        image_1_339 <= io_pixelVal_in_1_5;
      end else if (10'h153 == _T_28[9:0]) begin
        image_1_339 <= io_pixelVal_in_1_4;
      end else if (10'h153 == _T_25[9:0]) begin
        image_1_339 <= io_pixelVal_in_1_3;
      end else if (10'h153 == _T_22[9:0]) begin
        image_1_339 <= io_pixelVal_in_1_2;
      end else if (10'h153 == _T_19[9:0]) begin
        image_1_339 <= io_pixelVal_in_1_1;
      end else if (10'h153 == _T_15[9:0]) begin
        image_1_339 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_340 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h154 == _T_37[9:0]) begin
        image_1_340 <= io_pixelVal_in_1_7;
      end else if (10'h154 == _T_34[9:0]) begin
        image_1_340 <= io_pixelVal_in_1_6;
      end else if (10'h154 == _T_31[9:0]) begin
        image_1_340 <= io_pixelVal_in_1_5;
      end else if (10'h154 == _T_28[9:0]) begin
        image_1_340 <= io_pixelVal_in_1_4;
      end else if (10'h154 == _T_25[9:0]) begin
        image_1_340 <= io_pixelVal_in_1_3;
      end else if (10'h154 == _T_22[9:0]) begin
        image_1_340 <= io_pixelVal_in_1_2;
      end else if (10'h154 == _T_19[9:0]) begin
        image_1_340 <= io_pixelVal_in_1_1;
      end else if (10'h154 == _T_15[9:0]) begin
        image_1_340 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_341 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h155 == _T_37[9:0]) begin
        image_1_341 <= io_pixelVal_in_1_7;
      end else if (10'h155 == _T_34[9:0]) begin
        image_1_341 <= io_pixelVal_in_1_6;
      end else if (10'h155 == _T_31[9:0]) begin
        image_1_341 <= io_pixelVal_in_1_5;
      end else if (10'h155 == _T_28[9:0]) begin
        image_1_341 <= io_pixelVal_in_1_4;
      end else if (10'h155 == _T_25[9:0]) begin
        image_1_341 <= io_pixelVal_in_1_3;
      end else if (10'h155 == _T_22[9:0]) begin
        image_1_341 <= io_pixelVal_in_1_2;
      end else if (10'h155 == _T_19[9:0]) begin
        image_1_341 <= io_pixelVal_in_1_1;
      end else if (10'h155 == _T_15[9:0]) begin
        image_1_341 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_342 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h156 == _T_37[9:0]) begin
        image_1_342 <= io_pixelVal_in_1_7;
      end else if (10'h156 == _T_34[9:0]) begin
        image_1_342 <= io_pixelVal_in_1_6;
      end else if (10'h156 == _T_31[9:0]) begin
        image_1_342 <= io_pixelVal_in_1_5;
      end else if (10'h156 == _T_28[9:0]) begin
        image_1_342 <= io_pixelVal_in_1_4;
      end else if (10'h156 == _T_25[9:0]) begin
        image_1_342 <= io_pixelVal_in_1_3;
      end else if (10'h156 == _T_22[9:0]) begin
        image_1_342 <= io_pixelVal_in_1_2;
      end else if (10'h156 == _T_19[9:0]) begin
        image_1_342 <= io_pixelVal_in_1_1;
      end else if (10'h156 == _T_15[9:0]) begin
        image_1_342 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_343 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h157 == _T_37[9:0]) begin
        image_1_343 <= io_pixelVal_in_1_7;
      end else if (10'h157 == _T_34[9:0]) begin
        image_1_343 <= io_pixelVal_in_1_6;
      end else if (10'h157 == _T_31[9:0]) begin
        image_1_343 <= io_pixelVal_in_1_5;
      end else if (10'h157 == _T_28[9:0]) begin
        image_1_343 <= io_pixelVal_in_1_4;
      end else if (10'h157 == _T_25[9:0]) begin
        image_1_343 <= io_pixelVal_in_1_3;
      end else if (10'h157 == _T_22[9:0]) begin
        image_1_343 <= io_pixelVal_in_1_2;
      end else if (10'h157 == _T_19[9:0]) begin
        image_1_343 <= io_pixelVal_in_1_1;
      end else if (10'h157 == _T_15[9:0]) begin
        image_1_343 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_344 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h158 == _T_37[9:0]) begin
        image_1_344 <= io_pixelVal_in_1_7;
      end else if (10'h158 == _T_34[9:0]) begin
        image_1_344 <= io_pixelVal_in_1_6;
      end else if (10'h158 == _T_31[9:0]) begin
        image_1_344 <= io_pixelVal_in_1_5;
      end else if (10'h158 == _T_28[9:0]) begin
        image_1_344 <= io_pixelVal_in_1_4;
      end else if (10'h158 == _T_25[9:0]) begin
        image_1_344 <= io_pixelVal_in_1_3;
      end else if (10'h158 == _T_22[9:0]) begin
        image_1_344 <= io_pixelVal_in_1_2;
      end else if (10'h158 == _T_19[9:0]) begin
        image_1_344 <= io_pixelVal_in_1_1;
      end else if (10'h158 == _T_15[9:0]) begin
        image_1_344 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_345 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h159 == _T_37[9:0]) begin
        image_1_345 <= io_pixelVal_in_1_7;
      end else if (10'h159 == _T_34[9:0]) begin
        image_1_345 <= io_pixelVal_in_1_6;
      end else if (10'h159 == _T_31[9:0]) begin
        image_1_345 <= io_pixelVal_in_1_5;
      end else if (10'h159 == _T_28[9:0]) begin
        image_1_345 <= io_pixelVal_in_1_4;
      end else if (10'h159 == _T_25[9:0]) begin
        image_1_345 <= io_pixelVal_in_1_3;
      end else if (10'h159 == _T_22[9:0]) begin
        image_1_345 <= io_pixelVal_in_1_2;
      end else if (10'h159 == _T_19[9:0]) begin
        image_1_345 <= io_pixelVal_in_1_1;
      end else if (10'h159 == _T_15[9:0]) begin
        image_1_345 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_346 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h15a == _T_37[9:0]) begin
        image_1_346 <= io_pixelVal_in_1_7;
      end else if (10'h15a == _T_34[9:0]) begin
        image_1_346 <= io_pixelVal_in_1_6;
      end else if (10'h15a == _T_31[9:0]) begin
        image_1_346 <= io_pixelVal_in_1_5;
      end else if (10'h15a == _T_28[9:0]) begin
        image_1_346 <= io_pixelVal_in_1_4;
      end else if (10'h15a == _T_25[9:0]) begin
        image_1_346 <= io_pixelVal_in_1_3;
      end else if (10'h15a == _T_22[9:0]) begin
        image_1_346 <= io_pixelVal_in_1_2;
      end else if (10'h15a == _T_19[9:0]) begin
        image_1_346 <= io_pixelVal_in_1_1;
      end else if (10'h15a == _T_15[9:0]) begin
        image_1_346 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_347 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h15b == _T_37[9:0]) begin
        image_1_347 <= io_pixelVal_in_1_7;
      end else if (10'h15b == _T_34[9:0]) begin
        image_1_347 <= io_pixelVal_in_1_6;
      end else if (10'h15b == _T_31[9:0]) begin
        image_1_347 <= io_pixelVal_in_1_5;
      end else if (10'h15b == _T_28[9:0]) begin
        image_1_347 <= io_pixelVal_in_1_4;
      end else if (10'h15b == _T_25[9:0]) begin
        image_1_347 <= io_pixelVal_in_1_3;
      end else if (10'h15b == _T_22[9:0]) begin
        image_1_347 <= io_pixelVal_in_1_2;
      end else if (10'h15b == _T_19[9:0]) begin
        image_1_347 <= io_pixelVal_in_1_1;
      end else if (10'h15b == _T_15[9:0]) begin
        image_1_347 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_348 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h15c == _T_37[9:0]) begin
        image_1_348 <= io_pixelVal_in_1_7;
      end else if (10'h15c == _T_34[9:0]) begin
        image_1_348 <= io_pixelVal_in_1_6;
      end else if (10'h15c == _T_31[9:0]) begin
        image_1_348 <= io_pixelVal_in_1_5;
      end else if (10'h15c == _T_28[9:0]) begin
        image_1_348 <= io_pixelVal_in_1_4;
      end else if (10'h15c == _T_25[9:0]) begin
        image_1_348 <= io_pixelVal_in_1_3;
      end else if (10'h15c == _T_22[9:0]) begin
        image_1_348 <= io_pixelVal_in_1_2;
      end else if (10'h15c == _T_19[9:0]) begin
        image_1_348 <= io_pixelVal_in_1_1;
      end else if (10'h15c == _T_15[9:0]) begin
        image_1_348 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_349 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h15d == _T_37[9:0]) begin
        image_1_349 <= io_pixelVal_in_1_7;
      end else if (10'h15d == _T_34[9:0]) begin
        image_1_349 <= io_pixelVal_in_1_6;
      end else if (10'h15d == _T_31[9:0]) begin
        image_1_349 <= io_pixelVal_in_1_5;
      end else if (10'h15d == _T_28[9:0]) begin
        image_1_349 <= io_pixelVal_in_1_4;
      end else if (10'h15d == _T_25[9:0]) begin
        image_1_349 <= io_pixelVal_in_1_3;
      end else if (10'h15d == _T_22[9:0]) begin
        image_1_349 <= io_pixelVal_in_1_2;
      end else if (10'h15d == _T_19[9:0]) begin
        image_1_349 <= io_pixelVal_in_1_1;
      end else if (10'h15d == _T_15[9:0]) begin
        image_1_349 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_350 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h15e == _T_37[9:0]) begin
        image_1_350 <= io_pixelVal_in_1_7;
      end else if (10'h15e == _T_34[9:0]) begin
        image_1_350 <= io_pixelVal_in_1_6;
      end else if (10'h15e == _T_31[9:0]) begin
        image_1_350 <= io_pixelVal_in_1_5;
      end else if (10'h15e == _T_28[9:0]) begin
        image_1_350 <= io_pixelVal_in_1_4;
      end else if (10'h15e == _T_25[9:0]) begin
        image_1_350 <= io_pixelVal_in_1_3;
      end else if (10'h15e == _T_22[9:0]) begin
        image_1_350 <= io_pixelVal_in_1_2;
      end else if (10'h15e == _T_19[9:0]) begin
        image_1_350 <= io_pixelVal_in_1_1;
      end else if (10'h15e == _T_15[9:0]) begin
        image_1_350 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_351 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h15f == _T_37[9:0]) begin
        image_1_351 <= io_pixelVal_in_1_7;
      end else if (10'h15f == _T_34[9:0]) begin
        image_1_351 <= io_pixelVal_in_1_6;
      end else if (10'h15f == _T_31[9:0]) begin
        image_1_351 <= io_pixelVal_in_1_5;
      end else if (10'h15f == _T_28[9:0]) begin
        image_1_351 <= io_pixelVal_in_1_4;
      end else if (10'h15f == _T_25[9:0]) begin
        image_1_351 <= io_pixelVal_in_1_3;
      end else if (10'h15f == _T_22[9:0]) begin
        image_1_351 <= io_pixelVal_in_1_2;
      end else if (10'h15f == _T_19[9:0]) begin
        image_1_351 <= io_pixelVal_in_1_1;
      end else if (10'h15f == _T_15[9:0]) begin
        image_1_351 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_352 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h160 == _T_37[9:0]) begin
        image_1_352 <= io_pixelVal_in_1_7;
      end else if (10'h160 == _T_34[9:0]) begin
        image_1_352 <= io_pixelVal_in_1_6;
      end else if (10'h160 == _T_31[9:0]) begin
        image_1_352 <= io_pixelVal_in_1_5;
      end else if (10'h160 == _T_28[9:0]) begin
        image_1_352 <= io_pixelVal_in_1_4;
      end else if (10'h160 == _T_25[9:0]) begin
        image_1_352 <= io_pixelVal_in_1_3;
      end else if (10'h160 == _T_22[9:0]) begin
        image_1_352 <= io_pixelVal_in_1_2;
      end else if (10'h160 == _T_19[9:0]) begin
        image_1_352 <= io_pixelVal_in_1_1;
      end else if (10'h160 == _T_15[9:0]) begin
        image_1_352 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_353 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h161 == _T_37[9:0]) begin
        image_1_353 <= io_pixelVal_in_1_7;
      end else if (10'h161 == _T_34[9:0]) begin
        image_1_353 <= io_pixelVal_in_1_6;
      end else if (10'h161 == _T_31[9:0]) begin
        image_1_353 <= io_pixelVal_in_1_5;
      end else if (10'h161 == _T_28[9:0]) begin
        image_1_353 <= io_pixelVal_in_1_4;
      end else if (10'h161 == _T_25[9:0]) begin
        image_1_353 <= io_pixelVal_in_1_3;
      end else if (10'h161 == _T_22[9:0]) begin
        image_1_353 <= io_pixelVal_in_1_2;
      end else if (10'h161 == _T_19[9:0]) begin
        image_1_353 <= io_pixelVal_in_1_1;
      end else if (10'h161 == _T_15[9:0]) begin
        image_1_353 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_354 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h162 == _T_37[9:0]) begin
        image_1_354 <= io_pixelVal_in_1_7;
      end else if (10'h162 == _T_34[9:0]) begin
        image_1_354 <= io_pixelVal_in_1_6;
      end else if (10'h162 == _T_31[9:0]) begin
        image_1_354 <= io_pixelVal_in_1_5;
      end else if (10'h162 == _T_28[9:0]) begin
        image_1_354 <= io_pixelVal_in_1_4;
      end else if (10'h162 == _T_25[9:0]) begin
        image_1_354 <= io_pixelVal_in_1_3;
      end else if (10'h162 == _T_22[9:0]) begin
        image_1_354 <= io_pixelVal_in_1_2;
      end else if (10'h162 == _T_19[9:0]) begin
        image_1_354 <= io_pixelVal_in_1_1;
      end else if (10'h162 == _T_15[9:0]) begin
        image_1_354 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_355 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h163 == _T_37[9:0]) begin
        image_1_355 <= io_pixelVal_in_1_7;
      end else if (10'h163 == _T_34[9:0]) begin
        image_1_355 <= io_pixelVal_in_1_6;
      end else if (10'h163 == _T_31[9:0]) begin
        image_1_355 <= io_pixelVal_in_1_5;
      end else if (10'h163 == _T_28[9:0]) begin
        image_1_355 <= io_pixelVal_in_1_4;
      end else if (10'h163 == _T_25[9:0]) begin
        image_1_355 <= io_pixelVal_in_1_3;
      end else if (10'h163 == _T_22[9:0]) begin
        image_1_355 <= io_pixelVal_in_1_2;
      end else if (10'h163 == _T_19[9:0]) begin
        image_1_355 <= io_pixelVal_in_1_1;
      end else if (10'h163 == _T_15[9:0]) begin
        image_1_355 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_356 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h164 == _T_37[9:0]) begin
        image_1_356 <= io_pixelVal_in_1_7;
      end else if (10'h164 == _T_34[9:0]) begin
        image_1_356 <= io_pixelVal_in_1_6;
      end else if (10'h164 == _T_31[9:0]) begin
        image_1_356 <= io_pixelVal_in_1_5;
      end else if (10'h164 == _T_28[9:0]) begin
        image_1_356 <= io_pixelVal_in_1_4;
      end else if (10'h164 == _T_25[9:0]) begin
        image_1_356 <= io_pixelVal_in_1_3;
      end else if (10'h164 == _T_22[9:0]) begin
        image_1_356 <= io_pixelVal_in_1_2;
      end else if (10'h164 == _T_19[9:0]) begin
        image_1_356 <= io_pixelVal_in_1_1;
      end else if (10'h164 == _T_15[9:0]) begin
        image_1_356 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_357 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h165 == _T_37[9:0]) begin
        image_1_357 <= io_pixelVal_in_1_7;
      end else if (10'h165 == _T_34[9:0]) begin
        image_1_357 <= io_pixelVal_in_1_6;
      end else if (10'h165 == _T_31[9:0]) begin
        image_1_357 <= io_pixelVal_in_1_5;
      end else if (10'h165 == _T_28[9:0]) begin
        image_1_357 <= io_pixelVal_in_1_4;
      end else if (10'h165 == _T_25[9:0]) begin
        image_1_357 <= io_pixelVal_in_1_3;
      end else if (10'h165 == _T_22[9:0]) begin
        image_1_357 <= io_pixelVal_in_1_2;
      end else if (10'h165 == _T_19[9:0]) begin
        image_1_357 <= io_pixelVal_in_1_1;
      end else if (10'h165 == _T_15[9:0]) begin
        image_1_357 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_358 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h166 == _T_37[9:0]) begin
        image_1_358 <= io_pixelVal_in_1_7;
      end else if (10'h166 == _T_34[9:0]) begin
        image_1_358 <= io_pixelVal_in_1_6;
      end else if (10'h166 == _T_31[9:0]) begin
        image_1_358 <= io_pixelVal_in_1_5;
      end else if (10'h166 == _T_28[9:0]) begin
        image_1_358 <= io_pixelVal_in_1_4;
      end else if (10'h166 == _T_25[9:0]) begin
        image_1_358 <= io_pixelVal_in_1_3;
      end else if (10'h166 == _T_22[9:0]) begin
        image_1_358 <= io_pixelVal_in_1_2;
      end else if (10'h166 == _T_19[9:0]) begin
        image_1_358 <= io_pixelVal_in_1_1;
      end else if (10'h166 == _T_15[9:0]) begin
        image_1_358 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_359 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h167 == _T_37[9:0]) begin
        image_1_359 <= io_pixelVal_in_1_7;
      end else if (10'h167 == _T_34[9:0]) begin
        image_1_359 <= io_pixelVal_in_1_6;
      end else if (10'h167 == _T_31[9:0]) begin
        image_1_359 <= io_pixelVal_in_1_5;
      end else if (10'h167 == _T_28[9:0]) begin
        image_1_359 <= io_pixelVal_in_1_4;
      end else if (10'h167 == _T_25[9:0]) begin
        image_1_359 <= io_pixelVal_in_1_3;
      end else if (10'h167 == _T_22[9:0]) begin
        image_1_359 <= io_pixelVal_in_1_2;
      end else if (10'h167 == _T_19[9:0]) begin
        image_1_359 <= io_pixelVal_in_1_1;
      end else if (10'h167 == _T_15[9:0]) begin
        image_1_359 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_360 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h168 == _T_37[9:0]) begin
        image_1_360 <= io_pixelVal_in_1_7;
      end else if (10'h168 == _T_34[9:0]) begin
        image_1_360 <= io_pixelVal_in_1_6;
      end else if (10'h168 == _T_31[9:0]) begin
        image_1_360 <= io_pixelVal_in_1_5;
      end else if (10'h168 == _T_28[9:0]) begin
        image_1_360 <= io_pixelVal_in_1_4;
      end else if (10'h168 == _T_25[9:0]) begin
        image_1_360 <= io_pixelVal_in_1_3;
      end else if (10'h168 == _T_22[9:0]) begin
        image_1_360 <= io_pixelVal_in_1_2;
      end else if (10'h168 == _T_19[9:0]) begin
        image_1_360 <= io_pixelVal_in_1_1;
      end else if (10'h168 == _T_15[9:0]) begin
        image_1_360 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_361 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h169 == _T_37[9:0]) begin
        image_1_361 <= io_pixelVal_in_1_7;
      end else if (10'h169 == _T_34[9:0]) begin
        image_1_361 <= io_pixelVal_in_1_6;
      end else if (10'h169 == _T_31[9:0]) begin
        image_1_361 <= io_pixelVal_in_1_5;
      end else if (10'h169 == _T_28[9:0]) begin
        image_1_361 <= io_pixelVal_in_1_4;
      end else if (10'h169 == _T_25[9:0]) begin
        image_1_361 <= io_pixelVal_in_1_3;
      end else if (10'h169 == _T_22[9:0]) begin
        image_1_361 <= io_pixelVal_in_1_2;
      end else if (10'h169 == _T_19[9:0]) begin
        image_1_361 <= io_pixelVal_in_1_1;
      end else if (10'h169 == _T_15[9:0]) begin
        image_1_361 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_362 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h16a == _T_37[9:0]) begin
        image_1_362 <= io_pixelVal_in_1_7;
      end else if (10'h16a == _T_34[9:0]) begin
        image_1_362 <= io_pixelVal_in_1_6;
      end else if (10'h16a == _T_31[9:0]) begin
        image_1_362 <= io_pixelVal_in_1_5;
      end else if (10'h16a == _T_28[9:0]) begin
        image_1_362 <= io_pixelVal_in_1_4;
      end else if (10'h16a == _T_25[9:0]) begin
        image_1_362 <= io_pixelVal_in_1_3;
      end else if (10'h16a == _T_22[9:0]) begin
        image_1_362 <= io_pixelVal_in_1_2;
      end else if (10'h16a == _T_19[9:0]) begin
        image_1_362 <= io_pixelVal_in_1_1;
      end else if (10'h16a == _T_15[9:0]) begin
        image_1_362 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_363 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h16b == _T_37[9:0]) begin
        image_1_363 <= io_pixelVal_in_1_7;
      end else if (10'h16b == _T_34[9:0]) begin
        image_1_363 <= io_pixelVal_in_1_6;
      end else if (10'h16b == _T_31[9:0]) begin
        image_1_363 <= io_pixelVal_in_1_5;
      end else if (10'h16b == _T_28[9:0]) begin
        image_1_363 <= io_pixelVal_in_1_4;
      end else if (10'h16b == _T_25[9:0]) begin
        image_1_363 <= io_pixelVal_in_1_3;
      end else if (10'h16b == _T_22[9:0]) begin
        image_1_363 <= io_pixelVal_in_1_2;
      end else if (10'h16b == _T_19[9:0]) begin
        image_1_363 <= io_pixelVal_in_1_1;
      end else if (10'h16b == _T_15[9:0]) begin
        image_1_363 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_364 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h16c == _T_37[9:0]) begin
        image_1_364 <= io_pixelVal_in_1_7;
      end else if (10'h16c == _T_34[9:0]) begin
        image_1_364 <= io_pixelVal_in_1_6;
      end else if (10'h16c == _T_31[9:0]) begin
        image_1_364 <= io_pixelVal_in_1_5;
      end else if (10'h16c == _T_28[9:0]) begin
        image_1_364 <= io_pixelVal_in_1_4;
      end else if (10'h16c == _T_25[9:0]) begin
        image_1_364 <= io_pixelVal_in_1_3;
      end else if (10'h16c == _T_22[9:0]) begin
        image_1_364 <= io_pixelVal_in_1_2;
      end else if (10'h16c == _T_19[9:0]) begin
        image_1_364 <= io_pixelVal_in_1_1;
      end else if (10'h16c == _T_15[9:0]) begin
        image_1_364 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_365 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h16d == _T_37[9:0]) begin
        image_1_365 <= io_pixelVal_in_1_7;
      end else if (10'h16d == _T_34[9:0]) begin
        image_1_365 <= io_pixelVal_in_1_6;
      end else if (10'h16d == _T_31[9:0]) begin
        image_1_365 <= io_pixelVal_in_1_5;
      end else if (10'h16d == _T_28[9:0]) begin
        image_1_365 <= io_pixelVal_in_1_4;
      end else if (10'h16d == _T_25[9:0]) begin
        image_1_365 <= io_pixelVal_in_1_3;
      end else if (10'h16d == _T_22[9:0]) begin
        image_1_365 <= io_pixelVal_in_1_2;
      end else if (10'h16d == _T_19[9:0]) begin
        image_1_365 <= io_pixelVal_in_1_1;
      end else if (10'h16d == _T_15[9:0]) begin
        image_1_365 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_366 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h16e == _T_37[9:0]) begin
        image_1_366 <= io_pixelVal_in_1_7;
      end else if (10'h16e == _T_34[9:0]) begin
        image_1_366 <= io_pixelVal_in_1_6;
      end else if (10'h16e == _T_31[9:0]) begin
        image_1_366 <= io_pixelVal_in_1_5;
      end else if (10'h16e == _T_28[9:0]) begin
        image_1_366 <= io_pixelVal_in_1_4;
      end else if (10'h16e == _T_25[9:0]) begin
        image_1_366 <= io_pixelVal_in_1_3;
      end else if (10'h16e == _T_22[9:0]) begin
        image_1_366 <= io_pixelVal_in_1_2;
      end else if (10'h16e == _T_19[9:0]) begin
        image_1_366 <= io_pixelVal_in_1_1;
      end else if (10'h16e == _T_15[9:0]) begin
        image_1_366 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_367 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h16f == _T_37[9:0]) begin
        image_1_367 <= io_pixelVal_in_1_7;
      end else if (10'h16f == _T_34[9:0]) begin
        image_1_367 <= io_pixelVal_in_1_6;
      end else if (10'h16f == _T_31[9:0]) begin
        image_1_367 <= io_pixelVal_in_1_5;
      end else if (10'h16f == _T_28[9:0]) begin
        image_1_367 <= io_pixelVal_in_1_4;
      end else if (10'h16f == _T_25[9:0]) begin
        image_1_367 <= io_pixelVal_in_1_3;
      end else if (10'h16f == _T_22[9:0]) begin
        image_1_367 <= io_pixelVal_in_1_2;
      end else if (10'h16f == _T_19[9:0]) begin
        image_1_367 <= io_pixelVal_in_1_1;
      end else if (10'h16f == _T_15[9:0]) begin
        image_1_367 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_368 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h170 == _T_37[9:0]) begin
        image_1_368 <= io_pixelVal_in_1_7;
      end else if (10'h170 == _T_34[9:0]) begin
        image_1_368 <= io_pixelVal_in_1_6;
      end else if (10'h170 == _T_31[9:0]) begin
        image_1_368 <= io_pixelVal_in_1_5;
      end else if (10'h170 == _T_28[9:0]) begin
        image_1_368 <= io_pixelVal_in_1_4;
      end else if (10'h170 == _T_25[9:0]) begin
        image_1_368 <= io_pixelVal_in_1_3;
      end else if (10'h170 == _T_22[9:0]) begin
        image_1_368 <= io_pixelVal_in_1_2;
      end else if (10'h170 == _T_19[9:0]) begin
        image_1_368 <= io_pixelVal_in_1_1;
      end else if (10'h170 == _T_15[9:0]) begin
        image_1_368 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_369 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h171 == _T_37[9:0]) begin
        image_1_369 <= io_pixelVal_in_1_7;
      end else if (10'h171 == _T_34[9:0]) begin
        image_1_369 <= io_pixelVal_in_1_6;
      end else if (10'h171 == _T_31[9:0]) begin
        image_1_369 <= io_pixelVal_in_1_5;
      end else if (10'h171 == _T_28[9:0]) begin
        image_1_369 <= io_pixelVal_in_1_4;
      end else if (10'h171 == _T_25[9:0]) begin
        image_1_369 <= io_pixelVal_in_1_3;
      end else if (10'h171 == _T_22[9:0]) begin
        image_1_369 <= io_pixelVal_in_1_2;
      end else if (10'h171 == _T_19[9:0]) begin
        image_1_369 <= io_pixelVal_in_1_1;
      end else if (10'h171 == _T_15[9:0]) begin
        image_1_369 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_370 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h172 == _T_37[9:0]) begin
        image_1_370 <= io_pixelVal_in_1_7;
      end else if (10'h172 == _T_34[9:0]) begin
        image_1_370 <= io_pixelVal_in_1_6;
      end else if (10'h172 == _T_31[9:0]) begin
        image_1_370 <= io_pixelVal_in_1_5;
      end else if (10'h172 == _T_28[9:0]) begin
        image_1_370 <= io_pixelVal_in_1_4;
      end else if (10'h172 == _T_25[9:0]) begin
        image_1_370 <= io_pixelVal_in_1_3;
      end else if (10'h172 == _T_22[9:0]) begin
        image_1_370 <= io_pixelVal_in_1_2;
      end else if (10'h172 == _T_19[9:0]) begin
        image_1_370 <= io_pixelVal_in_1_1;
      end else if (10'h172 == _T_15[9:0]) begin
        image_1_370 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_371 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h173 == _T_37[9:0]) begin
        image_1_371 <= io_pixelVal_in_1_7;
      end else if (10'h173 == _T_34[9:0]) begin
        image_1_371 <= io_pixelVal_in_1_6;
      end else if (10'h173 == _T_31[9:0]) begin
        image_1_371 <= io_pixelVal_in_1_5;
      end else if (10'h173 == _T_28[9:0]) begin
        image_1_371 <= io_pixelVal_in_1_4;
      end else if (10'h173 == _T_25[9:0]) begin
        image_1_371 <= io_pixelVal_in_1_3;
      end else if (10'h173 == _T_22[9:0]) begin
        image_1_371 <= io_pixelVal_in_1_2;
      end else if (10'h173 == _T_19[9:0]) begin
        image_1_371 <= io_pixelVal_in_1_1;
      end else if (10'h173 == _T_15[9:0]) begin
        image_1_371 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_372 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h174 == _T_37[9:0]) begin
        image_1_372 <= io_pixelVal_in_1_7;
      end else if (10'h174 == _T_34[9:0]) begin
        image_1_372 <= io_pixelVal_in_1_6;
      end else if (10'h174 == _T_31[9:0]) begin
        image_1_372 <= io_pixelVal_in_1_5;
      end else if (10'h174 == _T_28[9:0]) begin
        image_1_372 <= io_pixelVal_in_1_4;
      end else if (10'h174 == _T_25[9:0]) begin
        image_1_372 <= io_pixelVal_in_1_3;
      end else if (10'h174 == _T_22[9:0]) begin
        image_1_372 <= io_pixelVal_in_1_2;
      end else if (10'h174 == _T_19[9:0]) begin
        image_1_372 <= io_pixelVal_in_1_1;
      end else if (10'h174 == _T_15[9:0]) begin
        image_1_372 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_373 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h175 == _T_37[9:0]) begin
        image_1_373 <= io_pixelVal_in_1_7;
      end else if (10'h175 == _T_34[9:0]) begin
        image_1_373 <= io_pixelVal_in_1_6;
      end else if (10'h175 == _T_31[9:0]) begin
        image_1_373 <= io_pixelVal_in_1_5;
      end else if (10'h175 == _T_28[9:0]) begin
        image_1_373 <= io_pixelVal_in_1_4;
      end else if (10'h175 == _T_25[9:0]) begin
        image_1_373 <= io_pixelVal_in_1_3;
      end else if (10'h175 == _T_22[9:0]) begin
        image_1_373 <= io_pixelVal_in_1_2;
      end else if (10'h175 == _T_19[9:0]) begin
        image_1_373 <= io_pixelVal_in_1_1;
      end else if (10'h175 == _T_15[9:0]) begin
        image_1_373 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_374 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h176 == _T_37[9:0]) begin
        image_1_374 <= io_pixelVal_in_1_7;
      end else if (10'h176 == _T_34[9:0]) begin
        image_1_374 <= io_pixelVal_in_1_6;
      end else if (10'h176 == _T_31[9:0]) begin
        image_1_374 <= io_pixelVal_in_1_5;
      end else if (10'h176 == _T_28[9:0]) begin
        image_1_374 <= io_pixelVal_in_1_4;
      end else if (10'h176 == _T_25[9:0]) begin
        image_1_374 <= io_pixelVal_in_1_3;
      end else if (10'h176 == _T_22[9:0]) begin
        image_1_374 <= io_pixelVal_in_1_2;
      end else if (10'h176 == _T_19[9:0]) begin
        image_1_374 <= io_pixelVal_in_1_1;
      end else if (10'h176 == _T_15[9:0]) begin
        image_1_374 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_375 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h177 == _T_37[9:0]) begin
        image_1_375 <= io_pixelVal_in_1_7;
      end else if (10'h177 == _T_34[9:0]) begin
        image_1_375 <= io_pixelVal_in_1_6;
      end else if (10'h177 == _T_31[9:0]) begin
        image_1_375 <= io_pixelVal_in_1_5;
      end else if (10'h177 == _T_28[9:0]) begin
        image_1_375 <= io_pixelVal_in_1_4;
      end else if (10'h177 == _T_25[9:0]) begin
        image_1_375 <= io_pixelVal_in_1_3;
      end else if (10'h177 == _T_22[9:0]) begin
        image_1_375 <= io_pixelVal_in_1_2;
      end else if (10'h177 == _T_19[9:0]) begin
        image_1_375 <= io_pixelVal_in_1_1;
      end else if (10'h177 == _T_15[9:0]) begin
        image_1_375 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_376 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h178 == _T_37[9:0]) begin
        image_1_376 <= io_pixelVal_in_1_7;
      end else if (10'h178 == _T_34[9:0]) begin
        image_1_376 <= io_pixelVal_in_1_6;
      end else if (10'h178 == _T_31[9:0]) begin
        image_1_376 <= io_pixelVal_in_1_5;
      end else if (10'h178 == _T_28[9:0]) begin
        image_1_376 <= io_pixelVal_in_1_4;
      end else if (10'h178 == _T_25[9:0]) begin
        image_1_376 <= io_pixelVal_in_1_3;
      end else if (10'h178 == _T_22[9:0]) begin
        image_1_376 <= io_pixelVal_in_1_2;
      end else if (10'h178 == _T_19[9:0]) begin
        image_1_376 <= io_pixelVal_in_1_1;
      end else if (10'h178 == _T_15[9:0]) begin
        image_1_376 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_377 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h179 == _T_37[9:0]) begin
        image_1_377 <= io_pixelVal_in_1_7;
      end else if (10'h179 == _T_34[9:0]) begin
        image_1_377 <= io_pixelVal_in_1_6;
      end else if (10'h179 == _T_31[9:0]) begin
        image_1_377 <= io_pixelVal_in_1_5;
      end else if (10'h179 == _T_28[9:0]) begin
        image_1_377 <= io_pixelVal_in_1_4;
      end else if (10'h179 == _T_25[9:0]) begin
        image_1_377 <= io_pixelVal_in_1_3;
      end else if (10'h179 == _T_22[9:0]) begin
        image_1_377 <= io_pixelVal_in_1_2;
      end else if (10'h179 == _T_19[9:0]) begin
        image_1_377 <= io_pixelVal_in_1_1;
      end else if (10'h179 == _T_15[9:0]) begin
        image_1_377 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_378 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h17a == _T_37[9:0]) begin
        image_1_378 <= io_pixelVal_in_1_7;
      end else if (10'h17a == _T_34[9:0]) begin
        image_1_378 <= io_pixelVal_in_1_6;
      end else if (10'h17a == _T_31[9:0]) begin
        image_1_378 <= io_pixelVal_in_1_5;
      end else if (10'h17a == _T_28[9:0]) begin
        image_1_378 <= io_pixelVal_in_1_4;
      end else if (10'h17a == _T_25[9:0]) begin
        image_1_378 <= io_pixelVal_in_1_3;
      end else if (10'h17a == _T_22[9:0]) begin
        image_1_378 <= io_pixelVal_in_1_2;
      end else if (10'h17a == _T_19[9:0]) begin
        image_1_378 <= io_pixelVal_in_1_1;
      end else if (10'h17a == _T_15[9:0]) begin
        image_1_378 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_379 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h17b == _T_37[9:0]) begin
        image_1_379 <= io_pixelVal_in_1_7;
      end else if (10'h17b == _T_34[9:0]) begin
        image_1_379 <= io_pixelVal_in_1_6;
      end else if (10'h17b == _T_31[9:0]) begin
        image_1_379 <= io_pixelVal_in_1_5;
      end else if (10'h17b == _T_28[9:0]) begin
        image_1_379 <= io_pixelVal_in_1_4;
      end else if (10'h17b == _T_25[9:0]) begin
        image_1_379 <= io_pixelVal_in_1_3;
      end else if (10'h17b == _T_22[9:0]) begin
        image_1_379 <= io_pixelVal_in_1_2;
      end else if (10'h17b == _T_19[9:0]) begin
        image_1_379 <= io_pixelVal_in_1_1;
      end else if (10'h17b == _T_15[9:0]) begin
        image_1_379 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_380 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h17c == _T_37[9:0]) begin
        image_1_380 <= io_pixelVal_in_1_7;
      end else if (10'h17c == _T_34[9:0]) begin
        image_1_380 <= io_pixelVal_in_1_6;
      end else if (10'h17c == _T_31[9:0]) begin
        image_1_380 <= io_pixelVal_in_1_5;
      end else if (10'h17c == _T_28[9:0]) begin
        image_1_380 <= io_pixelVal_in_1_4;
      end else if (10'h17c == _T_25[9:0]) begin
        image_1_380 <= io_pixelVal_in_1_3;
      end else if (10'h17c == _T_22[9:0]) begin
        image_1_380 <= io_pixelVal_in_1_2;
      end else if (10'h17c == _T_19[9:0]) begin
        image_1_380 <= io_pixelVal_in_1_1;
      end else if (10'h17c == _T_15[9:0]) begin
        image_1_380 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_381 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h17d == _T_37[9:0]) begin
        image_1_381 <= io_pixelVal_in_1_7;
      end else if (10'h17d == _T_34[9:0]) begin
        image_1_381 <= io_pixelVal_in_1_6;
      end else if (10'h17d == _T_31[9:0]) begin
        image_1_381 <= io_pixelVal_in_1_5;
      end else if (10'h17d == _T_28[9:0]) begin
        image_1_381 <= io_pixelVal_in_1_4;
      end else if (10'h17d == _T_25[9:0]) begin
        image_1_381 <= io_pixelVal_in_1_3;
      end else if (10'h17d == _T_22[9:0]) begin
        image_1_381 <= io_pixelVal_in_1_2;
      end else if (10'h17d == _T_19[9:0]) begin
        image_1_381 <= io_pixelVal_in_1_1;
      end else if (10'h17d == _T_15[9:0]) begin
        image_1_381 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_382 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h17e == _T_37[9:0]) begin
        image_1_382 <= io_pixelVal_in_1_7;
      end else if (10'h17e == _T_34[9:0]) begin
        image_1_382 <= io_pixelVal_in_1_6;
      end else if (10'h17e == _T_31[9:0]) begin
        image_1_382 <= io_pixelVal_in_1_5;
      end else if (10'h17e == _T_28[9:0]) begin
        image_1_382 <= io_pixelVal_in_1_4;
      end else if (10'h17e == _T_25[9:0]) begin
        image_1_382 <= io_pixelVal_in_1_3;
      end else if (10'h17e == _T_22[9:0]) begin
        image_1_382 <= io_pixelVal_in_1_2;
      end else if (10'h17e == _T_19[9:0]) begin
        image_1_382 <= io_pixelVal_in_1_1;
      end else if (10'h17e == _T_15[9:0]) begin
        image_1_382 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_383 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h17f == _T_37[9:0]) begin
        image_1_383 <= io_pixelVal_in_1_7;
      end else if (10'h17f == _T_34[9:0]) begin
        image_1_383 <= io_pixelVal_in_1_6;
      end else if (10'h17f == _T_31[9:0]) begin
        image_1_383 <= io_pixelVal_in_1_5;
      end else if (10'h17f == _T_28[9:0]) begin
        image_1_383 <= io_pixelVal_in_1_4;
      end else if (10'h17f == _T_25[9:0]) begin
        image_1_383 <= io_pixelVal_in_1_3;
      end else if (10'h17f == _T_22[9:0]) begin
        image_1_383 <= io_pixelVal_in_1_2;
      end else if (10'h17f == _T_19[9:0]) begin
        image_1_383 <= io_pixelVal_in_1_1;
      end else if (10'h17f == _T_15[9:0]) begin
        image_1_383 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_384 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h180 == _T_37[9:0]) begin
        image_1_384 <= io_pixelVal_in_1_7;
      end else if (10'h180 == _T_34[9:0]) begin
        image_1_384 <= io_pixelVal_in_1_6;
      end else if (10'h180 == _T_31[9:0]) begin
        image_1_384 <= io_pixelVal_in_1_5;
      end else if (10'h180 == _T_28[9:0]) begin
        image_1_384 <= io_pixelVal_in_1_4;
      end else if (10'h180 == _T_25[9:0]) begin
        image_1_384 <= io_pixelVal_in_1_3;
      end else if (10'h180 == _T_22[9:0]) begin
        image_1_384 <= io_pixelVal_in_1_2;
      end else if (10'h180 == _T_19[9:0]) begin
        image_1_384 <= io_pixelVal_in_1_1;
      end else if (10'h180 == _T_15[9:0]) begin
        image_1_384 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_385 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h181 == _T_37[9:0]) begin
        image_1_385 <= io_pixelVal_in_1_7;
      end else if (10'h181 == _T_34[9:0]) begin
        image_1_385 <= io_pixelVal_in_1_6;
      end else if (10'h181 == _T_31[9:0]) begin
        image_1_385 <= io_pixelVal_in_1_5;
      end else if (10'h181 == _T_28[9:0]) begin
        image_1_385 <= io_pixelVal_in_1_4;
      end else if (10'h181 == _T_25[9:0]) begin
        image_1_385 <= io_pixelVal_in_1_3;
      end else if (10'h181 == _T_22[9:0]) begin
        image_1_385 <= io_pixelVal_in_1_2;
      end else if (10'h181 == _T_19[9:0]) begin
        image_1_385 <= io_pixelVal_in_1_1;
      end else if (10'h181 == _T_15[9:0]) begin
        image_1_385 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_386 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h182 == _T_37[9:0]) begin
        image_1_386 <= io_pixelVal_in_1_7;
      end else if (10'h182 == _T_34[9:0]) begin
        image_1_386 <= io_pixelVal_in_1_6;
      end else if (10'h182 == _T_31[9:0]) begin
        image_1_386 <= io_pixelVal_in_1_5;
      end else if (10'h182 == _T_28[9:0]) begin
        image_1_386 <= io_pixelVal_in_1_4;
      end else if (10'h182 == _T_25[9:0]) begin
        image_1_386 <= io_pixelVal_in_1_3;
      end else if (10'h182 == _T_22[9:0]) begin
        image_1_386 <= io_pixelVal_in_1_2;
      end else if (10'h182 == _T_19[9:0]) begin
        image_1_386 <= io_pixelVal_in_1_1;
      end else if (10'h182 == _T_15[9:0]) begin
        image_1_386 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_387 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h183 == _T_37[9:0]) begin
        image_1_387 <= io_pixelVal_in_1_7;
      end else if (10'h183 == _T_34[9:0]) begin
        image_1_387 <= io_pixelVal_in_1_6;
      end else if (10'h183 == _T_31[9:0]) begin
        image_1_387 <= io_pixelVal_in_1_5;
      end else if (10'h183 == _T_28[9:0]) begin
        image_1_387 <= io_pixelVal_in_1_4;
      end else if (10'h183 == _T_25[9:0]) begin
        image_1_387 <= io_pixelVal_in_1_3;
      end else if (10'h183 == _T_22[9:0]) begin
        image_1_387 <= io_pixelVal_in_1_2;
      end else if (10'h183 == _T_19[9:0]) begin
        image_1_387 <= io_pixelVal_in_1_1;
      end else if (10'h183 == _T_15[9:0]) begin
        image_1_387 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_388 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h184 == _T_37[9:0]) begin
        image_1_388 <= io_pixelVal_in_1_7;
      end else if (10'h184 == _T_34[9:0]) begin
        image_1_388 <= io_pixelVal_in_1_6;
      end else if (10'h184 == _T_31[9:0]) begin
        image_1_388 <= io_pixelVal_in_1_5;
      end else if (10'h184 == _T_28[9:0]) begin
        image_1_388 <= io_pixelVal_in_1_4;
      end else if (10'h184 == _T_25[9:0]) begin
        image_1_388 <= io_pixelVal_in_1_3;
      end else if (10'h184 == _T_22[9:0]) begin
        image_1_388 <= io_pixelVal_in_1_2;
      end else if (10'h184 == _T_19[9:0]) begin
        image_1_388 <= io_pixelVal_in_1_1;
      end else if (10'h184 == _T_15[9:0]) begin
        image_1_388 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_389 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h185 == _T_37[9:0]) begin
        image_1_389 <= io_pixelVal_in_1_7;
      end else if (10'h185 == _T_34[9:0]) begin
        image_1_389 <= io_pixelVal_in_1_6;
      end else if (10'h185 == _T_31[9:0]) begin
        image_1_389 <= io_pixelVal_in_1_5;
      end else if (10'h185 == _T_28[9:0]) begin
        image_1_389 <= io_pixelVal_in_1_4;
      end else if (10'h185 == _T_25[9:0]) begin
        image_1_389 <= io_pixelVal_in_1_3;
      end else if (10'h185 == _T_22[9:0]) begin
        image_1_389 <= io_pixelVal_in_1_2;
      end else if (10'h185 == _T_19[9:0]) begin
        image_1_389 <= io_pixelVal_in_1_1;
      end else if (10'h185 == _T_15[9:0]) begin
        image_1_389 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_390 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h186 == _T_37[9:0]) begin
        image_1_390 <= io_pixelVal_in_1_7;
      end else if (10'h186 == _T_34[9:0]) begin
        image_1_390 <= io_pixelVal_in_1_6;
      end else if (10'h186 == _T_31[9:0]) begin
        image_1_390 <= io_pixelVal_in_1_5;
      end else if (10'h186 == _T_28[9:0]) begin
        image_1_390 <= io_pixelVal_in_1_4;
      end else if (10'h186 == _T_25[9:0]) begin
        image_1_390 <= io_pixelVal_in_1_3;
      end else if (10'h186 == _T_22[9:0]) begin
        image_1_390 <= io_pixelVal_in_1_2;
      end else if (10'h186 == _T_19[9:0]) begin
        image_1_390 <= io_pixelVal_in_1_1;
      end else if (10'h186 == _T_15[9:0]) begin
        image_1_390 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_391 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h187 == _T_37[9:0]) begin
        image_1_391 <= io_pixelVal_in_1_7;
      end else if (10'h187 == _T_34[9:0]) begin
        image_1_391 <= io_pixelVal_in_1_6;
      end else if (10'h187 == _T_31[9:0]) begin
        image_1_391 <= io_pixelVal_in_1_5;
      end else if (10'h187 == _T_28[9:0]) begin
        image_1_391 <= io_pixelVal_in_1_4;
      end else if (10'h187 == _T_25[9:0]) begin
        image_1_391 <= io_pixelVal_in_1_3;
      end else if (10'h187 == _T_22[9:0]) begin
        image_1_391 <= io_pixelVal_in_1_2;
      end else if (10'h187 == _T_19[9:0]) begin
        image_1_391 <= io_pixelVal_in_1_1;
      end else if (10'h187 == _T_15[9:0]) begin
        image_1_391 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_392 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h188 == _T_37[9:0]) begin
        image_1_392 <= io_pixelVal_in_1_7;
      end else if (10'h188 == _T_34[9:0]) begin
        image_1_392 <= io_pixelVal_in_1_6;
      end else if (10'h188 == _T_31[9:0]) begin
        image_1_392 <= io_pixelVal_in_1_5;
      end else if (10'h188 == _T_28[9:0]) begin
        image_1_392 <= io_pixelVal_in_1_4;
      end else if (10'h188 == _T_25[9:0]) begin
        image_1_392 <= io_pixelVal_in_1_3;
      end else if (10'h188 == _T_22[9:0]) begin
        image_1_392 <= io_pixelVal_in_1_2;
      end else if (10'h188 == _T_19[9:0]) begin
        image_1_392 <= io_pixelVal_in_1_1;
      end else if (10'h188 == _T_15[9:0]) begin
        image_1_392 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_393 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h189 == _T_37[9:0]) begin
        image_1_393 <= io_pixelVal_in_1_7;
      end else if (10'h189 == _T_34[9:0]) begin
        image_1_393 <= io_pixelVal_in_1_6;
      end else if (10'h189 == _T_31[9:0]) begin
        image_1_393 <= io_pixelVal_in_1_5;
      end else if (10'h189 == _T_28[9:0]) begin
        image_1_393 <= io_pixelVal_in_1_4;
      end else if (10'h189 == _T_25[9:0]) begin
        image_1_393 <= io_pixelVal_in_1_3;
      end else if (10'h189 == _T_22[9:0]) begin
        image_1_393 <= io_pixelVal_in_1_2;
      end else if (10'h189 == _T_19[9:0]) begin
        image_1_393 <= io_pixelVal_in_1_1;
      end else if (10'h189 == _T_15[9:0]) begin
        image_1_393 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_394 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h18a == _T_37[9:0]) begin
        image_1_394 <= io_pixelVal_in_1_7;
      end else if (10'h18a == _T_34[9:0]) begin
        image_1_394 <= io_pixelVal_in_1_6;
      end else if (10'h18a == _T_31[9:0]) begin
        image_1_394 <= io_pixelVal_in_1_5;
      end else if (10'h18a == _T_28[9:0]) begin
        image_1_394 <= io_pixelVal_in_1_4;
      end else if (10'h18a == _T_25[9:0]) begin
        image_1_394 <= io_pixelVal_in_1_3;
      end else if (10'h18a == _T_22[9:0]) begin
        image_1_394 <= io_pixelVal_in_1_2;
      end else if (10'h18a == _T_19[9:0]) begin
        image_1_394 <= io_pixelVal_in_1_1;
      end else if (10'h18a == _T_15[9:0]) begin
        image_1_394 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_395 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h18b == _T_37[9:0]) begin
        image_1_395 <= io_pixelVal_in_1_7;
      end else if (10'h18b == _T_34[9:0]) begin
        image_1_395 <= io_pixelVal_in_1_6;
      end else if (10'h18b == _T_31[9:0]) begin
        image_1_395 <= io_pixelVal_in_1_5;
      end else if (10'h18b == _T_28[9:0]) begin
        image_1_395 <= io_pixelVal_in_1_4;
      end else if (10'h18b == _T_25[9:0]) begin
        image_1_395 <= io_pixelVal_in_1_3;
      end else if (10'h18b == _T_22[9:0]) begin
        image_1_395 <= io_pixelVal_in_1_2;
      end else if (10'h18b == _T_19[9:0]) begin
        image_1_395 <= io_pixelVal_in_1_1;
      end else if (10'h18b == _T_15[9:0]) begin
        image_1_395 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_396 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h18c == _T_37[9:0]) begin
        image_1_396 <= io_pixelVal_in_1_7;
      end else if (10'h18c == _T_34[9:0]) begin
        image_1_396 <= io_pixelVal_in_1_6;
      end else if (10'h18c == _T_31[9:0]) begin
        image_1_396 <= io_pixelVal_in_1_5;
      end else if (10'h18c == _T_28[9:0]) begin
        image_1_396 <= io_pixelVal_in_1_4;
      end else if (10'h18c == _T_25[9:0]) begin
        image_1_396 <= io_pixelVal_in_1_3;
      end else if (10'h18c == _T_22[9:0]) begin
        image_1_396 <= io_pixelVal_in_1_2;
      end else if (10'h18c == _T_19[9:0]) begin
        image_1_396 <= io_pixelVal_in_1_1;
      end else if (10'h18c == _T_15[9:0]) begin
        image_1_396 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_397 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h18d == _T_37[9:0]) begin
        image_1_397 <= io_pixelVal_in_1_7;
      end else if (10'h18d == _T_34[9:0]) begin
        image_1_397 <= io_pixelVal_in_1_6;
      end else if (10'h18d == _T_31[9:0]) begin
        image_1_397 <= io_pixelVal_in_1_5;
      end else if (10'h18d == _T_28[9:0]) begin
        image_1_397 <= io_pixelVal_in_1_4;
      end else if (10'h18d == _T_25[9:0]) begin
        image_1_397 <= io_pixelVal_in_1_3;
      end else if (10'h18d == _T_22[9:0]) begin
        image_1_397 <= io_pixelVal_in_1_2;
      end else if (10'h18d == _T_19[9:0]) begin
        image_1_397 <= io_pixelVal_in_1_1;
      end else if (10'h18d == _T_15[9:0]) begin
        image_1_397 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_398 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h18e == _T_37[9:0]) begin
        image_1_398 <= io_pixelVal_in_1_7;
      end else if (10'h18e == _T_34[9:0]) begin
        image_1_398 <= io_pixelVal_in_1_6;
      end else if (10'h18e == _T_31[9:0]) begin
        image_1_398 <= io_pixelVal_in_1_5;
      end else if (10'h18e == _T_28[9:0]) begin
        image_1_398 <= io_pixelVal_in_1_4;
      end else if (10'h18e == _T_25[9:0]) begin
        image_1_398 <= io_pixelVal_in_1_3;
      end else if (10'h18e == _T_22[9:0]) begin
        image_1_398 <= io_pixelVal_in_1_2;
      end else if (10'h18e == _T_19[9:0]) begin
        image_1_398 <= io_pixelVal_in_1_1;
      end else if (10'h18e == _T_15[9:0]) begin
        image_1_398 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_399 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h18f == _T_37[9:0]) begin
        image_1_399 <= io_pixelVal_in_1_7;
      end else if (10'h18f == _T_34[9:0]) begin
        image_1_399 <= io_pixelVal_in_1_6;
      end else if (10'h18f == _T_31[9:0]) begin
        image_1_399 <= io_pixelVal_in_1_5;
      end else if (10'h18f == _T_28[9:0]) begin
        image_1_399 <= io_pixelVal_in_1_4;
      end else if (10'h18f == _T_25[9:0]) begin
        image_1_399 <= io_pixelVal_in_1_3;
      end else if (10'h18f == _T_22[9:0]) begin
        image_1_399 <= io_pixelVal_in_1_2;
      end else if (10'h18f == _T_19[9:0]) begin
        image_1_399 <= io_pixelVal_in_1_1;
      end else if (10'h18f == _T_15[9:0]) begin
        image_1_399 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_400 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h190 == _T_37[9:0]) begin
        image_1_400 <= io_pixelVal_in_1_7;
      end else if (10'h190 == _T_34[9:0]) begin
        image_1_400 <= io_pixelVal_in_1_6;
      end else if (10'h190 == _T_31[9:0]) begin
        image_1_400 <= io_pixelVal_in_1_5;
      end else if (10'h190 == _T_28[9:0]) begin
        image_1_400 <= io_pixelVal_in_1_4;
      end else if (10'h190 == _T_25[9:0]) begin
        image_1_400 <= io_pixelVal_in_1_3;
      end else if (10'h190 == _T_22[9:0]) begin
        image_1_400 <= io_pixelVal_in_1_2;
      end else if (10'h190 == _T_19[9:0]) begin
        image_1_400 <= io_pixelVal_in_1_1;
      end else if (10'h190 == _T_15[9:0]) begin
        image_1_400 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_401 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h191 == _T_37[9:0]) begin
        image_1_401 <= io_pixelVal_in_1_7;
      end else if (10'h191 == _T_34[9:0]) begin
        image_1_401 <= io_pixelVal_in_1_6;
      end else if (10'h191 == _T_31[9:0]) begin
        image_1_401 <= io_pixelVal_in_1_5;
      end else if (10'h191 == _T_28[9:0]) begin
        image_1_401 <= io_pixelVal_in_1_4;
      end else if (10'h191 == _T_25[9:0]) begin
        image_1_401 <= io_pixelVal_in_1_3;
      end else if (10'h191 == _T_22[9:0]) begin
        image_1_401 <= io_pixelVal_in_1_2;
      end else if (10'h191 == _T_19[9:0]) begin
        image_1_401 <= io_pixelVal_in_1_1;
      end else if (10'h191 == _T_15[9:0]) begin
        image_1_401 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_402 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h192 == _T_37[9:0]) begin
        image_1_402 <= io_pixelVal_in_1_7;
      end else if (10'h192 == _T_34[9:0]) begin
        image_1_402 <= io_pixelVal_in_1_6;
      end else if (10'h192 == _T_31[9:0]) begin
        image_1_402 <= io_pixelVal_in_1_5;
      end else if (10'h192 == _T_28[9:0]) begin
        image_1_402 <= io_pixelVal_in_1_4;
      end else if (10'h192 == _T_25[9:0]) begin
        image_1_402 <= io_pixelVal_in_1_3;
      end else if (10'h192 == _T_22[9:0]) begin
        image_1_402 <= io_pixelVal_in_1_2;
      end else if (10'h192 == _T_19[9:0]) begin
        image_1_402 <= io_pixelVal_in_1_1;
      end else if (10'h192 == _T_15[9:0]) begin
        image_1_402 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_403 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h193 == _T_37[9:0]) begin
        image_1_403 <= io_pixelVal_in_1_7;
      end else if (10'h193 == _T_34[9:0]) begin
        image_1_403 <= io_pixelVal_in_1_6;
      end else if (10'h193 == _T_31[9:0]) begin
        image_1_403 <= io_pixelVal_in_1_5;
      end else if (10'h193 == _T_28[9:0]) begin
        image_1_403 <= io_pixelVal_in_1_4;
      end else if (10'h193 == _T_25[9:0]) begin
        image_1_403 <= io_pixelVal_in_1_3;
      end else if (10'h193 == _T_22[9:0]) begin
        image_1_403 <= io_pixelVal_in_1_2;
      end else if (10'h193 == _T_19[9:0]) begin
        image_1_403 <= io_pixelVal_in_1_1;
      end else if (10'h193 == _T_15[9:0]) begin
        image_1_403 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_404 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h194 == _T_37[9:0]) begin
        image_1_404 <= io_pixelVal_in_1_7;
      end else if (10'h194 == _T_34[9:0]) begin
        image_1_404 <= io_pixelVal_in_1_6;
      end else if (10'h194 == _T_31[9:0]) begin
        image_1_404 <= io_pixelVal_in_1_5;
      end else if (10'h194 == _T_28[9:0]) begin
        image_1_404 <= io_pixelVal_in_1_4;
      end else if (10'h194 == _T_25[9:0]) begin
        image_1_404 <= io_pixelVal_in_1_3;
      end else if (10'h194 == _T_22[9:0]) begin
        image_1_404 <= io_pixelVal_in_1_2;
      end else if (10'h194 == _T_19[9:0]) begin
        image_1_404 <= io_pixelVal_in_1_1;
      end else if (10'h194 == _T_15[9:0]) begin
        image_1_404 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_405 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h195 == _T_37[9:0]) begin
        image_1_405 <= io_pixelVal_in_1_7;
      end else if (10'h195 == _T_34[9:0]) begin
        image_1_405 <= io_pixelVal_in_1_6;
      end else if (10'h195 == _T_31[9:0]) begin
        image_1_405 <= io_pixelVal_in_1_5;
      end else if (10'h195 == _T_28[9:0]) begin
        image_1_405 <= io_pixelVal_in_1_4;
      end else if (10'h195 == _T_25[9:0]) begin
        image_1_405 <= io_pixelVal_in_1_3;
      end else if (10'h195 == _T_22[9:0]) begin
        image_1_405 <= io_pixelVal_in_1_2;
      end else if (10'h195 == _T_19[9:0]) begin
        image_1_405 <= io_pixelVal_in_1_1;
      end else if (10'h195 == _T_15[9:0]) begin
        image_1_405 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_406 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h196 == _T_37[9:0]) begin
        image_1_406 <= io_pixelVal_in_1_7;
      end else if (10'h196 == _T_34[9:0]) begin
        image_1_406 <= io_pixelVal_in_1_6;
      end else if (10'h196 == _T_31[9:0]) begin
        image_1_406 <= io_pixelVal_in_1_5;
      end else if (10'h196 == _T_28[9:0]) begin
        image_1_406 <= io_pixelVal_in_1_4;
      end else if (10'h196 == _T_25[9:0]) begin
        image_1_406 <= io_pixelVal_in_1_3;
      end else if (10'h196 == _T_22[9:0]) begin
        image_1_406 <= io_pixelVal_in_1_2;
      end else if (10'h196 == _T_19[9:0]) begin
        image_1_406 <= io_pixelVal_in_1_1;
      end else if (10'h196 == _T_15[9:0]) begin
        image_1_406 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_407 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h197 == _T_37[9:0]) begin
        image_1_407 <= io_pixelVal_in_1_7;
      end else if (10'h197 == _T_34[9:0]) begin
        image_1_407 <= io_pixelVal_in_1_6;
      end else if (10'h197 == _T_31[9:0]) begin
        image_1_407 <= io_pixelVal_in_1_5;
      end else if (10'h197 == _T_28[9:0]) begin
        image_1_407 <= io_pixelVal_in_1_4;
      end else if (10'h197 == _T_25[9:0]) begin
        image_1_407 <= io_pixelVal_in_1_3;
      end else if (10'h197 == _T_22[9:0]) begin
        image_1_407 <= io_pixelVal_in_1_2;
      end else if (10'h197 == _T_19[9:0]) begin
        image_1_407 <= io_pixelVal_in_1_1;
      end else if (10'h197 == _T_15[9:0]) begin
        image_1_407 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_408 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h198 == _T_37[9:0]) begin
        image_1_408 <= io_pixelVal_in_1_7;
      end else if (10'h198 == _T_34[9:0]) begin
        image_1_408 <= io_pixelVal_in_1_6;
      end else if (10'h198 == _T_31[9:0]) begin
        image_1_408 <= io_pixelVal_in_1_5;
      end else if (10'h198 == _T_28[9:0]) begin
        image_1_408 <= io_pixelVal_in_1_4;
      end else if (10'h198 == _T_25[9:0]) begin
        image_1_408 <= io_pixelVal_in_1_3;
      end else if (10'h198 == _T_22[9:0]) begin
        image_1_408 <= io_pixelVal_in_1_2;
      end else if (10'h198 == _T_19[9:0]) begin
        image_1_408 <= io_pixelVal_in_1_1;
      end else if (10'h198 == _T_15[9:0]) begin
        image_1_408 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_409 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h199 == _T_37[9:0]) begin
        image_1_409 <= io_pixelVal_in_1_7;
      end else if (10'h199 == _T_34[9:0]) begin
        image_1_409 <= io_pixelVal_in_1_6;
      end else if (10'h199 == _T_31[9:0]) begin
        image_1_409 <= io_pixelVal_in_1_5;
      end else if (10'h199 == _T_28[9:0]) begin
        image_1_409 <= io_pixelVal_in_1_4;
      end else if (10'h199 == _T_25[9:0]) begin
        image_1_409 <= io_pixelVal_in_1_3;
      end else if (10'h199 == _T_22[9:0]) begin
        image_1_409 <= io_pixelVal_in_1_2;
      end else if (10'h199 == _T_19[9:0]) begin
        image_1_409 <= io_pixelVal_in_1_1;
      end else if (10'h199 == _T_15[9:0]) begin
        image_1_409 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_410 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h19a == _T_37[9:0]) begin
        image_1_410 <= io_pixelVal_in_1_7;
      end else if (10'h19a == _T_34[9:0]) begin
        image_1_410 <= io_pixelVal_in_1_6;
      end else if (10'h19a == _T_31[9:0]) begin
        image_1_410 <= io_pixelVal_in_1_5;
      end else if (10'h19a == _T_28[9:0]) begin
        image_1_410 <= io_pixelVal_in_1_4;
      end else if (10'h19a == _T_25[9:0]) begin
        image_1_410 <= io_pixelVal_in_1_3;
      end else if (10'h19a == _T_22[9:0]) begin
        image_1_410 <= io_pixelVal_in_1_2;
      end else if (10'h19a == _T_19[9:0]) begin
        image_1_410 <= io_pixelVal_in_1_1;
      end else if (10'h19a == _T_15[9:0]) begin
        image_1_410 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_411 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h19b == _T_37[9:0]) begin
        image_1_411 <= io_pixelVal_in_1_7;
      end else if (10'h19b == _T_34[9:0]) begin
        image_1_411 <= io_pixelVal_in_1_6;
      end else if (10'h19b == _T_31[9:0]) begin
        image_1_411 <= io_pixelVal_in_1_5;
      end else if (10'h19b == _T_28[9:0]) begin
        image_1_411 <= io_pixelVal_in_1_4;
      end else if (10'h19b == _T_25[9:0]) begin
        image_1_411 <= io_pixelVal_in_1_3;
      end else if (10'h19b == _T_22[9:0]) begin
        image_1_411 <= io_pixelVal_in_1_2;
      end else if (10'h19b == _T_19[9:0]) begin
        image_1_411 <= io_pixelVal_in_1_1;
      end else if (10'h19b == _T_15[9:0]) begin
        image_1_411 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_412 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h19c == _T_37[9:0]) begin
        image_1_412 <= io_pixelVal_in_1_7;
      end else if (10'h19c == _T_34[9:0]) begin
        image_1_412 <= io_pixelVal_in_1_6;
      end else if (10'h19c == _T_31[9:0]) begin
        image_1_412 <= io_pixelVal_in_1_5;
      end else if (10'h19c == _T_28[9:0]) begin
        image_1_412 <= io_pixelVal_in_1_4;
      end else if (10'h19c == _T_25[9:0]) begin
        image_1_412 <= io_pixelVal_in_1_3;
      end else if (10'h19c == _T_22[9:0]) begin
        image_1_412 <= io_pixelVal_in_1_2;
      end else if (10'h19c == _T_19[9:0]) begin
        image_1_412 <= io_pixelVal_in_1_1;
      end else if (10'h19c == _T_15[9:0]) begin
        image_1_412 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_413 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h19d == _T_37[9:0]) begin
        image_1_413 <= io_pixelVal_in_1_7;
      end else if (10'h19d == _T_34[9:0]) begin
        image_1_413 <= io_pixelVal_in_1_6;
      end else if (10'h19d == _T_31[9:0]) begin
        image_1_413 <= io_pixelVal_in_1_5;
      end else if (10'h19d == _T_28[9:0]) begin
        image_1_413 <= io_pixelVal_in_1_4;
      end else if (10'h19d == _T_25[9:0]) begin
        image_1_413 <= io_pixelVal_in_1_3;
      end else if (10'h19d == _T_22[9:0]) begin
        image_1_413 <= io_pixelVal_in_1_2;
      end else if (10'h19d == _T_19[9:0]) begin
        image_1_413 <= io_pixelVal_in_1_1;
      end else if (10'h19d == _T_15[9:0]) begin
        image_1_413 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_414 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h19e == _T_37[9:0]) begin
        image_1_414 <= io_pixelVal_in_1_7;
      end else if (10'h19e == _T_34[9:0]) begin
        image_1_414 <= io_pixelVal_in_1_6;
      end else if (10'h19e == _T_31[9:0]) begin
        image_1_414 <= io_pixelVal_in_1_5;
      end else if (10'h19e == _T_28[9:0]) begin
        image_1_414 <= io_pixelVal_in_1_4;
      end else if (10'h19e == _T_25[9:0]) begin
        image_1_414 <= io_pixelVal_in_1_3;
      end else if (10'h19e == _T_22[9:0]) begin
        image_1_414 <= io_pixelVal_in_1_2;
      end else if (10'h19e == _T_19[9:0]) begin
        image_1_414 <= io_pixelVal_in_1_1;
      end else if (10'h19e == _T_15[9:0]) begin
        image_1_414 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_415 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h19f == _T_37[9:0]) begin
        image_1_415 <= io_pixelVal_in_1_7;
      end else if (10'h19f == _T_34[9:0]) begin
        image_1_415 <= io_pixelVal_in_1_6;
      end else if (10'h19f == _T_31[9:0]) begin
        image_1_415 <= io_pixelVal_in_1_5;
      end else if (10'h19f == _T_28[9:0]) begin
        image_1_415 <= io_pixelVal_in_1_4;
      end else if (10'h19f == _T_25[9:0]) begin
        image_1_415 <= io_pixelVal_in_1_3;
      end else if (10'h19f == _T_22[9:0]) begin
        image_1_415 <= io_pixelVal_in_1_2;
      end else if (10'h19f == _T_19[9:0]) begin
        image_1_415 <= io_pixelVal_in_1_1;
      end else if (10'h19f == _T_15[9:0]) begin
        image_1_415 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_416 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a0 == _T_37[9:0]) begin
        image_1_416 <= io_pixelVal_in_1_7;
      end else if (10'h1a0 == _T_34[9:0]) begin
        image_1_416 <= io_pixelVal_in_1_6;
      end else if (10'h1a0 == _T_31[9:0]) begin
        image_1_416 <= io_pixelVal_in_1_5;
      end else if (10'h1a0 == _T_28[9:0]) begin
        image_1_416 <= io_pixelVal_in_1_4;
      end else if (10'h1a0 == _T_25[9:0]) begin
        image_1_416 <= io_pixelVal_in_1_3;
      end else if (10'h1a0 == _T_22[9:0]) begin
        image_1_416 <= io_pixelVal_in_1_2;
      end else if (10'h1a0 == _T_19[9:0]) begin
        image_1_416 <= io_pixelVal_in_1_1;
      end else if (10'h1a0 == _T_15[9:0]) begin
        image_1_416 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_417 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a1 == _T_37[9:0]) begin
        image_1_417 <= io_pixelVal_in_1_7;
      end else if (10'h1a1 == _T_34[9:0]) begin
        image_1_417 <= io_pixelVal_in_1_6;
      end else if (10'h1a1 == _T_31[9:0]) begin
        image_1_417 <= io_pixelVal_in_1_5;
      end else if (10'h1a1 == _T_28[9:0]) begin
        image_1_417 <= io_pixelVal_in_1_4;
      end else if (10'h1a1 == _T_25[9:0]) begin
        image_1_417 <= io_pixelVal_in_1_3;
      end else if (10'h1a1 == _T_22[9:0]) begin
        image_1_417 <= io_pixelVal_in_1_2;
      end else if (10'h1a1 == _T_19[9:0]) begin
        image_1_417 <= io_pixelVal_in_1_1;
      end else if (10'h1a1 == _T_15[9:0]) begin
        image_1_417 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_418 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a2 == _T_37[9:0]) begin
        image_1_418 <= io_pixelVal_in_1_7;
      end else if (10'h1a2 == _T_34[9:0]) begin
        image_1_418 <= io_pixelVal_in_1_6;
      end else if (10'h1a2 == _T_31[9:0]) begin
        image_1_418 <= io_pixelVal_in_1_5;
      end else if (10'h1a2 == _T_28[9:0]) begin
        image_1_418 <= io_pixelVal_in_1_4;
      end else if (10'h1a2 == _T_25[9:0]) begin
        image_1_418 <= io_pixelVal_in_1_3;
      end else if (10'h1a2 == _T_22[9:0]) begin
        image_1_418 <= io_pixelVal_in_1_2;
      end else if (10'h1a2 == _T_19[9:0]) begin
        image_1_418 <= io_pixelVal_in_1_1;
      end else if (10'h1a2 == _T_15[9:0]) begin
        image_1_418 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_419 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a3 == _T_37[9:0]) begin
        image_1_419 <= io_pixelVal_in_1_7;
      end else if (10'h1a3 == _T_34[9:0]) begin
        image_1_419 <= io_pixelVal_in_1_6;
      end else if (10'h1a3 == _T_31[9:0]) begin
        image_1_419 <= io_pixelVal_in_1_5;
      end else if (10'h1a3 == _T_28[9:0]) begin
        image_1_419 <= io_pixelVal_in_1_4;
      end else if (10'h1a3 == _T_25[9:0]) begin
        image_1_419 <= io_pixelVal_in_1_3;
      end else if (10'h1a3 == _T_22[9:0]) begin
        image_1_419 <= io_pixelVal_in_1_2;
      end else if (10'h1a3 == _T_19[9:0]) begin
        image_1_419 <= io_pixelVal_in_1_1;
      end else if (10'h1a3 == _T_15[9:0]) begin
        image_1_419 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_420 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a4 == _T_37[9:0]) begin
        image_1_420 <= io_pixelVal_in_1_7;
      end else if (10'h1a4 == _T_34[9:0]) begin
        image_1_420 <= io_pixelVal_in_1_6;
      end else if (10'h1a4 == _T_31[9:0]) begin
        image_1_420 <= io_pixelVal_in_1_5;
      end else if (10'h1a4 == _T_28[9:0]) begin
        image_1_420 <= io_pixelVal_in_1_4;
      end else if (10'h1a4 == _T_25[9:0]) begin
        image_1_420 <= io_pixelVal_in_1_3;
      end else if (10'h1a4 == _T_22[9:0]) begin
        image_1_420 <= io_pixelVal_in_1_2;
      end else if (10'h1a4 == _T_19[9:0]) begin
        image_1_420 <= io_pixelVal_in_1_1;
      end else if (10'h1a4 == _T_15[9:0]) begin
        image_1_420 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_421 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a5 == _T_37[9:0]) begin
        image_1_421 <= io_pixelVal_in_1_7;
      end else if (10'h1a5 == _T_34[9:0]) begin
        image_1_421 <= io_pixelVal_in_1_6;
      end else if (10'h1a5 == _T_31[9:0]) begin
        image_1_421 <= io_pixelVal_in_1_5;
      end else if (10'h1a5 == _T_28[9:0]) begin
        image_1_421 <= io_pixelVal_in_1_4;
      end else if (10'h1a5 == _T_25[9:0]) begin
        image_1_421 <= io_pixelVal_in_1_3;
      end else if (10'h1a5 == _T_22[9:0]) begin
        image_1_421 <= io_pixelVal_in_1_2;
      end else if (10'h1a5 == _T_19[9:0]) begin
        image_1_421 <= io_pixelVal_in_1_1;
      end else if (10'h1a5 == _T_15[9:0]) begin
        image_1_421 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_422 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a6 == _T_37[9:0]) begin
        image_1_422 <= io_pixelVal_in_1_7;
      end else if (10'h1a6 == _T_34[9:0]) begin
        image_1_422 <= io_pixelVal_in_1_6;
      end else if (10'h1a6 == _T_31[9:0]) begin
        image_1_422 <= io_pixelVal_in_1_5;
      end else if (10'h1a6 == _T_28[9:0]) begin
        image_1_422 <= io_pixelVal_in_1_4;
      end else if (10'h1a6 == _T_25[9:0]) begin
        image_1_422 <= io_pixelVal_in_1_3;
      end else if (10'h1a6 == _T_22[9:0]) begin
        image_1_422 <= io_pixelVal_in_1_2;
      end else if (10'h1a6 == _T_19[9:0]) begin
        image_1_422 <= io_pixelVal_in_1_1;
      end else if (10'h1a6 == _T_15[9:0]) begin
        image_1_422 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_423 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a7 == _T_37[9:0]) begin
        image_1_423 <= io_pixelVal_in_1_7;
      end else if (10'h1a7 == _T_34[9:0]) begin
        image_1_423 <= io_pixelVal_in_1_6;
      end else if (10'h1a7 == _T_31[9:0]) begin
        image_1_423 <= io_pixelVal_in_1_5;
      end else if (10'h1a7 == _T_28[9:0]) begin
        image_1_423 <= io_pixelVal_in_1_4;
      end else if (10'h1a7 == _T_25[9:0]) begin
        image_1_423 <= io_pixelVal_in_1_3;
      end else if (10'h1a7 == _T_22[9:0]) begin
        image_1_423 <= io_pixelVal_in_1_2;
      end else if (10'h1a7 == _T_19[9:0]) begin
        image_1_423 <= io_pixelVal_in_1_1;
      end else if (10'h1a7 == _T_15[9:0]) begin
        image_1_423 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_424 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a8 == _T_37[9:0]) begin
        image_1_424 <= io_pixelVal_in_1_7;
      end else if (10'h1a8 == _T_34[9:0]) begin
        image_1_424 <= io_pixelVal_in_1_6;
      end else if (10'h1a8 == _T_31[9:0]) begin
        image_1_424 <= io_pixelVal_in_1_5;
      end else if (10'h1a8 == _T_28[9:0]) begin
        image_1_424 <= io_pixelVal_in_1_4;
      end else if (10'h1a8 == _T_25[9:0]) begin
        image_1_424 <= io_pixelVal_in_1_3;
      end else if (10'h1a8 == _T_22[9:0]) begin
        image_1_424 <= io_pixelVal_in_1_2;
      end else if (10'h1a8 == _T_19[9:0]) begin
        image_1_424 <= io_pixelVal_in_1_1;
      end else if (10'h1a8 == _T_15[9:0]) begin
        image_1_424 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_425 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a9 == _T_37[9:0]) begin
        image_1_425 <= io_pixelVal_in_1_7;
      end else if (10'h1a9 == _T_34[9:0]) begin
        image_1_425 <= io_pixelVal_in_1_6;
      end else if (10'h1a9 == _T_31[9:0]) begin
        image_1_425 <= io_pixelVal_in_1_5;
      end else if (10'h1a9 == _T_28[9:0]) begin
        image_1_425 <= io_pixelVal_in_1_4;
      end else if (10'h1a9 == _T_25[9:0]) begin
        image_1_425 <= io_pixelVal_in_1_3;
      end else if (10'h1a9 == _T_22[9:0]) begin
        image_1_425 <= io_pixelVal_in_1_2;
      end else if (10'h1a9 == _T_19[9:0]) begin
        image_1_425 <= io_pixelVal_in_1_1;
      end else if (10'h1a9 == _T_15[9:0]) begin
        image_1_425 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_426 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1aa == _T_37[9:0]) begin
        image_1_426 <= io_pixelVal_in_1_7;
      end else if (10'h1aa == _T_34[9:0]) begin
        image_1_426 <= io_pixelVal_in_1_6;
      end else if (10'h1aa == _T_31[9:0]) begin
        image_1_426 <= io_pixelVal_in_1_5;
      end else if (10'h1aa == _T_28[9:0]) begin
        image_1_426 <= io_pixelVal_in_1_4;
      end else if (10'h1aa == _T_25[9:0]) begin
        image_1_426 <= io_pixelVal_in_1_3;
      end else if (10'h1aa == _T_22[9:0]) begin
        image_1_426 <= io_pixelVal_in_1_2;
      end else if (10'h1aa == _T_19[9:0]) begin
        image_1_426 <= io_pixelVal_in_1_1;
      end else if (10'h1aa == _T_15[9:0]) begin
        image_1_426 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_427 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ab == _T_37[9:0]) begin
        image_1_427 <= io_pixelVal_in_1_7;
      end else if (10'h1ab == _T_34[9:0]) begin
        image_1_427 <= io_pixelVal_in_1_6;
      end else if (10'h1ab == _T_31[9:0]) begin
        image_1_427 <= io_pixelVal_in_1_5;
      end else if (10'h1ab == _T_28[9:0]) begin
        image_1_427 <= io_pixelVal_in_1_4;
      end else if (10'h1ab == _T_25[9:0]) begin
        image_1_427 <= io_pixelVal_in_1_3;
      end else if (10'h1ab == _T_22[9:0]) begin
        image_1_427 <= io_pixelVal_in_1_2;
      end else if (10'h1ab == _T_19[9:0]) begin
        image_1_427 <= io_pixelVal_in_1_1;
      end else if (10'h1ab == _T_15[9:0]) begin
        image_1_427 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_428 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ac == _T_37[9:0]) begin
        image_1_428 <= io_pixelVal_in_1_7;
      end else if (10'h1ac == _T_34[9:0]) begin
        image_1_428 <= io_pixelVal_in_1_6;
      end else if (10'h1ac == _T_31[9:0]) begin
        image_1_428 <= io_pixelVal_in_1_5;
      end else if (10'h1ac == _T_28[9:0]) begin
        image_1_428 <= io_pixelVal_in_1_4;
      end else if (10'h1ac == _T_25[9:0]) begin
        image_1_428 <= io_pixelVal_in_1_3;
      end else if (10'h1ac == _T_22[9:0]) begin
        image_1_428 <= io_pixelVal_in_1_2;
      end else if (10'h1ac == _T_19[9:0]) begin
        image_1_428 <= io_pixelVal_in_1_1;
      end else if (10'h1ac == _T_15[9:0]) begin
        image_1_428 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_429 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ad == _T_37[9:0]) begin
        image_1_429 <= io_pixelVal_in_1_7;
      end else if (10'h1ad == _T_34[9:0]) begin
        image_1_429 <= io_pixelVal_in_1_6;
      end else if (10'h1ad == _T_31[9:0]) begin
        image_1_429 <= io_pixelVal_in_1_5;
      end else if (10'h1ad == _T_28[9:0]) begin
        image_1_429 <= io_pixelVal_in_1_4;
      end else if (10'h1ad == _T_25[9:0]) begin
        image_1_429 <= io_pixelVal_in_1_3;
      end else if (10'h1ad == _T_22[9:0]) begin
        image_1_429 <= io_pixelVal_in_1_2;
      end else if (10'h1ad == _T_19[9:0]) begin
        image_1_429 <= io_pixelVal_in_1_1;
      end else if (10'h1ad == _T_15[9:0]) begin
        image_1_429 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_430 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ae == _T_37[9:0]) begin
        image_1_430 <= io_pixelVal_in_1_7;
      end else if (10'h1ae == _T_34[9:0]) begin
        image_1_430 <= io_pixelVal_in_1_6;
      end else if (10'h1ae == _T_31[9:0]) begin
        image_1_430 <= io_pixelVal_in_1_5;
      end else if (10'h1ae == _T_28[9:0]) begin
        image_1_430 <= io_pixelVal_in_1_4;
      end else if (10'h1ae == _T_25[9:0]) begin
        image_1_430 <= io_pixelVal_in_1_3;
      end else if (10'h1ae == _T_22[9:0]) begin
        image_1_430 <= io_pixelVal_in_1_2;
      end else if (10'h1ae == _T_19[9:0]) begin
        image_1_430 <= io_pixelVal_in_1_1;
      end else if (10'h1ae == _T_15[9:0]) begin
        image_1_430 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_431 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1af == _T_37[9:0]) begin
        image_1_431 <= io_pixelVal_in_1_7;
      end else if (10'h1af == _T_34[9:0]) begin
        image_1_431 <= io_pixelVal_in_1_6;
      end else if (10'h1af == _T_31[9:0]) begin
        image_1_431 <= io_pixelVal_in_1_5;
      end else if (10'h1af == _T_28[9:0]) begin
        image_1_431 <= io_pixelVal_in_1_4;
      end else if (10'h1af == _T_25[9:0]) begin
        image_1_431 <= io_pixelVal_in_1_3;
      end else if (10'h1af == _T_22[9:0]) begin
        image_1_431 <= io_pixelVal_in_1_2;
      end else if (10'h1af == _T_19[9:0]) begin
        image_1_431 <= io_pixelVal_in_1_1;
      end else if (10'h1af == _T_15[9:0]) begin
        image_1_431 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_432 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b0 == _T_37[9:0]) begin
        image_1_432 <= io_pixelVal_in_1_7;
      end else if (10'h1b0 == _T_34[9:0]) begin
        image_1_432 <= io_pixelVal_in_1_6;
      end else if (10'h1b0 == _T_31[9:0]) begin
        image_1_432 <= io_pixelVal_in_1_5;
      end else if (10'h1b0 == _T_28[9:0]) begin
        image_1_432 <= io_pixelVal_in_1_4;
      end else if (10'h1b0 == _T_25[9:0]) begin
        image_1_432 <= io_pixelVal_in_1_3;
      end else if (10'h1b0 == _T_22[9:0]) begin
        image_1_432 <= io_pixelVal_in_1_2;
      end else if (10'h1b0 == _T_19[9:0]) begin
        image_1_432 <= io_pixelVal_in_1_1;
      end else if (10'h1b0 == _T_15[9:0]) begin
        image_1_432 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_433 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b1 == _T_37[9:0]) begin
        image_1_433 <= io_pixelVal_in_1_7;
      end else if (10'h1b1 == _T_34[9:0]) begin
        image_1_433 <= io_pixelVal_in_1_6;
      end else if (10'h1b1 == _T_31[9:0]) begin
        image_1_433 <= io_pixelVal_in_1_5;
      end else if (10'h1b1 == _T_28[9:0]) begin
        image_1_433 <= io_pixelVal_in_1_4;
      end else if (10'h1b1 == _T_25[9:0]) begin
        image_1_433 <= io_pixelVal_in_1_3;
      end else if (10'h1b1 == _T_22[9:0]) begin
        image_1_433 <= io_pixelVal_in_1_2;
      end else if (10'h1b1 == _T_19[9:0]) begin
        image_1_433 <= io_pixelVal_in_1_1;
      end else if (10'h1b1 == _T_15[9:0]) begin
        image_1_433 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_434 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b2 == _T_37[9:0]) begin
        image_1_434 <= io_pixelVal_in_1_7;
      end else if (10'h1b2 == _T_34[9:0]) begin
        image_1_434 <= io_pixelVal_in_1_6;
      end else if (10'h1b2 == _T_31[9:0]) begin
        image_1_434 <= io_pixelVal_in_1_5;
      end else if (10'h1b2 == _T_28[9:0]) begin
        image_1_434 <= io_pixelVal_in_1_4;
      end else if (10'h1b2 == _T_25[9:0]) begin
        image_1_434 <= io_pixelVal_in_1_3;
      end else if (10'h1b2 == _T_22[9:0]) begin
        image_1_434 <= io_pixelVal_in_1_2;
      end else if (10'h1b2 == _T_19[9:0]) begin
        image_1_434 <= io_pixelVal_in_1_1;
      end else if (10'h1b2 == _T_15[9:0]) begin
        image_1_434 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_435 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b3 == _T_37[9:0]) begin
        image_1_435 <= io_pixelVal_in_1_7;
      end else if (10'h1b3 == _T_34[9:0]) begin
        image_1_435 <= io_pixelVal_in_1_6;
      end else if (10'h1b3 == _T_31[9:0]) begin
        image_1_435 <= io_pixelVal_in_1_5;
      end else if (10'h1b3 == _T_28[9:0]) begin
        image_1_435 <= io_pixelVal_in_1_4;
      end else if (10'h1b3 == _T_25[9:0]) begin
        image_1_435 <= io_pixelVal_in_1_3;
      end else if (10'h1b3 == _T_22[9:0]) begin
        image_1_435 <= io_pixelVal_in_1_2;
      end else if (10'h1b3 == _T_19[9:0]) begin
        image_1_435 <= io_pixelVal_in_1_1;
      end else if (10'h1b3 == _T_15[9:0]) begin
        image_1_435 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_436 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b4 == _T_37[9:0]) begin
        image_1_436 <= io_pixelVal_in_1_7;
      end else if (10'h1b4 == _T_34[9:0]) begin
        image_1_436 <= io_pixelVal_in_1_6;
      end else if (10'h1b4 == _T_31[9:0]) begin
        image_1_436 <= io_pixelVal_in_1_5;
      end else if (10'h1b4 == _T_28[9:0]) begin
        image_1_436 <= io_pixelVal_in_1_4;
      end else if (10'h1b4 == _T_25[9:0]) begin
        image_1_436 <= io_pixelVal_in_1_3;
      end else if (10'h1b4 == _T_22[9:0]) begin
        image_1_436 <= io_pixelVal_in_1_2;
      end else if (10'h1b4 == _T_19[9:0]) begin
        image_1_436 <= io_pixelVal_in_1_1;
      end else if (10'h1b4 == _T_15[9:0]) begin
        image_1_436 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_437 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b5 == _T_37[9:0]) begin
        image_1_437 <= io_pixelVal_in_1_7;
      end else if (10'h1b5 == _T_34[9:0]) begin
        image_1_437 <= io_pixelVal_in_1_6;
      end else if (10'h1b5 == _T_31[9:0]) begin
        image_1_437 <= io_pixelVal_in_1_5;
      end else if (10'h1b5 == _T_28[9:0]) begin
        image_1_437 <= io_pixelVal_in_1_4;
      end else if (10'h1b5 == _T_25[9:0]) begin
        image_1_437 <= io_pixelVal_in_1_3;
      end else if (10'h1b5 == _T_22[9:0]) begin
        image_1_437 <= io_pixelVal_in_1_2;
      end else if (10'h1b5 == _T_19[9:0]) begin
        image_1_437 <= io_pixelVal_in_1_1;
      end else if (10'h1b5 == _T_15[9:0]) begin
        image_1_437 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_438 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b6 == _T_37[9:0]) begin
        image_1_438 <= io_pixelVal_in_1_7;
      end else if (10'h1b6 == _T_34[9:0]) begin
        image_1_438 <= io_pixelVal_in_1_6;
      end else if (10'h1b6 == _T_31[9:0]) begin
        image_1_438 <= io_pixelVal_in_1_5;
      end else if (10'h1b6 == _T_28[9:0]) begin
        image_1_438 <= io_pixelVal_in_1_4;
      end else if (10'h1b6 == _T_25[9:0]) begin
        image_1_438 <= io_pixelVal_in_1_3;
      end else if (10'h1b6 == _T_22[9:0]) begin
        image_1_438 <= io_pixelVal_in_1_2;
      end else if (10'h1b6 == _T_19[9:0]) begin
        image_1_438 <= io_pixelVal_in_1_1;
      end else if (10'h1b6 == _T_15[9:0]) begin
        image_1_438 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_439 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b7 == _T_37[9:0]) begin
        image_1_439 <= io_pixelVal_in_1_7;
      end else if (10'h1b7 == _T_34[9:0]) begin
        image_1_439 <= io_pixelVal_in_1_6;
      end else if (10'h1b7 == _T_31[9:0]) begin
        image_1_439 <= io_pixelVal_in_1_5;
      end else if (10'h1b7 == _T_28[9:0]) begin
        image_1_439 <= io_pixelVal_in_1_4;
      end else if (10'h1b7 == _T_25[9:0]) begin
        image_1_439 <= io_pixelVal_in_1_3;
      end else if (10'h1b7 == _T_22[9:0]) begin
        image_1_439 <= io_pixelVal_in_1_2;
      end else if (10'h1b7 == _T_19[9:0]) begin
        image_1_439 <= io_pixelVal_in_1_1;
      end else if (10'h1b7 == _T_15[9:0]) begin
        image_1_439 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_440 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b8 == _T_37[9:0]) begin
        image_1_440 <= io_pixelVal_in_1_7;
      end else if (10'h1b8 == _T_34[9:0]) begin
        image_1_440 <= io_pixelVal_in_1_6;
      end else if (10'h1b8 == _T_31[9:0]) begin
        image_1_440 <= io_pixelVal_in_1_5;
      end else if (10'h1b8 == _T_28[9:0]) begin
        image_1_440 <= io_pixelVal_in_1_4;
      end else if (10'h1b8 == _T_25[9:0]) begin
        image_1_440 <= io_pixelVal_in_1_3;
      end else if (10'h1b8 == _T_22[9:0]) begin
        image_1_440 <= io_pixelVal_in_1_2;
      end else if (10'h1b8 == _T_19[9:0]) begin
        image_1_440 <= io_pixelVal_in_1_1;
      end else if (10'h1b8 == _T_15[9:0]) begin
        image_1_440 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_441 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b9 == _T_37[9:0]) begin
        image_1_441 <= io_pixelVal_in_1_7;
      end else if (10'h1b9 == _T_34[9:0]) begin
        image_1_441 <= io_pixelVal_in_1_6;
      end else if (10'h1b9 == _T_31[9:0]) begin
        image_1_441 <= io_pixelVal_in_1_5;
      end else if (10'h1b9 == _T_28[9:0]) begin
        image_1_441 <= io_pixelVal_in_1_4;
      end else if (10'h1b9 == _T_25[9:0]) begin
        image_1_441 <= io_pixelVal_in_1_3;
      end else if (10'h1b9 == _T_22[9:0]) begin
        image_1_441 <= io_pixelVal_in_1_2;
      end else if (10'h1b9 == _T_19[9:0]) begin
        image_1_441 <= io_pixelVal_in_1_1;
      end else if (10'h1b9 == _T_15[9:0]) begin
        image_1_441 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_442 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ba == _T_37[9:0]) begin
        image_1_442 <= io_pixelVal_in_1_7;
      end else if (10'h1ba == _T_34[9:0]) begin
        image_1_442 <= io_pixelVal_in_1_6;
      end else if (10'h1ba == _T_31[9:0]) begin
        image_1_442 <= io_pixelVal_in_1_5;
      end else if (10'h1ba == _T_28[9:0]) begin
        image_1_442 <= io_pixelVal_in_1_4;
      end else if (10'h1ba == _T_25[9:0]) begin
        image_1_442 <= io_pixelVal_in_1_3;
      end else if (10'h1ba == _T_22[9:0]) begin
        image_1_442 <= io_pixelVal_in_1_2;
      end else if (10'h1ba == _T_19[9:0]) begin
        image_1_442 <= io_pixelVal_in_1_1;
      end else if (10'h1ba == _T_15[9:0]) begin
        image_1_442 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_443 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1bb == _T_37[9:0]) begin
        image_1_443 <= io_pixelVal_in_1_7;
      end else if (10'h1bb == _T_34[9:0]) begin
        image_1_443 <= io_pixelVal_in_1_6;
      end else if (10'h1bb == _T_31[9:0]) begin
        image_1_443 <= io_pixelVal_in_1_5;
      end else if (10'h1bb == _T_28[9:0]) begin
        image_1_443 <= io_pixelVal_in_1_4;
      end else if (10'h1bb == _T_25[9:0]) begin
        image_1_443 <= io_pixelVal_in_1_3;
      end else if (10'h1bb == _T_22[9:0]) begin
        image_1_443 <= io_pixelVal_in_1_2;
      end else if (10'h1bb == _T_19[9:0]) begin
        image_1_443 <= io_pixelVal_in_1_1;
      end else if (10'h1bb == _T_15[9:0]) begin
        image_1_443 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_444 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1bc == _T_37[9:0]) begin
        image_1_444 <= io_pixelVal_in_1_7;
      end else if (10'h1bc == _T_34[9:0]) begin
        image_1_444 <= io_pixelVal_in_1_6;
      end else if (10'h1bc == _T_31[9:0]) begin
        image_1_444 <= io_pixelVal_in_1_5;
      end else if (10'h1bc == _T_28[9:0]) begin
        image_1_444 <= io_pixelVal_in_1_4;
      end else if (10'h1bc == _T_25[9:0]) begin
        image_1_444 <= io_pixelVal_in_1_3;
      end else if (10'h1bc == _T_22[9:0]) begin
        image_1_444 <= io_pixelVal_in_1_2;
      end else if (10'h1bc == _T_19[9:0]) begin
        image_1_444 <= io_pixelVal_in_1_1;
      end else if (10'h1bc == _T_15[9:0]) begin
        image_1_444 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_445 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1bd == _T_37[9:0]) begin
        image_1_445 <= io_pixelVal_in_1_7;
      end else if (10'h1bd == _T_34[9:0]) begin
        image_1_445 <= io_pixelVal_in_1_6;
      end else if (10'h1bd == _T_31[9:0]) begin
        image_1_445 <= io_pixelVal_in_1_5;
      end else if (10'h1bd == _T_28[9:0]) begin
        image_1_445 <= io_pixelVal_in_1_4;
      end else if (10'h1bd == _T_25[9:0]) begin
        image_1_445 <= io_pixelVal_in_1_3;
      end else if (10'h1bd == _T_22[9:0]) begin
        image_1_445 <= io_pixelVal_in_1_2;
      end else if (10'h1bd == _T_19[9:0]) begin
        image_1_445 <= io_pixelVal_in_1_1;
      end else if (10'h1bd == _T_15[9:0]) begin
        image_1_445 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_446 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1be == _T_37[9:0]) begin
        image_1_446 <= io_pixelVal_in_1_7;
      end else if (10'h1be == _T_34[9:0]) begin
        image_1_446 <= io_pixelVal_in_1_6;
      end else if (10'h1be == _T_31[9:0]) begin
        image_1_446 <= io_pixelVal_in_1_5;
      end else if (10'h1be == _T_28[9:0]) begin
        image_1_446 <= io_pixelVal_in_1_4;
      end else if (10'h1be == _T_25[9:0]) begin
        image_1_446 <= io_pixelVal_in_1_3;
      end else if (10'h1be == _T_22[9:0]) begin
        image_1_446 <= io_pixelVal_in_1_2;
      end else if (10'h1be == _T_19[9:0]) begin
        image_1_446 <= io_pixelVal_in_1_1;
      end else if (10'h1be == _T_15[9:0]) begin
        image_1_446 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_447 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1bf == _T_37[9:0]) begin
        image_1_447 <= io_pixelVal_in_1_7;
      end else if (10'h1bf == _T_34[9:0]) begin
        image_1_447 <= io_pixelVal_in_1_6;
      end else if (10'h1bf == _T_31[9:0]) begin
        image_1_447 <= io_pixelVal_in_1_5;
      end else if (10'h1bf == _T_28[9:0]) begin
        image_1_447 <= io_pixelVal_in_1_4;
      end else if (10'h1bf == _T_25[9:0]) begin
        image_1_447 <= io_pixelVal_in_1_3;
      end else if (10'h1bf == _T_22[9:0]) begin
        image_1_447 <= io_pixelVal_in_1_2;
      end else if (10'h1bf == _T_19[9:0]) begin
        image_1_447 <= io_pixelVal_in_1_1;
      end else if (10'h1bf == _T_15[9:0]) begin
        image_1_447 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_448 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c0 == _T_37[9:0]) begin
        image_1_448 <= io_pixelVal_in_1_7;
      end else if (10'h1c0 == _T_34[9:0]) begin
        image_1_448 <= io_pixelVal_in_1_6;
      end else if (10'h1c0 == _T_31[9:0]) begin
        image_1_448 <= io_pixelVal_in_1_5;
      end else if (10'h1c0 == _T_28[9:0]) begin
        image_1_448 <= io_pixelVal_in_1_4;
      end else if (10'h1c0 == _T_25[9:0]) begin
        image_1_448 <= io_pixelVal_in_1_3;
      end else if (10'h1c0 == _T_22[9:0]) begin
        image_1_448 <= io_pixelVal_in_1_2;
      end else if (10'h1c0 == _T_19[9:0]) begin
        image_1_448 <= io_pixelVal_in_1_1;
      end else if (10'h1c0 == _T_15[9:0]) begin
        image_1_448 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_449 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c1 == _T_37[9:0]) begin
        image_1_449 <= io_pixelVal_in_1_7;
      end else if (10'h1c1 == _T_34[9:0]) begin
        image_1_449 <= io_pixelVal_in_1_6;
      end else if (10'h1c1 == _T_31[9:0]) begin
        image_1_449 <= io_pixelVal_in_1_5;
      end else if (10'h1c1 == _T_28[9:0]) begin
        image_1_449 <= io_pixelVal_in_1_4;
      end else if (10'h1c1 == _T_25[9:0]) begin
        image_1_449 <= io_pixelVal_in_1_3;
      end else if (10'h1c1 == _T_22[9:0]) begin
        image_1_449 <= io_pixelVal_in_1_2;
      end else if (10'h1c1 == _T_19[9:0]) begin
        image_1_449 <= io_pixelVal_in_1_1;
      end else if (10'h1c1 == _T_15[9:0]) begin
        image_1_449 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_450 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c2 == _T_37[9:0]) begin
        image_1_450 <= io_pixelVal_in_1_7;
      end else if (10'h1c2 == _T_34[9:0]) begin
        image_1_450 <= io_pixelVal_in_1_6;
      end else if (10'h1c2 == _T_31[9:0]) begin
        image_1_450 <= io_pixelVal_in_1_5;
      end else if (10'h1c2 == _T_28[9:0]) begin
        image_1_450 <= io_pixelVal_in_1_4;
      end else if (10'h1c2 == _T_25[9:0]) begin
        image_1_450 <= io_pixelVal_in_1_3;
      end else if (10'h1c2 == _T_22[9:0]) begin
        image_1_450 <= io_pixelVal_in_1_2;
      end else if (10'h1c2 == _T_19[9:0]) begin
        image_1_450 <= io_pixelVal_in_1_1;
      end else if (10'h1c2 == _T_15[9:0]) begin
        image_1_450 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_451 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c3 == _T_37[9:0]) begin
        image_1_451 <= io_pixelVal_in_1_7;
      end else if (10'h1c3 == _T_34[9:0]) begin
        image_1_451 <= io_pixelVal_in_1_6;
      end else if (10'h1c3 == _T_31[9:0]) begin
        image_1_451 <= io_pixelVal_in_1_5;
      end else if (10'h1c3 == _T_28[9:0]) begin
        image_1_451 <= io_pixelVal_in_1_4;
      end else if (10'h1c3 == _T_25[9:0]) begin
        image_1_451 <= io_pixelVal_in_1_3;
      end else if (10'h1c3 == _T_22[9:0]) begin
        image_1_451 <= io_pixelVal_in_1_2;
      end else if (10'h1c3 == _T_19[9:0]) begin
        image_1_451 <= io_pixelVal_in_1_1;
      end else if (10'h1c3 == _T_15[9:0]) begin
        image_1_451 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_452 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c4 == _T_37[9:0]) begin
        image_1_452 <= io_pixelVal_in_1_7;
      end else if (10'h1c4 == _T_34[9:0]) begin
        image_1_452 <= io_pixelVal_in_1_6;
      end else if (10'h1c4 == _T_31[9:0]) begin
        image_1_452 <= io_pixelVal_in_1_5;
      end else if (10'h1c4 == _T_28[9:0]) begin
        image_1_452 <= io_pixelVal_in_1_4;
      end else if (10'h1c4 == _T_25[9:0]) begin
        image_1_452 <= io_pixelVal_in_1_3;
      end else if (10'h1c4 == _T_22[9:0]) begin
        image_1_452 <= io_pixelVal_in_1_2;
      end else if (10'h1c4 == _T_19[9:0]) begin
        image_1_452 <= io_pixelVal_in_1_1;
      end else if (10'h1c4 == _T_15[9:0]) begin
        image_1_452 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_453 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c5 == _T_37[9:0]) begin
        image_1_453 <= io_pixelVal_in_1_7;
      end else if (10'h1c5 == _T_34[9:0]) begin
        image_1_453 <= io_pixelVal_in_1_6;
      end else if (10'h1c5 == _T_31[9:0]) begin
        image_1_453 <= io_pixelVal_in_1_5;
      end else if (10'h1c5 == _T_28[9:0]) begin
        image_1_453 <= io_pixelVal_in_1_4;
      end else if (10'h1c5 == _T_25[9:0]) begin
        image_1_453 <= io_pixelVal_in_1_3;
      end else if (10'h1c5 == _T_22[9:0]) begin
        image_1_453 <= io_pixelVal_in_1_2;
      end else if (10'h1c5 == _T_19[9:0]) begin
        image_1_453 <= io_pixelVal_in_1_1;
      end else if (10'h1c5 == _T_15[9:0]) begin
        image_1_453 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_454 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c6 == _T_37[9:0]) begin
        image_1_454 <= io_pixelVal_in_1_7;
      end else if (10'h1c6 == _T_34[9:0]) begin
        image_1_454 <= io_pixelVal_in_1_6;
      end else if (10'h1c6 == _T_31[9:0]) begin
        image_1_454 <= io_pixelVal_in_1_5;
      end else if (10'h1c6 == _T_28[9:0]) begin
        image_1_454 <= io_pixelVal_in_1_4;
      end else if (10'h1c6 == _T_25[9:0]) begin
        image_1_454 <= io_pixelVal_in_1_3;
      end else if (10'h1c6 == _T_22[9:0]) begin
        image_1_454 <= io_pixelVal_in_1_2;
      end else if (10'h1c6 == _T_19[9:0]) begin
        image_1_454 <= io_pixelVal_in_1_1;
      end else if (10'h1c6 == _T_15[9:0]) begin
        image_1_454 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_455 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c7 == _T_37[9:0]) begin
        image_1_455 <= io_pixelVal_in_1_7;
      end else if (10'h1c7 == _T_34[9:0]) begin
        image_1_455 <= io_pixelVal_in_1_6;
      end else if (10'h1c7 == _T_31[9:0]) begin
        image_1_455 <= io_pixelVal_in_1_5;
      end else if (10'h1c7 == _T_28[9:0]) begin
        image_1_455 <= io_pixelVal_in_1_4;
      end else if (10'h1c7 == _T_25[9:0]) begin
        image_1_455 <= io_pixelVal_in_1_3;
      end else if (10'h1c7 == _T_22[9:0]) begin
        image_1_455 <= io_pixelVal_in_1_2;
      end else if (10'h1c7 == _T_19[9:0]) begin
        image_1_455 <= io_pixelVal_in_1_1;
      end else if (10'h1c7 == _T_15[9:0]) begin
        image_1_455 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_456 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c8 == _T_37[9:0]) begin
        image_1_456 <= io_pixelVal_in_1_7;
      end else if (10'h1c8 == _T_34[9:0]) begin
        image_1_456 <= io_pixelVal_in_1_6;
      end else if (10'h1c8 == _T_31[9:0]) begin
        image_1_456 <= io_pixelVal_in_1_5;
      end else if (10'h1c8 == _T_28[9:0]) begin
        image_1_456 <= io_pixelVal_in_1_4;
      end else if (10'h1c8 == _T_25[9:0]) begin
        image_1_456 <= io_pixelVal_in_1_3;
      end else if (10'h1c8 == _T_22[9:0]) begin
        image_1_456 <= io_pixelVal_in_1_2;
      end else if (10'h1c8 == _T_19[9:0]) begin
        image_1_456 <= io_pixelVal_in_1_1;
      end else if (10'h1c8 == _T_15[9:0]) begin
        image_1_456 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_457 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c9 == _T_37[9:0]) begin
        image_1_457 <= io_pixelVal_in_1_7;
      end else if (10'h1c9 == _T_34[9:0]) begin
        image_1_457 <= io_pixelVal_in_1_6;
      end else if (10'h1c9 == _T_31[9:0]) begin
        image_1_457 <= io_pixelVal_in_1_5;
      end else if (10'h1c9 == _T_28[9:0]) begin
        image_1_457 <= io_pixelVal_in_1_4;
      end else if (10'h1c9 == _T_25[9:0]) begin
        image_1_457 <= io_pixelVal_in_1_3;
      end else if (10'h1c9 == _T_22[9:0]) begin
        image_1_457 <= io_pixelVal_in_1_2;
      end else if (10'h1c9 == _T_19[9:0]) begin
        image_1_457 <= io_pixelVal_in_1_1;
      end else if (10'h1c9 == _T_15[9:0]) begin
        image_1_457 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_458 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ca == _T_37[9:0]) begin
        image_1_458 <= io_pixelVal_in_1_7;
      end else if (10'h1ca == _T_34[9:0]) begin
        image_1_458 <= io_pixelVal_in_1_6;
      end else if (10'h1ca == _T_31[9:0]) begin
        image_1_458 <= io_pixelVal_in_1_5;
      end else if (10'h1ca == _T_28[9:0]) begin
        image_1_458 <= io_pixelVal_in_1_4;
      end else if (10'h1ca == _T_25[9:0]) begin
        image_1_458 <= io_pixelVal_in_1_3;
      end else if (10'h1ca == _T_22[9:0]) begin
        image_1_458 <= io_pixelVal_in_1_2;
      end else if (10'h1ca == _T_19[9:0]) begin
        image_1_458 <= io_pixelVal_in_1_1;
      end else if (10'h1ca == _T_15[9:0]) begin
        image_1_458 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_459 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1cb == _T_37[9:0]) begin
        image_1_459 <= io_pixelVal_in_1_7;
      end else if (10'h1cb == _T_34[9:0]) begin
        image_1_459 <= io_pixelVal_in_1_6;
      end else if (10'h1cb == _T_31[9:0]) begin
        image_1_459 <= io_pixelVal_in_1_5;
      end else if (10'h1cb == _T_28[9:0]) begin
        image_1_459 <= io_pixelVal_in_1_4;
      end else if (10'h1cb == _T_25[9:0]) begin
        image_1_459 <= io_pixelVal_in_1_3;
      end else if (10'h1cb == _T_22[9:0]) begin
        image_1_459 <= io_pixelVal_in_1_2;
      end else if (10'h1cb == _T_19[9:0]) begin
        image_1_459 <= io_pixelVal_in_1_1;
      end else if (10'h1cb == _T_15[9:0]) begin
        image_1_459 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_460 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1cc == _T_37[9:0]) begin
        image_1_460 <= io_pixelVal_in_1_7;
      end else if (10'h1cc == _T_34[9:0]) begin
        image_1_460 <= io_pixelVal_in_1_6;
      end else if (10'h1cc == _T_31[9:0]) begin
        image_1_460 <= io_pixelVal_in_1_5;
      end else if (10'h1cc == _T_28[9:0]) begin
        image_1_460 <= io_pixelVal_in_1_4;
      end else if (10'h1cc == _T_25[9:0]) begin
        image_1_460 <= io_pixelVal_in_1_3;
      end else if (10'h1cc == _T_22[9:0]) begin
        image_1_460 <= io_pixelVal_in_1_2;
      end else if (10'h1cc == _T_19[9:0]) begin
        image_1_460 <= io_pixelVal_in_1_1;
      end else if (10'h1cc == _T_15[9:0]) begin
        image_1_460 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_461 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1cd == _T_37[9:0]) begin
        image_1_461 <= io_pixelVal_in_1_7;
      end else if (10'h1cd == _T_34[9:0]) begin
        image_1_461 <= io_pixelVal_in_1_6;
      end else if (10'h1cd == _T_31[9:0]) begin
        image_1_461 <= io_pixelVal_in_1_5;
      end else if (10'h1cd == _T_28[9:0]) begin
        image_1_461 <= io_pixelVal_in_1_4;
      end else if (10'h1cd == _T_25[9:0]) begin
        image_1_461 <= io_pixelVal_in_1_3;
      end else if (10'h1cd == _T_22[9:0]) begin
        image_1_461 <= io_pixelVal_in_1_2;
      end else if (10'h1cd == _T_19[9:0]) begin
        image_1_461 <= io_pixelVal_in_1_1;
      end else if (10'h1cd == _T_15[9:0]) begin
        image_1_461 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_462 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ce == _T_37[9:0]) begin
        image_1_462 <= io_pixelVal_in_1_7;
      end else if (10'h1ce == _T_34[9:0]) begin
        image_1_462 <= io_pixelVal_in_1_6;
      end else if (10'h1ce == _T_31[9:0]) begin
        image_1_462 <= io_pixelVal_in_1_5;
      end else if (10'h1ce == _T_28[9:0]) begin
        image_1_462 <= io_pixelVal_in_1_4;
      end else if (10'h1ce == _T_25[9:0]) begin
        image_1_462 <= io_pixelVal_in_1_3;
      end else if (10'h1ce == _T_22[9:0]) begin
        image_1_462 <= io_pixelVal_in_1_2;
      end else if (10'h1ce == _T_19[9:0]) begin
        image_1_462 <= io_pixelVal_in_1_1;
      end else if (10'h1ce == _T_15[9:0]) begin
        image_1_462 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_463 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1cf == _T_37[9:0]) begin
        image_1_463 <= io_pixelVal_in_1_7;
      end else if (10'h1cf == _T_34[9:0]) begin
        image_1_463 <= io_pixelVal_in_1_6;
      end else if (10'h1cf == _T_31[9:0]) begin
        image_1_463 <= io_pixelVal_in_1_5;
      end else if (10'h1cf == _T_28[9:0]) begin
        image_1_463 <= io_pixelVal_in_1_4;
      end else if (10'h1cf == _T_25[9:0]) begin
        image_1_463 <= io_pixelVal_in_1_3;
      end else if (10'h1cf == _T_22[9:0]) begin
        image_1_463 <= io_pixelVal_in_1_2;
      end else if (10'h1cf == _T_19[9:0]) begin
        image_1_463 <= io_pixelVal_in_1_1;
      end else if (10'h1cf == _T_15[9:0]) begin
        image_1_463 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_464 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d0 == _T_37[9:0]) begin
        image_1_464 <= io_pixelVal_in_1_7;
      end else if (10'h1d0 == _T_34[9:0]) begin
        image_1_464 <= io_pixelVal_in_1_6;
      end else if (10'h1d0 == _T_31[9:0]) begin
        image_1_464 <= io_pixelVal_in_1_5;
      end else if (10'h1d0 == _T_28[9:0]) begin
        image_1_464 <= io_pixelVal_in_1_4;
      end else if (10'h1d0 == _T_25[9:0]) begin
        image_1_464 <= io_pixelVal_in_1_3;
      end else if (10'h1d0 == _T_22[9:0]) begin
        image_1_464 <= io_pixelVal_in_1_2;
      end else if (10'h1d0 == _T_19[9:0]) begin
        image_1_464 <= io_pixelVal_in_1_1;
      end else if (10'h1d0 == _T_15[9:0]) begin
        image_1_464 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_465 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d1 == _T_37[9:0]) begin
        image_1_465 <= io_pixelVal_in_1_7;
      end else if (10'h1d1 == _T_34[9:0]) begin
        image_1_465 <= io_pixelVal_in_1_6;
      end else if (10'h1d1 == _T_31[9:0]) begin
        image_1_465 <= io_pixelVal_in_1_5;
      end else if (10'h1d1 == _T_28[9:0]) begin
        image_1_465 <= io_pixelVal_in_1_4;
      end else if (10'h1d1 == _T_25[9:0]) begin
        image_1_465 <= io_pixelVal_in_1_3;
      end else if (10'h1d1 == _T_22[9:0]) begin
        image_1_465 <= io_pixelVal_in_1_2;
      end else if (10'h1d1 == _T_19[9:0]) begin
        image_1_465 <= io_pixelVal_in_1_1;
      end else if (10'h1d1 == _T_15[9:0]) begin
        image_1_465 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_466 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d2 == _T_37[9:0]) begin
        image_1_466 <= io_pixelVal_in_1_7;
      end else if (10'h1d2 == _T_34[9:0]) begin
        image_1_466 <= io_pixelVal_in_1_6;
      end else if (10'h1d2 == _T_31[9:0]) begin
        image_1_466 <= io_pixelVal_in_1_5;
      end else if (10'h1d2 == _T_28[9:0]) begin
        image_1_466 <= io_pixelVal_in_1_4;
      end else if (10'h1d2 == _T_25[9:0]) begin
        image_1_466 <= io_pixelVal_in_1_3;
      end else if (10'h1d2 == _T_22[9:0]) begin
        image_1_466 <= io_pixelVal_in_1_2;
      end else if (10'h1d2 == _T_19[9:0]) begin
        image_1_466 <= io_pixelVal_in_1_1;
      end else if (10'h1d2 == _T_15[9:0]) begin
        image_1_466 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_467 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d3 == _T_37[9:0]) begin
        image_1_467 <= io_pixelVal_in_1_7;
      end else if (10'h1d3 == _T_34[9:0]) begin
        image_1_467 <= io_pixelVal_in_1_6;
      end else if (10'h1d3 == _T_31[9:0]) begin
        image_1_467 <= io_pixelVal_in_1_5;
      end else if (10'h1d3 == _T_28[9:0]) begin
        image_1_467 <= io_pixelVal_in_1_4;
      end else if (10'h1d3 == _T_25[9:0]) begin
        image_1_467 <= io_pixelVal_in_1_3;
      end else if (10'h1d3 == _T_22[9:0]) begin
        image_1_467 <= io_pixelVal_in_1_2;
      end else if (10'h1d3 == _T_19[9:0]) begin
        image_1_467 <= io_pixelVal_in_1_1;
      end else if (10'h1d3 == _T_15[9:0]) begin
        image_1_467 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_468 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d4 == _T_37[9:0]) begin
        image_1_468 <= io_pixelVal_in_1_7;
      end else if (10'h1d4 == _T_34[9:0]) begin
        image_1_468 <= io_pixelVal_in_1_6;
      end else if (10'h1d4 == _T_31[9:0]) begin
        image_1_468 <= io_pixelVal_in_1_5;
      end else if (10'h1d4 == _T_28[9:0]) begin
        image_1_468 <= io_pixelVal_in_1_4;
      end else if (10'h1d4 == _T_25[9:0]) begin
        image_1_468 <= io_pixelVal_in_1_3;
      end else if (10'h1d4 == _T_22[9:0]) begin
        image_1_468 <= io_pixelVal_in_1_2;
      end else if (10'h1d4 == _T_19[9:0]) begin
        image_1_468 <= io_pixelVal_in_1_1;
      end else if (10'h1d4 == _T_15[9:0]) begin
        image_1_468 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_469 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d5 == _T_37[9:0]) begin
        image_1_469 <= io_pixelVal_in_1_7;
      end else if (10'h1d5 == _T_34[9:0]) begin
        image_1_469 <= io_pixelVal_in_1_6;
      end else if (10'h1d5 == _T_31[9:0]) begin
        image_1_469 <= io_pixelVal_in_1_5;
      end else if (10'h1d5 == _T_28[9:0]) begin
        image_1_469 <= io_pixelVal_in_1_4;
      end else if (10'h1d5 == _T_25[9:0]) begin
        image_1_469 <= io_pixelVal_in_1_3;
      end else if (10'h1d5 == _T_22[9:0]) begin
        image_1_469 <= io_pixelVal_in_1_2;
      end else if (10'h1d5 == _T_19[9:0]) begin
        image_1_469 <= io_pixelVal_in_1_1;
      end else if (10'h1d5 == _T_15[9:0]) begin
        image_1_469 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_470 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d6 == _T_37[9:0]) begin
        image_1_470 <= io_pixelVal_in_1_7;
      end else if (10'h1d6 == _T_34[9:0]) begin
        image_1_470 <= io_pixelVal_in_1_6;
      end else if (10'h1d6 == _T_31[9:0]) begin
        image_1_470 <= io_pixelVal_in_1_5;
      end else if (10'h1d6 == _T_28[9:0]) begin
        image_1_470 <= io_pixelVal_in_1_4;
      end else if (10'h1d6 == _T_25[9:0]) begin
        image_1_470 <= io_pixelVal_in_1_3;
      end else if (10'h1d6 == _T_22[9:0]) begin
        image_1_470 <= io_pixelVal_in_1_2;
      end else if (10'h1d6 == _T_19[9:0]) begin
        image_1_470 <= io_pixelVal_in_1_1;
      end else if (10'h1d6 == _T_15[9:0]) begin
        image_1_470 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_471 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d7 == _T_37[9:0]) begin
        image_1_471 <= io_pixelVal_in_1_7;
      end else if (10'h1d7 == _T_34[9:0]) begin
        image_1_471 <= io_pixelVal_in_1_6;
      end else if (10'h1d7 == _T_31[9:0]) begin
        image_1_471 <= io_pixelVal_in_1_5;
      end else if (10'h1d7 == _T_28[9:0]) begin
        image_1_471 <= io_pixelVal_in_1_4;
      end else if (10'h1d7 == _T_25[9:0]) begin
        image_1_471 <= io_pixelVal_in_1_3;
      end else if (10'h1d7 == _T_22[9:0]) begin
        image_1_471 <= io_pixelVal_in_1_2;
      end else if (10'h1d7 == _T_19[9:0]) begin
        image_1_471 <= io_pixelVal_in_1_1;
      end else if (10'h1d7 == _T_15[9:0]) begin
        image_1_471 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_472 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d8 == _T_37[9:0]) begin
        image_1_472 <= io_pixelVal_in_1_7;
      end else if (10'h1d8 == _T_34[9:0]) begin
        image_1_472 <= io_pixelVal_in_1_6;
      end else if (10'h1d8 == _T_31[9:0]) begin
        image_1_472 <= io_pixelVal_in_1_5;
      end else if (10'h1d8 == _T_28[9:0]) begin
        image_1_472 <= io_pixelVal_in_1_4;
      end else if (10'h1d8 == _T_25[9:0]) begin
        image_1_472 <= io_pixelVal_in_1_3;
      end else if (10'h1d8 == _T_22[9:0]) begin
        image_1_472 <= io_pixelVal_in_1_2;
      end else if (10'h1d8 == _T_19[9:0]) begin
        image_1_472 <= io_pixelVal_in_1_1;
      end else if (10'h1d8 == _T_15[9:0]) begin
        image_1_472 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_473 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d9 == _T_37[9:0]) begin
        image_1_473 <= io_pixelVal_in_1_7;
      end else if (10'h1d9 == _T_34[9:0]) begin
        image_1_473 <= io_pixelVal_in_1_6;
      end else if (10'h1d9 == _T_31[9:0]) begin
        image_1_473 <= io_pixelVal_in_1_5;
      end else if (10'h1d9 == _T_28[9:0]) begin
        image_1_473 <= io_pixelVal_in_1_4;
      end else if (10'h1d9 == _T_25[9:0]) begin
        image_1_473 <= io_pixelVal_in_1_3;
      end else if (10'h1d9 == _T_22[9:0]) begin
        image_1_473 <= io_pixelVal_in_1_2;
      end else if (10'h1d9 == _T_19[9:0]) begin
        image_1_473 <= io_pixelVal_in_1_1;
      end else if (10'h1d9 == _T_15[9:0]) begin
        image_1_473 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_474 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1da == _T_37[9:0]) begin
        image_1_474 <= io_pixelVal_in_1_7;
      end else if (10'h1da == _T_34[9:0]) begin
        image_1_474 <= io_pixelVal_in_1_6;
      end else if (10'h1da == _T_31[9:0]) begin
        image_1_474 <= io_pixelVal_in_1_5;
      end else if (10'h1da == _T_28[9:0]) begin
        image_1_474 <= io_pixelVal_in_1_4;
      end else if (10'h1da == _T_25[9:0]) begin
        image_1_474 <= io_pixelVal_in_1_3;
      end else if (10'h1da == _T_22[9:0]) begin
        image_1_474 <= io_pixelVal_in_1_2;
      end else if (10'h1da == _T_19[9:0]) begin
        image_1_474 <= io_pixelVal_in_1_1;
      end else if (10'h1da == _T_15[9:0]) begin
        image_1_474 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_475 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1db == _T_37[9:0]) begin
        image_1_475 <= io_pixelVal_in_1_7;
      end else if (10'h1db == _T_34[9:0]) begin
        image_1_475 <= io_pixelVal_in_1_6;
      end else if (10'h1db == _T_31[9:0]) begin
        image_1_475 <= io_pixelVal_in_1_5;
      end else if (10'h1db == _T_28[9:0]) begin
        image_1_475 <= io_pixelVal_in_1_4;
      end else if (10'h1db == _T_25[9:0]) begin
        image_1_475 <= io_pixelVal_in_1_3;
      end else if (10'h1db == _T_22[9:0]) begin
        image_1_475 <= io_pixelVal_in_1_2;
      end else if (10'h1db == _T_19[9:0]) begin
        image_1_475 <= io_pixelVal_in_1_1;
      end else if (10'h1db == _T_15[9:0]) begin
        image_1_475 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_476 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1dc == _T_37[9:0]) begin
        image_1_476 <= io_pixelVal_in_1_7;
      end else if (10'h1dc == _T_34[9:0]) begin
        image_1_476 <= io_pixelVal_in_1_6;
      end else if (10'h1dc == _T_31[9:0]) begin
        image_1_476 <= io_pixelVal_in_1_5;
      end else if (10'h1dc == _T_28[9:0]) begin
        image_1_476 <= io_pixelVal_in_1_4;
      end else if (10'h1dc == _T_25[9:0]) begin
        image_1_476 <= io_pixelVal_in_1_3;
      end else if (10'h1dc == _T_22[9:0]) begin
        image_1_476 <= io_pixelVal_in_1_2;
      end else if (10'h1dc == _T_19[9:0]) begin
        image_1_476 <= io_pixelVal_in_1_1;
      end else if (10'h1dc == _T_15[9:0]) begin
        image_1_476 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_477 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1dd == _T_37[9:0]) begin
        image_1_477 <= io_pixelVal_in_1_7;
      end else if (10'h1dd == _T_34[9:0]) begin
        image_1_477 <= io_pixelVal_in_1_6;
      end else if (10'h1dd == _T_31[9:0]) begin
        image_1_477 <= io_pixelVal_in_1_5;
      end else if (10'h1dd == _T_28[9:0]) begin
        image_1_477 <= io_pixelVal_in_1_4;
      end else if (10'h1dd == _T_25[9:0]) begin
        image_1_477 <= io_pixelVal_in_1_3;
      end else if (10'h1dd == _T_22[9:0]) begin
        image_1_477 <= io_pixelVal_in_1_2;
      end else if (10'h1dd == _T_19[9:0]) begin
        image_1_477 <= io_pixelVal_in_1_1;
      end else if (10'h1dd == _T_15[9:0]) begin
        image_1_477 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_478 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1de == _T_37[9:0]) begin
        image_1_478 <= io_pixelVal_in_1_7;
      end else if (10'h1de == _T_34[9:0]) begin
        image_1_478 <= io_pixelVal_in_1_6;
      end else if (10'h1de == _T_31[9:0]) begin
        image_1_478 <= io_pixelVal_in_1_5;
      end else if (10'h1de == _T_28[9:0]) begin
        image_1_478 <= io_pixelVal_in_1_4;
      end else if (10'h1de == _T_25[9:0]) begin
        image_1_478 <= io_pixelVal_in_1_3;
      end else if (10'h1de == _T_22[9:0]) begin
        image_1_478 <= io_pixelVal_in_1_2;
      end else if (10'h1de == _T_19[9:0]) begin
        image_1_478 <= io_pixelVal_in_1_1;
      end else if (10'h1de == _T_15[9:0]) begin
        image_1_478 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_479 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1df == _T_37[9:0]) begin
        image_1_479 <= io_pixelVal_in_1_7;
      end else if (10'h1df == _T_34[9:0]) begin
        image_1_479 <= io_pixelVal_in_1_6;
      end else if (10'h1df == _T_31[9:0]) begin
        image_1_479 <= io_pixelVal_in_1_5;
      end else if (10'h1df == _T_28[9:0]) begin
        image_1_479 <= io_pixelVal_in_1_4;
      end else if (10'h1df == _T_25[9:0]) begin
        image_1_479 <= io_pixelVal_in_1_3;
      end else if (10'h1df == _T_22[9:0]) begin
        image_1_479 <= io_pixelVal_in_1_2;
      end else if (10'h1df == _T_19[9:0]) begin
        image_1_479 <= io_pixelVal_in_1_1;
      end else if (10'h1df == _T_15[9:0]) begin
        image_1_479 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_480 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e0 == _T_37[9:0]) begin
        image_1_480 <= io_pixelVal_in_1_7;
      end else if (10'h1e0 == _T_34[9:0]) begin
        image_1_480 <= io_pixelVal_in_1_6;
      end else if (10'h1e0 == _T_31[9:0]) begin
        image_1_480 <= io_pixelVal_in_1_5;
      end else if (10'h1e0 == _T_28[9:0]) begin
        image_1_480 <= io_pixelVal_in_1_4;
      end else if (10'h1e0 == _T_25[9:0]) begin
        image_1_480 <= io_pixelVal_in_1_3;
      end else if (10'h1e0 == _T_22[9:0]) begin
        image_1_480 <= io_pixelVal_in_1_2;
      end else if (10'h1e0 == _T_19[9:0]) begin
        image_1_480 <= io_pixelVal_in_1_1;
      end else if (10'h1e0 == _T_15[9:0]) begin
        image_1_480 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_481 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e1 == _T_37[9:0]) begin
        image_1_481 <= io_pixelVal_in_1_7;
      end else if (10'h1e1 == _T_34[9:0]) begin
        image_1_481 <= io_pixelVal_in_1_6;
      end else if (10'h1e1 == _T_31[9:0]) begin
        image_1_481 <= io_pixelVal_in_1_5;
      end else if (10'h1e1 == _T_28[9:0]) begin
        image_1_481 <= io_pixelVal_in_1_4;
      end else if (10'h1e1 == _T_25[9:0]) begin
        image_1_481 <= io_pixelVal_in_1_3;
      end else if (10'h1e1 == _T_22[9:0]) begin
        image_1_481 <= io_pixelVal_in_1_2;
      end else if (10'h1e1 == _T_19[9:0]) begin
        image_1_481 <= io_pixelVal_in_1_1;
      end else if (10'h1e1 == _T_15[9:0]) begin
        image_1_481 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_482 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e2 == _T_37[9:0]) begin
        image_1_482 <= io_pixelVal_in_1_7;
      end else if (10'h1e2 == _T_34[9:0]) begin
        image_1_482 <= io_pixelVal_in_1_6;
      end else if (10'h1e2 == _T_31[9:0]) begin
        image_1_482 <= io_pixelVal_in_1_5;
      end else if (10'h1e2 == _T_28[9:0]) begin
        image_1_482 <= io_pixelVal_in_1_4;
      end else if (10'h1e2 == _T_25[9:0]) begin
        image_1_482 <= io_pixelVal_in_1_3;
      end else if (10'h1e2 == _T_22[9:0]) begin
        image_1_482 <= io_pixelVal_in_1_2;
      end else if (10'h1e2 == _T_19[9:0]) begin
        image_1_482 <= io_pixelVal_in_1_1;
      end else if (10'h1e2 == _T_15[9:0]) begin
        image_1_482 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_483 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e3 == _T_37[9:0]) begin
        image_1_483 <= io_pixelVal_in_1_7;
      end else if (10'h1e3 == _T_34[9:0]) begin
        image_1_483 <= io_pixelVal_in_1_6;
      end else if (10'h1e3 == _T_31[9:0]) begin
        image_1_483 <= io_pixelVal_in_1_5;
      end else if (10'h1e3 == _T_28[9:0]) begin
        image_1_483 <= io_pixelVal_in_1_4;
      end else if (10'h1e3 == _T_25[9:0]) begin
        image_1_483 <= io_pixelVal_in_1_3;
      end else if (10'h1e3 == _T_22[9:0]) begin
        image_1_483 <= io_pixelVal_in_1_2;
      end else if (10'h1e3 == _T_19[9:0]) begin
        image_1_483 <= io_pixelVal_in_1_1;
      end else if (10'h1e3 == _T_15[9:0]) begin
        image_1_483 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_484 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e4 == _T_37[9:0]) begin
        image_1_484 <= io_pixelVal_in_1_7;
      end else if (10'h1e4 == _T_34[9:0]) begin
        image_1_484 <= io_pixelVal_in_1_6;
      end else if (10'h1e4 == _T_31[9:0]) begin
        image_1_484 <= io_pixelVal_in_1_5;
      end else if (10'h1e4 == _T_28[9:0]) begin
        image_1_484 <= io_pixelVal_in_1_4;
      end else if (10'h1e4 == _T_25[9:0]) begin
        image_1_484 <= io_pixelVal_in_1_3;
      end else if (10'h1e4 == _T_22[9:0]) begin
        image_1_484 <= io_pixelVal_in_1_2;
      end else if (10'h1e4 == _T_19[9:0]) begin
        image_1_484 <= io_pixelVal_in_1_1;
      end else if (10'h1e4 == _T_15[9:0]) begin
        image_1_484 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_485 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e5 == _T_37[9:0]) begin
        image_1_485 <= io_pixelVal_in_1_7;
      end else if (10'h1e5 == _T_34[9:0]) begin
        image_1_485 <= io_pixelVal_in_1_6;
      end else if (10'h1e5 == _T_31[9:0]) begin
        image_1_485 <= io_pixelVal_in_1_5;
      end else if (10'h1e5 == _T_28[9:0]) begin
        image_1_485 <= io_pixelVal_in_1_4;
      end else if (10'h1e5 == _T_25[9:0]) begin
        image_1_485 <= io_pixelVal_in_1_3;
      end else if (10'h1e5 == _T_22[9:0]) begin
        image_1_485 <= io_pixelVal_in_1_2;
      end else if (10'h1e5 == _T_19[9:0]) begin
        image_1_485 <= io_pixelVal_in_1_1;
      end else if (10'h1e5 == _T_15[9:0]) begin
        image_1_485 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_486 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e6 == _T_37[9:0]) begin
        image_1_486 <= io_pixelVal_in_1_7;
      end else if (10'h1e6 == _T_34[9:0]) begin
        image_1_486 <= io_pixelVal_in_1_6;
      end else if (10'h1e6 == _T_31[9:0]) begin
        image_1_486 <= io_pixelVal_in_1_5;
      end else if (10'h1e6 == _T_28[9:0]) begin
        image_1_486 <= io_pixelVal_in_1_4;
      end else if (10'h1e6 == _T_25[9:0]) begin
        image_1_486 <= io_pixelVal_in_1_3;
      end else if (10'h1e6 == _T_22[9:0]) begin
        image_1_486 <= io_pixelVal_in_1_2;
      end else if (10'h1e6 == _T_19[9:0]) begin
        image_1_486 <= io_pixelVal_in_1_1;
      end else if (10'h1e6 == _T_15[9:0]) begin
        image_1_486 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_487 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e7 == _T_37[9:0]) begin
        image_1_487 <= io_pixelVal_in_1_7;
      end else if (10'h1e7 == _T_34[9:0]) begin
        image_1_487 <= io_pixelVal_in_1_6;
      end else if (10'h1e7 == _T_31[9:0]) begin
        image_1_487 <= io_pixelVal_in_1_5;
      end else if (10'h1e7 == _T_28[9:0]) begin
        image_1_487 <= io_pixelVal_in_1_4;
      end else if (10'h1e7 == _T_25[9:0]) begin
        image_1_487 <= io_pixelVal_in_1_3;
      end else if (10'h1e7 == _T_22[9:0]) begin
        image_1_487 <= io_pixelVal_in_1_2;
      end else if (10'h1e7 == _T_19[9:0]) begin
        image_1_487 <= io_pixelVal_in_1_1;
      end else if (10'h1e7 == _T_15[9:0]) begin
        image_1_487 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_488 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e8 == _T_37[9:0]) begin
        image_1_488 <= io_pixelVal_in_1_7;
      end else if (10'h1e8 == _T_34[9:0]) begin
        image_1_488 <= io_pixelVal_in_1_6;
      end else if (10'h1e8 == _T_31[9:0]) begin
        image_1_488 <= io_pixelVal_in_1_5;
      end else if (10'h1e8 == _T_28[9:0]) begin
        image_1_488 <= io_pixelVal_in_1_4;
      end else if (10'h1e8 == _T_25[9:0]) begin
        image_1_488 <= io_pixelVal_in_1_3;
      end else if (10'h1e8 == _T_22[9:0]) begin
        image_1_488 <= io_pixelVal_in_1_2;
      end else if (10'h1e8 == _T_19[9:0]) begin
        image_1_488 <= io_pixelVal_in_1_1;
      end else if (10'h1e8 == _T_15[9:0]) begin
        image_1_488 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_489 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e9 == _T_37[9:0]) begin
        image_1_489 <= io_pixelVal_in_1_7;
      end else if (10'h1e9 == _T_34[9:0]) begin
        image_1_489 <= io_pixelVal_in_1_6;
      end else if (10'h1e9 == _T_31[9:0]) begin
        image_1_489 <= io_pixelVal_in_1_5;
      end else if (10'h1e9 == _T_28[9:0]) begin
        image_1_489 <= io_pixelVal_in_1_4;
      end else if (10'h1e9 == _T_25[9:0]) begin
        image_1_489 <= io_pixelVal_in_1_3;
      end else if (10'h1e9 == _T_22[9:0]) begin
        image_1_489 <= io_pixelVal_in_1_2;
      end else if (10'h1e9 == _T_19[9:0]) begin
        image_1_489 <= io_pixelVal_in_1_1;
      end else if (10'h1e9 == _T_15[9:0]) begin
        image_1_489 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_490 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ea == _T_37[9:0]) begin
        image_1_490 <= io_pixelVal_in_1_7;
      end else if (10'h1ea == _T_34[9:0]) begin
        image_1_490 <= io_pixelVal_in_1_6;
      end else if (10'h1ea == _T_31[9:0]) begin
        image_1_490 <= io_pixelVal_in_1_5;
      end else if (10'h1ea == _T_28[9:0]) begin
        image_1_490 <= io_pixelVal_in_1_4;
      end else if (10'h1ea == _T_25[9:0]) begin
        image_1_490 <= io_pixelVal_in_1_3;
      end else if (10'h1ea == _T_22[9:0]) begin
        image_1_490 <= io_pixelVal_in_1_2;
      end else if (10'h1ea == _T_19[9:0]) begin
        image_1_490 <= io_pixelVal_in_1_1;
      end else if (10'h1ea == _T_15[9:0]) begin
        image_1_490 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_491 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1eb == _T_37[9:0]) begin
        image_1_491 <= io_pixelVal_in_1_7;
      end else if (10'h1eb == _T_34[9:0]) begin
        image_1_491 <= io_pixelVal_in_1_6;
      end else if (10'h1eb == _T_31[9:0]) begin
        image_1_491 <= io_pixelVal_in_1_5;
      end else if (10'h1eb == _T_28[9:0]) begin
        image_1_491 <= io_pixelVal_in_1_4;
      end else if (10'h1eb == _T_25[9:0]) begin
        image_1_491 <= io_pixelVal_in_1_3;
      end else if (10'h1eb == _T_22[9:0]) begin
        image_1_491 <= io_pixelVal_in_1_2;
      end else if (10'h1eb == _T_19[9:0]) begin
        image_1_491 <= io_pixelVal_in_1_1;
      end else if (10'h1eb == _T_15[9:0]) begin
        image_1_491 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_492 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ec == _T_37[9:0]) begin
        image_1_492 <= io_pixelVal_in_1_7;
      end else if (10'h1ec == _T_34[9:0]) begin
        image_1_492 <= io_pixelVal_in_1_6;
      end else if (10'h1ec == _T_31[9:0]) begin
        image_1_492 <= io_pixelVal_in_1_5;
      end else if (10'h1ec == _T_28[9:0]) begin
        image_1_492 <= io_pixelVal_in_1_4;
      end else if (10'h1ec == _T_25[9:0]) begin
        image_1_492 <= io_pixelVal_in_1_3;
      end else if (10'h1ec == _T_22[9:0]) begin
        image_1_492 <= io_pixelVal_in_1_2;
      end else if (10'h1ec == _T_19[9:0]) begin
        image_1_492 <= io_pixelVal_in_1_1;
      end else if (10'h1ec == _T_15[9:0]) begin
        image_1_492 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_493 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ed == _T_37[9:0]) begin
        image_1_493 <= io_pixelVal_in_1_7;
      end else if (10'h1ed == _T_34[9:0]) begin
        image_1_493 <= io_pixelVal_in_1_6;
      end else if (10'h1ed == _T_31[9:0]) begin
        image_1_493 <= io_pixelVal_in_1_5;
      end else if (10'h1ed == _T_28[9:0]) begin
        image_1_493 <= io_pixelVal_in_1_4;
      end else if (10'h1ed == _T_25[9:0]) begin
        image_1_493 <= io_pixelVal_in_1_3;
      end else if (10'h1ed == _T_22[9:0]) begin
        image_1_493 <= io_pixelVal_in_1_2;
      end else if (10'h1ed == _T_19[9:0]) begin
        image_1_493 <= io_pixelVal_in_1_1;
      end else if (10'h1ed == _T_15[9:0]) begin
        image_1_493 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_494 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ee == _T_37[9:0]) begin
        image_1_494 <= io_pixelVal_in_1_7;
      end else if (10'h1ee == _T_34[9:0]) begin
        image_1_494 <= io_pixelVal_in_1_6;
      end else if (10'h1ee == _T_31[9:0]) begin
        image_1_494 <= io_pixelVal_in_1_5;
      end else if (10'h1ee == _T_28[9:0]) begin
        image_1_494 <= io_pixelVal_in_1_4;
      end else if (10'h1ee == _T_25[9:0]) begin
        image_1_494 <= io_pixelVal_in_1_3;
      end else if (10'h1ee == _T_22[9:0]) begin
        image_1_494 <= io_pixelVal_in_1_2;
      end else if (10'h1ee == _T_19[9:0]) begin
        image_1_494 <= io_pixelVal_in_1_1;
      end else if (10'h1ee == _T_15[9:0]) begin
        image_1_494 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_495 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ef == _T_37[9:0]) begin
        image_1_495 <= io_pixelVal_in_1_7;
      end else if (10'h1ef == _T_34[9:0]) begin
        image_1_495 <= io_pixelVal_in_1_6;
      end else if (10'h1ef == _T_31[9:0]) begin
        image_1_495 <= io_pixelVal_in_1_5;
      end else if (10'h1ef == _T_28[9:0]) begin
        image_1_495 <= io_pixelVal_in_1_4;
      end else if (10'h1ef == _T_25[9:0]) begin
        image_1_495 <= io_pixelVal_in_1_3;
      end else if (10'h1ef == _T_22[9:0]) begin
        image_1_495 <= io_pixelVal_in_1_2;
      end else if (10'h1ef == _T_19[9:0]) begin
        image_1_495 <= io_pixelVal_in_1_1;
      end else if (10'h1ef == _T_15[9:0]) begin
        image_1_495 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_496 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f0 == _T_37[9:0]) begin
        image_1_496 <= io_pixelVal_in_1_7;
      end else if (10'h1f0 == _T_34[9:0]) begin
        image_1_496 <= io_pixelVal_in_1_6;
      end else if (10'h1f0 == _T_31[9:0]) begin
        image_1_496 <= io_pixelVal_in_1_5;
      end else if (10'h1f0 == _T_28[9:0]) begin
        image_1_496 <= io_pixelVal_in_1_4;
      end else if (10'h1f0 == _T_25[9:0]) begin
        image_1_496 <= io_pixelVal_in_1_3;
      end else if (10'h1f0 == _T_22[9:0]) begin
        image_1_496 <= io_pixelVal_in_1_2;
      end else if (10'h1f0 == _T_19[9:0]) begin
        image_1_496 <= io_pixelVal_in_1_1;
      end else if (10'h1f0 == _T_15[9:0]) begin
        image_1_496 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_497 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f1 == _T_37[9:0]) begin
        image_1_497 <= io_pixelVal_in_1_7;
      end else if (10'h1f1 == _T_34[9:0]) begin
        image_1_497 <= io_pixelVal_in_1_6;
      end else if (10'h1f1 == _T_31[9:0]) begin
        image_1_497 <= io_pixelVal_in_1_5;
      end else if (10'h1f1 == _T_28[9:0]) begin
        image_1_497 <= io_pixelVal_in_1_4;
      end else if (10'h1f1 == _T_25[9:0]) begin
        image_1_497 <= io_pixelVal_in_1_3;
      end else if (10'h1f1 == _T_22[9:0]) begin
        image_1_497 <= io_pixelVal_in_1_2;
      end else if (10'h1f1 == _T_19[9:0]) begin
        image_1_497 <= io_pixelVal_in_1_1;
      end else if (10'h1f1 == _T_15[9:0]) begin
        image_1_497 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_498 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f2 == _T_37[9:0]) begin
        image_1_498 <= io_pixelVal_in_1_7;
      end else if (10'h1f2 == _T_34[9:0]) begin
        image_1_498 <= io_pixelVal_in_1_6;
      end else if (10'h1f2 == _T_31[9:0]) begin
        image_1_498 <= io_pixelVal_in_1_5;
      end else if (10'h1f2 == _T_28[9:0]) begin
        image_1_498 <= io_pixelVal_in_1_4;
      end else if (10'h1f2 == _T_25[9:0]) begin
        image_1_498 <= io_pixelVal_in_1_3;
      end else if (10'h1f2 == _T_22[9:0]) begin
        image_1_498 <= io_pixelVal_in_1_2;
      end else if (10'h1f2 == _T_19[9:0]) begin
        image_1_498 <= io_pixelVal_in_1_1;
      end else if (10'h1f2 == _T_15[9:0]) begin
        image_1_498 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_499 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f3 == _T_37[9:0]) begin
        image_1_499 <= io_pixelVal_in_1_7;
      end else if (10'h1f3 == _T_34[9:0]) begin
        image_1_499 <= io_pixelVal_in_1_6;
      end else if (10'h1f3 == _T_31[9:0]) begin
        image_1_499 <= io_pixelVal_in_1_5;
      end else if (10'h1f3 == _T_28[9:0]) begin
        image_1_499 <= io_pixelVal_in_1_4;
      end else if (10'h1f3 == _T_25[9:0]) begin
        image_1_499 <= io_pixelVal_in_1_3;
      end else if (10'h1f3 == _T_22[9:0]) begin
        image_1_499 <= io_pixelVal_in_1_2;
      end else if (10'h1f3 == _T_19[9:0]) begin
        image_1_499 <= io_pixelVal_in_1_1;
      end else if (10'h1f3 == _T_15[9:0]) begin
        image_1_499 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_500 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f4 == _T_37[9:0]) begin
        image_1_500 <= io_pixelVal_in_1_7;
      end else if (10'h1f4 == _T_34[9:0]) begin
        image_1_500 <= io_pixelVal_in_1_6;
      end else if (10'h1f4 == _T_31[9:0]) begin
        image_1_500 <= io_pixelVal_in_1_5;
      end else if (10'h1f4 == _T_28[9:0]) begin
        image_1_500 <= io_pixelVal_in_1_4;
      end else if (10'h1f4 == _T_25[9:0]) begin
        image_1_500 <= io_pixelVal_in_1_3;
      end else if (10'h1f4 == _T_22[9:0]) begin
        image_1_500 <= io_pixelVal_in_1_2;
      end else if (10'h1f4 == _T_19[9:0]) begin
        image_1_500 <= io_pixelVal_in_1_1;
      end else if (10'h1f4 == _T_15[9:0]) begin
        image_1_500 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_501 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f5 == _T_37[9:0]) begin
        image_1_501 <= io_pixelVal_in_1_7;
      end else if (10'h1f5 == _T_34[9:0]) begin
        image_1_501 <= io_pixelVal_in_1_6;
      end else if (10'h1f5 == _T_31[9:0]) begin
        image_1_501 <= io_pixelVal_in_1_5;
      end else if (10'h1f5 == _T_28[9:0]) begin
        image_1_501 <= io_pixelVal_in_1_4;
      end else if (10'h1f5 == _T_25[9:0]) begin
        image_1_501 <= io_pixelVal_in_1_3;
      end else if (10'h1f5 == _T_22[9:0]) begin
        image_1_501 <= io_pixelVal_in_1_2;
      end else if (10'h1f5 == _T_19[9:0]) begin
        image_1_501 <= io_pixelVal_in_1_1;
      end else if (10'h1f5 == _T_15[9:0]) begin
        image_1_501 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_502 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f6 == _T_37[9:0]) begin
        image_1_502 <= io_pixelVal_in_1_7;
      end else if (10'h1f6 == _T_34[9:0]) begin
        image_1_502 <= io_pixelVal_in_1_6;
      end else if (10'h1f6 == _T_31[9:0]) begin
        image_1_502 <= io_pixelVal_in_1_5;
      end else if (10'h1f6 == _T_28[9:0]) begin
        image_1_502 <= io_pixelVal_in_1_4;
      end else if (10'h1f6 == _T_25[9:0]) begin
        image_1_502 <= io_pixelVal_in_1_3;
      end else if (10'h1f6 == _T_22[9:0]) begin
        image_1_502 <= io_pixelVal_in_1_2;
      end else if (10'h1f6 == _T_19[9:0]) begin
        image_1_502 <= io_pixelVal_in_1_1;
      end else if (10'h1f6 == _T_15[9:0]) begin
        image_1_502 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_503 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f7 == _T_37[9:0]) begin
        image_1_503 <= io_pixelVal_in_1_7;
      end else if (10'h1f7 == _T_34[9:0]) begin
        image_1_503 <= io_pixelVal_in_1_6;
      end else if (10'h1f7 == _T_31[9:0]) begin
        image_1_503 <= io_pixelVal_in_1_5;
      end else if (10'h1f7 == _T_28[9:0]) begin
        image_1_503 <= io_pixelVal_in_1_4;
      end else if (10'h1f7 == _T_25[9:0]) begin
        image_1_503 <= io_pixelVal_in_1_3;
      end else if (10'h1f7 == _T_22[9:0]) begin
        image_1_503 <= io_pixelVal_in_1_2;
      end else if (10'h1f7 == _T_19[9:0]) begin
        image_1_503 <= io_pixelVal_in_1_1;
      end else if (10'h1f7 == _T_15[9:0]) begin
        image_1_503 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_504 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f8 == _T_37[9:0]) begin
        image_1_504 <= io_pixelVal_in_1_7;
      end else if (10'h1f8 == _T_34[9:0]) begin
        image_1_504 <= io_pixelVal_in_1_6;
      end else if (10'h1f8 == _T_31[9:0]) begin
        image_1_504 <= io_pixelVal_in_1_5;
      end else if (10'h1f8 == _T_28[9:0]) begin
        image_1_504 <= io_pixelVal_in_1_4;
      end else if (10'h1f8 == _T_25[9:0]) begin
        image_1_504 <= io_pixelVal_in_1_3;
      end else if (10'h1f8 == _T_22[9:0]) begin
        image_1_504 <= io_pixelVal_in_1_2;
      end else if (10'h1f8 == _T_19[9:0]) begin
        image_1_504 <= io_pixelVal_in_1_1;
      end else if (10'h1f8 == _T_15[9:0]) begin
        image_1_504 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_505 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f9 == _T_37[9:0]) begin
        image_1_505 <= io_pixelVal_in_1_7;
      end else if (10'h1f9 == _T_34[9:0]) begin
        image_1_505 <= io_pixelVal_in_1_6;
      end else if (10'h1f9 == _T_31[9:0]) begin
        image_1_505 <= io_pixelVal_in_1_5;
      end else if (10'h1f9 == _T_28[9:0]) begin
        image_1_505 <= io_pixelVal_in_1_4;
      end else if (10'h1f9 == _T_25[9:0]) begin
        image_1_505 <= io_pixelVal_in_1_3;
      end else if (10'h1f9 == _T_22[9:0]) begin
        image_1_505 <= io_pixelVal_in_1_2;
      end else if (10'h1f9 == _T_19[9:0]) begin
        image_1_505 <= io_pixelVal_in_1_1;
      end else if (10'h1f9 == _T_15[9:0]) begin
        image_1_505 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_506 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1fa == _T_37[9:0]) begin
        image_1_506 <= io_pixelVal_in_1_7;
      end else if (10'h1fa == _T_34[9:0]) begin
        image_1_506 <= io_pixelVal_in_1_6;
      end else if (10'h1fa == _T_31[9:0]) begin
        image_1_506 <= io_pixelVal_in_1_5;
      end else if (10'h1fa == _T_28[9:0]) begin
        image_1_506 <= io_pixelVal_in_1_4;
      end else if (10'h1fa == _T_25[9:0]) begin
        image_1_506 <= io_pixelVal_in_1_3;
      end else if (10'h1fa == _T_22[9:0]) begin
        image_1_506 <= io_pixelVal_in_1_2;
      end else if (10'h1fa == _T_19[9:0]) begin
        image_1_506 <= io_pixelVal_in_1_1;
      end else if (10'h1fa == _T_15[9:0]) begin
        image_1_506 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_507 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1fb == _T_37[9:0]) begin
        image_1_507 <= io_pixelVal_in_1_7;
      end else if (10'h1fb == _T_34[9:0]) begin
        image_1_507 <= io_pixelVal_in_1_6;
      end else if (10'h1fb == _T_31[9:0]) begin
        image_1_507 <= io_pixelVal_in_1_5;
      end else if (10'h1fb == _T_28[9:0]) begin
        image_1_507 <= io_pixelVal_in_1_4;
      end else if (10'h1fb == _T_25[9:0]) begin
        image_1_507 <= io_pixelVal_in_1_3;
      end else if (10'h1fb == _T_22[9:0]) begin
        image_1_507 <= io_pixelVal_in_1_2;
      end else if (10'h1fb == _T_19[9:0]) begin
        image_1_507 <= io_pixelVal_in_1_1;
      end else if (10'h1fb == _T_15[9:0]) begin
        image_1_507 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_508 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1fc == _T_37[9:0]) begin
        image_1_508 <= io_pixelVal_in_1_7;
      end else if (10'h1fc == _T_34[9:0]) begin
        image_1_508 <= io_pixelVal_in_1_6;
      end else if (10'h1fc == _T_31[9:0]) begin
        image_1_508 <= io_pixelVal_in_1_5;
      end else if (10'h1fc == _T_28[9:0]) begin
        image_1_508 <= io_pixelVal_in_1_4;
      end else if (10'h1fc == _T_25[9:0]) begin
        image_1_508 <= io_pixelVal_in_1_3;
      end else if (10'h1fc == _T_22[9:0]) begin
        image_1_508 <= io_pixelVal_in_1_2;
      end else if (10'h1fc == _T_19[9:0]) begin
        image_1_508 <= io_pixelVal_in_1_1;
      end else if (10'h1fc == _T_15[9:0]) begin
        image_1_508 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_509 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1fd == _T_37[9:0]) begin
        image_1_509 <= io_pixelVal_in_1_7;
      end else if (10'h1fd == _T_34[9:0]) begin
        image_1_509 <= io_pixelVal_in_1_6;
      end else if (10'h1fd == _T_31[9:0]) begin
        image_1_509 <= io_pixelVal_in_1_5;
      end else if (10'h1fd == _T_28[9:0]) begin
        image_1_509 <= io_pixelVal_in_1_4;
      end else if (10'h1fd == _T_25[9:0]) begin
        image_1_509 <= io_pixelVal_in_1_3;
      end else if (10'h1fd == _T_22[9:0]) begin
        image_1_509 <= io_pixelVal_in_1_2;
      end else if (10'h1fd == _T_19[9:0]) begin
        image_1_509 <= io_pixelVal_in_1_1;
      end else if (10'h1fd == _T_15[9:0]) begin
        image_1_509 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_510 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1fe == _T_37[9:0]) begin
        image_1_510 <= io_pixelVal_in_1_7;
      end else if (10'h1fe == _T_34[9:0]) begin
        image_1_510 <= io_pixelVal_in_1_6;
      end else if (10'h1fe == _T_31[9:0]) begin
        image_1_510 <= io_pixelVal_in_1_5;
      end else if (10'h1fe == _T_28[9:0]) begin
        image_1_510 <= io_pixelVal_in_1_4;
      end else if (10'h1fe == _T_25[9:0]) begin
        image_1_510 <= io_pixelVal_in_1_3;
      end else if (10'h1fe == _T_22[9:0]) begin
        image_1_510 <= io_pixelVal_in_1_2;
      end else if (10'h1fe == _T_19[9:0]) begin
        image_1_510 <= io_pixelVal_in_1_1;
      end else if (10'h1fe == _T_15[9:0]) begin
        image_1_510 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_511 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ff == _T_37[9:0]) begin
        image_1_511 <= io_pixelVal_in_1_7;
      end else if (10'h1ff == _T_34[9:0]) begin
        image_1_511 <= io_pixelVal_in_1_6;
      end else if (10'h1ff == _T_31[9:0]) begin
        image_1_511 <= io_pixelVal_in_1_5;
      end else if (10'h1ff == _T_28[9:0]) begin
        image_1_511 <= io_pixelVal_in_1_4;
      end else if (10'h1ff == _T_25[9:0]) begin
        image_1_511 <= io_pixelVal_in_1_3;
      end else if (10'h1ff == _T_22[9:0]) begin
        image_1_511 <= io_pixelVal_in_1_2;
      end else if (10'h1ff == _T_19[9:0]) begin
        image_1_511 <= io_pixelVal_in_1_1;
      end else if (10'h1ff == _T_15[9:0]) begin
        image_1_511 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_512 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h200 == _T_37[9:0]) begin
        image_1_512 <= io_pixelVal_in_1_7;
      end else if (10'h200 == _T_34[9:0]) begin
        image_1_512 <= io_pixelVal_in_1_6;
      end else if (10'h200 == _T_31[9:0]) begin
        image_1_512 <= io_pixelVal_in_1_5;
      end else if (10'h200 == _T_28[9:0]) begin
        image_1_512 <= io_pixelVal_in_1_4;
      end else if (10'h200 == _T_25[9:0]) begin
        image_1_512 <= io_pixelVal_in_1_3;
      end else if (10'h200 == _T_22[9:0]) begin
        image_1_512 <= io_pixelVal_in_1_2;
      end else if (10'h200 == _T_19[9:0]) begin
        image_1_512 <= io_pixelVal_in_1_1;
      end else if (10'h200 == _T_15[9:0]) begin
        image_1_512 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_513 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h201 == _T_37[9:0]) begin
        image_1_513 <= io_pixelVal_in_1_7;
      end else if (10'h201 == _T_34[9:0]) begin
        image_1_513 <= io_pixelVal_in_1_6;
      end else if (10'h201 == _T_31[9:0]) begin
        image_1_513 <= io_pixelVal_in_1_5;
      end else if (10'h201 == _T_28[9:0]) begin
        image_1_513 <= io_pixelVal_in_1_4;
      end else if (10'h201 == _T_25[9:0]) begin
        image_1_513 <= io_pixelVal_in_1_3;
      end else if (10'h201 == _T_22[9:0]) begin
        image_1_513 <= io_pixelVal_in_1_2;
      end else if (10'h201 == _T_19[9:0]) begin
        image_1_513 <= io_pixelVal_in_1_1;
      end else if (10'h201 == _T_15[9:0]) begin
        image_1_513 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_514 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h202 == _T_37[9:0]) begin
        image_1_514 <= io_pixelVal_in_1_7;
      end else if (10'h202 == _T_34[9:0]) begin
        image_1_514 <= io_pixelVal_in_1_6;
      end else if (10'h202 == _T_31[9:0]) begin
        image_1_514 <= io_pixelVal_in_1_5;
      end else if (10'h202 == _T_28[9:0]) begin
        image_1_514 <= io_pixelVal_in_1_4;
      end else if (10'h202 == _T_25[9:0]) begin
        image_1_514 <= io_pixelVal_in_1_3;
      end else if (10'h202 == _T_22[9:0]) begin
        image_1_514 <= io_pixelVal_in_1_2;
      end else if (10'h202 == _T_19[9:0]) begin
        image_1_514 <= io_pixelVal_in_1_1;
      end else if (10'h202 == _T_15[9:0]) begin
        image_1_514 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_515 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h203 == _T_37[9:0]) begin
        image_1_515 <= io_pixelVal_in_1_7;
      end else if (10'h203 == _T_34[9:0]) begin
        image_1_515 <= io_pixelVal_in_1_6;
      end else if (10'h203 == _T_31[9:0]) begin
        image_1_515 <= io_pixelVal_in_1_5;
      end else if (10'h203 == _T_28[9:0]) begin
        image_1_515 <= io_pixelVal_in_1_4;
      end else if (10'h203 == _T_25[9:0]) begin
        image_1_515 <= io_pixelVal_in_1_3;
      end else if (10'h203 == _T_22[9:0]) begin
        image_1_515 <= io_pixelVal_in_1_2;
      end else if (10'h203 == _T_19[9:0]) begin
        image_1_515 <= io_pixelVal_in_1_1;
      end else if (10'h203 == _T_15[9:0]) begin
        image_1_515 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_516 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h204 == _T_37[9:0]) begin
        image_1_516 <= io_pixelVal_in_1_7;
      end else if (10'h204 == _T_34[9:0]) begin
        image_1_516 <= io_pixelVal_in_1_6;
      end else if (10'h204 == _T_31[9:0]) begin
        image_1_516 <= io_pixelVal_in_1_5;
      end else if (10'h204 == _T_28[9:0]) begin
        image_1_516 <= io_pixelVal_in_1_4;
      end else if (10'h204 == _T_25[9:0]) begin
        image_1_516 <= io_pixelVal_in_1_3;
      end else if (10'h204 == _T_22[9:0]) begin
        image_1_516 <= io_pixelVal_in_1_2;
      end else if (10'h204 == _T_19[9:0]) begin
        image_1_516 <= io_pixelVal_in_1_1;
      end else if (10'h204 == _T_15[9:0]) begin
        image_1_516 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_517 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h205 == _T_37[9:0]) begin
        image_1_517 <= io_pixelVal_in_1_7;
      end else if (10'h205 == _T_34[9:0]) begin
        image_1_517 <= io_pixelVal_in_1_6;
      end else if (10'h205 == _T_31[9:0]) begin
        image_1_517 <= io_pixelVal_in_1_5;
      end else if (10'h205 == _T_28[9:0]) begin
        image_1_517 <= io_pixelVal_in_1_4;
      end else if (10'h205 == _T_25[9:0]) begin
        image_1_517 <= io_pixelVal_in_1_3;
      end else if (10'h205 == _T_22[9:0]) begin
        image_1_517 <= io_pixelVal_in_1_2;
      end else if (10'h205 == _T_19[9:0]) begin
        image_1_517 <= io_pixelVal_in_1_1;
      end else if (10'h205 == _T_15[9:0]) begin
        image_1_517 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_518 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h206 == _T_37[9:0]) begin
        image_1_518 <= io_pixelVal_in_1_7;
      end else if (10'h206 == _T_34[9:0]) begin
        image_1_518 <= io_pixelVal_in_1_6;
      end else if (10'h206 == _T_31[9:0]) begin
        image_1_518 <= io_pixelVal_in_1_5;
      end else if (10'h206 == _T_28[9:0]) begin
        image_1_518 <= io_pixelVal_in_1_4;
      end else if (10'h206 == _T_25[9:0]) begin
        image_1_518 <= io_pixelVal_in_1_3;
      end else if (10'h206 == _T_22[9:0]) begin
        image_1_518 <= io_pixelVal_in_1_2;
      end else if (10'h206 == _T_19[9:0]) begin
        image_1_518 <= io_pixelVal_in_1_1;
      end else if (10'h206 == _T_15[9:0]) begin
        image_1_518 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_519 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h207 == _T_37[9:0]) begin
        image_1_519 <= io_pixelVal_in_1_7;
      end else if (10'h207 == _T_34[9:0]) begin
        image_1_519 <= io_pixelVal_in_1_6;
      end else if (10'h207 == _T_31[9:0]) begin
        image_1_519 <= io_pixelVal_in_1_5;
      end else if (10'h207 == _T_28[9:0]) begin
        image_1_519 <= io_pixelVal_in_1_4;
      end else if (10'h207 == _T_25[9:0]) begin
        image_1_519 <= io_pixelVal_in_1_3;
      end else if (10'h207 == _T_22[9:0]) begin
        image_1_519 <= io_pixelVal_in_1_2;
      end else if (10'h207 == _T_19[9:0]) begin
        image_1_519 <= io_pixelVal_in_1_1;
      end else if (10'h207 == _T_15[9:0]) begin
        image_1_519 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_520 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h208 == _T_37[9:0]) begin
        image_1_520 <= io_pixelVal_in_1_7;
      end else if (10'h208 == _T_34[9:0]) begin
        image_1_520 <= io_pixelVal_in_1_6;
      end else if (10'h208 == _T_31[9:0]) begin
        image_1_520 <= io_pixelVal_in_1_5;
      end else if (10'h208 == _T_28[9:0]) begin
        image_1_520 <= io_pixelVal_in_1_4;
      end else if (10'h208 == _T_25[9:0]) begin
        image_1_520 <= io_pixelVal_in_1_3;
      end else if (10'h208 == _T_22[9:0]) begin
        image_1_520 <= io_pixelVal_in_1_2;
      end else if (10'h208 == _T_19[9:0]) begin
        image_1_520 <= io_pixelVal_in_1_1;
      end else if (10'h208 == _T_15[9:0]) begin
        image_1_520 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_521 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h209 == _T_37[9:0]) begin
        image_1_521 <= io_pixelVal_in_1_7;
      end else if (10'h209 == _T_34[9:0]) begin
        image_1_521 <= io_pixelVal_in_1_6;
      end else if (10'h209 == _T_31[9:0]) begin
        image_1_521 <= io_pixelVal_in_1_5;
      end else if (10'h209 == _T_28[9:0]) begin
        image_1_521 <= io_pixelVal_in_1_4;
      end else if (10'h209 == _T_25[9:0]) begin
        image_1_521 <= io_pixelVal_in_1_3;
      end else if (10'h209 == _T_22[9:0]) begin
        image_1_521 <= io_pixelVal_in_1_2;
      end else if (10'h209 == _T_19[9:0]) begin
        image_1_521 <= io_pixelVal_in_1_1;
      end else if (10'h209 == _T_15[9:0]) begin
        image_1_521 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_522 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h20a == _T_37[9:0]) begin
        image_1_522 <= io_pixelVal_in_1_7;
      end else if (10'h20a == _T_34[9:0]) begin
        image_1_522 <= io_pixelVal_in_1_6;
      end else if (10'h20a == _T_31[9:0]) begin
        image_1_522 <= io_pixelVal_in_1_5;
      end else if (10'h20a == _T_28[9:0]) begin
        image_1_522 <= io_pixelVal_in_1_4;
      end else if (10'h20a == _T_25[9:0]) begin
        image_1_522 <= io_pixelVal_in_1_3;
      end else if (10'h20a == _T_22[9:0]) begin
        image_1_522 <= io_pixelVal_in_1_2;
      end else if (10'h20a == _T_19[9:0]) begin
        image_1_522 <= io_pixelVal_in_1_1;
      end else if (10'h20a == _T_15[9:0]) begin
        image_1_522 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_523 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h20b == _T_37[9:0]) begin
        image_1_523 <= io_pixelVal_in_1_7;
      end else if (10'h20b == _T_34[9:0]) begin
        image_1_523 <= io_pixelVal_in_1_6;
      end else if (10'h20b == _T_31[9:0]) begin
        image_1_523 <= io_pixelVal_in_1_5;
      end else if (10'h20b == _T_28[9:0]) begin
        image_1_523 <= io_pixelVal_in_1_4;
      end else if (10'h20b == _T_25[9:0]) begin
        image_1_523 <= io_pixelVal_in_1_3;
      end else if (10'h20b == _T_22[9:0]) begin
        image_1_523 <= io_pixelVal_in_1_2;
      end else if (10'h20b == _T_19[9:0]) begin
        image_1_523 <= io_pixelVal_in_1_1;
      end else if (10'h20b == _T_15[9:0]) begin
        image_1_523 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_524 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h20c == _T_37[9:0]) begin
        image_1_524 <= io_pixelVal_in_1_7;
      end else if (10'h20c == _T_34[9:0]) begin
        image_1_524 <= io_pixelVal_in_1_6;
      end else if (10'h20c == _T_31[9:0]) begin
        image_1_524 <= io_pixelVal_in_1_5;
      end else if (10'h20c == _T_28[9:0]) begin
        image_1_524 <= io_pixelVal_in_1_4;
      end else if (10'h20c == _T_25[9:0]) begin
        image_1_524 <= io_pixelVal_in_1_3;
      end else if (10'h20c == _T_22[9:0]) begin
        image_1_524 <= io_pixelVal_in_1_2;
      end else if (10'h20c == _T_19[9:0]) begin
        image_1_524 <= io_pixelVal_in_1_1;
      end else if (10'h20c == _T_15[9:0]) begin
        image_1_524 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_525 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h20d == _T_37[9:0]) begin
        image_1_525 <= io_pixelVal_in_1_7;
      end else if (10'h20d == _T_34[9:0]) begin
        image_1_525 <= io_pixelVal_in_1_6;
      end else if (10'h20d == _T_31[9:0]) begin
        image_1_525 <= io_pixelVal_in_1_5;
      end else if (10'h20d == _T_28[9:0]) begin
        image_1_525 <= io_pixelVal_in_1_4;
      end else if (10'h20d == _T_25[9:0]) begin
        image_1_525 <= io_pixelVal_in_1_3;
      end else if (10'h20d == _T_22[9:0]) begin
        image_1_525 <= io_pixelVal_in_1_2;
      end else if (10'h20d == _T_19[9:0]) begin
        image_1_525 <= io_pixelVal_in_1_1;
      end else if (10'h20d == _T_15[9:0]) begin
        image_1_525 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_526 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h20e == _T_37[9:0]) begin
        image_1_526 <= io_pixelVal_in_1_7;
      end else if (10'h20e == _T_34[9:0]) begin
        image_1_526 <= io_pixelVal_in_1_6;
      end else if (10'h20e == _T_31[9:0]) begin
        image_1_526 <= io_pixelVal_in_1_5;
      end else if (10'h20e == _T_28[9:0]) begin
        image_1_526 <= io_pixelVal_in_1_4;
      end else if (10'h20e == _T_25[9:0]) begin
        image_1_526 <= io_pixelVal_in_1_3;
      end else if (10'h20e == _T_22[9:0]) begin
        image_1_526 <= io_pixelVal_in_1_2;
      end else if (10'h20e == _T_19[9:0]) begin
        image_1_526 <= io_pixelVal_in_1_1;
      end else if (10'h20e == _T_15[9:0]) begin
        image_1_526 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_527 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h20f == _T_37[9:0]) begin
        image_1_527 <= io_pixelVal_in_1_7;
      end else if (10'h20f == _T_34[9:0]) begin
        image_1_527 <= io_pixelVal_in_1_6;
      end else if (10'h20f == _T_31[9:0]) begin
        image_1_527 <= io_pixelVal_in_1_5;
      end else if (10'h20f == _T_28[9:0]) begin
        image_1_527 <= io_pixelVal_in_1_4;
      end else if (10'h20f == _T_25[9:0]) begin
        image_1_527 <= io_pixelVal_in_1_3;
      end else if (10'h20f == _T_22[9:0]) begin
        image_1_527 <= io_pixelVal_in_1_2;
      end else if (10'h20f == _T_19[9:0]) begin
        image_1_527 <= io_pixelVal_in_1_1;
      end else if (10'h20f == _T_15[9:0]) begin
        image_1_527 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_528 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h210 == _T_37[9:0]) begin
        image_1_528 <= io_pixelVal_in_1_7;
      end else if (10'h210 == _T_34[9:0]) begin
        image_1_528 <= io_pixelVal_in_1_6;
      end else if (10'h210 == _T_31[9:0]) begin
        image_1_528 <= io_pixelVal_in_1_5;
      end else if (10'h210 == _T_28[9:0]) begin
        image_1_528 <= io_pixelVal_in_1_4;
      end else if (10'h210 == _T_25[9:0]) begin
        image_1_528 <= io_pixelVal_in_1_3;
      end else if (10'h210 == _T_22[9:0]) begin
        image_1_528 <= io_pixelVal_in_1_2;
      end else if (10'h210 == _T_19[9:0]) begin
        image_1_528 <= io_pixelVal_in_1_1;
      end else if (10'h210 == _T_15[9:0]) begin
        image_1_528 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_529 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h211 == _T_37[9:0]) begin
        image_1_529 <= io_pixelVal_in_1_7;
      end else if (10'h211 == _T_34[9:0]) begin
        image_1_529 <= io_pixelVal_in_1_6;
      end else if (10'h211 == _T_31[9:0]) begin
        image_1_529 <= io_pixelVal_in_1_5;
      end else if (10'h211 == _T_28[9:0]) begin
        image_1_529 <= io_pixelVal_in_1_4;
      end else if (10'h211 == _T_25[9:0]) begin
        image_1_529 <= io_pixelVal_in_1_3;
      end else if (10'h211 == _T_22[9:0]) begin
        image_1_529 <= io_pixelVal_in_1_2;
      end else if (10'h211 == _T_19[9:0]) begin
        image_1_529 <= io_pixelVal_in_1_1;
      end else if (10'h211 == _T_15[9:0]) begin
        image_1_529 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_530 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h212 == _T_37[9:0]) begin
        image_1_530 <= io_pixelVal_in_1_7;
      end else if (10'h212 == _T_34[9:0]) begin
        image_1_530 <= io_pixelVal_in_1_6;
      end else if (10'h212 == _T_31[9:0]) begin
        image_1_530 <= io_pixelVal_in_1_5;
      end else if (10'h212 == _T_28[9:0]) begin
        image_1_530 <= io_pixelVal_in_1_4;
      end else if (10'h212 == _T_25[9:0]) begin
        image_1_530 <= io_pixelVal_in_1_3;
      end else if (10'h212 == _T_22[9:0]) begin
        image_1_530 <= io_pixelVal_in_1_2;
      end else if (10'h212 == _T_19[9:0]) begin
        image_1_530 <= io_pixelVal_in_1_1;
      end else if (10'h212 == _T_15[9:0]) begin
        image_1_530 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_531 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h213 == _T_37[9:0]) begin
        image_1_531 <= io_pixelVal_in_1_7;
      end else if (10'h213 == _T_34[9:0]) begin
        image_1_531 <= io_pixelVal_in_1_6;
      end else if (10'h213 == _T_31[9:0]) begin
        image_1_531 <= io_pixelVal_in_1_5;
      end else if (10'h213 == _T_28[9:0]) begin
        image_1_531 <= io_pixelVal_in_1_4;
      end else if (10'h213 == _T_25[9:0]) begin
        image_1_531 <= io_pixelVal_in_1_3;
      end else if (10'h213 == _T_22[9:0]) begin
        image_1_531 <= io_pixelVal_in_1_2;
      end else if (10'h213 == _T_19[9:0]) begin
        image_1_531 <= io_pixelVal_in_1_1;
      end else if (10'h213 == _T_15[9:0]) begin
        image_1_531 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_532 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h214 == _T_37[9:0]) begin
        image_1_532 <= io_pixelVal_in_1_7;
      end else if (10'h214 == _T_34[9:0]) begin
        image_1_532 <= io_pixelVal_in_1_6;
      end else if (10'h214 == _T_31[9:0]) begin
        image_1_532 <= io_pixelVal_in_1_5;
      end else if (10'h214 == _T_28[9:0]) begin
        image_1_532 <= io_pixelVal_in_1_4;
      end else if (10'h214 == _T_25[9:0]) begin
        image_1_532 <= io_pixelVal_in_1_3;
      end else if (10'h214 == _T_22[9:0]) begin
        image_1_532 <= io_pixelVal_in_1_2;
      end else if (10'h214 == _T_19[9:0]) begin
        image_1_532 <= io_pixelVal_in_1_1;
      end else if (10'h214 == _T_15[9:0]) begin
        image_1_532 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_533 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h215 == _T_37[9:0]) begin
        image_1_533 <= io_pixelVal_in_1_7;
      end else if (10'h215 == _T_34[9:0]) begin
        image_1_533 <= io_pixelVal_in_1_6;
      end else if (10'h215 == _T_31[9:0]) begin
        image_1_533 <= io_pixelVal_in_1_5;
      end else if (10'h215 == _T_28[9:0]) begin
        image_1_533 <= io_pixelVal_in_1_4;
      end else if (10'h215 == _T_25[9:0]) begin
        image_1_533 <= io_pixelVal_in_1_3;
      end else if (10'h215 == _T_22[9:0]) begin
        image_1_533 <= io_pixelVal_in_1_2;
      end else if (10'h215 == _T_19[9:0]) begin
        image_1_533 <= io_pixelVal_in_1_1;
      end else if (10'h215 == _T_15[9:0]) begin
        image_1_533 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_534 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h216 == _T_37[9:0]) begin
        image_1_534 <= io_pixelVal_in_1_7;
      end else if (10'h216 == _T_34[9:0]) begin
        image_1_534 <= io_pixelVal_in_1_6;
      end else if (10'h216 == _T_31[9:0]) begin
        image_1_534 <= io_pixelVal_in_1_5;
      end else if (10'h216 == _T_28[9:0]) begin
        image_1_534 <= io_pixelVal_in_1_4;
      end else if (10'h216 == _T_25[9:0]) begin
        image_1_534 <= io_pixelVal_in_1_3;
      end else if (10'h216 == _T_22[9:0]) begin
        image_1_534 <= io_pixelVal_in_1_2;
      end else if (10'h216 == _T_19[9:0]) begin
        image_1_534 <= io_pixelVal_in_1_1;
      end else if (10'h216 == _T_15[9:0]) begin
        image_1_534 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_535 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h217 == _T_37[9:0]) begin
        image_1_535 <= io_pixelVal_in_1_7;
      end else if (10'h217 == _T_34[9:0]) begin
        image_1_535 <= io_pixelVal_in_1_6;
      end else if (10'h217 == _T_31[9:0]) begin
        image_1_535 <= io_pixelVal_in_1_5;
      end else if (10'h217 == _T_28[9:0]) begin
        image_1_535 <= io_pixelVal_in_1_4;
      end else if (10'h217 == _T_25[9:0]) begin
        image_1_535 <= io_pixelVal_in_1_3;
      end else if (10'h217 == _T_22[9:0]) begin
        image_1_535 <= io_pixelVal_in_1_2;
      end else if (10'h217 == _T_19[9:0]) begin
        image_1_535 <= io_pixelVal_in_1_1;
      end else if (10'h217 == _T_15[9:0]) begin
        image_1_535 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_536 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h218 == _T_37[9:0]) begin
        image_1_536 <= io_pixelVal_in_1_7;
      end else if (10'h218 == _T_34[9:0]) begin
        image_1_536 <= io_pixelVal_in_1_6;
      end else if (10'h218 == _T_31[9:0]) begin
        image_1_536 <= io_pixelVal_in_1_5;
      end else if (10'h218 == _T_28[9:0]) begin
        image_1_536 <= io_pixelVal_in_1_4;
      end else if (10'h218 == _T_25[9:0]) begin
        image_1_536 <= io_pixelVal_in_1_3;
      end else if (10'h218 == _T_22[9:0]) begin
        image_1_536 <= io_pixelVal_in_1_2;
      end else if (10'h218 == _T_19[9:0]) begin
        image_1_536 <= io_pixelVal_in_1_1;
      end else if (10'h218 == _T_15[9:0]) begin
        image_1_536 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_537 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h219 == _T_37[9:0]) begin
        image_1_537 <= io_pixelVal_in_1_7;
      end else if (10'h219 == _T_34[9:0]) begin
        image_1_537 <= io_pixelVal_in_1_6;
      end else if (10'h219 == _T_31[9:0]) begin
        image_1_537 <= io_pixelVal_in_1_5;
      end else if (10'h219 == _T_28[9:0]) begin
        image_1_537 <= io_pixelVal_in_1_4;
      end else if (10'h219 == _T_25[9:0]) begin
        image_1_537 <= io_pixelVal_in_1_3;
      end else if (10'h219 == _T_22[9:0]) begin
        image_1_537 <= io_pixelVal_in_1_2;
      end else if (10'h219 == _T_19[9:0]) begin
        image_1_537 <= io_pixelVal_in_1_1;
      end else if (10'h219 == _T_15[9:0]) begin
        image_1_537 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_538 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h21a == _T_37[9:0]) begin
        image_1_538 <= io_pixelVal_in_1_7;
      end else if (10'h21a == _T_34[9:0]) begin
        image_1_538 <= io_pixelVal_in_1_6;
      end else if (10'h21a == _T_31[9:0]) begin
        image_1_538 <= io_pixelVal_in_1_5;
      end else if (10'h21a == _T_28[9:0]) begin
        image_1_538 <= io_pixelVal_in_1_4;
      end else if (10'h21a == _T_25[9:0]) begin
        image_1_538 <= io_pixelVal_in_1_3;
      end else if (10'h21a == _T_22[9:0]) begin
        image_1_538 <= io_pixelVal_in_1_2;
      end else if (10'h21a == _T_19[9:0]) begin
        image_1_538 <= io_pixelVal_in_1_1;
      end else if (10'h21a == _T_15[9:0]) begin
        image_1_538 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_539 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h21b == _T_37[9:0]) begin
        image_1_539 <= io_pixelVal_in_1_7;
      end else if (10'h21b == _T_34[9:0]) begin
        image_1_539 <= io_pixelVal_in_1_6;
      end else if (10'h21b == _T_31[9:0]) begin
        image_1_539 <= io_pixelVal_in_1_5;
      end else if (10'h21b == _T_28[9:0]) begin
        image_1_539 <= io_pixelVal_in_1_4;
      end else if (10'h21b == _T_25[9:0]) begin
        image_1_539 <= io_pixelVal_in_1_3;
      end else if (10'h21b == _T_22[9:0]) begin
        image_1_539 <= io_pixelVal_in_1_2;
      end else if (10'h21b == _T_19[9:0]) begin
        image_1_539 <= io_pixelVal_in_1_1;
      end else if (10'h21b == _T_15[9:0]) begin
        image_1_539 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_540 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h21c == _T_37[9:0]) begin
        image_1_540 <= io_pixelVal_in_1_7;
      end else if (10'h21c == _T_34[9:0]) begin
        image_1_540 <= io_pixelVal_in_1_6;
      end else if (10'h21c == _T_31[9:0]) begin
        image_1_540 <= io_pixelVal_in_1_5;
      end else if (10'h21c == _T_28[9:0]) begin
        image_1_540 <= io_pixelVal_in_1_4;
      end else if (10'h21c == _T_25[9:0]) begin
        image_1_540 <= io_pixelVal_in_1_3;
      end else if (10'h21c == _T_22[9:0]) begin
        image_1_540 <= io_pixelVal_in_1_2;
      end else if (10'h21c == _T_19[9:0]) begin
        image_1_540 <= io_pixelVal_in_1_1;
      end else if (10'h21c == _T_15[9:0]) begin
        image_1_540 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_541 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h21d == _T_37[9:0]) begin
        image_1_541 <= io_pixelVal_in_1_7;
      end else if (10'h21d == _T_34[9:0]) begin
        image_1_541 <= io_pixelVal_in_1_6;
      end else if (10'h21d == _T_31[9:0]) begin
        image_1_541 <= io_pixelVal_in_1_5;
      end else if (10'h21d == _T_28[9:0]) begin
        image_1_541 <= io_pixelVal_in_1_4;
      end else if (10'h21d == _T_25[9:0]) begin
        image_1_541 <= io_pixelVal_in_1_3;
      end else if (10'h21d == _T_22[9:0]) begin
        image_1_541 <= io_pixelVal_in_1_2;
      end else if (10'h21d == _T_19[9:0]) begin
        image_1_541 <= io_pixelVal_in_1_1;
      end else if (10'h21d == _T_15[9:0]) begin
        image_1_541 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_542 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h21e == _T_37[9:0]) begin
        image_1_542 <= io_pixelVal_in_1_7;
      end else if (10'h21e == _T_34[9:0]) begin
        image_1_542 <= io_pixelVal_in_1_6;
      end else if (10'h21e == _T_31[9:0]) begin
        image_1_542 <= io_pixelVal_in_1_5;
      end else if (10'h21e == _T_28[9:0]) begin
        image_1_542 <= io_pixelVal_in_1_4;
      end else if (10'h21e == _T_25[9:0]) begin
        image_1_542 <= io_pixelVal_in_1_3;
      end else if (10'h21e == _T_22[9:0]) begin
        image_1_542 <= io_pixelVal_in_1_2;
      end else if (10'h21e == _T_19[9:0]) begin
        image_1_542 <= io_pixelVal_in_1_1;
      end else if (10'h21e == _T_15[9:0]) begin
        image_1_542 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_543 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h21f == _T_37[9:0]) begin
        image_1_543 <= io_pixelVal_in_1_7;
      end else if (10'h21f == _T_34[9:0]) begin
        image_1_543 <= io_pixelVal_in_1_6;
      end else if (10'h21f == _T_31[9:0]) begin
        image_1_543 <= io_pixelVal_in_1_5;
      end else if (10'h21f == _T_28[9:0]) begin
        image_1_543 <= io_pixelVal_in_1_4;
      end else if (10'h21f == _T_25[9:0]) begin
        image_1_543 <= io_pixelVal_in_1_3;
      end else if (10'h21f == _T_22[9:0]) begin
        image_1_543 <= io_pixelVal_in_1_2;
      end else if (10'h21f == _T_19[9:0]) begin
        image_1_543 <= io_pixelVal_in_1_1;
      end else if (10'h21f == _T_15[9:0]) begin
        image_1_543 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_544 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h220 == _T_37[9:0]) begin
        image_1_544 <= io_pixelVal_in_1_7;
      end else if (10'h220 == _T_34[9:0]) begin
        image_1_544 <= io_pixelVal_in_1_6;
      end else if (10'h220 == _T_31[9:0]) begin
        image_1_544 <= io_pixelVal_in_1_5;
      end else if (10'h220 == _T_28[9:0]) begin
        image_1_544 <= io_pixelVal_in_1_4;
      end else if (10'h220 == _T_25[9:0]) begin
        image_1_544 <= io_pixelVal_in_1_3;
      end else if (10'h220 == _T_22[9:0]) begin
        image_1_544 <= io_pixelVal_in_1_2;
      end else if (10'h220 == _T_19[9:0]) begin
        image_1_544 <= io_pixelVal_in_1_1;
      end else if (10'h220 == _T_15[9:0]) begin
        image_1_544 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_545 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h221 == _T_37[9:0]) begin
        image_1_545 <= io_pixelVal_in_1_7;
      end else if (10'h221 == _T_34[9:0]) begin
        image_1_545 <= io_pixelVal_in_1_6;
      end else if (10'h221 == _T_31[9:0]) begin
        image_1_545 <= io_pixelVal_in_1_5;
      end else if (10'h221 == _T_28[9:0]) begin
        image_1_545 <= io_pixelVal_in_1_4;
      end else if (10'h221 == _T_25[9:0]) begin
        image_1_545 <= io_pixelVal_in_1_3;
      end else if (10'h221 == _T_22[9:0]) begin
        image_1_545 <= io_pixelVal_in_1_2;
      end else if (10'h221 == _T_19[9:0]) begin
        image_1_545 <= io_pixelVal_in_1_1;
      end else if (10'h221 == _T_15[9:0]) begin
        image_1_545 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_546 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h222 == _T_37[9:0]) begin
        image_1_546 <= io_pixelVal_in_1_7;
      end else if (10'h222 == _T_34[9:0]) begin
        image_1_546 <= io_pixelVal_in_1_6;
      end else if (10'h222 == _T_31[9:0]) begin
        image_1_546 <= io_pixelVal_in_1_5;
      end else if (10'h222 == _T_28[9:0]) begin
        image_1_546 <= io_pixelVal_in_1_4;
      end else if (10'h222 == _T_25[9:0]) begin
        image_1_546 <= io_pixelVal_in_1_3;
      end else if (10'h222 == _T_22[9:0]) begin
        image_1_546 <= io_pixelVal_in_1_2;
      end else if (10'h222 == _T_19[9:0]) begin
        image_1_546 <= io_pixelVal_in_1_1;
      end else if (10'h222 == _T_15[9:0]) begin
        image_1_546 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_547 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h223 == _T_37[9:0]) begin
        image_1_547 <= io_pixelVal_in_1_7;
      end else if (10'h223 == _T_34[9:0]) begin
        image_1_547 <= io_pixelVal_in_1_6;
      end else if (10'h223 == _T_31[9:0]) begin
        image_1_547 <= io_pixelVal_in_1_5;
      end else if (10'h223 == _T_28[9:0]) begin
        image_1_547 <= io_pixelVal_in_1_4;
      end else if (10'h223 == _T_25[9:0]) begin
        image_1_547 <= io_pixelVal_in_1_3;
      end else if (10'h223 == _T_22[9:0]) begin
        image_1_547 <= io_pixelVal_in_1_2;
      end else if (10'h223 == _T_19[9:0]) begin
        image_1_547 <= io_pixelVal_in_1_1;
      end else if (10'h223 == _T_15[9:0]) begin
        image_1_547 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_548 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h224 == _T_37[9:0]) begin
        image_1_548 <= io_pixelVal_in_1_7;
      end else if (10'h224 == _T_34[9:0]) begin
        image_1_548 <= io_pixelVal_in_1_6;
      end else if (10'h224 == _T_31[9:0]) begin
        image_1_548 <= io_pixelVal_in_1_5;
      end else if (10'h224 == _T_28[9:0]) begin
        image_1_548 <= io_pixelVal_in_1_4;
      end else if (10'h224 == _T_25[9:0]) begin
        image_1_548 <= io_pixelVal_in_1_3;
      end else if (10'h224 == _T_22[9:0]) begin
        image_1_548 <= io_pixelVal_in_1_2;
      end else if (10'h224 == _T_19[9:0]) begin
        image_1_548 <= io_pixelVal_in_1_1;
      end else if (10'h224 == _T_15[9:0]) begin
        image_1_548 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_549 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h225 == _T_37[9:0]) begin
        image_1_549 <= io_pixelVal_in_1_7;
      end else if (10'h225 == _T_34[9:0]) begin
        image_1_549 <= io_pixelVal_in_1_6;
      end else if (10'h225 == _T_31[9:0]) begin
        image_1_549 <= io_pixelVal_in_1_5;
      end else if (10'h225 == _T_28[9:0]) begin
        image_1_549 <= io_pixelVal_in_1_4;
      end else if (10'h225 == _T_25[9:0]) begin
        image_1_549 <= io_pixelVal_in_1_3;
      end else if (10'h225 == _T_22[9:0]) begin
        image_1_549 <= io_pixelVal_in_1_2;
      end else if (10'h225 == _T_19[9:0]) begin
        image_1_549 <= io_pixelVal_in_1_1;
      end else if (10'h225 == _T_15[9:0]) begin
        image_1_549 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_550 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h226 == _T_37[9:0]) begin
        image_1_550 <= io_pixelVal_in_1_7;
      end else if (10'h226 == _T_34[9:0]) begin
        image_1_550 <= io_pixelVal_in_1_6;
      end else if (10'h226 == _T_31[9:0]) begin
        image_1_550 <= io_pixelVal_in_1_5;
      end else if (10'h226 == _T_28[9:0]) begin
        image_1_550 <= io_pixelVal_in_1_4;
      end else if (10'h226 == _T_25[9:0]) begin
        image_1_550 <= io_pixelVal_in_1_3;
      end else if (10'h226 == _T_22[9:0]) begin
        image_1_550 <= io_pixelVal_in_1_2;
      end else if (10'h226 == _T_19[9:0]) begin
        image_1_550 <= io_pixelVal_in_1_1;
      end else if (10'h226 == _T_15[9:0]) begin
        image_1_550 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_551 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h227 == _T_37[9:0]) begin
        image_1_551 <= io_pixelVal_in_1_7;
      end else if (10'h227 == _T_34[9:0]) begin
        image_1_551 <= io_pixelVal_in_1_6;
      end else if (10'h227 == _T_31[9:0]) begin
        image_1_551 <= io_pixelVal_in_1_5;
      end else if (10'h227 == _T_28[9:0]) begin
        image_1_551 <= io_pixelVal_in_1_4;
      end else if (10'h227 == _T_25[9:0]) begin
        image_1_551 <= io_pixelVal_in_1_3;
      end else if (10'h227 == _T_22[9:0]) begin
        image_1_551 <= io_pixelVal_in_1_2;
      end else if (10'h227 == _T_19[9:0]) begin
        image_1_551 <= io_pixelVal_in_1_1;
      end else if (10'h227 == _T_15[9:0]) begin
        image_1_551 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_552 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h228 == _T_37[9:0]) begin
        image_1_552 <= io_pixelVal_in_1_7;
      end else if (10'h228 == _T_34[9:0]) begin
        image_1_552 <= io_pixelVal_in_1_6;
      end else if (10'h228 == _T_31[9:0]) begin
        image_1_552 <= io_pixelVal_in_1_5;
      end else if (10'h228 == _T_28[9:0]) begin
        image_1_552 <= io_pixelVal_in_1_4;
      end else if (10'h228 == _T_25[9:0]) begin
        image_1_552 <= io_pixelVal_in_1_3;
      end else if (10'h228 == _T_22[9:0]) begin
        image_1_552 <= io_pixelVal_in_1_2;
      end else if (10'h228 == _T_19[9:0]) begin
        image_1_552 <= io_pixelVal_in_1_1;
      end else if (10'h228 == _T_15[9:0]) begin
        image_1_552 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_553 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h229 == _T_37[9:0]) begin
        image_1_553 <= io_pixelVal_in_1_7;
      end else if (10'h229 == _T_34[9:0]) begin
        image_1_553 <= io_pixelVal_in_1_6;
      end else if (10'h229 == _T_31[9:0]) begin
        image_1_553 <= io_pixelVal_in_1_5;
      end else if (10'h229 == _T_28[9:0]) begin
        image_1_553 <= io_pixelVal_in_1_4;
      end else if (10'h229 == _T_25[9:0]) begin
        image_1_553 <= io_pixelVal_in_1_3;
      end else if (10'h229 == _T_22[9:0]) begin
        image_1_553 <= io_pixelVal_in_1_2;
      end else if (10'h229 == _T_19[9:0]) begin
        image_1_553 <= io_pixelVal_in_1_1;
      end else if (10'h229 == _T_15[9:0]) begin
        image_1_553 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_554 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h22a == _T_37[9:0]) begin
        image_1_554 <= io_pixelVal_in_1_7;
      end else if (10'h22a == _T_34[9:0]) begin
        image_1_554 <= io_pixelVal_in_1_6;
      end else if (10'h22a == _T_31[9:0]) begin
        image_1_554 <= io_pixelVal_in_1_5;
      end else if (10'h22a == _T_28[9:0]) begin
        image_1_554 <= io_pixelVal_in_1_4;
      end else if (10'h22a == _T_25[9:0]) begin
        image_1_554 <= io_pixelVal_in_1_3;
      end else if (10'h22a == _T_22[9:0]) begin
        image_1_554 <= io_pixelVal_in_1_2;
      end else if (10'h22a == _T_19[9:0]) begin
        image_1_554 <= io_pixelVal_in_1_1;
      end else if (10'h22a == _T_15[9:0]) begin
        image_1_554 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_555 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h22b == _T_37[9:0]) begin
        image_1_555 <= io_pixelVal_in_1_7;
      end else if (10'h22b == _T_34[9:0]) begin
        image_1_555 <= io_pixelVal_in_1_6;
      end else if (10'h22b == _T_31[9:0]) begin
        image_1_555 <= io_pixelVal_in_1_5;
      end else if (10'h22b == _T_28[9:0]) begin
        image_1_555 <= io_pixelVal_in_1_4;
      end else if (10'h22b == _T_25[9:0]) begin
        image_1_555 <= io_pixelVal_in_1_3;
      end else if (10'h22b == _T_22[9:0]) begin
        image_1_555 <= io_pixelVal_in_1_2;
      end else if (10'h22b == _T_19[9:0]) begin
        image_1_555 <= io_pixelVal_in_1_1;
      end else if (10'h22b == _T_15[9:0]) begin
        image_1_555 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_556 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h22c == _T_37[9:0]) begin
        image_1_556 <= io_pixelVal_in_1_7;
      end else if (10'h22c == _T_34[9:0]) begin
        image_1_556 <= io_pixelVal_in_1_6;
      end else if (10'h22c == _T_31[9:0]) begin
        image_1_556 <= io_pixelVal_in_1_5;
      end else if (10'h22c == _T_28[9:0]) begin
        image_1_556 <= io_pixelVal_in_1_4;
      end else if (10'h22c == _T_25[9:0]) begin
        image_1_556 <= io_pixelVal_in_1_3;
      end else if (10'h22c == _T_22[9:0]) begin
        image_1_556 <= io_pixelVal_in_1_2;
      end else if (10'h22c == _T_19[9:0]) begin
        image_1_556 <= io_pixelVal_in_1_1;
      end else if (10'h22c == _T_15[9:0]) begin
        image_1_556 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_557 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h22d == _T_37[9:0]) begin
        image_1_557 <= io_pixelVal_in_1_7;
      end else if (10'h22d == _T_34[9:0]) begin
        image_1_557 <= io_pixelVal_in_1_6;
      end else if (10'h22d == _T_31[9:0]) begin
        image_1_557 <= io_pixelVal_in_1_5;
      end else if (10'h22d == _T_28[9:0]) begin
        image_1_557 <= io_pixelVal_in_1_4;
      end else if (10'h22d == _T_25[9:0]) begin
        image_1_557 <= io_pixelVal_in_1_3;
      end else if (10'h22d == _T_22[9:0]) begin
        image_1_557 <= io_pixelVal_in_1_2;
      end else if (10'h22d == _T_19[9:0]) begin
        image_1_557 <= io_pixelVal_in_1_1;
      end else if (10'h22d == _T_15[9:0]) begin
        image_1_557 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_558 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h22e == _T_37[9:0]) begin
        image_1_558 <= io_pixelVal_in_1_7;
      end else if (10'h22e == _T_34[9:0]) begin
        image_1_558 <= io_pixelVal_in_1_6;
      end else if (10'h22e == _T_31[9:0]) begin
        image_1_558 <= io_pixelVal_in_1_5;
      end else if (10'h22e == _T_28[9:0]) begin
        image_1_558 <= io_pixelVal_in_1_4;
      end else if (10'h22e == _T_25[9:0]) begin
        image_1_558 <= io_pixelVal_in_1_3;
      end else if (10'h22e == _T_22[9:0]) begin
        image_1_558 <= io_pixelVal_in_1_2;
      end else if (10'h22e == _T_19[9:0]) begin
        image_1_558 <= io_pixelVal_in_1_1;
      end else if (10'h22e == _T_15[9:0]) begin
        image_1_558 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_559 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h22f == _T_37[9:0]) begin
        image_1_559 <= io_pixelVal_in_1_7;
      end else if (10'h22f == _T_34[9:0]) begin
        image_1_559 <= io_pixelVal_in_1_6;
      end else if (10'h22f == _T_31[9:0]) begin
        image_1_559 <= io_pixelVal_in_1_5;
      end else if (10'h22f == _T_28[9:0]) begin
        image_1_559 <= io_pixelVal_in_1_4;
      end else if (10'h22f == _T_25[9:0]) begin
        image_1_559 <= io_pixelVal_in_1_3;
      end else if (10'h22f == _T_22[9:0]) begin
        image_1_559 <= io_pixelVal_in_1_2;
      end else if (10'h22f == _T_19[9:0]) begin
        image_1_559 <= io_pixelVal_in_1_1;
      end else if (10'h22f == _T_15[9:0]) begin
        image_1_559 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_560 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h230 == _T_37[9:0]) begin
        image_1_560 <= io_pixelVal_in_1_7;
      end else if (10'h230 == _T_34[9:0]) begin
        image_1_560 <= io_pixelVal_in_1_6;
      end else if (10'h230 == _T_31[9:0]) begin
        image_1_560 <= io_pixelVal_in_1_5;
      end else if (10'h230 == _T_28[9:0]) begin
        image_1_560 <= io_pixelVal_in_1_4;
      end else if (10'h230 == _T_25[9:0]) begin
        image_1_560 <= io_pixelVal_in_1_3;
      end else if (10'h230 == _T_22[9:0]) begin
        image_1_560 <= io_pixelVal_in_1_2;
      end else if (10'h230 == _T_19[9:0]) begin
        image_1_560 <= io_pixelVal_in_1_1;
      end else if (10'h230 == _T_15[9:0]) begin
        image_1_560 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_561 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h231 == _T_37[9:0]) begin
        image_1_561 <= io_pixelVal_in_1_7;
      end else if (10'h231 == _T_34[9:0]) begin
        image_1_561 <= io_pixelVal_in_1_6;
      end else if (10'h231 == _T_31[9:0]) begin
        image_1_561 <= io_pixelVal_in_1_5;
      end else if (10'h231 == _T_28[9:0]) begin
        image_1_561 <= io_pixelVal_in_1_4;
      end else if (10'h231 == _T_25[9:0]) begin
        image_1_561 <= io_pixelVal_in_1_3;
      end else if (10'h231 == _T_22[9:0]) begin
        image_1_561 <= io_pixelVal_in_1_2;
      end else if (10'h231 == _T_19[9:0]) begin
        image_1_561 <= io_pixelVal_in_1_1;
      end else if (10'h231 == _T_15[9:0]) begin
        image_1_561 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_562 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h232 == _T_37[9:0]) begin
        image_1_562 <= io_pixelVal_in_1_7;
      end else if (10'h232 == _T_34[9:0]) begin
        image_1_562 <= io_pixelVal_in_1_6;
      end else if (10'h232 == _T_31[9:0]) begin
        image_1_562 <= io_pixelVal_in_1_5;
      end else if (10'h232 == _T_28[9:0]) begin
        image_1_562 <= io_pixelVal_in_1_4;
      end else if (10'h232 == _T_25[9:0]) begin
        image_1_562 <= io_pixelVal_in_1_3;
      end else if (10'h232 == _T_22[9:0]) begin
        image_1_562 <= io_pixelVal_in_1_2;
      end else if (10'h232 == _T_19[9:0]) begin
        image_1_562 <= io_pixelVal_in_1_1;
      end else if (10'h232 == _T_15[9:0]) begin
        image_1_562 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_563 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h233 == _T_37[9:0]) begin
        image_1_563 <= io_pixelVal_in_1_7;
      end else if (10'h233 == _T_34[9:0]) begin
        image_1_563 <= io_pixelVal_in_1_6;
      end else if (10'h233 == _T_31[9:0]) begin
        image_1_563 <= io_pixelVal_in_1_5;
      end else if (10'h233 == _T_28[9:0]) begin
        image_1_563 <= io_pixelVal_in_1_4;
      end else if (10'h233 == _T_25[9:0]) begin
        image_1_563 <= io_pixelVal_in_1_3;
      end else if (10'h233 == _T_22[9:0]) begin
        image_1_563 <= io_pixelVal_in_1_2;
      end else if (10'h233 == _T_19[9:0]) begin
        image_1_563 <= io_pixelVal_in_1_1;
      end else if (10'h233 == _T_15[9:0]) begin
        image_1_563 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_564 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h234 == _T_37[9:0]) begin
        image_1_564 <= io_pixelVal_in_1_7;
      end else if (10'h234 == _T_34[9:0]) begin
        image_1_564 <= io_pixelVal_in_1_6;
      end else if (10'h234 == _T_31[9:0]) begin
        image_1_564 <= io_pixelVal_in_1_5;
      end else if (10'h234 == _T_28[9:0]) begin
        image_1_564 <= io_pixelVal_in_1_4;
      end else if (10'h234 == _T_25[9:0]) begin
        image_1_564 <= io_pixelVal_in_1_3;
      end else if (10'h234 == _T_22[9:0]) begin
        image_1_564 <= io_pixelVal_in_1_2;
      end else if (10'h234 == _T_19[9:0]) begin
        image_1_564 <= io_pixelVal_in_1_1;
      end else if (10'h234 == _T_15[9:0]) begin
        image_1_564 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_565 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h235 == _T_37[9:0]) begin
        image_1_565 <= io_pixelVal_in_1_7;
      end else if (10'h235 == _T_34[9:0]) begin
        image_1_565 <= io_pixelVal_in_1_6;
      end else if (10'h235 == _T_31[9:0]) begin
        image_1_565 <= io_pixelVal_in_1_5;
      end else if (10'h235 == _T_28[9:0]) begin
        image_1_565 <= io_pixelVal_in_1_4;
      end else if (10'h235 == _T_25[9:0]) begin
        image_1_565 <= io_pixelVal_in_1_3;
      end else if (10'h235 == _T_22[9:0]) begin
        image_1_565 <= io_pixelVal_in_1_2;
      end else if (10'h235 == _T_19[9:0]) begin
        image_1_565 <= io_pixelVal_in_1_1;
      end else if (10'h235 == _T_15[9:0]) begin
        image_1_565 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_566 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h236 == _T_37[9:0]) begin
        image_1_566 <= io_pixelVal_in_1_7;
      end else if (10'h236 == _T_34[9:0]) begin
        image_1_566 <= io_pixelVal_in_1_6;
      end else if (10'h236 == _T_31[9:0]) begin
        image_1_566 <= io_pixelVal_in_1_5;
      end else if (10'h236 == _T_28[9:0]) begin
        image_1_566 <= io_pixelVal_in_1_4;
      end else if (10'h236 == _T_25[9:0]) begin
        image_1_566 <= io_pixelVal_in_1_3;
      end else if (10'h236 == _T_22[9:0]) begin
        image_1_566 <= io_pixelVal_in_1_2;
      end else if (10'h236 == _T_19[9:0]) begin
        image_1_566 <= io_pixelVal_in_1_1;
      end else if (10'h236 == _T_15[9:0]) begin
        image_1_566 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_567 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h237 == _T_37[9:0]) begin
        image_1_567 <= io_pixelVal_in_1_7;
      end else if (10'h237 == _T_34[9:0]) begin
        image_1_567 <= io_pixelVal_in_1_6;
      end else if (10'h237 == _T_31[9:0]) begin
        image_1_567 <= io_pixelVal_in_1_5;
      end else if (10'h237 == _T_28[9:0]) begin
        image_1_567 <= io_pixelVal_in_1_4;
      end else if (10'h237 == _T_25[9:0]) begin
        image_1_567 <= io_pixelVal_in_1_3;
      end else if (10'h237 == _T_22[9:0]) begin
        image_1_567 <= io_pixelVal_in_1_2;
      end else if (10'h237 == _T_19[9:0]) begin
        image_1_567 <= io_pixelVal_in_1_1;
      end else if (10'h237 == _T_15[9:0]) begin
        image_1_567 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_568 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h238 == _T_37[9:0]) begin
        image_1_568 <= io_pixelVal_in_1_7;
      end else if (10'h238 == _T_34[9:0]) begin
        image_1_568 <= io_pixelVal_in_1_6;
      end else if (10'h238 == _T_31[9:0]) begin
        image_1_568 <= io_pixelVal_in_1_5;
      end else if (10'h238 == _T_28[9:0]) begin
        image_1_568 <= io_pixelVal_in_1_4;
      end else if (10'h238 == _T_25[9:0]) begin
        image_1_568 <= io_pixelVal_in_1_3;
      end else if (10'h238 == _T_22[9:0]) begin
        image_1_568 <= io_pixelVal_in_1_2;
      end else if (10'h238 == _T_19[9:0]) begin
        image_1_568 <= io_pixelVal_in_1_1;
      end else if (10'h238 == _T_15[9:0]) begin
        image_1_568 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_569 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h239 == _T_37[9:0]) begin
        image_1_569 <= io_pixelVal_in_1_7;
      end else if (10'h239 == _T_34[9:0]) begin
        image_1_569 <= io_pixelVal_in_1_6;
      end else if (10'h239 == _T_31[9:0]) begin
        image_1_569 <= io_pixelVal_in_1_5;
      end else if (10'h239 == _T_28[9:0]) begin
        image_1_569 <= io_pixelVal_in_1_4;
      end else if (10'h239 == _T_25[9:0]) begin
        image_1_569 <= io_pixelVal_in_1_3;
      end else if (10'h239 == _T_22[9:0]) begin
        image_1_569 <= io_pixelVal_in_1_2;
      end else if (10'h239 == _T_19[9:0]) begin
        image_1_569 <= io_pixelVal_in_1_1;
      end else if (10'h239 == _T_15[9:0]) begin
        image_1_569 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_570 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h23a == _T_37[9:0]) begin
        image_1_570 <= io_pixelVal_in_1_7;
      end else if (10'h23a == _T_34[9:0]) begin
        image_1_570 <= io_pixelVal_in_1_6;
      end else if (10'h23a == _T_31[9:0]) begin
        image_1_570 <= io_pixelVal_in_1_5;
      end else if (10'h23a == _T_28[9:0]) begin
        image_1_570 <= io_pixelVal_in_1_4;
      end else if (10'h23a == _T_25[9:0]) begin
        image_1_570 <= io_pixelVal_in_1_3;
      end else if (10'h23a == _T_22[9:0]) begin
        image_1_570 <= io_pixelVal_in_1_2;
      end else if (10'h23a == _T_19[9:0]) begin
        image_1_570 <= io_pixelVal_in_1_1;
      end else if (10'h23a == _T_15[9:0]) begin
        image_1_570 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_571 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h23b == _T_37[9:0]) begin
        image_1_571 <= io_pixelVal_in_1_7;
      end else if (10'h23b == _T_34[9:0]) begin
        image_1_571 <= io_pixelVal_in_1_6;
      end else if (10'h23b == _T_31[9:0]) begin
        image_1_571 <= io_pixelVal_in_1_5;
      end else if (10'h23b == _T_28[9:0]) begin
        image_1_571 <= io_pixelVal_in_1_4;
      end else if (10'h23b == _T_25[9:0]) begin
        image_1_571 <= io_pixelVal_in_1_3;
      end else if (10'h23b == _T_22[9:0]) begin
        image_1_571 <= io_pixelVal_in_1_2;
      end else if (10'h23b == _T_19[9:0]) begin
        image_1_571 <= io_pixelVal_in_1_1;
      end else if (10'h23b == _T_15[9:0]) begin
        image_1_571 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_572 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h23c == _T_37[9:0]) begin
        image_1_572 <= io_pixelVal_in_1_7;
      end else if (10'h23c == _T_34[9:0]) begin
        image_1_572 <= io_pixelVal_in_1_6;
      end else if (10'h23c == _T_31[9:0]) begin
        image_1_572 <= io_pixelVal_in_1_5;
      end else if (10'h23c == _T_28[9:0]) begin
        image_1_572 <= io_pixelVal_in_1_4;
      end else if (10'h23c == _T_25[9:0]) begin
        image_1_572 <= io_pixelVal_in_1_3;
      end else if (10'h23c == _T_22[9:0]) begin
        image_1_572 <= io_pixelVal_in_1_2;
      end else if (10'h23c == _T_19[9:0]) begin
        image_1_572 <= io_pixelVal_in_1_1;
      end else if (10'h23c == _T_15[9:0]) begin
        image_1_572 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_573 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h23d == _T_37[9:0]) begin
        image_1_573 <= io_pixelVal_in_1_7;
      end else if (10'h23d == _T_34[9:0]) begin
        image_1_573 <= io_pixelVal_in_1_6;
      end else if (10'h23d == _T_31[9:0]) begin
        image_1_573 <= io_pixelVal_in_1_5;
      end else if (10'h23d == _T_28[9:0]) begin
        image_1_573 <= io_pixelVal_in_1_4;
      end else if (10'h23d == _T_25[9:0]) begin
        image_1_573 <= io_pixelVal_in_1_3;
      end else if (10'h23d == _T_22[9:0]) begin
        image_1_573 <= io_pixelVal_in_1_2;
      end else if (10'h23d == _T_19[9:0]) begin
        image_1_573 <= io_pixelVal_in_1_1;
      end else if (10'h23d == _T_15[9:0]) begin
        image_1_573 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_574 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h23e == _T_37[9:0]) begin
        image_1_574 <= io_pixelVal_in_1_7;
      end else if (10'h23e == _T_34[9:0]) begin
        image_1_574 <= io_pixelVal_in_1_6;
      end else if (10'h23e == _T_31[9:0]) begin
        image_1_574 <= io_pixelVal_in_1_5;
      end else if (10'h23e == _T_28[9:0]) begin
        image_1_574 <= io_pixelVal_in_1_4;
      end else if (10'h23e == _T_25[9:0]) begin
        image_1_574 <= io_pixelVal_in_1_3;
      end else if (10'h23e == _T_22[9:0]) begin
        image_1_574 <= io_pixelVal_in_1_2;
      end else if (10'h23e == _T_19[9:0]) begin
        image_1_574 <= io_pixelVal_in_1_1;
      end else if (10'h23e == _T_15[9:0]) begin
        image_1_574 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_1_575 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h23f == _T_37[9:0]) begin
        image_1_575 <= io_pixelVal_in_1_7;
      end else if (10'h23f == _T_34[9:0]) begin
        image_1_575 <= io_pixelVal_in_1_6;
      end else if (10'h23f == _T_31[9:0]) begin
        image_1_575 <= io_pixelVal_in_1_5;
      end else if (10'h23f == _T_28[9:0]) begin
        image_1_575 <= io_pixelVal_in_1_4;
      end else if (10'h23f == _T_25[9:0]) begin
        image_1_575 <= io_pixelVal_in_1_3;
      end else if (10'h23f == _T_22[9:0]) begin
        image_1_575 <= io_pixelVal_in_1_2;
      end else if (10'h23f == _T_19[9:0]) begin
        image_1_575 <= io_pixelVal_in_1_1;
      end else if (10'h23f == _T_15[9:0]) begin
        image_1_575 <= io_pixelVal_in_1_0;
      end
    end
    if (reset) begin
      image_2_0 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h0 == _T_37[9:0]) begin
        image_2_0 <= io_pixelVal_in_2_7;
      end else if (10'h0 == _T_34[9:0]) begin
        image_2_0 <= io_pixelVal_in_2_6;
      end else if (10'h0 == _T_31[9:0]) begin
        image_2_0 <= io_pixelVal_in_2_5;
      end else if (10'h0 == _T_28[9:0]) begin
        image_2_0 <= io_pixelVal_in_2_4;
      end else if (10'h0 == _T_25[9:0]) begin
        image_2_0 <= io_pixelVal_in_2_3;
      end else if (10'h0 == _T_22[9:0]) begin
        image_2_0 <= io_pixelVal_in_2_2;
      end else if (10'h0 == _T_19[9:0]) begin
        image_2_0 <= io_pixelVal_in_2_1;
      end else if (10'h0 == _T_15[9:0]) begin
        image_2_0 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_1 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1 == _T_37[9:0]) begin
        image_2_1 <= io_pixelVal_in_2_7;
      end else if (10'h1 == _T_34[9:0]) begin
        image_2_1 <= io_pixelVal_in_2_6;
      end else if (10'h1 == _T_31[9:0]) begin
        image_2_1 <= io_pixelVal_in_2_5;
      end else if (10'h1 == _T_28[9:0]) begin
        image_2_1 <= io_pixelVal_in_2_4;
      end else if (10'h1 == _T_25[9:0]) begin
        image_2_1 <= io_pixelVal_in_2_3;
      end else if (10'h1 == _T_22[9:0]) begin
        image_2_1 <= io_pixelVal_in_2_2;
      end else if (10'h1 == _T_19[9:0]) begin
        image_2_1 <= io_pixelVal_in_2_1;
      end else if (10'h1 == _T_15[9:0]) begin
        image_2_1 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_2 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h2 == _T_37[9:0]) begin
        image_2_2 <= io_pixelVal_in_2_7;
      end else if (10'h2 == _T_34[9:0]) begin
        image_2_2 <= io_pixelVal_in_2_6;
      end else if (10'h2 == _T_31[9:0]) begin
        image_2_2 <= io_pixelVal_in_2_5;
      end else if (10'h2 == _T_28[9:0]) begin
        image_2_2 <= io_pixelVal_in_2_4;
      end else if (10'h2 == _T_25[9:0]) begin
        image_2_2 <= io_pixelVal_in_2_3;
      end else if (10'h2 == _T_22[9:0]) begin
        image_2_2 <= io_pixelVal_in_2_2;
      end else if (10'h2 == _T_19[9:0]) begin
        image_2_2 <= io_pixelVal_in_2_1;
      end else if (10'h2 == _T_15[9:0]) begin
        image_2_2 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_3 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h3 == _T_37[9:0]) begin
        image_2_3 <= io_pixelVal_in_2_7;
      end else if (10'h3 == _T_34[9:0]) begin
        image_2_3 <= io_pixelVal_in_2_6;
      end else if (10'h3 == _T_31[9:0]) begin
        image_2_3 <= io_pixelVal_in_2_5;
      end else if (10'h3 == _T_28[9:0]) begin
        image_2_3 <= io_pixelVal_in_2_4;
      end else if (10'h3 == _T_25[9:0]) begin
        image_2_3 <= io_pixelVal_in_2_3;
      end else if (10'h3 == _T_22[9:0]) begin
        image_2_3 <= io_pixelVal_in_2_2;
      end else if (10'h3 == _T_19[9:0]) begin
        image_2_3 <= io_pixelVal_in_2_1;
      end else if (10'h3 == _T_15[9:0]) begin
        image_2_3 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_4 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h4 == _T_37[9:0]) begin
        image_2_4 <= io_pixelVal_in_2_7;
      end else if (10'h4 == _T_34[9:0]) begin
        image_2_4 <= io_pixelVal_in_2_6;
      end else if (10'h4 == _T_31[9:0]) begin
        image_2_4 <= io_pixelVal_in_2_5;
      end else if (10'h4 == _T_28[9:0]) begin
        image_2_4 <= io_pixelVal_in_2_4;
      end else if (10'h4 == _T_25[9:0]) begin
        image_2_4 <= io_pixelVal_in_2_3;
      end else if (10'h4 == _T_22[9:0]) begin
        image_2_4 <= io_pixelVal_in_2_2;
      end else if (10'h4 == _T_19[9:0]) begin
        image_2_4 <= io_pixelVal_in_2_1;
      end else if (10'h4 == _T_15[9:0]) begin
        image_2_4 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_5 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h5 == _T_37[9:0]) begin
        image_2_5 <= io_pixelVal_in_2_7;
      end else if (10'h5 == _T_34[9:0]) begin
        image_2_5 <= io_pixelVal_in_2_6;
      end else if (10'h5 == _T_31[9:0]) begin
        image_2_5 <= io_pixelVal_in_2_5;
      end else if (10'h5 == _T_28[9:0]) begin
        image_2_5 <= io_pixelVal_in_2_4;
      end else if (10'h5 == _T_25[9:0]) begin
        image_2_5 <= io_pixelVal_in_2_3;
      end else if (10'h5 == _T_22[9:0]) begin
        image_2_5 <= io_pixelVal_in_2_2;
      end else if (10'h5 == _T_19[9:0]) begin
        image_2_5 <= io_pixelVal_in_2_1;
      end else if (10'h5 == _T_15[9:0]) begin
        image_2_5 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_6 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h6 == _T_37[9:0]) begin
        image_2_6 <= io_pixelVal_in_2_7;
      end else if (10'h6 == _T_34[9:0]) begin
        image_2_6 <= io_pixelVal_in_2_6;
      end else if (10'h6 == _T_31[9:0]) begin
        image_2_6 <= io_pixelVal_in_2_5;
      end else if (10'h6 == _T_28[9:0]) begin
        image_2_6 <= io_pixelVal_in_2_4;
      end else if (10'h6 == _T_25[9:0]) begin
        image_2_6 <= io_pixelVal_in_2_3;
      end else if (10'h6 == _T_22[9:0]) begin
        image_2_6 <= io_pixelVal_in_2_2;
      end else if (10'h6 == _T_19[9:0]) begin
        image_2_6 <= io_pixelVal_in_2_1;
      end else if (10'h6 == _T_15[9:0]) begin
        image_2_6 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_7 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h7 == _T_37[9:0]) begin
        image_2_7 <= io_pixelVal_in_2_7;
      end else if (10'h7 == _T_34[9:0]) begin
        image_2_7 <= io_pixelVal_in_2_6;
      end else if (10'h7 == _T_31[9:0]) begin
        image_2_7 <= io_pixelVal_in_2_5;
      end else if (10'h7 == _T_28[9:0]) begin
        image_2_7 <= io_pixelVal_in_2_4;
      end else if (10'h7 == _T_25[9:0]) begin
        image_2_7 <= io_pixelVal_in_2_3;
      end else if (10'h7 == _T_22[9:0]) begin
        image_2_7 <= io_pixelVal_in_2_2;
      end else if (10'h7 == _T_19[9:0]) begin
        image_2_7 <= io_pixelVal_in_2_1;
      end else if (10'h7 == _T_15[9:0]) begin
        image_2_7 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_8 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h8 == _T_37[9:0]) begin
        image_2_8 <= io_pixelVal_in_2_7;
      end else if (10'h8 == _T_34[9:0]) begin
        image_2_8 <= io_pixelVal_in_2_6;
      end else if (10'h8 == _T_31[9:0]) begin
        image_2_8 <= io_pixelVal_in_2_5;
      end else if (10'h8 == _T_28[9:0]) begin
        image_2_8 <= io_pixelVal_in_2_4;
      end else if (10'h8 == _T_25[9:0]) begin
        image_2_8 <= io_pixelVal_in_2_3;
      end else if (10'h8 == _T_22[9:0]) begin
        image_2_8 <= io_pixelVal_in_2_2;
      end else if (10'h8 == _T_19[9:0]) begin
        image_2_8 <= io_pixelVal_in_2_1;
      end else if (10'h8 == _T_15[9:0]) begin
        image_2_8 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_9 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h9 == _T_37[9:0]) begin
        image_2_9 <= io_pixelVal_in_2_7;
      end else if (10'h9 == _T_34[9:0]) begin
        image_2_9 <= io_pixelVal_in_2_6;
      end else if (10'h9 == _T_31[9:0]) begin
        image_2_9 <= io_pixelVal_in_2_5;
      end else if (10'h9 == _T_28[9:0]) begin
        image_2_9 <= io_pixelVal_in_2_4;
      end else if (10'h9 == _T_25[9:0]) begin
        image_2_9 <= io_pixelVal_in_2_3;
      end else if (10'h9 == _T_22[9:0]) begin
        image_2_9 <= io_pixelVal_in_2_2;
      end else if (10'h9 == _T_19[9:0]) begin
        image_2_9 <= io_pixelVal_in_2_1;
      end else if (10'h9 == _T_15[9:0]) begin
        image_2_9 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_10 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha == _T_37[9:0]) begin
        image_2_10 <= io_pixelVal_in_2_7;
      end else if (10'ha == _T_34[9:0]) begin
        image_2_10 <= io_pixelVal_in_2_6;
      end else if (10'ha == _T_31[9:0]) begin
        image_2_10 <= io_pixelVal_in_2_5;
      end else if (10'ha == _T_28[9:0]) begin
        image_2_10 <= io_pixelVal_in_2_4;
      end else if (10'ha == _T_25[9:0]) begin
        image_2_10 <= io_pixelVal_in_2_3;
      end else if (10'ha == _T_22[9:0]) begin
        image_2_10 <= io_pixelVal_in_2_2;
      end else if (10'ha == _T_19[9:0]) begin
        image_2_10 <= io_pixelVal_in_2_1;
      end else if (10'ha == _T_15[9:0]) begin
        image_2_10 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_11 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb == _T_37[9:0]) begin
        image_2_11 <= io_pixelVal_in_2_7;
      end else if (10'hb == _T_34[9:0]) begin
        image_2_11 <= io_pixelVal_in_2_6;
      end else if (10'hb == _T_31[9:0]) begin
        image_2_11 <= io_pixelVal_in_2_5;
      end else if (10'hb == _T_28[9:0]) begin
        image_2_11 <= io_pixelVal_in_2_4;
      end else if (10'hb == _T_25[9:0]) begin
        image_2_11 <= io_pixelVal_in_2_3;
      end else if (10'hb == _T_22[9:0]) begin
        image_2_11 <= io_pixelVal_in_2_2;
      end else if (10'hb == _T_19[9:0]) begin
        image_2_11 <= io_pixelVal_in_2_1;
      end else if (10'hb == _T_15[9:0]) begin
        image_2_11 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_12 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc == _T_37[9:0]) begin
        image_2_12 <= io_pixelVal_in_2_7;
      end else if (10'hc == _T_34[9:0]) begin
        image_2_12 <= io_pixelVal_in_2_6;
      end else if (10'hc == _T_31[9:0]) begin
        image_2_12 <= io_pixelVal_in_2_5;
      end else if (10'hc == _T_28[9:0]) begin
        image_2_12 <= io_pixelVal_in_2_4;
      end else if (10'hc == _T_25[9:0]) begin
        image_2_12 <= io_pixelVal_in_2_3;
      end else if (10'hc == _T_22[9:0]) begin
        image_2_12 <= io_pixelVal_in_2_2;
      end else if (10'hc == _T_19[9:0]) begin
        image_2_12 <= io_pixelVal_in_2_1;
      end else if (10'hc == _T_15[9:0]) begin
        image_2_12 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_13 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd == _T_37[9:0]) begin
        image_2_13 <= io_pixelVal_in_2_7;
      end else if (10'hd == _T_34[9:0]) begin
        image_2_13 <= io_pixelVal_in_2_6;
      end else if (10'hd == _T_31[9:0]) begin
        image_2_13 <= io_pixelVal_in_2_5;
      end else if (10'hd == _T_28[9:0]) begin
        image_2_13 <= io_pixelVal_in_2_4;
      end else if (10'hd == _T_25[9:0]) begin
        image_2_13 <= io_pixelVal_in_2_3;
      end else if (10'hd == _T_22[9:0]) begin
        image_2_13 <= io_pixelVal_in_2_2;
      end else if (10'hd == _T_19[9:0]) begin
        image_2_13 <= io_pixelVal_in_2_1;
      end else if (10'hd == _T_15[9:0]) begin
        image_2_13 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_14 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he == _T_37[9:0]) begin
        image_2_14 <= io_pixelVal_in_2_7;
      end else if (10'he == _T_34[9:0]) begin
        image_2_14 <= io_pixelVal_in_2_6;
      end else if (10'he == _T_31[9:0]) begin
        image_2_14 <= io_pixelVal_in_2_5;
      end else if (10'he == _T_28[9:0]) begin
        image_2_14 <= io_pixelVal_in_2_4;
      end else if (10'he == _T_25[9:0]) begin
        image_2_14 <= io_pixelVal_in_2_3;
      end else if (10'he == _T_22[9:0]) begin
        image_2_14 <= io_pixelVal_in_2_2;
      end else if (10'he == _T_19[9:0]) begin
        image_2_14 <= io_pixelVal_in_2_1;
      end else if (10'he == _T_15[9:0]) begin
        image_2_14 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_15 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf == _T_37[9:0]) begin
        image_2_15 <= io_pixelVal_in_2_7;
      end else if (10'hf == _T_34[9:0]) begin
        image_2_15 <= io_pixelVal_in_2_6;
      end else if (10'hf == _T_31[9:0]) begin
        image_2_15 <= io_pixelVal_in_2_5;
      end else if (10'hf == _T_28[9:0]) begin
        image_2_15 <= io_pixelVal_in_2_4;
      end else if (10'hf == _T_25[9:0]) begin
        image_2_15 <= io_pixelVal_in_2_3;
      end else if (10'hf == _T_22[9:0]) begin
        image_2_15 <= io_pixelVal_in_2_2;
      end else if (10'hf == _T_19[9:0]) begin
        image_2_15 <= io_pixelVal_in_2_1;
      end else if (10'hf == _T_15[9:0]) begin
        image_2_15 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_16 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h10 == _T_37[9:0]) begin
        image_2_16 <= io_pixelVal_in_2_7;
      end else if (10'h10 == _T_34[9:0]) begin
        image_2_16 <= io_pixelVal_in_2_6;
      end else if (10'h10 == _T_31[9:0]) begin
        image_2_16 <= io_pixelVal_in_2_5;
      end else if (10'h10 == _T_28[9:0]) begin
        image_2_16 <= io_pixelVal_in_2_4;
      end else if (10'h10 == _T_25[9:0]) begin
        image_2_16 <= io_pixelVal_in_2_3;
      end else if (10'h10 == _T_22[9:0]) begin
        image_2_16 <= io_pixelVal_in_2_2;
      end else if (10'h10 == _T_19[9:0]) begin
        image_2_16 <= io_pixelVal_in_2_1;
      end else if (10'h10 == _T_15[9:0]) begin
        image_2_16 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_17 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h11 == _T_37[9:0]) begin
        image_2_17 <= io_pixelVal_in_2_7;
      end else if (10'h11 == _T_34[9:0]) begin
        image_2_17 <= io_pixelVal_in_2_6;
      end else if (10'h11 == _T_31[9:0]) begin
        image_2_17 <= io_pixelVal_in_2_5;
      end else if (10'h11 == _T_28[9:0]) begin
        image_2_17 <= io_pixelVal_in_2_4;
      end else if (10'h11 == _T_25[9:0]) begin
        image_2_17 <= io_pixelVal_in_2_3;
      end else if (10'h11 == _T_22[9:0]) begin
        image_2_17 <= io_pixelVal_in_2_2;
      end else if (10'h11 == _T_19[9:0]) begin
        image_2_17 <= io_pixelVal_in_2_1;
      end else if (10'h11 == _T_15[9:0]) begin
        image_2_17 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_18 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h12 == _T_37[9:0]) begin
        image_2_18 <= io_pixelVal_in_2_7;
      end else if (10'h12 == _T_34[9:0]) begin
        image_2_18 <= io_pixelVal_in_2_6;
      end else if (10'h12 == _T_31[9:0]) begin
        image_2_18 <= io_pixelVal_in_2_5;
      end else if (10'h12 == _T_28[9:0]) begin
        image_2_18 <= io_pixelVal_in_2_4;
      end else if (10'h12 == _T_25[9:0]) begin
        image_2_18 <= io_pixelVal_in_2_3;
      end else if (10'h12 == _T_22[9:0]) begin
        image_2_18 <= io_pixelVal_in_2_2;
      end else if (10'h12 == _T_19[9:0]) begin
        image_2_18 <= io_pixelVal_in_2_1;
      end else if (10'h12 == _T_15[9:0]) begin
        image_2_18 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_19 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h13 == _T_37[9:0]) begin
        image_2_19 <= io_pixelVal_in_2_7;
      end else if (10'h13 == _T_34[9:0]) begin
        image_2_19 <= io_pixelVal_in_2_6;
      end else if (10'h13 == _T_31[9:0]) begin
        image_2_19 <= io_pixelVal_in_2_5;
      end else if (10'h13 == _T_28[9:0]) begin
        image_2_19 <= io_pixelVal_in_2_4;
      end else if (10'h13 == _T_25[9:0]) begin
        image_2_19 <= io_pixelVal_in_2_3;
      end else if (10'h13 == _T_22[9:0]) begin
        image_2_19 <= io_pixelVal_in_2_2;
      end else if (10'h13 == _T_19[9:0]) begin
        image_2_19 <= io_pixelVal_in_2_1;
      end else if (10'h13 == _T_15[9:0]) begin
        image_2_19 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_20 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h14 == _T_37[9:0]) begin
        image_2_20 <= io_pixelVal_in_2_7;
      end else if (10'h14 == _T_34[9:0]) begin
        image_2_20 <= io_pixelVal_in_2_6;
      end else if (10'h14 == _T_31[9:0]) begin
        image_2_20 <= io_pixelVal_in_2_5;
      end else if (10'h14 == _T_28[9:0]) begin
        image_2_20 <= io_pixelVal_in_2_4;
      end else if (10'h14 == _T_25[9:0]) begin
        image_2_20 <= io_pixelVal_in_2_3;
      end else if (10'h14 == _T_22[9:0]) begin
        image_2_20 <= io_pixelVal_in_2_2;
      end else if (10'h14 == _T_19[9:0]) begin
        image_2_20 <= io_pixelVal_in_2_1;
      end else if (10'h14 == _T_15[9:0]) begin
        image_2_20 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_21 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h15 == _T_37[9:0]) begin
        image_2_21 <= io_pixelVal_in_2_7;
      end else if (10'h15 == _T_34[9:0]) begin
        image_2_21 <= io_pixelVal_in_2_6;
      end else if (10'h15 == _T_31[9:0]) begin
        image_2_21 <= io_pixelVal_in_2_5;
      end else if (10'h15 == _T_28[9:0]) begin
        image_2_21 <= io_pixelVal_in_2_4;
      end else if (10'h15 == _T_25[9:0]) begin
        image_2_21 <= io_pixelVal_in_2_3;
      end else if (10'h15 == _T_22[9:0]) begin
        image_2_21 <= io_pixelVal_in_2_2;
      end else if (10'h15 == _T_19[9:0]) begin
        image_2_21 <= io_pixelVal_in_2_1;
      end else if (10'h15 == _T_15[9:0]) begin
        image_2_21 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_22 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h16 == _T_37[9:0]) begin
        image_2_22 <= io_pixelVal_in_2_7;
      end else if (10'h16 == _T_34[9:0]) begin
        image_2_22 <= io_pixelVal_in_2_6;
      end else if (10'h16 == _T_31[9:0]) begin
        image_2_22 <= io_pixelVal_in_2_5;
      end else if (10'h16 == _T_28[9:0]) begin
        image_2_22 <= io_pixelVal_in_2_4;
      end else if (10'h16 == _T_25[9:0]) begin
        image_2_22 <= io_pixelVal_in_2_3;
      end else if (10'h16 == _T_22[9:0]) begin
        image_2_22 <= io_pixelVal_in_2_2;
      end else if (10'h16 == _T_19[9:0]) begin
        image_2_22 <= io_pixelVal_in_2_1;
      end else if (10'h16 == _T_15[9:0]) begin
        image_2_22 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_23 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h17 == _T_37[9:0]) begin
        image_2_23 <= io_pixelVal_in_2_7;
      end else if (10'h17 == _T_34[9:0]) begin
        image_2_23 <= io_pixelVal_in_2_6;
      end else if (10'h17 == _T_31[9:0]) begin
        image_2_23 <= io_pixelVal_in_2_5;
      end else if (10'h17 == _T_28[9:0]) begin
        image_2_23 <= io_pixelVal_in_2_4;
      end else if (10'h17 == _T_25[9:0]) begin
        image_2_23 <= io_pixelVal_in_2_3;
      end else if (10'h17 == _T_22[9:0]) begin
        image_2_23 <= io_pixelVal_in_2_2;
      end else if (10'h17 == _T_19[9:0]) begin
        image_2_23 <= io_pixelVal_in_2_1;
      end else if (10'h17 == _T_15[9:0]) begin
        image_2_23 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_24 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h18 == _T_37[9:0]) begin
        image_2_24 <= io_pixelVal_in_2_7;
      end else if (10'h18 == _T_34[9:0]) begin
        image_2_24 <= io_pixelVal_in_2_6;
      end else if (10'h18 == _T_31[9:0]) begin
        image_2_24 <= io_pixelVal_in_2_5;
      end else if (10'h18 == _T_28[9:0]) begin
        image_2_24 <= io_pixelVal_in_2_4;
      end else if (10'h18 == _T_25[9:0]) begin
        image_2_24 <= io_pixelVal_in_2_3;
      end else if (10'h18 == _T_22[9:0]) begin
        image_2_24 <= io_pixelVal_in_2_2;
      end else if (10'h18 == _T_19[9:0]) begin
        image_2_24 <= io_pixelVal_in_2_1;
      end else if (10'h18 == _T_15[9:0]) begin
        image_2_24 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_25 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h19 == _T_37[9:0]) begin
        image_2_25 <= io_pixelVal_in_2_7;
      end else if (10'h19 == _T_34[9:0]) begin
        image_2_25 <= io_pixelVal_in_2_6;
      end else if (10'h19 == _T_31[9:0]) begin
        image_2_25 <= io_pixelVal_in_2_5;
      end else if (10'h19 == _T_28[9:0]) begin
        image_2_25 <= io_pixelVal_in_2_4;
      end else if (10'h19 == _T_25[9:0]) begin
        image_2_25 <= io_pixelVal_in_2_3;
      end else if (10'h19 == _T_22[9:0]) begin
        image_2_25 <= io_pixelVal_in_2_2;
      end else if (10'h19 == _T_19[9:0]) begin
        image_2_25 <= io_pixelVal_in_2_1;
      end else if (10'h19 == _T_15[9:0]) begin
        image_2_25 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_26 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a == _T_37[9:0]) begin
        image_2_26 <= io_pixelVal_in_2_7;
      end else if (10'h1a == _T_34[9:0]) begin
        image_2_26 <= io_pixelVal_in_2_6;
      end else if (10'h1a == _T_31[9:0]) begin
        image_2_26 <= io_pixelVal_in_2_5;
      end else if (10'h1a == _T_28[9:0]) begin
        image_2_26 <= io_pixelVal_in_2_4;
      end else if (10'h1a == _T_25[9:0]) begin
        image_2_26 <= io_pixelVal_in_2_3;
      end else if (10'h1a == _T_22[9:0]) begin
        image_2_26 <= io_pixelVal_in_2_2;
      end else if (10'h1a == _T_19[9:0]) begin
        image_2_26 <= io_pixelVal_in_2_1;
      end else if (10'h1a == _T_15[9:0]) begin
        image_2_26 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_27 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b == _T_37[9:0]) begin
        image_2_27 <= io_pixelVal_in_2_7;
      end else if (10'h1b == _T_34[9:0]) begin
        image_2_27 <= io_pixelVal_in_2_6;
      end else if (10'h1b == _T_31[9:0]) begin
        image_2_27 <= io_pixelVal_in_2_5;
      end else if (10'h1b == _T_28[9:0]) begin
        image_2_27 <= io_pixelVal_in_2_4;
      end else if (10'h1b == _T_25[9:0]) begin
        image_2_27 <= io_pixelVal_in_2_3;
      end else if (10'h1b == _T_22[9:0]) begin
        image_2_27 <= io_pixelVal_in_2_2;
      end else if (10'h1b == _T_19[9:0]) begin
        image_2_27 <= io_pixelVal_in_2_1;
      end else if (10'h1b == _T_15[9:0]) begin
        image_2_27 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_28 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c == _T_37[9:0]) begin
        image_2_28 <= io_pixelVal_in_2_7;
      end else if (10'h1c == _T_34[9:0]) begin
        image_2_28 <= io_pixelVal_in_2_6;
      end else if (10'h1c == _T_31[9:0]) begin
        image_2_28 <= io_pixelVal_in_2_5;
      end else if (10'h1c == _T_28[9:0]) begin
        image_2_28 <= io_pixelVal_in_2_4;
      end else if (10'h1c == _T_25[9:0]) begin
        image_2_28 <= io_pixelVal_in_2_3;
      end else if (10'h1c == _T_22[9:0]) begin
        image_2_28 <= io_pixelVal_in_2_2;
      end else if (10'h1c == _T_19[9:0]) begin
        image_2_28 <= io_pixelVal_in_2_1;
      end else if (10'h1c == _T_15[9:0]) begin
        image_2_28 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_29 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d == _T_37[9:0]) begin
        image_2_29 <= io_pixelVal_in_2_7;
      end else if (10'h1d == _T_34[9:0]) begin
        image_2_29 <= io_pixelVal_in_2_6;
      end else if (10'h1d == _T_31[9:0]) begin
        image_2_29 <= io_pixelVal_in_2_5;
      end else if (10'h1d == _T_28[9:0]) begin
        image_2_29 <= io_pixelVal_in_2_4;
      end else if (10'h1d == _T_25[9:0]) begin
        image_2_29 <= io_pixelVal_in_2_3;
      end else if (10'h1d == _T_22[9:0]) begin
        image_2_29 <= io_pixelVal_in_2_2;
      end else if (10'h1d == _T_19[9:0]) begin
        image_2_29 <= io_pixelVal_in_2_1;
      end else if (10'h1d == _T_15[9:0]) begin
        image_2_29 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_30 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e == _T_37[9:0]) begin
        image_2_30 <= io_pixelVal_in_2_7;
      end else if (10'h1e == _T_34[9:0]) begin
        image_2_30 <= io_pixelVal_in_2_6;
      end else if (10'h1e == _T_31[9:0]) begin
        image_2_30 <= io_pixelVal_in_2_5;
      end else if (10'h1e == _T_28[9:0]) begin
        image_2_30 <= io_pixelVal_in_2_4;
      end else if (10'h1e == _T_25[9:0]) begin
        image_2_30 <= io_pixelVal_in_2_3;
      end else if (10'h1e == _T_22[9:0]) begin
        image_2_30 <= io_pixelVal_in_2_2;
      end else if (10'h1e == _T_19[9:0]) begin
        image_2_30 <= io_pixelVal_in_2_1;
      end else if (10'h1e == _T_15[9:0]) begin
        image_2_30 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_31 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f == _T_37[9:0]) begin
        image_2_31 <= io_pixelVal_in_2_7;
      end else if (10'h1f == _T_34[9:0]) begin
        image_2_31 <= io_pixelVal_in_2_6;
      end else if (10'h1f == _T_31[9:0]) begin
        image_2_31 <= io_pixelVal_in_2_5;
      end else if (10'h1f == _T_28[9:0]) begin
        image_2_31 <= io_pixelVal_in_2_4;
      end else if (10'h1f == _T_25[9:0]) begin
        image_2_31 <= io_pixelVal_in_2_3;
      end else if (10'h1f == _T_22[9:0]) begin
        image_2_31 <= io_pixelVal_in_2_2;
      end else if (10'h1f == _T_19[9:0]) begin
        image_2_31 <= io_pixelVal_in_2_1;
      end else if (10'h1f == _T_15[9:0]) begin
        image_2_31 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_32 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h20 == _T_37[9:0]) begin
        image_2_32 <= io_pixelVal_in_2_7;
      end else if (10'h20 == _T_34[9:0]) begin
        image_2_32 <= io_pixelVal_in_2_6;
      end else if (10'h20 == _T_31[9:0]) begin
        image_2_32 <= io_pixelVal_in_2_5;
      end else if (10'h20 == _T_28[9:0]) begin
        image_2_32 <= io_pixelVal_in_2_4;
      end else if (10'h20 == _T_25[9:0]) begin
        image_2_32 <= io_pixelVal_in_2_3;
      end else if (10'h20 == _T_22[9:0]) begin
        image_2_32 <= io_pixelVal_in_2_2;
      end else if (10'h20 == _T_19[9:0]) begin
        image_2_32 <= io_pixelVal_in_2_1;
      end else if (10'h20 == _T_15[9:0]) begin
        image_2_32 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_33 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h21 == _T_37[9:0]) begin
        image_2_33 <= io_pixelVal_in_2_7;
      end else if (10'h21 == _T_34[9:0]) begin
        image_2_33 <= io_pixelVal_in_2_6;
      end else if (10'h21 == _T_31[9:0]) begin
        image_2_33 <= io_pixelVal_in_2_5;
      end else if (10'h21 == _T_28[9:0]) begin
        image_2_33 <= io_pixelVal_in_2_4;
      end else if (10'h21 == _T_25[9:0]) begin
        image_2_33 <= io_pixelVal_in_2_3;
      end else if (10'h21 == _T_22[9:0]) begin
        image_2_33 <= io_pixelVal_in_2_2;
      end else if (10'h21 == _T_19[9:0]) begin
        image_2_33 <= io_pixelVal_in_2_1;
      end else if (10'h21 == _T_15[9:0]) begin
        image_2_33 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_34 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h22 == _T_37[9:0]) begin
        image_2_34 <= io_pixelVal_in_2_7;
      end else if (10'h22 == _T_34[9:0]) begin
        image_2_34 <= io_pixelVal_in_2_6;
      end else if (10'h22 == _T_31[9:0]) begin
        image_2_34 <= io_pixelVal_in_2_5;
      end else if (10'h22 == _T_28[9:0]) begin
        image_2_34 <= io_pixelVal_in_2_4;
      end else if (10'h22 == _T_25[9:0]) begin
        image_2_34 <= io_pixelVal_in_2_3;
      end else if (10'h22 == _T_22[9:0]) begin
        image_2_34 <= io_pixelVal_in_2_2;
      end else if (10'h22 == _T_19[9:0]) begin
        image_2_34 <= io_pixelVal_in_2_1;
      end else if (10'h22 == _T_15[9:0]) begin
        image_2_34 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_35 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h23 == _T_37[9:0]) begin
        image_2_35 <= io_pixelVal_in_2_7;
      end else if (10'h23 == _T_34[9:0]) begin
        image_2_35 <= io_pixelVal_in_2_6;
      end else if (10'h23 == _T_31[9:0]) begin
        image_2_35 <= io_pixelVal_in_2_5;
      end else if (10'h23 == _T_28[9:0]) begin
        image_2_35 <= io_pixelVal_in_2_4;
      end else if (10'h23 == _T_25[9:0]) begin
        image_2_35 <= io_pixelVal_in_2_3;
      end else if (10'h23 == _T_22[9:0]) begin
        image_2_35 <= io_pixelVal_in_2_2;
      end else if (10'h23 == _T_19[9:0]) begin
        image_2_35 <= io_pixelVal_in_2_1;
      end else if (10'h23 == _T_15[9:0]) begin
        image_2_35 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_36 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h24 == _T_37[9:0]) begin
        image_2_36 <= io_pixelVal_in_2_7;
      end else if (10'h24 == _T_34[9:0]) begin
        image_2_36 <= io_pixelVal_in_2_6;
      end else if (10'h24 == _T_31[9:0]) begin
        image_2_36 <= io_pixelVal_in_2_5;
      end else if (10'h24 == _T_28[9:0]) begin
        image_2_36 <= io_pixelVal_in_2_4;
      end else if (10'h24 == _T_25[9:0]) begin
        image_2_36 <= io_pixelVal_in_2_3;
      end else if (10'h24 == _T_22[9:0]) begin
        image_2_36 <= io_pixelVal_in_2_2;
      end else if (10'h24 == _T_19[9:0]) begin
        image_2_36 <= io_pixelVal_in_2_1;
      end else if (10'h24 == _T_15[9:0]) begin
        image_2_36 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_37 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h25 == _T_37[9:0]) begin
        image_2_37 <= io_pixelVal_in_2_7;
      end else if (10'h25 == _T_34[9:0]) begin
        image_2_37 <= io_pixelVal_in_2_6;
      end else if (10'h25 == _T_31[9:0]) begin
        image_2_37 <= io_pixelVal_in_2_5;
      end else if (10'h25 == _T_28[9:0]) begin
        image_2_37 <= io_pixelVal_in_2_4;
      end else if (10'h25 == _T_25[9:0]) begin
        image_2_37 <= io_pixelVal_in_2_3;
      end else if (10'h25 == _T_22[9:0]) begin
        image_2_37 <= io_pixelVal_in_2_2;
      end else if (10'h25 == _T_19[9:0]) begin
        image_2_37 <= io_pixelVal_in_2_1;
      end else if (10'h25 == _T_15[9:0]) begin
        image_2_37 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_38 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h26 == _T_37[9:0]) begin
        image_2_38 <= io_pixelVal_in_2_7;
      end else if (10'h26 == _T_34[9:0]) begin
        image_2_38 <= io_pixelVal_in_2_6;
      end else if (10'h26 == _T_31[9:0]) begin
        image_2_38 <= io_pixelVal_in_2_5;
      end else if (10'h26 == _T_28[9:0]) begin
        image_2_38 <= io_pixelVal_in_2_4;
      end else if (10'h26 == _T_25[9:0]) begin
        image_2_38 <= io_pixelVal_in_2_3;
      end else if (10'h26 == _T_22[9:0]) begin
        image_2_38 <= io_pixelVal_in_2_2;
      end else if (10'h26 == _T_19[9:0]) begin
        image_2_38 <= io_pixelVal_in_2_1;
      end else if (10'h26 == _T_15[9:0]) begin
        image_2_38 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_39 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h27 == _T_37[9:0]) begin
        image_2_39 <= io_pixelVal_in_2_7;
      end else if (10'h27 == _T_34[9:0]) begin
        image_2_39 <= io_pixelVal_in_2_6;
      end else if (10'h27 == _T_31[9:0]) begin
        image_2_39 <= io_pixelVal_in_2_5;
      end else if (10'h27 == _T_28[9:0]) begin
        image_2_39 <= io_pixelVal_in_2_4;
      end else if (10'h27 == _T_25[9:0]) begin
        image_2_39 <= io_pixelVal_in_2_3;
      end else if (10'h27 == _T_22[9:0]) begin
        image_2_39 <= io_pixelVal_in_2_2;
      end else if (10'h27 == _T_19[9:0]) begin
        image_2_39 <= io_pixelVal_in_2_1;
      end else if (10'h27 == _T_15[9:0]) begin
        image_2_39 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_40 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h28 == _T_37[9:0]) begin
        image_2_40 <= io_pixelVal_in_2_7;
      end else if (10'h28 == _T_34[9:0]) begin
        image_2_40 <= io_pixelVal_in_2_6;
      end else if (10'h28 == _T_31[9:0]) begin
        image_2_40 <= io_pixelVal_in_2_5;
      end else if (10'h28 == _T_28[9:0]) begin
        image_2_40 <= io_pixelVal_in_2_4;
      end else if (10'h28 == _T_25[9:0]) begin
        image_2_40 <= io_pixelVal_in_2_3;
      end else if (10'h28 == _T_22[9:0]) begin
        image_2_40 <= io_pixelVal_in_2_2;
      end else if (10'h28 == _T_19[9:0]) begin
        image_2_40 <= io_pixelVal_in_2_1;
      end else if (10'h28 == _T_15[9:0]) begin
        image_2_40 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_41 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h29 == _T_37[9:0]) begin
        image_2_41 <= io_pixelVal_in_2_7;
      end else if (10'h29 == _T_34[9:0]) begin
        image_2_41 <= io_pixelVal_in_2_6;
      end else if (10'h29 == _T_31[9:0]) begin
        image_2_41 <= io_pixelVal_in_2_5;
      end else if (10'h29 == _T_28[9:0]) begin
        image_2_41 <= io_pixelVal_in_2_4;
      end else if (10'h29 == _T_25[9:0]) begin
        image_2_41 <= io_pixelVal_in_2_3;
      end else if (10'h29 == _T_22[9:0]) begin
        image_2_41 <= io_pixelVal_in_2_2;
      end else if (10'h29 == _T_19[9:0]) begin
        image_2_41 <= io_pixelVal_in_2_1;
      end else if (10'h29 == _T_15[9:0]) begin
        image_2_41 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_42 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h2a == _T_37[9:0]) begin
        image_2_42 <= io_pixelVal_in_2_7;
      end else if (10'h2a == _T_34[9:0]) begin
        image_2_42 <= io_pixelVal_in_2_6;
      end else if (10'h2a == _T_31[9:0]) begin
        image_2_42 <= io_pixelVal_in_2_5;
      end else if (10'h2a == _T_28[9:0]) begin
        image_2_42 <= io_pixelVal_in_2_4;
      end else if (10'h2a == _T_25[9:0]) begin
        image_2_42 <= io_pixelVal_in_2_3;
      end else if (10'h2a == _T_22[9:0]) begin
        image_2_42 <= io_pixelVal_in_2_2;
      end else if (10'h2a == _T_19[9:0]) begin
        image_2_42 <= io_pixelVal_in_2_1;
      end else if (10'h2a == _T_15[9:0]) begin
        image_2_42 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_43 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h2b == _T_37[9:0]) begin
        image_2_43 <= io_pixelVal_in_2_7;
      end else if (10'h2b == _T_34[9:0]) begin
        image_2_43 <= io_pixelVal_in_2_6;
      end else if (10'h2b == _T_31[9:0]) begin
        image_2_43 <= io_pixelVal_in_2_5;
      end else if (10'h2b == _T_28[9:0]) begin
        image_2_43 <= io_pixelVal_in_2_4;
      end else if (10'h2b == _T_25[9:0]) begin
        image_2_43 <= io_pixelVal_in_2_3;
      end else if (10'h2b == _T_22[9:0]) begin
        image_2_43 <= io_pixelVal_in_2_2;
      end else if (10'h2b == _T_19[9:0]) begin
        image_2_43 <= io_pixelVal_in_2_1;
      end else if (10'h2b == _T_15[9:0]) begin
        image_2_43 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_44 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h2c == _T_37[9:0]) begin
        image_2_44 <= io_pixelVal_in_2_7;
      end else if (10'h2c == _T_34[9:0]) begin
        image_2_44 <= io_pixelVal_in_2_6;
      end else if (10'h2c == _T_31[9:0]) begin
        image_2_44 <= io_pixelVal_in_2_5;
      end else if (10'h2c == _T_28[9:0]) begin
        image_2_44 <= io_pixelVal_in_2_4;
      end else if (10'h2c == _T_25[9:0]) begin
        image_2_44 <= io_pixelVal_in_2_3;
      end else if (10'h2c == _T_22[9:0]) begin
        image_2_44 <= io_pixelVal_in_2_2;
      end else if (10'h2c == _T_19[9:0]) begin
        image_2_44 <= io_pixelVal_in_2_1;
      end else if (10'h2c == _T_15[9:0]) begin
        image_2_44 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_45 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h2d == _T_37[9:0]) begin
        image_2_45 <= io_pixelVal_in_2_7;
      end else if (10'h2d == _T_34[9:0]) begin
        image_2_45 <= io_pixelVal_in_2_6;
      end else if (10'h2d == _T_31[9:0]) begin
        image_2_45 <= io_pixelVal_in_2_5;
      end else if (10'h2d == _T_28[9:0]) begin
        image_2_45 <= io_pixelVal_in_2_4;
      end else if (10'h2d == _T_25[9:0]) begin
        image_2_45 <= io_pixelVal_in_2_3;
      end else if (10'h2d == _T_22[9:0]) begin
        image_2_45 <= io_pixelVal_in_2_2;
      end else if (10'h2d == _T_19[9:0]) begin
        image_2_45 <= io_pixelVal_in_2_1;
      end else if (10'h2d == _T_15[9:0]) begin
        image_2_45 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_46 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h2e == _T_37[9:0]) begin
        image_2_46 <= io_pixelVal_in_2_7;
      end else if (10'h2e == _T_34[9:0]) begin
        image_2_46 <= io_pixelVal_in_2_6;
      end else if (10'h2e == _T_31[9:0]) begin
        image_2_46 <= io_pixelVal_in_2_5;
      end else if (10'h2e == _T_28[9:0]) begin
        image_2_46 <= io_pixelVal_in_2_4;
      end else if (10'h2e == _T_25[9:0]) begin
        image_2_46 <= io_pixelVal_in_2_3;
      end else if (10'h2e == _T_22[9:0]) begin
        image_2_46 <= io_pixelVal_in_2_2;
      end else if (10'h2e == _T_19[9:0]) begin
        image_2_46 <= io_pixelVal_in_2_1;
      end else if (10'h2e == _T_15[9:0]) begin
        image_2_46 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_47 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h2f == _T_37[9:0]) begin
        image_2_47 <= io_pixelVal_in_2_7;
      end else if (10'h2f == _T_34[9:0]) begin
        image_2_47 <= io_pixelVal_in_2_6;
      end else if (10'h2f == _T_31[9:0]) begin
        image_2_47 <= io_pixelVal_in_2_5;
      end else if (10'h2f == _T_28[9:0]) begin
        image_2_47 <= io_pixelVal_in_2_4;
      end else if (10'h2f == _T_25[9:0]) begin
        image_2_47 <= io_pixelVal_in_2_3;
      end else if (10'h2f == _T_22[9:0]) begin
        image_2_47 <= io_pixelVal_in_2_2;
      end else if (10'h2f == _T_19[9:0]) begin
        image_2_47 <= io_pixelVal_in_2_1;
      end else if (10'h2f == _T_15[9:0]) begin
        image_2_47 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_48 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h30 == _T_37[9:0]) begin
        image_2_48 <= io_pixelVal_in_2_7;
      end else if (10'h30 == _T_34[9:0]) begin
        image_2_48 <= io_pixelVal_in_2_6;
      end else if (10'h30 == _T_31[9:0]) begin
        image_2_48 <= io_pixelVal_in_2_5;
      end else if (10'h30 == _T_28[9:0]) begin
        image_2_48 <= io_pixelVal_in_2_4;
      end else if (10'h30 == _T_25[9:0]) begin
        image_2_48 <= io_pixelVal_in_2_3;
      end else if (10'h30 == _T_22[9:0]) begin
        image_2_48 <= io_pixelVal_in_2_2;
      end else if (10'h30 == _T_19[9:0]) begin
        image_2_48 <= io_pixelVal_in_2_1;
      end else if (10'h30 == _T_15[9:0]) begin
        image_2_48 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_49 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h31 == _T_37[9:0]) begin
        image_2_49 <= io_pixelVal_in_2_7;
      end else if (10'h31 == _T_34[9:0]) begin
        image_2_49 <= io_pixelVal_in_2_6;
      end else if (10'h31 == _T_31[9:0]) begin
        image_2_49 <= io_pixelVal_in_2_5;
      end else if (10'h31 == _T_28[9:0]) begin
        image_2_49 <= io_pixelVal_in_2_4;
      end else if (10'h31 == _T_25[9:0]) begin
        image_2_49 <= io_pixelVal_in_2_3;
      end else if (10'h31 == _T_22[9:0]) begin
        image_2_49 <= io_pixelVal_in_2_2;
      end else if (10'h31 == _T_19[9:0]) begin
        image_2_49 <= io_pixelVal_in_2_1;
      end else if (10'h31 == _T_15[9:0]) begin
        image_2_49 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_50 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h32 == _T_37[9:0]) begin
        image_2_50 <= io_pixelVal_in_2_7;
      end else if (10'h32 == _T_34[9:0]) begin
        image_2_50 <= io_pixelVal_in_2_6;
      end else if (10'h32 == _T_31[9:0]) begin
        image_2_50 <= io_pixelVal_in_2_5;
      end else if (10'h32 == _T_28[9:0]) begin
        image_2_50 <= io_pixelVal_in_2_4;
      end else if (10'h32 == _T_25[9:0]) begin
        image_2_50 <= io_pixelVal_in_2_3;
      end else if (10'h32 == _T_22[9:0]) begin
        image_2_50 <= io_pixelVal_in_2_2;
      end else if (10'h32 == _T_19[9:0]) begin
        image_2_50 <= io_pixelVal_in_2_1;
      end else if (10'h32 == _T_15[9:0]) begin
        image_2_50 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_51 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h33 == _T_37[9:0]) begin
        image_2_51 <= io_pixelVal_in_2_7;
      end else if (10'h33 == _T_34[9:0]) begin
        image_2_51 <= io_pixelVal_in_2_6;
      end else if (10'h33 == _T_31[9:0]) begin
        image_2_51 <= io_pixelVal_in_2_5;
      end else if (10'h33 == _T_28[9:0]) begin
        image_2_51 <= io_pixelVal_in_2_4;
      end else if (10'h33 == _T_25[9:0]) begin
        image_2_51 <= io_pixelVal_in_2_3;
      end else if (10'h33 == _T_22[9:0]) begin
        image_2_51 <= io_pixelVal_in_2_2;
      end else if (10'h33 == _T_19[9:0]) begin
        image_2_51 <= io_pixelVal_in_2_1;
      end else if (10'h33 == _T_15[9:0]) begin
        image_2_51 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_52 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h34 == _T_37[9:0]) begin
        image_2_52 <= io_pixelVal_in_2_7;
      end else if (10'h34 == _T_34[9:0]) begin
        image_2_52 <= io_pixelVal_in_2_6;
      end else if (10'h34 == _T_31[9:0]) begin
        image_2_52 <= io_pixelVal_in_2_5;
      end else if (10'h34 == _T_28[9:0]) begin
        image_2_52 <= io_pixelVal_in_2_4;
      end else if (10'h34 == _T_25[9:0]) begin
        image_2_52 <= io_pixelVal_in_2_3;
      end else if (10'h34 == _T_22[9:0]) begin
        image_2_52 <= io_pixelVal_in_2_2;
      end else if (10'h34 == _T_19[9:0]) begin
        image_2_52 <= io_pixelVal_in_2_1;
      end else if (10'h34 == _T_15[9:0]) begin
        image_2_52 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_53 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h35 == _T_37[9:0]) begin
        image_2_53 <= io_pixelVal_in_2_7;
      end else if (10'h35 == _T_34[9:0]) begin
        image_2_53 <= io_pixelVal_in_2_6;
      end else if (10'h35 == _T_31[9:0]) begin
        image_2_53 <= io_pixelVal_in_2_5;
      end else if (10'h35 == _T_28[9:0]) begin
        image_2_53 <= io_pixelVal_in_2_4;
      end else if (10'h35 == _T_25[9:0]) begin
        image_2_53 <= io_pixelVal_in_2_3;
      end else if (10'h35 == _T_22[9:0]) begin
        image_2_53 <= io_pixelVal_in_2_2;
      end else if (10'h35 == _T_19[9:0]) begin
        image_2_53 <= io_pixelVal_in_2_1;
      end else if (10'h35 == _T_15[9:0]) begin
        image_2_53 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_54 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h36 == _T_37[9:0]) begin
        image_2_54 <= io_pixelVal_in_2_7;
      end else if (10'h36 == _T_34[9:0]) begin
        image_2_54 <= io_pixelVal_in_2_6;
      end else if (10'h36 == _T_31[9:0]) begin
        image_2_54 <= io_pixelVal_in_2_5;
      end else if (10'h36 == _T_28[9:0]) begin
        image_2_54 <= io_pixelVal_in_2_4;
      end else if (10'h36 == _T_25[9:0]) begin
        image_2_54 <= io_pixelVal_in_2_3;
      end else if (10'h36 == _T_22[9:0]) begin
        image_2_54 <= io_pixelVal_in_2_2;
      end else if (10'h36 == _T_19[9:0]) begin
        image_2_54 <= io_pixelVal_in_2_1;
      end else if (10'h36 == _T_15[9:0]) begin
        image_2_54 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_55 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h37 == _T_37[9:0]) begin
        image_2_55 <= io_pixelVal_in_2_7;
      end else if (10'h37 == _T_34[9:0]) begin
        image_2_55 <= io_pixelVal_in_2_6;
      end else if (10'h37 == _T_31[9:0]) begin
        image_2_55 <= io_pixelVal_in_2_5;
      end else if (10'h37 == _T_28[9:0]) begin
        image_2_55 <= io_pixelVal_in_2_4;
      end else if (10'h37 == _T_25[9:0]) begin
        image_2_55 <= io_pixelVal_in_2_3;
      end else if (10'h37 == _T_22[9:0]) begin
        image_2_55 <= io_pixelVal_in_2_2;
      end else if (10'h37 == _T_19[9:0]) begin
        image_2_55 <= io_pixelVal_in_2_1;
      end else if (10'h37 == _T_15[9:0]) begin
        image_2_55 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_56 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h38 == _T_37[9:0]) begin
        image_2_56 <= io_pixelVal_in_2_7;
      end else if (10'h38 == _T_34[9:0]) begin
        image_2_56 <= io_pixelVal_in_2_6;
      end else if (10'h38 == _T_31[9:0]) begin
        image_2_56 <= io_pixelVal_in_2_5;
      end else if (10'h38 == _T_28[9:0]) begin
        image_2_56 <= io_pixelVal_in_2_4;
      end else if (10'h38 == _T_25[9:0]) begin
        image_2_56 <= io_pixelVal_in_2_3;
      end else if (10'h38 == _T_22[9:0]) begin
        image_2_56 <= io_pixelVal_in_2_2;
      end else if (10'h38 == _T_19[9:0]) begin
        image_2_56 <= io_pixelVal_in_2_1;
      end else if (10'h38 == _T_15[9:0]) begin
        image_2_56 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_57 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h39 == _T_37[9:0]) begin
        image_2_57 <= io_pixelVal_in_2_7;
      end else if (10'h39 == _T_34[9:0]) begin
        image_2_57 <= io_pixelVal_in_2_6;
      end else if (10'h39 == _T_31[9:0]) begin
        image_2_57 <= io_pixelVal_in_2_5;
      end else if (10'h39 == _T_28[9:0]) begin
        image_2_57 <= io_pixelVal_in_2_4;
      end else if (10'h39 == _T_25[9:0]) begin
        image_2_57 <= io_pixelVal_in_2_3;
      end else if (10'h39 == _T_22[9:0]) begin
        image_2_57 <= io_pixelVal_in_2_2;
      end else if (10'h39 == _T_19[9:0]) begin
        image_2_57 <= io_pixelVal_in_2_1;
      end else if (10'h39 == _T_15[9:0]) begin
        image_2_57 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_58 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h3a == _T_37[9:0]) begin
        image_2_58 <= io_pixelVal_in_2_7;
      end else if (10'h3a == _T_34[9:0]) begin
        image_2_58 <= io_pixelVal_in_2_6;
      end else if (10'h3a == _T_31[9:0]) begin
        image_2_58 <= io_pixelVal_in_2_5;
      end else if (10'h3a == _T_28[9:0]) begin
        image_2_58 <= io_pixelVal_in_2_4;
      end else if (10'h3a == _T_25[9:0]) begin
        image_2_58 <= io_pixelVal_in_2_3;
      end else if (10'h3a == _T_22[9:0]) begin
        image_2_58 <= io_pixelVal_in_2_2;
      end else if (10'h3a == _T_19[9:0]) begin
        image_2_58 <= io_pixelVal_in_2_1;
      end else if (10'h3a == _T_15[9:0]) begin
        image_2_58 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_59 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h3b == _T_37[9:0]) begin
        image_2_59 <= io_pixelVal_in_2_7;
      end else if (10'h3b == _T_34[9:0]) begin
        image_2_59 <= io_pixelVal_in_2_6;
      end else if (10'h3b == _T_31[9:0]) begin
        image_2_59 <= io_pixelVal_in_2_5;
      end else if (10'h3b == _T_28[9:0]) begin
        image_2_59 <= io_pixelVal_in_2_4;
      end else if (10'h3b == _T_25[9:0]) begin
        image_2_59 <= io_pixelVal_in_2_3;
      end else if (10'h3b == _T_22[9:0]) begin
        image_2_59 <= io_pixelVal_in_2_2;
      end else if (10'h3b == _T_19[9:0]) begin
        image_2_59 <= io_pixelVal_in_2_1;
      end else if (10'h3b == _T_15[9:0]) begin
        image_2_59 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_60 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h3c == _T_37[9:0]) begin
        image_2_60 <= io_pixelVal_in_2_7;
      end else if (10'h3c == _T_34[9:0]) begin
        image_2_60 <= io_pixelVal_in_2_6;
      end else if (10'h3c == _T_31[9:0]) begin
        image_2_60 <= io_pixelVal_in_2_5;
      end else if (10'h3c == _T_28[9:0]) begin
        image_2_60 <= io_pixelVal_in_2_4;
      end else if (10'h3c == _T_25[9:0]) begin
        image_2_60 <= io_pixelVal_in_2_3;
      end else if (10'h3c == _T_22[9:0]) begin
        image_2_60 <= io_pixelVal_in_2_2;
      end else if (10'h3c == _T_19[9:0]) begin
        image_2_60 <= io_pixelVal_in_2_1;
      end else if (10'h3c == _T_15[9:0]) begin
        image_2_60 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_61 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h3d == _T_37[9:0]) begin
        image_2_61 <= io_pixelVal_in_2_7;
      end else if (10'h3d == _T_34[9:0]) begin
        image_2_61 <= io_pixelVal_in_2_6;
      end else if (10'h3d == _T_31[9:0]) begin
        image_2_61 <= io_pixelVal_in_2_5;
      end else if (10'h3d == _T_28[9:0]) begin
        image_2_61 <= io_pixelVal_in_2_4;
      end else if (10'h3d == _T_25[9:0]) begin
        image_2_61 <= io_pixelVal_in_2_3;
      end else if (10'h3d == _T_22[9:0]) begin
        image_2_61 <= io_pixelVal_in_2_2;
      end else if (10'h3d == _T_19[9:0]) begin
        image_2_61 <= io_pixelVal_in_2_1;
      end else if (10'h3d == _T_15[9:0]) begin
        image_2_61 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_62 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h3e == _T_37[9:0]) begin
        image_2_62 <= io_pixelVal_in_2_7;
      end else if (10'h3e == _T_34[9:0]) begin
        image_2_62 <= io_pixelVal_in_2_6;
      end else if (10'h3e == _T_31[9:0]) begin
        image_2_62 <= io_pixelVal_in_2_5;
      end else if (10'h3e == _T_28[9:0]) begin
        image_2_62 <= io_pixelVal_in_2_4;
      end else if (10'h3e == _T_25[9:0]) begin
        image_2_62 <= io_pixelVal_in_2_3;
      end else if (10'h3e == _T_22[9:0]) begin
        image_2_62 <= io_pixelVal_in_2_2;
      end else if (10'h3e == _T_19[9:0]) begin
        image_2_62 <= io_pixelVal_in_2_1;
      end else if (10'h3e == _T_15[9:0]) begin
        image_2_62 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_63 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h3f == _T_37[9:0]) begin
        image_2_63 <= io_pixelVal_in_2_7;
      end else if (10'h3f == _T_34[9:0]) begin
        image_2_63 <= io_pixelVal_in_2_6;
      end else if (10'h3f == _T_31[9:0]) begin
        image_2_63 <= io_pixelVal_in_2_5;
      end else if (10'h3f == _T_28[9:0]) begin
        image_2_63 <= io_pixelVal_in_2_4;
      end else if (10'h3f == _T_25[9:0]) begin
        image_2_63 <= io_pixelVal_in_2_3;
      end else if (10'h3f == _T_22[9:0]) begin
        image_2_63 <= io_pixelVal_in_2_2;
      end else if (10'h3f == _T_19[9:0]) begin
        image_2_63 <= io_pixelVal_in_2_1;
      end else if (10'h3f == _T_15[9:0]) begin
        image_2_63 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_64 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h40 == _T_37[9:0]) begin
        image_2_64 <= io_pixelVal_in_2_7;
      end else if (10'h40 == _T_34[9:0]) begin
        image_2_64 <= io_pixelVal_in_2_6;
      end else if (10'h40 == _T_31[9:0]) begin
        image_2_64 <= io_pixelVal_in_2_5;
      end else if (10'h40 == _T_28[9:0]) begin
        image_2_64 <= io_pixelVal_in_2_4;
      end else if (10'h40 == _T_25[9:0]) begin
        image_2_64 <= io_pixelVal_in_2_3;
      end else if (10'h40 == _T_22[9:0]) begin
        image_2_64 <= io_pixelVal_in_2_2;
      end else if (10'h40 == _T_19[9:0]) begin
        image_2_64 <= io_pixelVal_in_2_1;
      end else if (10'h40 == _T_15[9:0]) begin
        image_2_64 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_65 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h41 == _T_37[9:0]) begin
        image_2_65 <= io_pixelVal_in_2_7;
      end else if (10'h41 == _T_34[9:0]) begin
        image_2_65 <= io_pixelVal_in_2_6;
      end else if (10'h41 == _T_31[9:0]) begin
        image_2_65 <= io_pixelVal_in_2_5;
      end else if (10'h41 == _T_28[9:0]) begin
        image_2_65 <= io_pixelVal_in_2_4;
      end else if (10'h41 == _T_25[9:0]) begin
        image_2_65 <= io_pixelVal_in_2_3;
      end else if (10'h41 == _T_22[9:0]) begin
        image_2_65 <= io_pixelVal_in_2_2;
      end else if (10'h41 == _T_19[9:0]) begin
        image_2_65 <= io_pixelVal_in_2_1;
      end else if (10'h41 == _T_15[9:0]) begin
        image_2_65 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_66 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h42 == _T_37[9:0]) begin
        image_2_66 <= io_pixelVal_in_2_7;
      end else if (10'h42 == _T_34[9:0]) begin
        image_2_66 <= io_pixelVal_in_2_6;
      end else if (10'h42 == _T_31[9:0]) begin
        image_2_66 <= io_pixelVal_in_2_5;
      end else if (10'h42 == _T_28[9:0]) begin
        image_2_66 <= io_pixelVal_in_2_4;
      end else if (10'h42 == _T_25[9:0]) begin
        image_2_66 <= io_pixelVal_in_2_3;
      end else if (10'h42 == _T_22[9:0]) begin
        image_2_66 <= io_pixelVal_in_2_2;
      end else if (10'h42 == _T_19[9:0]) begin
        image_2_66 <= io_pixelVal_in_2_1;
      end else if (10'h42 == _T_15[9:0]) begin
        image_2_66 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_67 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h43 == _T_37[9:0]) begin
        image_2_67 <= io_pixelVal_in_2_7;
      end else if (10'h43 == _T_34[9:0]) begin
        image_2_67 <= io_pixelVal_in_2_6;
      end else if (10'h43 == _T_31[9:0]) begin
        image_2_67 <= io_pixelVal_in_2_5;
      end else if (10'h43 == _T_28[9:0]) begin
        image_2_67 <= io_pixelVal_in_2_4;
      end else if (10'h43 == _T_25[9:0]) begin
        image_2_67 <= io_pixelVal_in_2_3;
      end else if (10'h43 == _T_22[9:0]) begin
        image_2_67 <= io_pixelVal_in_2_2;
      end else if (10'h43 == _T_19[9:0]) begin
        image_2_67 <= io_pixelVal_in_2_1;
      end else if (10'h43 == _T_15[9:0]) begin
        image_2_67 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_68 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h44 == _T_37[9:0]) begin
        image_2_68 <= io_pixelVal_in_2_7;
      end else if (10'h44 == _T_34[9:0]) begin
        image_2_68 <= io_pixelVal_in_2_6;
      end else if (10'h44 == _T_31[9:0]) begin
        image_2_68 <= io_pixelVal_in_2_5;
      end else if (10'h44 == _T_28[9:0]) begin
        image_2_68 <= io_pixelVal_in_2_4;
      end else if (10'h44 == _T_25[9:0]) begin
        image_2_68 <= io_pixelVal_in_2_3;
      end else if (10'h44 == _T_22[9:0]) begin
        image_2_68 <= io_pixelVal_in_2_2;
      end else if (10'h44 == _T_19[9:0]) begin
        image_2_68 <= io_pixelVal_in_2_1;
      end else if (10'h44 == _T_15[9:0]) begin
        image_2_68 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_69 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h45 == _T_37[9:0]) begin
        image_2_69 <= io_pixelVal_in_2_7;
      end else if (10'h45 == _T_34[9:0]) begin
        image_2_69 <= io_pixelVal_in_2_6;
      end else if (10'h45 == _T_31[9:0]) begin
        image_2_69 <= io_pixelVal_in_2_5;
      end else if (10'h45 == _T_28[9:0]) begin
        image_2_69 <= io_pixelVal_in_2_4;
      end else if (10'h45 == _T_25[9:0]) begin
        image_2_69 <= io_pixelVal_in_2_3;
      end else if (10'h45 == _T_22[9:0]) begin
        image_2_69 <= io_pixelVal_in_2_2;
      end else if (10'h45 == _T_19[9:0]) begin
        image_2_69 <= io_pixelVal_in_2_1;
      end else if (10'h45 == _T_15[9:0]) begin
        image_2_69 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_70 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h46 == _T_37[9:0]) begin
        image_2_70 <= io_pixelVal_in_2_7;
      end else if (10'h46 == _T_34[9:0]) begin
        image_2_70 <= io_pixelVal_in_2_6;
      end else if (10'h46 == _T_31[9:0]) begin
        image_2_70 <= io_pixelVal_in_2_5;
      end else if (10'h46 == _T_28[9:0]) begin
        image_2_70 <= io_pixelVal_in_2_4;
      end else if (10'h46 == _T_25[9:0]) begin
        image_2_70 <= io_pixelVal_in_2_3;
      end else if (10'h46 == _T_22[9:0]) begin
        image_2_70 <= io_pixelVal_in_2_2;
      end else if (10'h46 == _T_19[9:0]) begin
        image_2_70 <= io_pixelVal_in_2_1;
      end else if (10'h46 == _T_15[9:0]) begin
        image_2_70 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_71 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h47 == _T_37[9:0]) begin
        image_2_71 <= io_pixelVal_in_2_7;
      end else if (10'h47 == _T_34[9:0]) begin
        image_2_71 <= io_pixelVal_in_2_6;
      end else if (10'h47 == _T_31[9:0]) begin
        image_2_71 <= io_pixelVal_in_2_5;
      end else if (10'h47 == _T_28[9:0]) begin
        image_2_71 <= io_pixelVal_in_2_4;
      end else if (10'h47 == _T_25[9:0]) begin
        image_2_71 <= io_pixelVal_in_2_3;
      end else if (10'h47 == _T_22[9:0]) begin
        image_2_71 <= io_pixelVal_in_2_2;
      end else if (10'h47 == _T_19[9:0]) begin
        image_2_71 <= io_pixelVal_in_2_1;
      end else if (10'h47 == _T_15[9:0]) begin
        image_2_71 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_72 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h48 == _T_37[9:0]) begin
        image_2_72 <= io_pixelVal_in_2_7;
      end else if (10'h48 == _T_34[9:0]) begin
        image_2_72 <= io_pixelVal_in_2_6;
      end else if (10'h48 == _T_31[9:0]) begin
        image_2_72 <= io_pixelVal_in_2_5;
      end else if (10'h48 == _T_28[9:0]) begin
        image_2_72 <= io_pixelVal_in_2_4;
      end else if (10'h48 == _T_25[9:0]) begin
        image_2_72 <= io_pixelVal_in_2_3;
      end else if (10'h48 == _T_22[9:0]) begin
        image_2_72 <= io_pixelVal_in_2_2;
      end else if (10'h48 == _T_19[9:0]) begin
        image_2_72 <= io_pixelVal_in_2_1;
      end else if (10'h48 == _T_15[9:0]) begin
        image_2_72 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_73 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h49 == _T_37[9:0]) begin
        image_2_73 <= io_pixelVal_in_2_7;
      end else if (10'h49 == _T_34[9:0]) begin
        image_2_73 <= io_pixelVal_in_2_6;
      end else if (10'h49 == _T_31[9:0]) begin
        image_2_73 <= io_pixelVal_in_2_5;
      end else if (10'h49 == _T_28[9:0]) begin
        image_2_73 <= io_pixelVal_in_2_4;
      end else if (10'h49 == _T_25[9:0]) begin
        image_2_73 <= io_pixelVal_in_2_3;
      end else if (10'h49 == _T_22[9:0]) begin
        image_2_73 <= io_pixelVal_in_2_2;
      end else if (10'h49 == _T_19[9:0]) begin
        image_2_73 <= io_pixelVal_in_2_1;
      end else if (10'h49 == _T_15[9:0]) begin
        image_2_73 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_74 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h4a == _T_37[9:0]) begin
        image_2_74 <= io_pixelVal_in_2_7;
      end else if (10'h4a == _T_34[9:0]) begin
        image_2_74 <= io_pixelVal_in_2_6;
      end else if (10'h4a == _T_31[9:0]) begin
        image_2_74 <= io_pixelVal_in_2_5;
      end else if (10'h4a == _T_28[9:0]) begin
        image_2_74 <= io_pixelVal_in_2_4;
      end else if (10'h4a == _T_25[9:0]) begin
        image_2_74 <= io_pixelVal_in_2_3;
      end else if (10'h4a == _T_22[9:0]) begin
        image_2_74 <= io_pixelVal_in_2_2;
      end else if (10'h4a == _T_19[9:0]) begin
        image_2_74 <= io_pixelVal_in_2_1;
      end else if (10'h4a == _T_15[9:0]) begin
        image_2_74 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_75 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h4b == _T_37[9:0]) begin
        image_2_75 <= io_pixelVal_in_2_7;
      end else if (10'h4b == _T_34[9:0]) begin
        image_2_75 <= io_pixelVal_in_2_6;
      end else if (10'h4b == _T_31[9:0]) begin
        image_2_75 <= io_pixelVal_in_2_5;
      end else if (10'h4b == _T_28[9:0]) begin
        image_2_75 <= io_pixelVal_in_2_4;
      end else if (10'h4b == _T_25[9:0]) begin
        image_2_75 <= io_pixelVal_in_2_3;
      end else if (10'h4b == _T_22[9:0]) begin
        image_2_75 <= io_pixelVal_in_2_2;
      end else if (10'h4b == _T_19[9:0]) begin
        image_2_75 <= io_pixelVal_in_2_1;
      end else if (10'h4b == _T_15[9:0]) begin
        image_2_75 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_76 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h4c == _T_37[9:0]) begin
        image_2_76 <= io_pixelVal_in_2_7;
      end else if (10'h4c == _T_34[9:0]) begin
        image_2_76 <= io_pixelVal_in_2_6;
      end else if (10'h4c == _T_31[9:0]) begin
        image_2_76 <= io_pixelVal_in_2_5;
      end else if (10'h4c == _T_28[9:0]) begin
        image_2_76 <= io_pixelVal_in_2_4;
      end else if (10'h4c == _T_25[9:0]) begin
        image_2_76 <= io_pixelVal_in_2_3;
      end else if (10'h4c == _T_22[9:0]) begin
        image_2_76 <= io_pixelVal_in_2_2;
      end else if (10'h4c == _T_19[9:0]) begin
        image_2_76 <= io_pixelVal_in_2_1;
      end else if (10'h4c == _T_15[9:0]) begin
        image_2_76 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_77 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h4d == _T_37[9:0]) begin
        image_2_77 <= io_pixelVal_in_2_7;
      end else if (10'h4d == _T_34[9:0]) begin
        image_2_77 <= io_pixelVal_in_2_6;
      end else if (10'h4d == _T_31[9:0]) begin
        image_2_77 <= io_pixelVal_in_2_5;
      end else if (10'h4d == _T_28[9:0]) begin
        image_2_77 <= io_pixelVal_in_2_4;
      end else if (10'h4d == _T_25[9:0]) begin
        image_2_77 <= io_pixelVal_in_2_3;
      end else if (10'h4d == _T_22[9:0]) begin
        image_2_77 <= io_pixelVal_in_2_2;
      end else if (10'h4d == _T_19[9:0]) begin
        image_2_77 <= io_pixelVal_in_2_1;
      end else if (10'h4d == _T_15[9:0]) begin
        image_2_77 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_78 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h4e == _T_37[9:0]) begin
        image_2_78 <= io_pixelVal_in_2_7;
      end else if (10'h4e == _T_34[9:0]) begin
        image_2_78 <= io_pixelVal_in_2_6;
      end else if (10'h4e == _T_31[9:0]) begin
        image_2_78 <= io_pixelVal_in_2_5;
      end else if (10'h4e == _T_28[9:0]) begin
        image_2_78 <= io_pixelVal_in_2_4;
      end else if (10'h4e == _T_25[9:0]) begin
        image_2_78 <= io_pixelVal_in_2_3;
      end else if (10'h4e == _T_22[9:0]) begin
        image_2_78 <= io_pixelVal_in_2_2;
      end else if (10'h4e == _T_19[9:0]) begin
        image_2_78 <= io_pixelVal_in_2_1;
      end else if (10'h4e == _T_15[9:0]) begin
        image_2_78 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_79 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h4f == _T_37[9:0]) begin
        image_2_79 <= io_pixelVal_in_2_7;
      end else if (10'h4f == _T_34[9:0]) begin
        image_2_79 <= io_pixelVal_in_2_6;
      end else if (10'h4f == _T_31[9:0]) begin
        image_2_79 <= io_pixelVal_in_2_5;
      end else if (10'h4f == _T_28[9:0]) begin
        image_2_79 <= io_pixelVal_in_2_4;
      end else if (10'h4f == _T_25[9:0]) begin
        image_2_79 <= io_pixelVal_in_2_3;
      end else if (10'h4f == _T_22[9:0]) begin
        image_2_79 <= io_pixelVal_in_2_2;
      end else if (10'h4f == _T_19[9:0]) begin
        image_2_79 <= io_pixelVal_in_2_1;
      end else if (10'h4f == _T_15[9:0]) begin
        image_2_79 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_80 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h50 == _T_37[9:0]) begin
        image_2_80 <= io_pixelVal_in_2_7;
      end else if (10'h50 == _T_34[9:0]) begin
        image_2_80 <= io_pixelVal_in_2_6;
      end else if (10'h50 == _T_31[9:0]) begin
        image_2_80 <= io_pixelVal_in_2_5;
      end else if (10'h50 == _T_28[9:0]) begin
        image_2_80 <= io_pixelVal_in_2_4;
      end else if (10'h50 == _T_25[9:0]) begin
        image_2_80 <= io_pixelVal_in_2_3;
      end else if (10'h50 == _T_22[9:0]) begin
        image_2_80 <= io_pixelVal_in_2_2;
      end else if (10'h50 == _T_19[9:0]) begin
        image_2_80 <= io_pixelVal_in_2_1;
      end else if (10'h50 == _T_15[9:0]) begin
        image_2_80 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_81 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h51 == _T_37[9:0]) begin
        image_2_81 <= io_pixelVal_in_2_7;
      end else if (10'h51 == _T_34[9:0]) begin
        image_2_81 <= io_pixelVal_in_2_6;
      end else if (10'h51 == _T_31[9:0]) begin
        image_2_81 <= io_pixelVal_in_2_5;
      end else if (10'h51 == _T_28[9:0]) begin
        image_2_81 <= io_pixelVal_in_2_4;
      end else if (10'h51 == _T_25[9:0]) begin
        image_2_81 <= io_pixelVal_in_2_3;
      end else if (10'h51 == _T_22[9:0]) begin
        image_2_81 <= io_pixelVal_in_2_2;
      end else if (10'h51 == _T_19[9:0]) begin
        image_2_81 <= io_pixelVal_in_2_1;
      end else if (10'h51 == _T_15[9:0]) begin
        image_2_81 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_82 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h52 == _T_37[9:0]) begin
        image_2_82 <= io_pixelVal_in_2_7;
      end else if (10'h52 == _T_34[9:0]) begin
        image_2_82 <= io_pixelVal_in_2_6;
      end else if (10'h52 == _T_31[9:0]) begin
        image_2_82 <= io_pixelVal_in_2_5;
      end else if (10'h52 == _T_28[9:0]) begin
        image_2_82 <= io_pixelVal_in_2_4;
      end else if (10'h52 == _T_25[9:0]) begin
        image_2_82 <= io_pixelVal_in_2_3;
      end else if (10'h52 == _T_22[9:0]) begin
        image_2_82 <= io_pixelVal_in_2_2;
      end else if (10'h52 == _T_19[9:0]) begin
        image_2_82 <= io_pixelVal_in_2_1;
      end else if (10'h52 == _T_15[9:0]) begin
        image_2_82 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_83 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h53 == _T_37[9:0]) begin
        image_2_83 <= io_pixelVal_in_2_7;
      end else if (10'h53 == _T_34[9:0]) begin
        image_2_83 <= io_pixelVal_in_2_6;
      end else if (10'h53 == _T_31[9:0]) begin
        image_2_83 <= io_pixelVal_in_2_5;
      end else if (10'h53 == _T_28[9:0]) begin
        image_2_83 <= io_pixelVal_in_2_4;
      end else if (10'h53 == _T_25[9:0]) begin
        image_2_83 <= io_pixelVal_in_2_3;
      end else if (10'h53 == _T_22[9:0]) begin
        image_2_83 <= io_pixelVal_in_2_2;
      end else if (10'h53 == _T_19[9:0]) begin
        image_2_83 <= io_pixelVal_in_2_1;
      end else if (10'h53 == _T_15[9:0]) begin
        image_2_83 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_84 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h54 == _T_37[9:0]) begin
        image_2_84 <= io_pixelVal_in_2_7;
      end else if (10'h54 == _T_34[9:0]) begin
        image_2_84 <= io_pixelVal_in_2_6;
      end else if (10'h54 == _T_31[9:0]) begin
        image_2_84 <= io_pixelVal_in_2_5;
      end else if (10'h54 == _T_28[9:0]) begin
        image_2_84 <= io_pixelVal_in_2_4;
      end else if (10'h54 == _T_25[9:0]) begin
        image_2_84 <= io_pixelVal_in_2_3;
      end else if (10'h54 == _T_22[9:0]) begin
        image_2_84 <= io_pixelVal_in_2_2;
      end else if (10'h54 == _T_19[9:0]) begin
        image_2_84 <= io_pixelVal_in_2_1;
      end else if (10'h54 == _T_15[9:0]) begin
        image_2_84 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_85 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h55 == _T_37[9:0]) begin
        image_2_85 <= io_pixelVal_in_2_7;
      end else if (10'h55 == _T_34[9:0]) begin
        image_2_85 <= io_pixelVal_in_2_6;
      end else if (10'h55 == _T_31[9:0]) begin
        image_2_85 <= io_pixelVal_in_2_5;
      end else if (10'h55 == _T_28[9:0]) begin
        image_2_85 <= io_pixelVal_in_2_4;
      end else if (10'h55 == _T_25[9:0]) begin
        image_2_85 <= io_pixelVal_in_2_3;
      end else if (10'h55 == _T_22[9:0]) begin
        image_2_85 <= io_pixelVal_in_2_2;
      end else if (10'h55 == _T_19[9:0]) begin
        image_2_85 <= io_pixelVal_in_2_1;
      end else if (10'h55 == _T_15[9:0]) begin
        image_2_85 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_86 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h56 == _T_37[9:0]) begin
        image_2_86 <= io_pixelVal_in_2_7;
      end else if (10'h56 == _T_34[9:0]) begin
        image_2_86 <= io_pixelVal_in_2_6;
      end else if (10'h56 == _T_31[9:0]) begin
        image_2_86 <= io_pixelVal_in_2_5;
      end else if (10'h56 == _T_28[9:0]) begin
        image_2_86 <= io_pixelVal_in_2_4;
      end else if (10'h56 == _T_25[9:0]) begin
        image_2_86 <= io_pixelVal_in_2_3;
      end else if (10'h56 == _T_22[9:0]) begin
        image_2_86 <= io_pixelVal_in_2_2;
      end else if (10'h56 == _T_19[9:0]) begin
        image_2_86 <= io_pixelVal_in_2_1;
      end else if (10'h56 == _T_15[9:0]) begin
        image_2_86 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_87 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h57 == _T_37[9:0]) begin
        image_2_87 <= io_pixelVal_in_2_7;
      end else if (10'h57 == _T_34[9:0]) begin
        image_2_87 <= io_pixelVal_in_2_6;
      end else if (10'h57 == _T_31[9:0]) begin
        image_2_87 <= io_pixelVal_in_2_5;
      end else if (10'h57 == _T_28[9:0]) begin
        image_2_87 <= io_pixelVal_in_2_4;
      end else if (10'h57 == _T_25[9:0]) begin
        image_2_87 <= io_pixelVal_in_2_3;
      end else if (10'h57 == _T_22[9:0]) begin
        image_2_87 <= io_pixelVal_in_2_2;
      end else if (10'h57 == _T_19[9:0]) begin
        image_2_87 <= io_pixelVal_in_2_1;
      end else if (10'h57 == _T_15[9:0]) begin
        image_2_87 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_88 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h58 == _T_37[9:0]) begin
        image_2_88 <= io_pixelVal_in_2_7;
      end else if (10'h58 == _T_34[9:0]) begin
        image_2_88 <= io_pixelVal_in_2_6;
      end else if (10'h58 == _T_31[9:0]) begin
        image_2_88 <= io_pixelVal_in_2_5;
      end else if (10'h58 == _T_28[9:0]) begin
        image_2_88 <= io_pixelVal_in_2_4;
      end else if (10'h58 == _T_25[9:0]) begin
        image_2_88 <= io_pixelVal_in_2_3;
      end else if (10'h58 == _T_22[9:0]) begin
        image_2_88 <= io_pixelVal_in_2_2;
      end else if (10'h58 == _T_19[9:0]) begin
        image_2_88 <= io_pixelVal_in_2_1;
      end else if (10'h58 == _T_15[9:0]) begin
        image_2_88 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_89 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h59 == _T_37[9:0]) begin
        image_2_89 <= io_pixelVal_in_2_7;
      end else if (10'h59 == _T_34[9:0]) begin
        image_2_89 <= io_pixelVal_in_2_6;
      end else if (10'h59 == _T_31[9:0]) begin
        image_2_89 <= io_pixelVal_in_2_5;
      end else if (10'h59 == _T_28[9:0]) begin
        image_2_89 <= io_pixelVal_in_2_4;
      end else if (10'h59 == _T_25[9:0]) begin
        image_2_89 <= io_pixelVal_in_2_3;
      end else if (10'h59 == _T_22[9:0]) begin
        image_2_89 <= io_pixelVal_in_2_2;
      end else if (10'h59 == _T_19[9:0]) begin
        image_2_89 <= io_pixelVal_in_2_1;
      end else if (10'h59 == _T_15[9:0]) begin
        image_2_89 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_90 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h5a == _T_37[9:0]) begin
        image_2_90 <= io_pixelVal_in_2_7;
      end else if (10'h5a == _T_34[9:0]) begin
        image_2_90 <= io_pixelVal_in_2_6;
      end else if (10'h5a == _T_31[9:0]) begin
        image_2_90 <= io_pixelVal_in_2_5;
      end else if (10'h5a == _T_28[9:0]) begin
        image_2_90 <= io_pixelVal_in_2_4;
      end else if (10'h5a == _T_25[9:0]) begin
        image_2_90 <= io_pixelVal_in_2_3;
      end else if (10'h5a == _T_22[9:0]) begin
        image_2_90 <= io_pixelVal_in_2_2;
      end else if (10'h5a == _T_19[9:0]) begin
        image_2_90 <= io_pixelVal_in_2_1;
      end else if (10'h5a == _T_15[9:0]) begin
        image_2_90 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_91 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h5b == _T_37[9:0]) begin
        image_2_91 <= io_pixelVal_in_2_7;
      end else if (10'h5b == _T_34[9:0]) begin
        image_2_91 <= io_pixelVal_in_2_6;
      end else if (10'h5b == _T_31[9:0]) begin
        image_2_91 <= io_pixelVal_in_2_5;
      end else if (10'h5b == _T_28[9:0]) begin
        image_2_91 <= io_pixelVal_in_2_4;
      end else if (10'h5b == _T_25[9:0]) begin
        image_2_91 <= io_pixelVal_in_2_3;
      end else if (10'h5b == _T_22[9:0]) begin
        image_2_91 <= io_pixelVal_in_2_2;
      end else if (10'h5b == _T_19[9:0]) begin
        image_2_91 <= io_pixelVal_in_2_1;
      end else if (10'h5b == _T_15[9:0]) begin
        image_2_91 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_92 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h5c == _T_37[9:0]) begin
        image_2_92 <= io_pixelVal_in_2_7;
      end else if (10'h5c == _T_34[9:0]) begin
        image_2_92 <= io_pixelVal_in_2_6;
      end else if (10'h5c == _T_31[9:0]) begin
        image_2_92 <= io_pixelVal_in_2_5;
      end else if (10'h5c == _T_28[9:0]) begin
        image_2_92 <= io_pixelVal_in_2_4;
      end else if (10'h5c == _T_25[9:0]) begin
        image_2_92 <= io_pixelVal_in_2_3;
      end else if (10'h5c == _T_22[9:0]) begin
        image_2_92 <= io_pixelVal_in_2_2;
      end else if (10'h5c == _T_19[9:0]) begin
        image_2_92 <= io_pixelVal_in_2_1;
      end else if (10'h5c == _T_15[9:0]) begin
        image_2_92 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_93 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h5d == _T_37[9:0]) begin
        image_2_93 <= io_pixelVal_in_2_7;
      end else if (10'h5d == _T_34[9:0]) begin
        image_2_93 <= io_pixelVal_in_2_6;
      end else if (10'h5d == _T_31[9:0]) begin
        image_2_93 <= io_pixelVal_in_2_5;
      end else if (10'h5d == _T_28[9:0]) begin
        image_2_93 <= io_pixelVal_in_2_4;
      end else if (10'h5d == _T_25[9:0]) begin
        image_2_93 <= io_pixelVal_in_2_3;
      end else if (10'h5d == _T_22[9:0]) begin
        image_2_93 <= io_pixelVal_in_2_2;
      end else if (10'h5d == _T_19[9:0]) begin
        image_2_93 <= io_pixelVal_in_2_1;
      end else if (10'h5d == _T_15[9:0]) begin
        image_2_93 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_94 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h5e == _T_37[9:0]) begin
        image_2_94 <= io_pixelVal_in_2_7;
      end else if (10'h5e == _T_34[9:0]) begin
        image_2_94 <= io_pixelVal_in_2_6;
      end else if (10'h5e == _T_31[9:0]) begin
        image_2_94 <= io_pixelVal_in_2_5;
      end else if (10'h5e == _T_28[9:0]) begin
        image_2_94 <= io_pixelVal_in_2_4;
      end else if (10'h5e == _T_25[9:0]) begin
        image_2_94 <= io_pixelVal_in_2_3;
      end else if (10'h5e == _T_22[9:0]) begin
        image_2_94 <= io_pixelVal_in_2_2;
      end else if (10'h5e == _T_19[9:0]) begin
        image_2_94 <= io_pixelVal_in_2_1;
      end else if (10'h5e == _T_15[9:0]) begin
        image_2_94 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_95 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h5f == _T_37[9:0]) begin
        image_2_95 <= io_pixelVal_in_2_7;
      end else if (10'h5f == _T_34[9:0]) begin
        image_2_95 <= io_pixelVal_in_2_6;
      end else if (10'h5f == _T_31[9:0]) begin
        image_2_95 <= io_pixelVal_in_2_5;
      end else if (10'h5f == _T_28[9:0]) begin
        image_2_95 <= io_pixelVal_in_2_4;
      end else if (10'h5f == _T_25[9:0]) begin
        image_2_95 <= io_pixelVal_in_2_3;
      end else if (10'h5f == _T_22[9:0]) begin
        image_2_95 <= io_pixelVal_in_2_2;
      end else if (10'h5f == _T_19[9:0]) begin
        image_2_95 <= io_pixelVal_in_2_1;
      end else if (10'h5f == _T_15[9:0]) begin
        image_2_95 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_96 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h60 == _T_37[9:0]) begin
        image_2_96 <= io_pixelVal_in_2_7;
      end else if (10'h60 == _T_34[9:0]) begin
        image_2_96 <= io_pixelVal_in_2_6;
      end else if (10'h60 == _T_31[9:0]) begin
        image_2_96 <= io_pixelVal_in_2_5;
      end else if (10'h60 == _T_28[9:0]) begin
        image_2_96 <= io_pixelVal_in_2_4;
      end else if (10'h60 == _T_25[9:0]) begin
        image_2_96 <= io_pixelVal_in_2_3;
      end else if (10'h60 == _T_22[9:0]) begin
        image_2_96 <= io_pixelVal_in_2_2;
      end else if (10'h60 == _T_19[9:0]) begin
        image_2_96 <= io_pixelVal_in_2_1;
      end else if (10'h60 == _T_15[9:0]) begin
        image_2_96 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_97 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h61 == _T_37[9:0]) begin
        image_2_97 <= io_pixelVal_in_2_7;
      end else if (10'h61 == _T_34[9:0]) begin
        image_2_97 <= io_pixelVal_in_2_6;
      end else if (10'h61 == _T_31[9:0]) begin
        image_2_97 <= io_pixelVal_in_2_5;
      end else if (10'h61 == _T_28[9:0]) begin
        image_2_97 <= io_pixelVal_in_2_4;
      end else if (10'h61 == _T_25[9:0]) begin
        image_2_97 <= io_pixelVal_in_2_3;
      end else if (10'h61 == _T_22[9:0]) begin
        image_2_97 <= io_pixelVal_in_2_2;
      end else if (10'h61 == _T_19[9:0]) begin
        image_2_97 <= io_pixelVal_in_2_1;
      end else if (10'h61 == _T_15[9:0]) begin
        image_2_97 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_98 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h62 == _T_37[9:0]) begin
        image_2_98 <= io_pixelVal_in_2_7;
      end else if (10'h62 == _T_34[9:0]) begin
        image_2_98 <= io_pixelVal_in_2_6;
      end else if (10'h62 == _T_31[9:0]) begin
        image_2_98 <= io_pixelVal_in_2_5;
      end else if (10'h62 == _T_28[9:0]) begin
        image_2_98 <= io_pixelVal_in_2_4;
      end else if (10'h62 == _T_25[9:0]) begin
        image_2_98 <= io_pixelVal_in_2_3;
      end else if (10'h62 == _T_22[9:0]) begin
        image_2_98 <= io_pixelVal_in_2_2;
      end else if (10'h62 == _T_19[9:0]) begin
        image_2_98 <= io_pixelVal_in_2_1;
      end else if (10'h62 == _T_15[9:0]) begin
        image_2_98 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_99 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h63 == _T_37[9:0]) begin
        image_2_99 <= io_pixelVal_in_2_7;
      end else if (10'h63 == _T_34[9:0]) begin
        image_2_99 <= io_pixelVal_in_2_6;
      end else if (10'h63 == _T_31[9:0]) begin
        image_2_99 <= io_pixelVal_in_2_5;
      end else if (10'h63 == _T_28[9:0]) begin
        image_2_99 <= io_pixelVal_in_2_4;
      end else if (10'h63 == _T_25[9:0]) begin
        image_2_99 <= io_pixelVal_in_2_3;
      end else if (10'h63 == _T_22[9:0]) begin
        image_2_99 <= io_pixelVal_in_2_2;
      end else if (10'h63 == _T_19[9:0]) begin
        image_2_99 <= io_pixelVal_in_2_1;
      end else if (10'h63 == _T_15[9:0]) begin
        image_2_99 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_100 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h64 == _T_37[9:0]) begin
        image_2_100 <= io_pixelVal_in_2_7;
      end else if (10'h64 == _T_34[9:0]) begin
        image_2_100 <= io_pixelVal_in_2_6;
      end else if (10'h64 == _T_31[9:0]) begin
        image_2_100 <= io_pixelVal_in_2_5;
      end else if (10'h64 == _T_28[9:0]) begin
        image_2_100 <= io_pixelVal_in_2_4;
      end else if (10'h64 == _T_25[9:0]) begin
        image_2_100 <= io_pixelVal_in_2_3;
      end else if (10'h64 == _T_22[9:0]) begin
        image_2_100 <= io_pixelVal_in_2_2;
      end else if (10'h64 == _T_19[9:0]) begin
        image_2_100 <= io_pixelVal_in_2_1;
      end else if (10'h64 == _T_15[9:0]) begin
        image_2_100 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_101 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h65 == _T_37[9:0]) begin
        image_2_101 <= io_pixelVal_in_2_7;
      end else if (10'h65 == _T_34[9:0]) begin
        image_2_101 <= io_pixelVal_in_2_6;
      end else if (10'h65 == _T_31[9:0]) begin
        image_2_101 <= io_pixelVal_in_2_5;
      end else if (10'h65 == _T_28[9:0]) begin
        image_2_101 <= io_pixelVal_in_2_4;
      end else if (10'h65 == _T_25[9:0]) begin
        image_2_101 <= io_pixelVal_in_2_3;
      end else if (10'h65 == _T_22[9:0]) begin
        image_2_101 <= io_pixelVal_in_2_2;
      end else if (10'h65 == _T_19[9:0]) begin
        image_2_101 <= io_pixelVal_in_2_1;
      end else if (10'h65 == _T_15[9:0]) begin
        image_2_101 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_102 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h66 == _T_37[9:0]) begin
        image_2_102 <= io_pixelVal_in_2_7;
      end else if (10'h66 == _T_34[9:0]) begin
        image_2_102 <= io_pixelVal_in_2_6;
      end else if (10'h66 == _T_31[9:0]) begin
        image_2_102 <= io_pixelVal_in_2_5;
      end else if (10'h66 == _T_28[9:0]) begin
        image_2_102 <= io_pixelVal_in_2_4;
      end else if (10'h66 == _T_25[9:0]) begin
        image_2_102 <= io_pixelVal_in_2_3;
      end else if (10'h66 == _T_22[9:0]) begin
        image_2_102 <= io_pixelVal_in_2_2;
      end else if (10'h66 == _T_19[9:0]) begin
        image_2_102 <= io_pixelVal_in_2_1;
      end else if (10'h66 == _T_15[9:0]) begin
        image_2_102 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_103 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h67 == _T_37[9:0]) begin
        image_2_103 <= io_pixelVal_in_2_7;
      end else if (10'h67 == _T_34[9:0]) begin
        image_2_103 <= io_pixelVal_in_2_6;
      end else if (10'h67 == _T_31[9:0]) begin
        image_2_103 <= io_pixelVal_in_2_5;
      end else if (10'h67 == _T_28[9:0]) begin
        image_2_103 <= io_pixelVal_in_2_4;
      end else if (10'h67 == _T_25[9:0]) begin
        image_2_103 <= io_pixelVal_in_2_3;
      end else if (10'h67 == _T_22[9:0]) begin
        image_2_103 <= io_pixelVal_in_2_2;
      end else if (10'h67 == _T_19[9:0]) begin
        image_2_103 <= io_pixelVal_in_2_1;
      end else if (10'h67 == _T_15[9:0]) begin
        image_2_103 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_104 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h68 == _T_37[9:0]) begin
        image_2_104 <= io_pixelVal_in_2_7;
      end else if (10'h68 == _T_34[9:0]) begin
        image_2_104 <= io_pixelVal_in_2_6;
      end else if (10'h68 == _T_31[9:0]) begin
        image_2_104 <= io_pixelVal_in_2_5;
      end else if (10'h68 == _T_28[9:0]) begin
        image_2_104 <= io_pixelVal_in_2_4;
      end else if (10'h68 == _T_25[9:0]) begin
        image_2_104 <= io_pixelVal_in_2_3;
      end else if (10'h68 == _T_22[9:0]) begin
        image_2_104 <= io_pixelVal_in_2_2;
      end else if (10'h68 == _T_19[9:0]) begin
        image_2_104 <= io_pixelVal_in_2_1;
      end else if (10'h68 == _T_15[9:0]) begin
        image_2_104 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_105 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h69 == _T_37[9:0]) begin
        image_2_105 <= io_pixelVal_in_2_7;
      end else if (10'h69 == _T_34[9:0]) begin
        image_2_105 <= io_pixelVal_in_2_6;
      end else if (10'h69 == _T_31[9:0]) begin
        image_2_105 <= io_pixelVal_in_2_5;
      end else if (10'h69 == _T_28[9:0]) begin
        image_2_105 <= io_pixelVal_in_2_4;
      end else if (10'h69 == _T_25[9:0]) begin
        image_2_105 <= io_pixelVal_in_2_3;
      end else if (10'h69 == _T_22[9:0]) begin
        image_2_105 <= io_pixelVal_in_2_2;
      end else if (10'h69 == _T_19[9:0]) begin
        image_2_105 <= io_pixelVal_in_2_1;
      end else if (10'h69 == _T_15[9:0]) begin
        image_2_105 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_106 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h6a == _T_37[9:0]) begin
        image_2_106 <= io_pixelVal_in_2_7;
      end else if (10'h6a == _T_34[9:0]) begin
        image_2_106 <= io_pixelVal_in_2_6;
      end else if (10'h6a == _T_31[9:0]) begin
        image_2_106 <= io_pixelVal_in_2_5;
      end else if (10'h6a == _T_28[9:0]) begin
        image_2_106 <= io_pixelVal_in_2_4;
      end else if (10'h6a == _T_25[9:0]) begin
        image_2_106 <= io_pixelVal_in_2_3;
      end else if (10'h6a == _T_22[9:0]) begin
        image_2_106 <= io_pixelVal_in_2_2;
      end else if (10'h6a == _T_19[9:0]) begin
        image_2_106 <= io_pixelVal_in_2_1;
      end else if (10'h6a == _T_15[9:0]) begin
        image_2_106 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_107 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h6b == _T_37[9:0]) begin
        image_2_107 <= io_pixelVal_in_2_7;
      end else if (10'h6b == _T_34[9:0]) begin
        image_2_107 <= io_pixelVal_in_2_6;
      end else if (10'h6b == _T_31[9:0]) begin
        image_2_107 <= io_pixelVal_in_2_5;
      end else if (10'h6b == _T_28[9:0]) begin
        image_2_107 <= io_pixelVal_in_2_4;
      end else if (10'h6b == _T_25[9:0]) begin
        image_2_107 <= io_pixelVal_in_2_3;
      end else if (10'h6b == _T_22[9:0]) begin
        image_2_107 <= io_pixelVal_in_2_2;
      end else if (10'h6b == _T_19[9:0]) begin
        image_2_107 <= io_pixelVal_in_2_1;
      end else if (10'h6b == _T_15[9:0]) begin
        image_2_107 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_108 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h6c == _T_37[9:0]) begin
        image_2_108 <= io_pixelVal_in_2_7;
      end else if (10'h6c == _T_34[9:0]) begin
        image_2_108 <= io_pixelVal_in_2_6;
      end else if (10'h6c == _T_31[9:0]) begin
        image_2_108 <= io_pixelVal_in_2_5;
      end else if (10'h6c == _T_28[9:0]) begin
        image_2_108 <= io_pixelVal_in_2_4;
      end else if (10'h6c == _T_25[9:0]) begin
        image_2_108 <= io_pixelVal_in_2_3;
      end else if (10'h6c == _T_22[9:0]) begin
        image_2_108 <= io_pixelVal_in_2_2;
      end else if (10'h6c == _T_19[9:0]) begin
        image_2_108 <= io_pixelVal_in_2_1;
      end else if (10'h6c == _T_15[9:0]) begin
        image_2_108 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_109 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h6d == _T_37[9:0]) begin
        image_2_109 <= io_pixelVal_in_2_7;
      end else if (10'h6d == _T_34[9:0]) begin
        image_2_109 <= io_pixelVal_in_2_6;
      end else if (10'h6d == _T_31[9:0]) begin
        image_2_109 <= io_pixelVal_in_2_5;
      end else if (10'h6d == _T_28[9:0]) begin
        image_2_109 <= io_pixelVal_in_2_4;
      end else if (10'h6d == _T_25[9:0]) begin
        image_2_109 <= io_pixelVal_in_2_3;
      end else if (10'h6d == _T_22[9:0]) begin
        image_2_109 <= io_pixelVal_in_2_2;
      end else if (10'h6d == _T_19[9:0]) begin
        image_2_109 <= io_pixelVal_in_2_1;
      end else if (10'h6d == _T_15[9:0]) begin
        image_2_109 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_110 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h6e == _T_37[9:0]) begin
        image_2_110 <= io_pixelVal_in_2_7;
      end else if (10'h6e == _T_34[9:0]) begin
        image_2_110 <= io_pixelVal_in_2_6;
      end else if (10'h6e == _T_31[9:0]) begin
        image_2_110 <= io_pixelVal_in_2_5;
      end else if (10'h6e == _T_28[9:0]) begin
        image_2_110 <= io_pixelVal_in_2_4;
      end else if (10'h6e == _T_25[9:0]) begin
        image_2_110 <= io_pixelVal_in_2_3;
      end else if (10'h6e == _T_22[9:0]) begin
        image_2_110 <= io_pixelVal_in_2_2;
      end else if (10'h6e == _T_19[9:0]) begin
        image_2_110 <= io_pixelVal_in_2_1;
      end else if (10'h6e == _T_15[9:0]) begin
        image_2_110 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_111 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h6f == _T_37[9:0]) begin
        image_2_111 <= io_pixelVal_in_2_7;
      end else if (10'h6f == _T_34[9:0]) begin
        image_2_111 <= io_pixelVal_in_2_6;
      end else if (10'h6f == _T_31[9:0]) begin
        image_2_111 <= io_pixelVal_in_2_5;
      end else if (10'h6f == _T_28[9:0]) begin
        image_2_111 <= io_pixelVal_in_2_4;
      end else if (10'h6f == _T_25[9:0]) begin
        image_2_111 <= io_pixelVal_in_2_3;
      end else if (10'h6f == _T_22[9:0]) begin
        image_2_111 <= io_pixelVal_in_2_2;
      end else if (10'h6f == _T_19[9:0]) begin
        image_2_111 <= io_pixelVal_in_2_1;
      end else if (10'h6f == _T_15[9:0]) begin
        image_2_111 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_112 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h70 == _T_37[9:0]) begin
        image_2_112 <= io_pixelVal_in_2_7;
      end else if (10'h70 == _T_34[9:0]) begin
        image_2_112 <= io_pixelVal_in_2_6;
      end else if (10'h70 == _T_31[9:0]) begin
        image_2_112 <= io_pixelVal_in_2_5;
      end else if (10'h70 == _T_28[9:0]) begin
        image_2_112 <= io_pixelVal_in_2_4;
      end else if (10'h70 == _T_25[9:0]) begin
        image_2_112 <= io_pixelVal_in_2_3;
      end else if (10'h70 == _T_22[9:0]) begin
        image_2_112 <= io_pixelVal_in_2_2;
      end else if (10'h70 == _T_19[9:0]) begin
        image_2_112 <= io_pixelVal_in_2_1;
      end else if (10'h70 == _T_15[9:0]) begin
        image_2_112 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_113 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h71 == _T_37[9:0]) begin
        image_2_113 <= io_pixelVal_in_2_7;
      end else if (10'h71 == _T_34[9:0]) begin
        image_2_113 <= io_pixelVal_in_2_6;
      end else if (10'h71 == _T_31[9:0]) begin
        image_2_113 <= io_pixelVal_in_2_5;
      end else if (10'h71 == _T_28[9:0]) begin
        image_2_113 <= io_pixelVal_in_2_4;
      end else if (10'h71 == _T_25[9:0]) begin
        image_2_113 <= io_pixelVal_in_2_3;
      end else if (10'h71 == _T_22[9:0]) begin
        image_2_113 <= io_pixelVal_in_2_2;
      end else if (10'h71 == _T_19[9:0]) begin
        image_2_113 <= io_pixelVal_in_2_1;
      end else if (10'h71 == _T_15[9:0]) begin
        image_2_113 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_114 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h72 == _T_37[9:0]) begin
        image_2_114 <= io_pixelVal_in_2_7;
      end else if (10'h72 == _T_34[9:0]) begin
        image_2_114 <= io_pixelVal_in_2_6;
      end else if (10'h72 == _T_31[9:0]) begin
        image_2_114 <= io_pixelVal_in_2_5;
      end else if (10'h72 == _T_28[9:0]) begin
        image_2_114 <= io_pixelVal_in_2_4;
      end else if (10'h72 == _T_25[9:0]) begin
        image_2_114 <= io_pixelVal_in_2_3;
      end else if (10'h72 == _T_22[9:0]) begin
        image_2_114 <= io_pixelVal_in_2_2;
      end else if (10'h72 == _T_19[9:0]) begin
        image_2_114 <= io_pixelVal_in_2_1;
      end else if (10'h72 == _T_15[9:0]) begin
        image_2_114 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_115 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h73 == _T_37[9:0]) begin
        image_2_115 <= io_pixelVal_in_2_7;
      end else if (10'h73 == _T_34[9:0]) begin
        image_2_115 <= io_pixelVal_in_2_6;
      end else if (10'h73 == _T_31[9:0]) begin
        image_2_115 <= io_pixelVal_in_2_5;
      end else if (10'h73 == _T_28[9:0]) begin
        image_2_115 <= io_pixelVal_in_2_4;
      end else if (10'h73 == _T_25[9:0]) begin
        image_2_115 <= io_pixelVal_in_2_3;
      end else if (10'h73 == _T_22[9:0]) begin
        image_2_115 <= io_pixelVal_in_2_2;
      end else if (10'h73 == _T_19[9:0]) begin
        image_2_115 <= io_pixelVal_in_2_1;
      end else if (10'h73 == _T_15[9:0]) begin
        image_2_115 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_116 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h74 == _T_37[9:0]) begin
        image_2_116 <= io_pixelVal_in_2_7;
      end else if (10'h74 == _T_34[9:0]) begin
        image_2_116 <= io_pixelVal_in_2_6;
      end else if (10'h74 == _T_31[9:0]) begin
        image_2_116 <= io_pixelVal_in_2_5;
      end else if (10'h74 == _T_28[9:0]) begin
        image_2_116 <= io_pixelVal_in_2_4;
      end else if (10'h74 == _T_25[9:0]) begin
        image_2_116 <= io_pixelVal_in_2_3;
      end else if (10'h74 == _T_22[9:0]) begin
        image_2_116 <= io_pixelVal_in_2_2;
      end else if (10'h74 == _T_19[9:0]) begin
        image_2_116 <= io_pixelVal_in_2_1;
      end else if (10'h74 == _T_15[9:0]) begin
        image_2_116 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_117 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h75 == _T_37[9:0]) begin
        image_2_117 <= io_pixelVal_in_2_7;
      end else if (10'h75 == _T_34[9:0]) begin
        image_2_117 <= io_pixelVal_in_2_6;
      end else if (10'h75 == _T_31[9:0]) begin
        image_2_117 <= io_pixelVal_in_2_5;
      end else if (10'h75 == _T_28[9:0]) begin
        image_2_117 <= io_pixelVal_in_2_4;
      end else if (10'h75 == _T_25[9:0]) begin
        image_2_117 <= io_pixelVal_in_2_3;
      end else if (10'h75 == _T_22[9:0]) begin
        image_2_117 <= io_pixelVal_in_2_2;
      end else if (10'h75 == _T_19[9:0]) begin
        image_2_117 <= io_pixelVal_in_2_1;
      end else if (10'h75 == _T_15[9:0]) begin
        image_2_117 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_118 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h76 == _T_37[9:0]) begin
        image_2_118 <= io_pixelVal_in_2_7;
      end else if (10'h76 == _T_34[9:0]) begin
        image_2_118 <= io_pixelVal_in_2_6;
      end else if (10'h76 == _T_31[9:0]) begin
        image_2_118 <= io_pixelVal_in_2_5;
      end else if (10'h76 == _T_28[9:0]) begin
        image_2_118 <= io_pixelVal_in_2_4;
      end else if (10'h76 == _T_25[9:0]) begin
        image_2_118 <= io_pixelVal_in_2_3;
      end else if (10'h76 == _T_22[9:0]) begin
        image_2_118 <= io_pixelVal_in_2_2;
      end else if (10'h76 == _T_19[9:0]) begin
        image_2_118 <= io_pixelVal_in_2_1;
      end else if (10'h76 == _T_15[9:0]) begin
        image_2_118 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_119 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h77 == _T_37[9:0]) begin
        image_2_119 <= io_pixelVal_in_2_7;
      end else if (10'h77 == _T_34[9:0]) begin
        image_2_119 <= io_pixelVal_in_2_6;
      end else if (10'h77 == _T_31[9:0]) begin
        image_2_119 <= io_pixelVal_in_2_5;
      end else if (10'h77 == _T_28[9:0]) begin
        image_2_119 <= io_pixelVal_in_2_4;
      end else if (10'h77 == _T_25[9:0]) begin
        image_2_119 <= io_pixelVal_in_2_3;
      end else if (10'h77 == _T_22[9:0]) begin
        image_2_119 <= io_pixelVal_in_2_2;
      end else if (10'h77 == _T_19[9:0]) begin
        image_2_119 <= io_pixelVal_in_2_1;
      end else if (10'h77 == _T_15[9:0]) begin
        image_2_119 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_120 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h78 == _T_37[9:0]) begin
        image_2_120 <= io_pixelVal_in_2_7;
      end else if (10'h78 == _T_34[9:0]) begin
        image_2_120 <= io_pixelVal_in_2_6;
      end else if (10'h78 == _T_31[9:0]) begin
        image_2_120 <= io_pixelVal_in_2_5;
      end else if (10'h78 == _T_28[9:0]) begin
        image_2_120 <= io_pixelVal_in_2_4;
      end else if (10'h78 == _T_25[9:0]) begin
        image_2_120 <= io_pixelVal_in_2_3;
      end else if (10'h78 == _T_22[9:0]) begin
        image_2_120 <= io_pixelVal_in_2_2;
      end else if (10'h78 == _T_19[9:0]) begin
        image_2_120 <= io_pixelVal_in_2_1;
      end else if (10'h78 == _T_15[9:0]) begin
        image_2_120 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_121 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h79 == _T_37[9:0]) begin
        image_2_121 <= io_pixelVal_in_2_7;
      end else if (10'h79 == _T_34[9:0]) begin
        image_2_121 <= io_pixelVal_in_2_6;
      end else if (10'h79 == _T_31[9:0]) begin
        image_2_121 <= io_pixelVal_in_2_5;
      end else if (10'h79 == _T_28[9:0]) begin
        image_2_121 <= io_pixelVal_in_2_4;
      end else if (10'h79 == _T_25[9:0]) begin
        image_2_121 <= io_pixelVal_in_2_3;
      end else if (10'h79 == _T_22[9:0]) begin
        image_2_121 <= io_pixelVal_in_2_2;
      end else if (10'h79 == _T_19[9:0]) begin
        image_2_121 <= io_pixelVal_in_2_1;
      end else if (10'h79 == _T_15[9:0]) begin
        image_2_121 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_122 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h7a == _T_37[9:0]) begin
        image_2_122 <= io_pixelVal_in_2_7;
      end else if (10'h7a == _T_34[9:0]) begin
        image_2_122 <= io_pixelVal_in_2_6;
      end else if (10'h7a == _T_31[9:0]) begin
        image_2_122 <= io_pixelVal_in_2_5;
      end else if (10'h7a == _T_28[9:0]) begin
        image_2_122 <= io_pixelVal_in_2_4;
      end else if (10'h7a == _T_25[9:0]) begin
        image_2_122 <= io_pixelVal_in_2_3;
      end else if (10'h7a == _T_22[9:0]) begin
        image_2_122 <= io_pixelVal_in_2_2;
      end else if (10'h7a == _T_19[9:0]) begin
        image_2_122 <= io_pixelVal_in_2_1;
      end else if (10'h7a == _T_15[9:0]) begin
        image_2_122 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_123 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h7b == _T_37[9:0]) begin
        image_2_123 <= io_pixelVal_in_2_7;
      end else if (10'h7b == _T_34[9:0]) begin
        image_2_123 <= io_pixelVal_in_2_6;
      end else if (10'h7b == _T_31[9:0]) begin
        image_2_123 <= io_pixelVal_in_2_5;
      end else if (10'h7b == _T_28[9:0]) begin
        image_2_123 <= io_pixelVal_in_2_4;
      end else if (10'h7b == _T_25[9:0]) begin
        image_2_123 <= io_pixelVal_in_2_3;
      end else if (10'h7b == _T_22[9:0]) begin
        image_2_123 <= io_pixelVal_in_2_2;
      end else if (10'h7b == _T_19[9:0]) begin
        image_2_123 <= io_pixelVal_in_2_1;
      end else if (10'h7b == _T_15[9:0]) begin
        image_2_123 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_124 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h7c == _T_37[9:0]) begin
        image_2_124 <= io_pixelVal_in_2_7;
      end else if (10'h7c == _T_34[9:0]) begin
        image_2_124 <= io_pixelVal_in_2_6;
      end else if (10'h7c == _T_31[9:0]) begin
        image_2_124 <= io_pixelVal_in_2_5;
      end else if (10'h7c == _T_28[9:0]) begin
        image_2_124 <= io_pixelVal_in_2_4;
      end else if (10'h7c == _T_25[9:0]) begin
        image_2_124 <= io_pixelVal_in_2_3;
      end else if (10'h7c == _T_22[9:0]) begin
        image_2_124 <= io_pixelVal_in_2_2;
      end else if (10'h7c == _T_19[9:0]) begin
        image_2_124 <= io_pixelVal_in_2_1;
      end else if (10'h7c == _T_15[9:0]) begin
        image_2_124 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_125 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h7d == _T_37[9:0]) begin
        image_2_125 <= io_pixelVal_in_2_7;
      end else if (10'h7d == _T_34[9:0]) begin
        image_2_125 <= io_pixelVal_in_2_6;
      end else if (10'h7d == _T_31[9:0]) begin
        image_2_125 <= io_pixelVal_in_2_5;
      end else if (10'h7d == _T_28[9:0]) begin
        image_2_125 <= io_pixelVal_in_2_4;
      end else if (10'h7d == _T_25[9:0]) begin
        image_2_125 <= io_pixelVal_in_2_3;
      end else if (10'h7d == _T_22[9:0]) begin
        image_2_125 <= io_pixelVal_in_2_2;
      end else if (10'h7d == _T_19[9:0]) begin
        image_2_125 <= io_pixelVal_in_2_1;
      end else if (10'h7d == _T_15[9:0]) begin
        image_2_125 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_126 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h7e == _T_37[9:0]) begin
        image_2_126 <= io_pixelVal_in_2_7;
      end else if (10'h7e == _T_34[9:0]) begin
        image_2_126 <= io_pixelVal_in_2_6;
      end else if (10'h7e == _T_31[9:0]) begin
        image_2_126 <= io_pixelVal_in_2_5;
      end else if (10'h7e == _T_28[9:0]) begin
        image_2_126 <= io_pixelVal_in_2_4;
      end else if (10'h7e == _T_25[9:0]) begin
        image_2_126 <= io_pixelVal_in_2_3;
      end else if (10'h7e == _T_22[9:0]) begin
        image_2_126 <= io_pixelVal_in_2_2;
      end else if (10'h7e == _T_19[9:0]) begin
        image_2_126 <= io_pixelVal_in_2_1;
      end else if (10'h7e == _T_15[9:0]) begin
        image_2_126 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_127 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h7f == _T_37[9:0]) begin
        image_2_127 <= io_pixelVal_in_2_7;
      end else if (10'h7f == _T_34[9:0]) begin
        image_2_127 <= io_pixelVal_in_2_6;
      end else if (10'h7f == _T_31[9:0]) begin
        image_2_127 <= io_pixelVal_in_2_5;
      end else if (10'h7f == _T_28[9:0]) begin
        image_2_127 <= io_pixelVal_in_2_4;
      end else if (10'h7f == _T_25[9:0]) begin
        image_2_127 <= io_pixelVal_in_2_3;
      end else if (10'h7f == _T_22[9:0]) begin
        image_2_127 <= io_pixelVal_in_2_2;
      end else if (10'h7f == _T_19[9:0]) begin
        image_2_127 <= io_pixelVal_in_2_1;
      end else if (10'h7f == _T_15[9:0]) begin
        image_2_127 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_128 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h80 == _T_37[9:0]) begin
        image_2_128 <= io_pixelVal_in_2_7;
      end else if (10'h80 == _T_34[9:0]) begin
        image_2_128 <= io_pixelVal_in_2_6;
      end else if (10'h80 == _T_31[9:0]) begin
        image_2_128 <= io_pixelVal_in_2_5;
      end else if (10'h80 == _T_28[9:0]) begin
        image_2_128 <= io_pixelVal_in_2_4;
      end else if (10'h80 == _T_25[9:0]) begin
        image_2_128 <= io_pixelVal_in_2_3;
      end else if (10'h80 == _T_22[9:0]) begin
        image_2_128 <= io_pixelVal_in_2_2;
      end else if (10'h80 == _T_19[9:0]) begin
        image_2_128 <= io_pixelVal_in_2_1;
      end else if (10'h80 == _T_15[9:0]) begin
        image_2_128 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_129 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h81 == _T_37[9:0]) begin
        image_2_129 <= io_pixelVal_in_2_7;
      end else if (10'h81 == _T_34[9:0]) begin
        image_2_129 <= io_pixelVal_in_2_6;
      end else if (10'h81 == _T_31[9:0]) begin
        image_2_129 <= io_pixelVal_in_2_5;
      end else if (10'h81 == _T_28[9:0]) begin
        image_2_129 <= io_pixelVal_in_2_4;
      end else if (10'h81 == _T_25[9:0]) begin
        image_2_129 <= io_pixelVal_in_2_3;
      end else if (10'h81 == _T_22[9:0]) begin
        image_2_129 <= io_pixelVal_in_2_2;
      end else if (10'h81 == _T_19[9:0]) begin
        image_2_129 <= io_pixelVal_in_2_1;
      end else if (10'h81 == _T_15[9:0]) begin
        image_2_129 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_130 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h82 == _T_37[9:0]) begin
        image_2_130 <= io_pixelVal_in_2_7;
      end else if (10'h82 == _T_34[9:0]) begin
        image_2_130 <= io_pixelVal_in_2_6;
      end else if (10'h82 == _T_31[9:0]) begin
        image_2_130 <= io_pixelVal_in_2_5;
      end else if (10'h82 == _T_28[9:0]) begin
        image_2_130 <= io_pixelVal_in_2_4;
      end else if (10'h82 == _T_25[9:0]) begin
        image_2_130 <= io_pixelVal_in_2_3;
      end else if (10'h82 == _T_22[9:0]) begin
        image_2_130 <= io_pixelVal_in_2_2;
      end else if (10'h82 == _T_19[9:0]) begin
        image_2_130 <= io_pixelVal_in_2_1;
      end else if (10'h82 == _T_15[9:0]) begin
        image_2_130 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_131 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h83 == _T_37[9:0]) begin
        image_2_131 <= io_pixelVal_in_2_7;
      end else if (10'h83 == _T_34[9:0]) begin
        image_2_131 <= io_pixelVal_in_2_6;
      end else if (10'h83 == _T_31[9:0]) begin
        image_2_131 <= io_pixelVal_in_2_5;
      end else if (10'h83 == _T_28[9:0]) begin
        image_2_131 <= io_pixelVal_in_2_4;
      end else if (10'h83 == _T_25[9:0]) begin
        image_2_131 <= io_pixelVal_in_2_3;
      end else if (10'h83 == _T_22[9:0]) begin
        image_2_131 <= io_pixelVal_in_2_2;
      end else if (10'h83 == _T_19[9:0]) begin
        image_2_131 <= io_pixelVal_in_2_1;
      end else if (10'h83 == _T_15[9:0]) begin
        image_2_131 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_132 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h84 == _T_37[9:0]) begin
        image_2_132 <= io_pixelVal_in_2_7;
      end else if (10'h84 == _T_34[9:0]) begin
        image_2_132 <= io_pixelVal_in_2_6;
      end else if (10'h84 == _T_31[9:0]) begin
        image_2_132 <= io_pixelVal_in_2_5;
      end else if (10'h84 == _T_28[9:0]) begin
        image_2_132 <= io_pixelVal_in_2_4;
      end else if (10'h84 == _T_25[9:0]) begin
        image_2_132 <= io_pixelVal_in_2_3;
      end else if (10'h84 == _T_22[9:0]) begin
        image_2_132 <= io_pixelVal_in_2_2;
      end else if (10'h84 == _T_19[9:0]) begin
        image_2_132 <= io_pixelVal_in_2_1;
      end else if (10'h84 == _T_15[9:0]) begin
        image_2_132 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_133 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h85 == _T_37[9:0]) begin
        image_2_133 <= io_pixelVal_in_2_7;
      end else if (10'h85 == _T_34[9:0]) begin
        image_2_133 <= io_pixelVal_in_2_6;
      end else if (10'h85 == _T_31[9:0]) begin
        image_2_133 <= io_pixelVal_in_2_5;
      end else if (10'h85 == _T_28[9:0]) begin
        image_2_133 <= io_pixelVal_in_2_4;
      end else if (10'h85 == _T_25[9:0]) begin
        image_2_133 <= io_pixelVal_in_2_3;
      end else if (10'h85 == _T_22[9:0]) begin
        image_2_133 <= io_pixelVal_in_2_2;
      end else if (10'h85 == _T_19[9:0]) begin
        image_2_133 <= io_pixelVal_in_2_1;
      end else if (10'h85 == _T_15[9:0]) begin
        image_2_133 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_134 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h86 == _T_37[9:0]) begin
        image_2_134 <= io_pixelVal_in_2_7;
      end else if (10'h86 == _T_34[9:0]) begin
        image_2_134 <= io_pixelVal_in_2_6;
      end else if (10'h86 == _T_31[9:0]) begin
        image_2_134 <= io_pixelVal_in_2_5;
      end else if (10'h86 == _T_28[9:0]) begin
        image_2_134 <= io_pixelVal_in_2_4;
      end else if (10'h86 == _T_25[9:0]) begin
        image_2_134 <= io_pixelVal_in_2_3;
      end else if (10'h86 == _T_22[9:0]) begin
        image_2_134 <= io_pixelVal_in_2_2;
      end else if (10'h86 == _T_19[9:0]) begin
        image_2_134 <= io_pixelVal_in_2_1;
      end else if (10'h86 == _T_15[9:0]) begin
        image_2_134 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_135 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h87 == _T_37[9:0]) begin
        image_2_135 <= io_pixelVal_in_2_7;
      end else if (10'h87 == _T_34[9:0]) begin
        image_2_135 <= io_pixelVal_in_2_6;
      end else if (10'h87 == _T_31[9:0]) begin
        image_2_135 <= io_pixelVal_in_2_5;
      end else if (10'h87 == _T_28[9:0]) begin
        image_2_135 <= io_pixelVal_in_2_4;
      end else if (10'h87 == _T_25[9:0]) begin
        image_2_135 <= io_pixelVal_in_2_3;
      end else if (10'h87 == _T_22[9:0]) begin
        image_2_135 <= io_pixelVal_in_2_2;
      end else if (10'h87 == _T_19[9:0]) begin
        image_2_135 <= io_pixelVal_in_2_1;
      end else if (10'h87 == _T_15[9:0]) begin
        image_2_135 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_136 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h88 == _T_37[9:0]) begin
        image_2_136 <= io_pixelVal_in_2_7;
      end else if (10'h88 == _T_34[9:0]) begin
        image_2_136 <= io_pixelVal_in_2_6;
      end else if (10'h88 == _T_31[9:0]) begin
        image_2_136 <= io_pixelVal_in_2_5;
      end else if (10'h88 == _T_28[9:0]) begin
        image_2_136 <= io_pixelVal_in_2_4;
      end else if (10'h88 == _T_25[9:0]) begin
        image_2_136 <= io_pixelVal_in_2_3;
      end else if (10'h88 == _T_22[9:0]) begin
        image_2_136 <= io_pixelVal_in_2_2;
      end else if (10'h88 == _T_19[9:0]) begin
        image_2_136 <= io_pixelVal_in_2_1;
      end else if (10'h88 == _T_15[9:0]) begin
        image_2_136 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_137 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h89 == _T_37[9:0]) begin
        image_2_137 <= io_pixelVal_in_2_7;
      end else if (10'h89 == _T_34[9:0]) begin
        image_2_137 <= io_pixelVal_in_2_6;
      end else if (10'h89 == _T_31[9:0]) begin
        image_2_137 <= io_pixelVal_in_2_5;
      end else if (10'h89 == _T_28[9:0]) begin
        image_2_137 <= io_pixelVal_in_2_4;
      end else if (10'h89 == _T_25[9:0]) begin
        image_2_137 <= io_pixelVal_in_2_3;
      end else if (10'h89 == _T_22[9:0]) begin
        image_2_137 <= io_pixelVal_in_2_2;
      end else if (10'h89 == _T_19[9:0]) begin
        image_2_137 <= io_pixelVal_in_2_1;
      end else if (10'h89 == _T_15[9:0]) begin
        image_2_137 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_138 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h8a == _T_37[9:0]) begin
        image_2_138 <= io_pixelVal_in_2_7;
      end else if (10'h8a == _T_34[9:0]) begin
        image_2_138 <= io_pixelVal_in_2_6;
      end else if (10'h8a == _T_31[9:0]) begin
        image_2_138 <= io_pixelVal_in_2_5;
      end else if (10'h8a == _T_28[9:0]) begin
        image_2_138 <= io_pixelVal_in_2_4;
      end else if (10'h8a == _T_25[9:0]) begin
        image_2_138 <= io_pixelVal_in_2_3;
      end else if (10'h8a == _T_22[9:0]) begin
        image_2_138 <= io_pixelVal_in_2_2;
      end else if (10'h8a == _T_19[9:0]) begin
        image_2_138 <= io_pixelVal_in_2_1;
      end else if (10'h8a == _T_15[9:0]) begin
        image_2_138 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_139 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h8b == _T_37[9:0]) begin
        image_2_139 <= io_pixelVal_in_2_7;
      end else if (10'h8b == _T_34[9:0]) begin
        image_2_139 <= io_pixelVal_in_2_6;
      end else if (10'h8b == _T_31[9:0]) begin
        image_2_139 <= io_pixelVal_in_2_5;
      end else if (10'h8b == _T_28[9:0]) begin
        image_2_139 <= io_pixelVal_in_2_4;
      end else if (10'h8b == _T_25[9:0]) begin
        image_2_139 <= io_pixelVal_in_2_3;
      end else if (10'h8b == _T_22[9:0]) begin
        image_2_139 <= io_pixelVal_in_2_2;
      end else if (10'h8b == _T_19[9:0]) begin
        image_2_139 <= io_pixelVal_in_2_1;
      end else if (10'h8b == _T_15[9:0]) begin
        image_2_139 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_140 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h8c == _T_37[9:0]) begin
        image_2_140 <= io_pixelVal_in_2_7;
      end else if (10'h8c == _T_34[9:0]) begin
        image_2_140 <= io_pixelVal_in_2_6;
      end else if (10'h8c == _T_31[9:0]) begin
        image_2_140 <= io_pixelVal_in_2_5;
      end else if (10'h8c == _T_28[9:0]) begin
        image_2_140 <= io_pixelVal_in_2_4;
      end else if (10'h8c == _T_25[9:0]) begin
        image_2_140 <= io_pixelVal_in_2_3;
      end else if (10'h8c == _T_22[9:0]) begin
        image_2_140 <= io_pixelVal_in_2_2;
      end else if (10'h8c == _T_19[9:0]) begin
        image_2_140 <= io_pixelVal_in_2_1;
      end else if (10'h8c == _T_15[9:0]) begin
        image_2_140 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_141 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h8d == _T_37[9:0]) begin
        image_2_141 <= io_pixelVal_in_2_7;
      end else if (10'h8d == _T_34[9:0]) begin
        image_2_141 <= io_pixelVal_in_2_6;
      end else if (10'h8d == _T_31[9:0]) begin
        image_2_141 <= io_pixelVal_in_2_5;
      end else if (10'h8d == _T_28[9:0]) begin
        image_2_141 <= io_pixelVal_in_2_4;
      end else if (10'h8d == _T_25[9:0]) begin
        image_2_141 <= io_pixelVal_in_2_3;
      end else if (10'h8d == _T_22[9:0]) begin
        image_2_141 <= io_pixelVal_in_2_2;
      end else if (10'h8d == _T_19[9:0]) begin
        image_2_141 <= io_pixelVal_in_2_1;
      end else if (10'h8d == _T_15[9:0]) begin
        image_2_141 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_142 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h8e == _T_37[9:0]) begin
        image_2_142 <= io_pixelVal_in_2_7;
      end else if (10'h8e == _T_34[9:0]) begin
        image_2_142 <= io_pixelVal_in_2_6;
      end else if (10'h8e == _T_31[9:0]) begin
        image_2_142 <= io_pixelVal_in_2_5;
      end else if (10'h8e == _T_28[9:0]) begin
        image_2_142 <= io_pixelVal_in_2_4;
      end else if (10'h8e == _T_25[9:0]) begin
        image_2_142 <= io_pixelVal_in_2_3;
      end else if (10'h8e == _T_22[9:0]) begin
        image_2_142 <= io_pixelVal_in_2_2;
      end else if (10'h8e == _T_19[9:0]) begin
        image_2_142 <= io_pixelVal_in_2_1;
      end else if (10'h8e == _T_15[9:0]) begin
        image_2_142 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_143 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h8f == _T_37[9:0]) begin
        image_2_143 <= io_pixelVal_in_2_7;
      end else if (10'h8f == _T_34[9:0]) begin
        image_2_143 <= io_pixelVal_in_2_6;
      end else if (10'h8f == _T_31[9:0]) begin
        image_2_143 <= io_pixelVal_in_2_5;
      end else if (10'h8f == _T_28[9:0]) begin
        image_2_143 <= io_pixelVal_in_2_4;
      end else if (10'h8f == _T_25[9:0]) begin
        image_2_143 <= io_pixelVal_in_2_3;
      end else if (10'h8f == _T_22[9:0]) begin
        image_2_143 <= io_pixelVal_in_2_2;
      end else if (10'h8f == _T_19[9:0]) begin
        image_2_143 <= io_pixelVal_in_2_1;
      end else if (10'h8f == _T_15[9:0]) begin
        image_2_143 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_144 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h90 == _T_37[9:0]) begin
        image_2_144 <= io_pixelVal_in_2_7;
      end else if (10'h90 == _T_34[9:0]) begin
        image_2_144 <= io_pixelVal_in_2_6;
      end else if (10'h90 == _T_31[9:0]) begin
        image_2_144 <= io_pixelVal_in_2_5;
      end else if (10'h90 == _T_28[9:0]) begin
        image_2_144 <= io_pixelVal_in_2_4;
      end else if (10'h90 == _T_25[9:0]) begin
        image_2_144 <= io_pixelVal_in_2_3;
      end else if (10'h90 == _T_22[9:0]) begin
        image_2_144 <= io_pixelVal_in_2_2;
      end else if (10'h90 == _T_19[9:0]) begin
        image_2_144 <= io_pixelVal_in_2_1;
      end else if (10'h90 == _T_15[9:0]) begin
        image_2_144 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_145 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h91 == _T_37[9:0]) begin
        image_2_145 <= io_pixelVal_in_2_7;
      end else if (10'h91 == _T_34[9:0]) begin
        image_2_145 <= io_pixelVal_in_2_6;
      end else if (10'h91 == _T_31[9:0]) begin
        image_2_145 <= io_pixelVal_in_2_5;
      end else if (10'h91 == _T_28[9:0]) begin
        image_2_145 <= io_pixelVal_in_2_4;
      end else if (10'h91 == _T_25[9:0]) begin
        image_2_145 <= io_pixelVal_in_2_3;
      end else if (10'h91 == _T_22[9:0]) begin
        image_2_145 <= io_pixelVal_in_2_2;
      end else if (10'h91 == _T_19[9:0]) begin
        image_2_145 <= io_pixelVal_in_2_1;
      end else if (10'h91 == _T_15[9:0]) begin
        image_2_145 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_146 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h92 == _T_37[9:0]) begin
        image_2_146 <= io_pixelVal_in_2_7;
      end else if (10'h92 == _T_34[9:0]) begin
        image_2_146 <= io_pixelVal_in_2_6;
      end else if (10'h92 == _T_31[9:0]) begin
        image_2_146 <= io_pixelVal_in_2_5;
      end else if (10'h92 == _T_28[9:0]) begin
        image_2_146 <= io_pixelVal_in_2_4;
      end else if (10'h92 == _T_25[9:0]) begin
        image_2_146 <= io_pixelVal_in_2_3;
      end else if (10'h92 == _T_22[9:0]) begin
        image_2_146 <= io_pixelVal_in_2_2;
      end else if (10'h92 == _T_19[9:0]) begin
        image_2_146 <= io_pixelVal_in_2_1;
      end else if (10'h92 == _T_15[9:0]) begin
        image_2_146 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_147 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h93 == _T_37[9:0]) begin
        image_2_147 <= io_pixelVal_in_2_7;
      end else if (10'h93 == _T_34[9:0]) begin
        image_2_147 <= io_pixelVal_in_2_6;
      end else if (10'h93 == _T_31[9:0]) begin
        image_2_147 <= io_pixelVal_in_2_5;
      end else if (10'h93 == _T_28[9:0]) begin
        image_2_147 <= io_pixelVal_in_2_4;
      end else if (10'h93 == _T_25[9:0]) begin
        image_2_147 <= io_pixelVal_in_2_3;
      end else if (10'h93 == _T_22[9:0]) begin
        image_2_147 <= io_pixelVal_in_2_2;
      end else if (10'h93 == _T_19[9:0]) begin
        image_2_147 <= io_pixelVal_in_2_1;
      end else if (10'h93 == _T_15[9:0]) begin
        image_2_147 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_148 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h94 == _T_37[9:0]) begin
        image_2_148 <= io_pixelVal_in_2_7;
      end else if (10'h94 == _T_34[9:0]) begin
        image_2_148 <= io_pixelVal_in_2_6;
      end else if (10'h94 == _T_31[9:0]) begin
        image_2_148 <= io_pixelVal_in_2_5;
      end else if (10'h94 == _T_28[9:0]) begin
        image_2_148 <= io_pixelVal_in_2_4;
      end else if (10'h94 == _T_25[9:0]) begin
        image_2_148 <= io_pixelVal_in_2_3;
      end else if (10'h94 == _T_22[9:0]) begin
        image_2_148 <= io_pixelVal_in_2_2;
      end else if (10'h94 == _T_19[9:0]) begin
        image_2_148 <= io_pixelVal_in_2_1;
      end else if (10'h94 == _T_15[9:0]) begin
        image_2_148 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_149 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h95 == _T_37[9:0]) begin
        image_2_149 <= io_pixelVal_in_2_7;
      end else if (10'h95 == _T_34[9:0]) begin
        image_2_149 <= io_pixelVal_in_2_6;
      end else if (10'h95 == _T_31[9:0]) begin
        image_2_149 <= io_pixelVal_in_2_5;
      end else if (10'h95 == _T_28[9:0]) begin
        image_2_149 <= io_pixelVal_in_2_4;
      end else if (10'h95 == _T_25[9:0]) begin
        image_2_149 <= io_pixelVal_in_2_3;
      end else if (10'h95 == _T_22[9:0]) begin
        image_2_149 <= io_pixelVal_in_2_2;
      end else if (10'h95 == _T_19[9:0]) begin
        image_2_149 <= io_pixelVal_in_2_1;
      end else if (10'h95 == _T_15[9:0]) begin
        image_2_149 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_150 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h96 == _T_37[9:0]) begin
        image_2_150 <= io_pixelVal_in_2_7;
      end else if (10'h96 == _T_34[9:0]) begin
        image_2_150 <= io_pixelVal_in_2_6;
      end else if (10'h96 == _T_31[9:0]) begin
        image_2_150 <= io_pixelVal_in_2_5;
      end else if (10'h96 == _T_28[9:0]) begin
        image_2_150 <= io_pixelVal_in_2_4;
      end else if (10'h96 == _T_25[9:0]) begin
        image_2_150 <= io_pixelVal_in_2_3;
      end else if (10'h96 == _T_22[9:0]) begin
        image_2_150 <= io_pixelVal_in_2_2;
      end else if (10'h96 == _T_19[9:0]) begin
        image_2_150 <= io_pixelVal_in_2_1;
      end else if (10'h96 == _T_15[9:0]) begin
        image_2_150 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_151 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h97 == _T_37[9:0]) begin
        image_2_151 <= io_pixelVal_in_2_7;
      end else if (10'h97 == _T_34[9:0]) begin
        image_2_151 <= io_pixelVal_in_2_6;
      end else if (10'h97 == _T_31[9:0]) begin
        image_2_151 <= io_pixelVal_in_2_5;
      end else if (10'h97 == _T_28[9:0]) begin
        image_2_151 <= io_pixelVal_in_2_4;
      end else if (10'h97 == _T_25[9:0]) begin
        image_2_151 <= io_pixelVal_in_2_3;
      end else if (10'h97 == _T_22[9:0]) begin
        image_2_151 <= io_pixelVal_in_2_2;
      end else if (10'h97 == _T_19[9:0]) begin
        image_2_151 <= io_pixelVal_in_2_1;
      end else if (10'h97 == _T_15[9:0]) begin
        image_2_151 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_152 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h98 == _T_37[9:0]) begin
        image_2_152 <= io_pixelVal_in_2_7;
      end else if (10'h98 == _T_34[9:0]) begin
        image_2_152 <= io_pixelVal_in_2_6;
      end else if (10'h98 == _T_31[9:0]) begin
        image_2_152 <= io_pixelVal_in_2_5;
      end else if (10'h98 == _T_28[9:0]) begin
        image_2_152 <= io_pixelVal_in_2_4;
      end else if (10'h98 == _T_25[9:0]) begin
        image_2_152 <= io_pixelVal_in_2_3;
      end else if (10'h98 == _T_22[9:0]) begin
        image_2_152 <= io_pixelVal_in_2_2;
      end else if (10'h98 == _T_19[9:0]) begin
        image_2_152 <= io_pixelVal_in_2_1;
      end else if (10'h98 == _T_15[9:0]) begin
        image_2_152 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_153 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h99 == _T_37[9:0]) begin
        image_2_153 <= io_pixelVal_in_2_7;
      end else if (10'h99 == _T_34[9:0]) begin
        image_2_153 <= io_pixelVal_in_2_6;
      end else if (10'h99 == _T_31[9:0]) begin
        image_2_153 <= io_pixelVal_in_2_5;
      end else if (10'h99 == _T_28[9:0]) begin
        image_2_153 <= io_pixelVal_in_2_4;
      end else if (10'h99 == _T_25[9:0]) begin
        image_2_153 <= io_pixelVal_in_2_3;
      end else if (10'h99 == _T_22[9:0]) begin
        image_2_153 <= io_pixelVal_in_2_2;
      end else if (10'h99 == _T_19[9:0]) begin
        image_2_153 <= io_pixelVal_in_2_1;
      end else if (10'h99 == _T_15[9:0]) begin
        image_2_153 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_154 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h9a == _T_37[9:0]) begin
        image_2_154 <= io_pixelVal_in_2_7;
      end else if (10'h9a == _T_34[9:0]) begin
        image_2_154 <= io_pixelVal_in_2_6;
      end else if (10'h9a == _T_31[9:0]) begin
        image_2_154 <= io_pixelVal_in_2_5;
      end else if (10'h9a == _T_28[9:0]) begin
        image_2_154 <= io_pixelVal_in_2_4;
      end else if (10'h9a == _T_25[9:0]) begin
        image_2_154 <= io_pixelVal_in_2_3;
      end else if (10'h9a == _T_22[9:0]) begin
        image_2_154 <= io_pixelVal_in_2_2;
      end else if (10'h9a == _T_19[9:0]) begin
        image_2_154 <= io_pixelVal_in_2_1;
      end else if (10'h9a == _T_15[9:0]) begin
        image_2_154 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_155 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h9b == _T_37[9:0]) begin
        image_2_155 <= io_pixelVal_in_2_7;
      end else if (10'h9b == _T_34[9:0]) begin
        image_2_155 <= io_pixelVal_in_2_6;
      end else if (10'h9b == _T_31[9:0]) begin
        image_2_155 <= io_pixelVal_in_2_5;
      end else if (10'h9b == _T_28[9:0]) begin
        image_2_155 <= io_pixelVal_in_2_4;
      end else if (10'h9b == _T_25[9:0]) begin
        image_2_155 <= io_pixelVal_in_2_3;
      end else if (10'h9b == _T_22[9:0]) begin
        image_2_155 <= io_pixelVal_in_2_2;
      end else if (10'h9b == _T_19[9:0]) begin
        image_2_155 <= io_pixelVal_in_2_1;
      end else if (10'h9b == _T_15[9:0]) begin
        image_2_155 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_156 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h9c == _T_37[9:0]) begin
        image_2_156 <= io_pixelVal_in_2_7;
      end else if (10'h9c == _T_34[9:0]) begin
        image_2_156 <= io_pixelVal_in_2_6;
      end else if (10'h9c == _T_31[9:0]) begin
        image_2_156 <= io_pixelVal_in_2_5;
      end else if (10'h9c == _T_28[9:0]) begin
        image_2_156 <= io_pixelVal_in_2_4;
      end else if (10'h9c == _T_25[9:0]) begin
        image_2_156 <= io_pixelVal_in_2_3;
      end else if (10'h9c == _T_22[9:0]) begin
        image_2_156 <= io_pixelVal_in_2_2;
      end else if (10'h9c == _T_19[9:0]) begin
        image_2_156 <= io_pixelVal_in_2_1;
      end else if (10'h9c == _T_15[9:0]) begin
        image_2_156 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_157 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h9d == _T_37[9:0]) begin
        image_2_157 <= io_pixelVal_in_2_7;
      end else if (10'h9d == _T_34[9:0]) begin
        image_2_157 <= io_pixelVal_in_2_6;
      end else if (10'h9d == _T_31[9:0]) begin
        image_2_157 <= io_pixelVal_in_2_5;
      end else if (10'h9d == _T_28[9:0]) begin
        image_2_157 <= io_pixelVal_in_2_4;
      end else if (10'h9d == _T_25[9:0]) begin
        image_2_157 <= io_pixelVal_in_2_3;
      end else if (10'h9d == _T_22[9:0]) begin
        image_2_157 <= io_pixelVal_in_2_2;
      end else if (10'h9d == _T_19[9:0]) begin
        image_2_157 <= io_pixelVal_in_2_1;
      end else if (10'h9d == _T_15[9:0]) begin
        image_2_157 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_158 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h9e == _T_37[9:0]) begin
        image_2_158 <= io_pixelVal_in_2_7;
      end else if (10'h9e == _T_34[9:0]) begin
        image_2_158 <= io_pixelVal_in_2_6;
      end else if (10'h9e == _T_31[9:0]) begin
        image_2_158 <= io_pixelVal_in_2_5;
      end else if (10'h9e == _T_28[9:0]) begin
        image_2_158 <= io_pixelVal_in_2_4;
      end else if (10'h9e == _T_25[9:0]) begin
        image_2_158 <= io_pixelVal_in_2_3;
      end else if (10'h9e == _T_22[9:0]) begin
        image_2_158 <= io_pixelVal_in_2_2;
      end else if (10'h9e == _T_19[9:0]) begin
        image_2_158 <= io_pixelVal_in_2_1;
      end else if (10'h9e == _T_15[9:0]) begin
        image_2_158 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_159 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h9f == _T_37[9:0]) begin
        image_2_159 <= io_pixelVal_in_2_7;
      end else if (10'h9f == _T_34[9:0]) begin
        image_2_159 <= io_pixelVal_in_2_6;
      end else if (10'h9f == _T_31[9:0]) begin
        image_2_159 <= io_pixelVal_in_2_5;
      end else if (10'h9f == _T_28[9:0]) begin
        image_2_159 <= io_pixelVal_in_2_4;
      end else if (10'h9f == _T_25[9:0]) begin
        image_2_159 <= io_pixelVal_in_2_3;
      end else if (10'h9f == _T_22[9:0]) begin
        image_2_159 <= io_pixelVal_in_2_2;
      end else if (10'h9f == _T_19[9:0]) begin
        image_2_159 <= io_pixelVal_in_2_1;
      end else if (10'h9f == _T_15[9:0]) begin
        image_2_159 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_160 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha0 == _T_37[9:0]) begin
        image_2_160 <= io_pixelVal_in_2_7;
      end else if (10'ha0 == _T_34[9:0]) begin
        image_2_160 <= io_pixelVal_in_2_6;
      end else if (10'ha0 == _T_31[9:0]) begin
        image_2_160 <= io_pixelVal_in_2_5;
      end else if (10'ha0 == _T_28[9:0]) begin
        image_2_160 <= io_pixelVal_in_2_4;
      end else if (10'ha0 == _T_25[9:0]) begin
        image_2_160 <= io_pixelVal_in_2_3;
      end else if (10'ha0 == _T_22[9:0]) begin
        image_2_160 <= io_pixelVal_in_2_2;
      end else if (10'ha0 == _T_19[9:0]) begin
        image_2_160 <= io_pixelVal_in_2_1;
      end else if (10'ha0 == _T_15[9:0]) begin
        image_2_160 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_161 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha1 == _T_37[9:0]) begin
        image_2_161 <= io_pixelVal_in_2_7;
      end else if (10'ha1 == _T_34[9:0]) begin
        image_2_161 <= io_pixelVal_in_2_6;
      end else if (10'ha1 == _T_31[9:0]) begin
        image_2_161 <= io_pixelVal_in_2_5;
      end else if (10'ha1 == _T_28[9:0]) begin
        image_2_161 <= io_pixelVal_in_2_4;
      end else if (10'ha1 == _T_25[9:0]) begin
        image_2_161 <= io_pixelVal_in_2_3;
      end else if (10'ha1 == _T_22[9:0]) begin
        image_2_161 <= io_pixelVal_in_2_2;
      end else if (10'ha1 == _T_19[9:0]) begin
        image_2_161 <= io_pixelVal_in_2_1;
      end else if (10'ha1 == _T_15[9:0]) begin
        image_2_161 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_162 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha2 == _T_37[9:0]) begin
        image_2_162 <= io_pixelVal_in_2_7;
      end else if (10'ha2 == _T_34[9:0]) begin
        image_2_162 <= io_pixelVal_in_2_6;
      end else if (10'ha2 == _T_31[9:0]) begin
        image_2_162 <= io_pixelVal_in_2_5;
      end else if (10'ha2 == _T_28[9:0]) begin
        image_2_162 <= io_pixelVal_in_2_4;
      end else if (10'ha2 == _T_25[9:0]) begin
        image_2_162 <= io_pixelVal_in_2_3;
      end else if (10'ha2 == _T_22[9:0]) begin
        image_2_162 <= io_pixelVal_in_2_2;
      end else if (10'ha2 == _T_19[9:0]) begin
        image_2_162 <= io_pixelVal_in_2_1;
      end else if (10'ha2 == _T_15[9:0]) begin
        image_2_162 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_163 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha3 == _T_37[9:0]) begin
        image_2_163 <= io_pixelVal_in_2_7;
      end else if (10'ha3 == _T_34[9:0]) begin
        image_2_163 <= io_pixelVal_in_2_6;
      end else if (10'ha3 == _T_31[9:0]) begin
        image_2_163 <= io_pixelVal_in_2_5;
      end else if (10'ha3 == _T_28[9:0]) begin
        image_2_163 <= io_pixelVal_in_2_4;
      end else if (10'ha3 == _T_25[9:0]) begin
        image_2_163 <= io_pixelVal_in_2_3;
      end else if (10'ha3 == _T_22[9:0]) begin
        image_2_163 <= io_pixelVal_in_2_2;
      end else if (10'ha3 == _T_19[9:0]) begin
        image_2_163 <= io_pixelVal_in_2_1;
      end else if (10'ha3 == _T_15[9:0]) begin
        image_2_163 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_164 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha4 == _T_37[9:0]) begin
        image_2_164 <= io_pixelVal_in_2_7;
      end else if (10'ha4 == _T_34[9:0]) begin
        image_2_164 <= io_pixelVal_in_2_6;
      end else if (10'ha4 == _T_31[9:0]) begin
        image_2_164 <= io_pixelVal_in_2_5;
      end else if (10'ha4 == _T_28[9:0]) begin
        image_2_164 <= io_pixelVal_in_2_4;
      end else if (10'ha4 == _T_25[9:0]) begin
        image_2_164 <= io_pixelVal_in_2_3;
      end else if (10'ha4 == _T_22[9:0]) begin
        image_2_164 <= io_pixelVal_in_2_2;
      end else if (10'ha4 == _T_19[9:0]) begin
        image_2_164 <= io_pixelVal_in_2_1;
      end else if (10'ha4 == _T_15[9:0]) begin
        image_2_164 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_165 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha5 == _T_37[9:0]) begin
        image_2_165 <= io_pixelVal_in_2_7;
      end else if (10'ha5 == _T_34[9:0]) begin
        image_2_165 <= io_pixelVal_in_2_6;
      end else if (10'ha5 == _T_31[9:0]) begin
        image_2_165 <= io_pixelVal_in_2_5;
      end else if (10'ha5 == _T_28[9:0]) begin
        image_2_165 <= io_pixelVal_in_2_4;
      end else if (10'ha5 == _T_25[9:0]) begin
        image_2_165 <= io_pixelVal_in_2_3;
      end else if (10'ha5 == _T_22[9:0]) begin
        image_2_165 <= io_pixelVal_in_2_2;
      end else if (10'ha5 == _T_19[9:0]) begin
        image_2_165 <= io_pixelVal_in_2_1;
      end else if (10'ha5 == _T_15[9:0]) begin
        image_2_165 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_166 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha6 == _T_37[9:0]) begin
        image_2_166 <= io_pixelVal_in_2_7;
      end else if (10'ha6 == _T_34[9:0]) begin
        image_2_166 <= io_pixelVal_in_2_6;
      end else if (10'ha6 == _T_31[9:0]) begin
        image_2_166 <= io_pixelVal_in_2_5;
      end else if (10'ha6 == _T_28[9:0]) begin
        image_2_166 <= io_pixelVal_in_2_4;
      end else if (10'ha6 == _T_25[9:0]) begin
        image_2_166 <= io_pixelVal_in_2_3;
      end else if (10'ha6 == _T_22[9:0]) begin
        image_2_166 <= io_pixelVal_in_2_2;
      end else if (10'ha6 == _T_19[9:0]) begin
        image_2_166 <= io_pixelVal_in_2_1;
      end else if (10'ha6 == _T_15[9:0]) begin
        image_2_166 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_167 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha7 == _T_37[9:0]) begin
        image_2_167 <= io_pixelVal_in_2_7;
      end else if (10'ha7 == _T_34[9:0]) begin
        image_2_167 <= io_pixelVal_in_2_6;
      end else if (10'ha7 == _T_31[9:0]) begin
        image_2_167 <= io_pixelVal_in_2_5;
      end else if (10'ha7 == _T_28[9:0]) begin
        image_2_167 <= io_pixelVal_in_2_4;
      end else if (10'ha7 == _T_25[9:0]) begin
        image_2_167 <= io_pixelVal_in_2_3;
      end else if (10'ha7 == _T_22[9:0]) begin
        image_2_167 <= io_pixelVal_in_2_2;
      end else if (10'ha7 == _T_19[9:0]) begin
        image_2_167 <= io_pixelVal_in_2_1;
      end else if (10'ha7 == _T_15[9:0]) begin
        image_2_167 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_168 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha8 == _T_37[9:0]) begin
        image_2_168 <= io_pixelVal_in_2_7;
      end else if (10'ha8 == _T_34[9:0]) begin
        image_2_168 <= io_pixelVal_in_2_6;
      end else if (10'ha8 == _T_31[9:0]) begin
        image_2_168 <= io_pixelVal_in_2_5;
      end else if (10'ha8 == _T_28[9:0]) begin
        image_2_168 <= io_pixelVal_in_2_4;
      end else if (10'ha8 == _T_25[9:0]) begin
        image_2_168 <= io_pixelVal_in_2_3;
      end else if (10'ha8 == _T_22[9:0]) begin
        image_2_168 <= io_pixelVal_in_2_2;
      end else if (10'ha8 == _T_19[9:0]) begin
        image_2_168 <= io_pixelVal_in_2_1;
      end else if (10'ha8 == _T_15[9:0]) begin
        image_2_168 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_169 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'ha9 == _T_37[9:0]) begin
        image_2_169 <= io_pixelVal_in_2_7;
      end else if (10'ha9 == _T_34[9:0]) begin
        image_2_169 <= io_pixelVal_in_2_6;
      end else if (10'ha9 == _T_31[9:0]) begin
        image_2_169 <= io_pixelVal_in_2_5;
      end else if (10'ha9 == _T_28[9:0]) begin
        image_2_169 <= io_pixelVal_in_2_4;
      end else if (10'ha9 == _T_25[9:0]) begin
        image_2_169 <= io_pixelVal_in_2_3;
      end else if (10'ha9 == _T_22[9:0]) begin
        image_2_169 <= io_pixelVal_in_2_2;
      end else if (10'ha9 == _T_19[9:0]) begin
        image_2_169 <= io_pixelVal_in_2_1;
      end else if (10'ha9 == _T_15[9:0]) begin
        image_2_169 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_170 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'haa == _T_37[9:0]) begin
        image_2_170 <= io_pixelVal_in_2_7;
      end else if (10'haa == _T_34[9:0]) begin
        image_2_170 <= io_pixelVal_in_2_6;
      end else if (10'haa == _T_31[9:0]) begin
        image_2_170 <= io_pixelVal_in_2_5;
      end else if (10'haa == _T_28[9:0]) begin
        image_2_170 <= io_pixelVal_in_2_4;
      end else if (10'haa == _T_25[9:0]) begin
        image_2_170 <= io_pixelVal_in_2_3;
      end else if (10'haa == _T_22[9:0]) begin
        image_2_170 <= io_pixelVal_in_2_2;
      end else if (10'haa == _T_19[9:0]) begin
        image_2_170 <= io_pixelVal_in_2_1;
      end else if (10'haa == _T_15[9:0]) begin
        image_2_170 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_171 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hab == _T_37[9:0]) begin
        image_2_171 <= io_pixelVal_in_2_7;
      end else if (10'hab == _T_34[9:0]) begin
        image_2_171 <= io_pixelVal_in_2_6;
      end else if (10'hab == _T_31[9:0]) begin
        image_2_171 <= io_pixelVal_in_2_5;
      end else if (10'hab == _T_28[9:0]) begin
        image_2_171 <= io_pixelVal_in_2_4;
      end else if (10'hab == _T_25[9:0]) begin
        image_2_171 <= io_pixelVal_in_2_3;
      end else if (10'hab == _T_22[9:0]) begin
        image_2_171 <= io_pixelVal_in_2_2;
      end else if (10'hab == _T_19[9:0]) begin
        image_2_171 <= io_pixelVal_in_2_1;
      end else if (10'hab == _T_15[9:0]) begin
        image_2_171 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_172 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hac == _T_37[9:0]) begin
        image_2_172 <= io_pixelVal_in_2_7;
      end else if (10'hac == _T_34[9:0]) begin
        image_2_172 <= io_pixelVal_in_2_6;
      end else if (10'hac == _T_31[9:0]) begin
        image_2_172 <= io_pixelVal_in_2_5;
      end else if (10'hac == _T_28[9:0]) begin
        image_2_172 <= io_pixelVal_in_2_4;
      end else if (10'hac == _T_25[9:0]) begin
        image_2_172 <= io_pixelVal_in_2_3;
      end else if (10'hac == _T_22[9:0]) begin
        image_2_172 <= io_pixelVal_in_2_2;
      end else if (10'hac == _T_19[9:0]) begin
        image_2_172 <= io_pixelVal_in_2_1;
      end else if (10'hac == _T_15[9:0]) begin
        image_2_172 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_173 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'had == _T_37[9:0]) begin
        image_2_173 <= io_pixelVal_in_2_7;
      end else if (10'had == _T_34[9:0]) begin
        image_2_173 <= io_pixelVal_in_2_6;
      end else if (10'had == _T_31[9:0]) begin
        image_2_173 <= io_pixelVal_in_2_5;
      end else if (10'had == _T_28[9:0]) begin
        image_2_173 <= io_pixelVal_in_2_4;
      end else if (10'had == _T_25[9:0]) begin
        image_2_173 <= io_pixelVal_in_2_3;
      end else if (10'had == _T_22[9:0]) begin
        image_2_173 <= io_pixelVal_in_2_2;
      end else if (10'had == _T_19[9:0]) begin
        image_2_173 <= io_pixelVal_in_2_1;
      end else if (10'had == _T_15[9:0]) begin
        image_2_173 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_174 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hae == _T_37[9:0]) begin
        image_2_174 <= io_pixelVal_in_2_7;
      end else if (10'hae == _T_34[9:0]) begin
        image_2_174 <= io_pixelVal_in_2_6;
      end else if (10'hae == _T_31[9:0]) begin
        image_2_174 <= io_pixelVal_in_2_5;
      end else if (10'hae == _T_28[9:0]) begin
        image_2_174 <= io_pixelVal_in_2_4;
      end else if (10'hae == _T_25[9:0]) begin
        image_2_174 <= io_pixelVal_in_2_3;
      end else if (10'hae == _T_22[9:0]) begin
        image_2_174 <= io_pixelVal_in_2_2;
      end else if (10'hae == _T_19[9:0]) begin
        image_2_174 <= io_pixelVal_in_2_1;
      end else if (10'hae == _T_15[9:0]) begin
        image_2_174 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_175 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'haf == _T_37[9:0]) begin
        image_2_175 <= io_pixelVal_in_2_7;
      end else if (10'haf == _T_34[9:0]) begin
        image_2_175 <= io_pixelVal_in_2_6;
      end else if (10'haf == _T_31[9:0]) begin
        image_2_175 <= io_pixelVal_in_2_5;
      end else if (10'haf == _T_28[9:0]) begin
        image_2_175 <= io_pixelVal_in_2_4;
      end else if (10'haf == _T_25[9:0]) begin
        image_2_175 <= io_pixelVal_in_2_3;
      end else if (10'haf == _T_22[9:0]) begin
        image_2_175 <= io_pixelVal_in_2_2;
      end else if (10'haf == _T_19[9:0]) begin
        image_2_175 <= io_pixelVal_in_2_1;
      end else if (10'haf == _T_15[9:0]) begin
        image_2_175 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_176 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb0 == _T_37[9:0]) begin
        image_2_176 <= io_pixelVal_in_2_7;
      end else if (10'hb0 == _T_34[9:0]) begin
        image_2_176 <= io_pixelVal_in_2_6;
      end else if (10'hb0 == _T_31[9:0]) begin
        image_2_176 <= io_pixelVal_in_2_5;
      end else if (10'hb0 == _T_28[9:0]) begin
        image_2_176 <= io_pixelVal_in_2_4;
      end else if (10'hb0 == _T_25[9:0]) begin
        image_2_176 <= io_pixelVal_in_2_3;
      end else if (10'hb0 == _T_22[9:0]) begin
        image_2_176 <= io_pixelVal_in_2_2;
      end else if (10'hb0 == _T_19[9:0]) begin
        image_2_176 <= io_pixelVal_in_2_1;
      end else if (10'hb0 == _T_15[9:0]) begin
        image_2_176 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_177 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb1 == _T_37[9:0]) begin
        image_2_177 <= io_pixelVal_in_2_7;
      end else if (10'hb1 == _T_34[9:0]) begin
        image_2_177 <= io_pixelVal_in_2_6;
      end else if (10'hb1 == _T_31[9:0]) begin
        image_2_177 <= io_pixelVal_in_2_5;
      end else if (10'hb1 == _T_28[9:0]) begin
        image_2_177 <= io_pixelVal_in_2_4;
      end else if (10'hb1 == _T_25[9:0]) begin
        image_2_177 <= io_pixelVal_in_2_3;
      end else if (10'hb1 == _T_22[9:0]) begin
        image_2_177 <= io_pixelVal_in_2_2;
      end else if (10'hb1 == _T_19[9:0]) begin
        image_2_177 <= io_pixelVal_in_2_1;
      end else if (10'hb1 == _T_15[9:0]) begin
        image_2_177 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_178 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb2 == _T_37[9:0]) begin
        image_2_178 <= io_pixelVal_in_2_7;
      end else if (10'hb2 == _T_34[9:0]) begin
        image_2_178 <= io_pixelVal_in_2_6;
      end else if (10'hb2 == _T_31[9:0]) begin
        image_2_178 <= io_pixelVal_in_2_5;
      end else if (10'hb2 == _T_28[9:0]) begin
        image_2_178 <= io_pixelVal_in_2_4;
      end else if (10'hb2 == _T_25[9:0]) begin
        image_2_178 <= io_pixelVal_in_2_3;
      end else if (10'hb2 == _T_22[9:0]) begin
        image_2_178 <= io_pixelVal_in_2_2;
      end else if (10'hb2 == _T_19[9:0]) begin
        image_2_178 <= io_pixelVal_in_2_1;
      end else if (10'hb2 == _T_15[9:0]) begin
        image_2_178 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_179 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb3 == _T_37[9:0]) begin
        image_2_179 <= io_pixelVal_in_2_7;
      end else if (10'hb3 == _T_34[9:0]) begin
        image_2_179 <= io_pixelVal_in_2_6;
      end else if (10'hb3 == _T_31[9:0]) begin
        image_2_179 <= io_pixelVal_in_2_5;
      end else if (10'hb3 == _T_28[9:0]) begin
        image_2_179 <= io_pixelVal_in_2_4;
      end else if (10'hb3 == _T_25[9:0]) begin
        image_2_179 <= io_pixelVal_in_2_3;
      end else if (10'hb3 == _T_22[9:0]) begin
        image_2_179 <= io_pixelVal_in_2_2;
      end else if (10'hb3 == _T_19[9:0]) begin
        image_2_179 <= io_pixelVal_in_2_1;
      end else if (10'hb3 == _T_15[9:0]) begin
        image_2_179 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_180 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb4 == _T_37[9:0]) begin
        image_2_180 <= io_pixelVal_in_2_7;
      end else if (10'hb4 == _T_34[9:0]) begin
        image_2_180 <= io_pixelVal_in_2_6;
      end else if (10'hb4 == _T_31[9:0]) begin
        image_2_180 <= io_pixelVal_in_2_5;
      end else if (10'hb4 == _T_28[9:0]) begin
        image_2_180 <= io_pixelVal_in_2_4;
      end else if (10'hb4 == _T_25[9:0]) begin
        image_2_180 <= io_pixelVal_in_2_3;
      end else if (10'hb4 == _T_22[9:0]) begin
        image_2_180 <= io_pixelVal_in_2_2;
      end else if (10'hb4 == _T_19[9:0]) begin
        image_2_180 <= io_pixelVal_in_2_1;
      end else if (10'hb4 == _T_15[9:0]) begin
        image_2_180 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_181 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb5 == _T_37[9:0]) begin
        image_2_181 <= io_pixelVal_in_2_7;
      end else if (10'hb5 == _T_34[9:0]) begin
        image_2_181 <= io_pixelVal_in_2_6;
      end else if (10'hb5 == _T_31[9:0]) begin
        image_2_181 <= io_pixelVal_in_2_5;
      end else if (10'hb5 == _T_28[9:0]) begin
        image_2_181 <= io_pixelVal_in_2_4;
      end else if (10'hb5 == _T_25[9:0]) begin
        image_2_181 <= io_pixelVal_in_2_3;
      end else if (10'hb5 == _T_22[9:0]) begin
        image_2_181 <= io_pixelVal_in_2_2;
      end else if (10'hb5 == _T_19[9:0]) begin
        image_2_181 <= io_pixelVal_in_2_1;
      end else if (10'hb5 == _T_15[9:0]) begin
        image_2_181 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_182 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb6 == _T_37[9:0]) begin
        image_2_182 <= io_pixelVal_in_2_7;
      end else if (10'hb6 == _T_34[9:0]) begin
        image_2_182 <= io_pixelVal_in_2_6;
      end else if (10'hb6 == _T_31[9:0]) begin
        image_2_182 <= io_pixelVal_in_2_5;
      end else if (10'hb6 == _T_28[9:0]) begin
        image_2_182 <= io_pixelVal_in_2_4;
      end else if (10'hb6 == _T_25[9:0]) begin
        image_2_182 <= io_pixelVal_in_2_3;
      end else if (10'hb6 == _T_22[9:0]) begin
        image_2_182 <= io_pixelVal_in_2_2;
      end else if (10'hb6 == _T_19[9:0]) begin
        image_2_182 <= io_pixelVal_in_2_1;
      end else if (10'hb6 == _T_15[9:0]) begin
        image_2_182 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_183 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb7 == _T_37[9:0]) begin
        image_2_183 <= io_pixelVal_in_2_7;
      end else if (10'hb7 == _T_34[9:0]) begin
        image_2_183 <= io_pixelVal_in_2_6;
      end else if (10'hb7 == _T_31[9:0]) begin
        image_2_183 <= io_pixelVal_in_2_5;
      end else if (10'hb7 == _T_28[9:0]) begin
        image_2_183 <= io_pixelVal_in_2_4;
      end else if (10'hb7 == _T_25[9:0]) begin
        image_2_183 <= io_pixelVal_in_2_3;
      end else if (10'hb7 == _T_22[9:0]) begin
        image_2_183 <= io_pixelVal_in_2_2;
      end else if (10'hb7 == _T_19[9:0]) begin
        image_2_183 <= io_pixelVal_in_2_1;
      end else if (10'hb7 == _T_15[9:0]) begin
        image_2_183 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_184 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb8 == _T_37[9:0]) begin
        image_2_184 <= io_pixelVal_in_2_7;
      end else if (10'hb8 == _T_34[9:0]) begin
        image_2_184 <= io_pixelVal_in_2_6;
      end else if (10'hb8 == _T_31[9:0]) begin
        image_2_184 <= io_pixelVal_in_2_5;
      end else if (10'hb8 == _T_28[9:0]) begin
        image_2_184 <= io_pixelVal_in_2_4;
      end else if (10'hb8 == _T_25[9:0]) begin
        image_2_184 <= io_pixelVal_in_2_3;
      end else if (10'hb8 == _T_22[9:0]) begin
        image_2_184 <= io_pixelVal_in_2_2;
      end else if (10'hb8 == _T_19[9:0]) begin
        image_2_184 <= io_pixelVal_in_2_1;
      end else if (10'hb8 == _T_15[9:0]) begin
        image_2_184 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_185 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hb9 == _T_37[9:0]) begin
        image_2_185 <= io_pixelVal_in_2_7;
      end else if (10'hb9 == _T_34[9:0]) begin
        image_2_185 <= io_pixelVal_in_2_6;
      end else if (10'hb9 == _T_31[9:0]) begin
        image_2_185 <= io_pixelVal_in_2_5;
      end else if (10'hb9 == _T_28[9:0]) begin
        image_2_185 <= io_pixelVal_in_2_4;
      end else if (10'hb9 == _T_25[9:0]) begin
        image_2_185 <= io_pixelVal_in_2_3;
      end else if (10'hb9 == _T_22[9:0]) begin
        image_2_185 <= io_pixelVal_in_2_2;
      end else if (10'hb9 == _T_19[9:0]) begin
        image_2_185 <= io_pixelVal_in_2_1;
      end else if (10'hb9 == _T_15[9:0]) begin
        image_2_185 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_186 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hba == _T_37[9:0]) begin
        image_2_186 <= io_pixelVal_in_2_7;
      end else if (10'hba == _T_34[9:0]) begin
        image_2_186 <= io_pixelVal_in_2_6;
      end else if (10'hba == _T_31[9:0]) begin
        image_2_186 <= io_pixelVal_in_2_5;
      end else if (10'hba == _T_28[9:0]) begin
        image_2_186 <= io_pixelVal_in_2_4;
      end else if (10'hba == _T_25[9:0]) begin
        image_2_186 <= io_pixelVal_in_2_3;
      end else if (10'hba == _T_22[9:0]) begin
        image_2_186 <= io_pixelVal_in_2_2;
      end else if (10'hba == _T_19[9:0]) begin
        image_2_186 <= io_pixelVal_in_2_1;
      end else if (10'hba == _T_15[9:0]) begin
        image_2_186 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_187 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hbb == _T_37[9:0]) begin
        image_2_187 <= io_pixelVal_in_2_7;
      end else if (10'hbb == _T_34[9:0]) begin
        image_2_187 <= io_pixelVal_in_2_6;
      end else if (10'hbb == _T_31[9:0]) begin
        image_2_187 <= io_pixelVal_in_2_5;
      end else if (10'hbb == _T_28[9:0]) begin
        image_2_187 <= io_pixelVal_in_2_4;
      end else if (10'hbb == _T_25[9:0]) begin
        image_2_187 <= io_pixelVal_in_2_3;
      end else if (10'hbb == _T_22[9:0]) begin
        image_2_187 <= io_pixelVal_in_2_2;
      end else if (10'hbb == _T_19[9:0]) begin
        image_2_187 <= io_pixelVal_in_2_1;
      end else if (10'hbb == _T_15[9:0]) begin
        image_2_187 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_188 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hbc == _T_37[9:0]) begin
        image_2_188 <= io_pixelVal_in_2_7;
      end else if (10'hbc == _T_34[9:0]) begin
        image_2_188 <= io_pixelVal_in_2_6;
      end else if (10'hbc == _T_31[9:0]) begin
        image_2_188 <= io_pixelVal_in_2_5;
      end else if (10'hbc == _T_28[9:0]) begin
        image_2_188 <= io_pixelVal_in_2_4;
      end else if (10'hbc == _T_25[9:0]) begin
        image_2_188 <= io_pixelVal_in_2_3;
      end else if (10'hbc == _T_22[9:0]) begin
        image_2_188 <= io_pixelVal_in_2_2;
      end else if (10'hbc == _T_19[9:0]) begin
        image_2_188 <= io_pixelVal_in_2_1;
      end else if (10'hbc == _T_15[9:0]) begin
        image_2_188 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_189 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hbd == _T_37[9:0]) begin
        image_2_189 <= io_pixelVal_in_2_7;
      end else if (10'hbd == _T_34[9:0]) begin
        image_2_189 <= io_pixelVal_in_2_6;
      end else if (10'hbd == _T_31[9:0]) begin
        image_2_189 <= io_pixelVal_in_2_5;
      end else if (10'hbd == _T_28[9:0]) begin
        image_2_189 <= io_pixelVal_in_2_4;
      end else if (10'hbd == _T_25[9:0]) begin
        image_2_189 <= io_pixelVal_in_2_3;
      end else if (10'hbd == _T_22[9:0]) begin
        image_2_189 <= io_pixelVal_in_2_2;
      end else if (10'hbd == _T_19[9:0]) begin
        image_2_189 <= io_pixelVal_in_2_1;
      end else if (10'hbd == _T_15[9:0]) begin
        image_2_189 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_190 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hbe == _T_37[9:0]) begin
        image_2_190 <= io_pixelVal_in_2_7;
      end else if (10'hbe == _T_34[9:0]) begin
        image_2_190 <= io_pixelVal_in_2_6;
      end else if (10'hbe == _T_31[9:0]) begin
        image_2_190 <= io_pixelVal_in_2_5;
      end else if (10'hbe == _T_28[9:0]) begin
        image_2_190 <= io_pixelVal_in_2_4;
      end else if (10'hbe == _T_25[9:0]) begin
        image_2_190 <= io_pixelVal_in_2_3;
      end else if (10'hbe == _T_22[9:0]) begin
        image_2_190 <= io_pixelVal_in_2_2;
      end else if (10'hbe == _T_19[9:0]) begin
        image_2_190 <= io_pixelVal_in_2_1;
      end else if (10'hbe == _T_15[9:0]) begin
        image_2_190 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_191 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hbf == _T_37[9:0]) begin
        image_2_191 <= io_pixelVal_in_2_7;
      end else if (10'hbf == _T_34[9:0]) begin
        image_2_191 <= io_pixelVal_in_2_6;
      end else if (10'hbf == _T_31[9:0]) begin
        image_2_191 <= io_pixelVal_in_2_5;
      end else if (10'hbf == _T_28[9:0]) begin
        image_2_191 <= io_pixelVal_in_2_4;
      end else if (10'hbf == _T_25[9:0]) begin
        image_2_191 <= io_pixelVal_in_2_3;
      end else if (10'hbf == _T_22[9:0]) begin
        image_2_191 <= io_pixelVal_in_2_2;
      end else if (10'hbf == _T_19[9:0]) begin
        image_2_191 <= io_pixelVal_in_2_1;
      end else if (10'hbf == _T_15[9:0]) begin
        image_2_191 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_192 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc0 == _T_37[9:0]) begin
        image_2_192 <= io_pixelVal_in_2_7;
      end else if (10'hc0 == _T_34[9:0]) begin
        image_2_192 <= io_pixelVal_in_2_6;
      end else if (10'hc0 == _T_31[9:0]) begin
        image_2_192 <= io_pixelVal_in_2_5;
      end else if (10'hc0 == _T_28[9:0]) begin
        image_2_192 <= io_pixelVal_in_2_4;
      end else if (10'hc0 == _T_25[9:0]) begin
        image_2_192 <= io_pixelVal_in_2_3;
      end else if (10'hc0 == _T_22[9:0]) begin
        image_2_192 <= io_pixelVal_in_2_2;
      end else if (10'hc0 == _T_19[9:0]) begin
        image_2_192 <= io_pixelVal_in_2_1;
      end else if (10'hc0 == _T_15[9:0]) begin
        image_2_192 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_193 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc1 == _T_37[9:0]) begin
        image_2_193 <= io_pixelVal_in_2_7;
      end else if (10'hc1 == _T_34[9:0]) begin
        image_2_193 <= io_pixelVal_in_2_6;
      end else if (10'hc1 == _T_31[9:0]) begin
        image_2_193 <= io_pixelVal_in_2_5;
      end else if (10'hc1 == _T_28[9:0]) begin
        image_2_193 <= io_pixelVal_in_2_4;
      end else if (10'hc1 == _T_25[9:0]) begin
        image_2_193 <= io_pixelVal_in_2_3;
      end else if (10'hc1 == _T_22[9:0]) begin
        image_2_193 <= io_pixelVal_in_2_2;
      end else if (10'hc1 == _T_19[9:0]) begin
        image_2_193 <= io_pixelVal_in_2_1;
      end else if (10'hc1 == _T_15[9:0]) begin
        image_2_193 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_194 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc2 == _T_37[9:0]) begin
        image_2_194 <= io_pixelVal_in_2_7;
      end else if (10'hc2 == _T_34[9:0]) begin
        image_2_194 <= io_pixelVal_in_2_6;
      end else if (10'hc2 == _T_31[9:0]) begin
        image_2_194 <= io_pixelVal_in_2_5;
      end else if (10'hc2 == _T_28[9:0]) begin
        image_2_194 <= io_pixelVal_in_2_4;
      end else if (10'hc2 == _T_25[9:0]) begin
        image_2_194 <= io_pixelVal_in_2_3;
      end else if (10'hc2 == _T_22[9:0]) begin
        image_2_194 <= io_pixelVal_in_2_2;
      end else if (10'hc2 == _T_19[9:0]) begin
        image_2_194 <= io_pixelVal_in_2_1;
      end else if (10'hc2 == _T_15[9:0]) begin
        image_2_194 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_195 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc3 == _T_37[9:0]) begin
        image_2_195 <= io_pixelVal_in_2_7;
      end else if (10'hc3 == _T_34[9:0]) begin
        image_2_195 <= io_pixelVal_in_2_6;
      end else if (10'hc3 == _T_31[9:0]) begin
        image_2_195 <= io_pixelVal_in_2_5;
      end else if (10'hc3 == _T_28[9:0]) begin
        image_2_195 <= io_pixelVal_in_2_4;
      end else if (10'hc3 == _T_25[9:0]) begin
        image_2_195 <= io_pixelVal_in_2_3;
      end else if (10'hc3 == _T_22[9:0]) begin
        image_2_195 <= io_pixelVal_in_2_2;
      end else if (10'hc3 == _T_19[9:0]) begin
        image_2_195 <= io_pixelVal_in_2_1;
      end else if (10'hc3 == _T_15[9:0]) begin
        image_2_195 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_196 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc4 == _T_37[9:0]) begin
        image_2_196 <= io_pixelVal_in_2_7;
      end else if (10'hc4 == _T_34[9:0]) begin
        image_2_196 <= io_pixelVal_in_2_6;
      end else if (10'hc4 == _T_31[9:0]) begin
        image_2_196 <= io_pixelVal_in_2_5;
      end else if (10'hc4 == _T_28[9:0]) begin
        image_2_196 <= io_pixelVal_in_2_4;
      end else if (10'hc4 == _T_25[9:0]) begin
        image_2_196 <= io_pixelVal_in_2_3;
      end else if (10'hc4 == _T_22[9:0]) begin
        image_2_196 <= io_pixelVal_in_2_2;
      end else if (10'hc4 == _T_19[9:0]) begin
        image_2_196 <= io_pixelVal_in_2_1;
      end else if (10'hc4 == _T_15[9:0]) begin
        image_2_196 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_197 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc5 == _T_37[9:0]) begin
        image_2_197 <= io_pixelVal_in_2_7;
      end else if (10'hc5 == _T_34[9:0]) begin
        image_2_197 <= io_pixelVal_in_2_6;
      end else if (10'hc5 == _T_31[9:0]) begin
        image_2_197 <= io_pixelVal_in_2_5;
      end else if (10'hc5 == _T_28[9:0]) begin
        image_2_197 <= io_pixelVal_in_2_4;
      end else if (10'hc5 == _T_25[9:0]) begin
        image_2_197 <= io_pixelVal_in_2_3;
      end else if (10'hc5 == _T_22[9:0]) begin
        image_2_197 <= io_pixelVal_in_2_2;
      end else if (10'hc5 == _T_19[9:0]) begin
        image_2_197 <= io_pixelVal_in_2_1;
      end else if (10'hc5 == _T_15[9:0]) begin
        image_2_197 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_198 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc6 == _T_37[9:0]) begin
        image_2_198 <= io_pixelVal_in_2_7;
      end else if (10'hc6 == _T_34[9:0]) begin
        image_2_198 <= io_pixelVal_in_2_6;
      end else if (10'hc6 == _T_31[9:0]) begin
        image_2_198 <= io_pixelVal_in_2_5;
      end else if (10'hc6 == _T_28[9:0]) begin
        image_2_198 <= io_pixelVal_in_2_4;
      end else if (10'hc6 == _T_25[9:0]) begin
        image_2_198 <= io_pixelVal_in_2_3;
      end else if (10'hc6 == _T_22[9:0]) begin
        image_2_198 <= io_pixelVal_in_2_2;
      end else if (10'hc6 == _T_19[9:0]) begin
        image_2_198 <= io_pixelVal_in_2_1;
      end else if (10'hc6 == _T_15[9:0]) begin
        image_2_198 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_199 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc7 == _T_37[9:0]) begin
        image_2_199 <= io_pixelVal_in_2_7;
      end else if (10'hc7 == _T_34[9:0]) begin
        image_2_199 <= io_pixelVal_in_2_6;
      end else if (10'hc7 == _T_31[9:0]) begin
        image_2_199 <= io_pixelVal_in_2_5;
      end else if (10'hc7 == _T_28[9:0]) begin
        image_2_199 <= io_pixelVal_in_2_4;
      end else if (10'hc7 == _T_25[9:0]) begin
        image_2_199 <= io_pixelVal_in_2_3;
      end else if (10'hc7 == _T_22[9:0]) begin
        image_2_199 <= io_pixelVal_in_2_2;
      end else if (10'hc7 == _T_19[9:0]) begin
        image_2_199 <= io_pixelVal_in_2_1;
      end else if (10'hc7 == _T_15[9:0]) begin
        image_2_199 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_200 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc8 == _T_37[9:0]) begin
        image_2_200 <= io_pixelVal_in_2_7;
      end else if (10'hc8 == _T_34[9:0]) begin
        image_2_200 <= io_pixelVal_in_2_6;
      end else if (10'hc8 == _T_31[9:0]) begin
        image_2_200 <= io_pixelVal_in_2_5;
      end else if (10'hc8 == _T_28[9:0]) begin
        image_2_200 <= io_pixelVal_in_2_4;
      end else if (10'hc8 == _T_25[9:0]) begin
        image_2_200 <= io_pixelVal_in_2_3;
      end else if (10'hc8 == _T_22[9:0]) begin
        image_2_200 <= io_pixelVal_in_2_2;
      end else if (10'hc8 == _T_19[9:0]) begin
        image_2_200 <= io_pixelVal_in_2_1;
      end else if (10'hc8 == _T_15[9:0]) begin
        image_2_200 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_201 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hc9 == _T_37[9:0]) begin
        image_2_201 <= io_pixelVal_in_2_7;
      end else if (10'hc9 == _T_34[9:0]) begin
        image_2_201 <= io_pixelVal_in_2_6;
      end else if (10'hc9 == _T_31[9:0]) begin
        image_2_201 <= io_pixelVal_in_2_5;
      end else if (10'hc9 == _T_28[9:0]) begin
        image_2_201 <= io_pixelVal_in_2_4;
      end else if (10'hc9 == _T_25[9:0]) begin
        image_2_201 <= io_pixelVal_in_2_3;
      end else if (10'hc9 == _T_22[9:0]) begin
        image_2_201 <= io_pixelVal_in_2_2;
      end else if (10'hc9 == _T_19[9:0]) begin
        image_2_201 <= io_pixelVal_in_2_1;
      end else if (10'hc9 == _T_15[9:0]) begin
        image_2_201 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_202 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hca == _T_37[9:0]) begin
        image_2_202 <= io_pixelVal_in_2_7;
      end else if (10'hca == _T_34[9:0]) begin
        image_2_202 <= io_pixelVal_in_2_6;
      end else if (10'hca == _T_31[9:0]) begin
        image_2_202 <= io_pixelVal_in_2_5;
      end else if (10'hca == _T_28[9:0]) begin
        image_2_202 <= io_pixelVal_in_2_4;
      end else if (10'hca == _T_25[9:0]) begin
        image_2_202 <= io_pixelVal_in_2_3;
      end else if (10'hca == _T_22[9:0]) begin
        image_2_202 <= io_pixelVal_in_2_2;
      end else if (10'hca == _T_19[9:0]) begin
        image_2_202 <= io_pixelVal_in_2_1;
      end else if (10'hca == _T_15[9:0]) begin
        image_2_202 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_203 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hcb == _T_37[9:0]) begin
        image_2_203 <= io_pixelVal_in_2_7;
      end else if (10'hcb == _T_34[9:0]) begin
        image_2_203 <= io_pixelVal_in_2_6;
      end else if (10'hcb == _T_31[9:0]) begin
        image_2_203 <= io_pixelVal_in_2_5;
      end else if (10'hcb == _T_28[9:0]) begin
        image_2_203 <= io_pixelVal_in_2_4;
      end else if (10'hcb == _T_25[9:0]) begin
        image_2_203 <= io_pixelVal_in_2_3;
      end else if (10'hcb == _T_22[9:0]) begin
        image_2_203 <= io_pixelVal_in_2_2;
      end else if (10'hcb == _T_19[9:0]) begin
        image_2_203 <= io_pixelVal_in_2_1;
      end else if (10'hcb == _T_15[9:0]) begin
        image_2_203 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_204 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hcc == _T_37[9:0]) begin
        image_2_204 <= io_pixelVal_in_2_7;
      end else if (10'hcc == _T_34[9:0]) begin
        image_2_204 <= io_pixelVal_in_2_6;
      end else if (10'hcc == _T_31[9:0]) begin
        image_2_204 <= io_pixelVal_in_2_5;
      end else if (10'hcc == _T_28[9:0]) begin
        image_2_204 <= io_pixelVal_in_2_4;
      end else if (10'hcc == _T_25[9:0]) begin
        image_2_204 <= io_pixelVal_in_2_3;
      end else if (10'hcc == _T_22[9:0]) begin
        image_2_204 <= io_pixelVal_in_2_2;
      end else if (10'hcc == _T_19[9:0]) begin
        image_2_204 <= io_pixelVal_in_2_1;
      end else if (10'hcc == _T_15[9:0]) begin
        image_2_204 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_205 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hcd == _T_37[9:0]) begin
        image_2_205 <= io_pixelVal_in_2_7;
      end else if (10'hcd == _T_34[9:0]) begin
        image_2_205 <= io_pixelVal_in_2_6;
      end else if (10'hcd == _T_31[9:0]) begin
        image_2_205 <= io_pixelVal_in_2_5;
      end else if (10'hcd == _T_28[9:0]) begin
        image_2_205 <= io_pixelVal_in_2_4;
      end else if (10'hcd == _T_25[9:0]) begin
        image_2_205 <= io_pixelVal_in_2_3;
      end else if (10'hcd == _T_22[9:0]) begin
        image_2_205 <= io_pixelVal_in_2_2;
      end else if (10'hcd == _T_19[9:0]) begin
        image_2_205 <= io_pixelVal_in_2_1;
      end else if (10'hcd == _T_15[9:0]) begin
        image_2_205 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_206 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hce == _T_37[9:0]) begin
        image_2_206 <= io_pixelVal_in_2_7;
      end else if (10'hce == _T_34[9:0]) begin
        image_2_206 <= io_pixelVal_in_2_6;
      end else if (10'hce == _T_31[9:0]) begin
        image_2_206 <= io_pixelVal_in_2_5;
      end else if (10'hce == _T_28[9:0]) begin
        image_2_206 <= io_pixelVal_in_2_4;
      end else if (10'hce == _T_25[9:0]) begin
        image_2_206 <= io_pixelVal_in_2_3;
      end else if (10'hce == _T_22[9:0]) begin
        image_2_206 <= io_pixelVal_in_2_2;
      end else if (10'hce == _T_19[9:0]) begin
        image_2_206 <= io_pixelVal_in_2_1;
      end else if (10'hce == _T_15[9:0]) begin
        image_2_206 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_207 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hcf == _T_37[9:0]) begin
        image_2_207 <= io_pixelVal_in_2_7;
      end else if (10'hcf == _T_34[9:0]) begin
        image_2_207 <= io_pixelVal_in_2_6;
      end else if (10'hcf == _T_31[9:0]) begin
        image_2_207 <= io_pixelVal_in_2_5;
      end else if (10'hcf == _T_28[9:0]) begin
        image_2_207 <= io_pixelVal_in_2_4;
      end else if (10'hcf == _T_25[9:0]) begin
        image_2_207 <= io_pixelVal_in_2_3;
      end else if (10'hcf == _T_22[9:0]) begin
        image_2_207 <= io_pixelVal_in_2_2;
      end else if (10'hcf == _T_19[9:0]) begin
        image_2_207 <= io_pixelVal_in_2_1;
      end else if (10'hcf == _T_15[9:0]) begin
        image_2_207 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_208 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd0 == _T_37[9:0]) begin
        image_2_208 <= io_pixelVal_in_2_7;
      end else if (10'hd0 == _T_34[9:0]) begin
        image_2_208 <= io_pixelVal_in_2_6;
      end else if (10'hd0 == _T_31[9:0]) begin
        image_2_208 <= io_pixelVal_in_2_5;
      end else if (10'hd0 == _T_28[9:0]) begin
        image_2_208 <= io_pixelVal_in_2_4;
      end else if (10'hd0 == _T_25[9:0]) begin
        image_2_208 <= io_pixelVal_in_2_3;
      end else if (10'hd0 == _T_22[9:0]) begin
        image_2_208 <= io_pixelVal_in_2_2;
      end else if (10'hd0 == _T_19[9:0]) begin
        image_2_208 <= io_pixelVal_in_2_1;
      end else if (10'hd0 == _T_15[9:0]) begin
        image_2_208 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_209 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd1 == _T_37[9:0]) begin
        image_2_209 <= io_pixelVal_in_2_7;
      end else if (10'hd1 == _T_34[9:0]) begin
        image_2_209 <= io_pixelVal_in_2_6;
      end else if (10'hd1 == _T_31[9:0]) begin
        image_2_209 <= io_pixelVal_in_2_5;
      end else if (10'hd1 == _T_28[9:0]) begin
        image_2_209 <= io_pixelVal_in_2_4;
      end else if (10'hd1 == _T_25[9:0]) begin
        image_2_209 <= io_pixelVal_in_2_3;
      end else if (10'hd1 == _T_22[9:0]) begin
        image_2_209 <= io_pixelVal_in_2_2;
      end else if (10'hd1 == _T_19[9:0]) begin
        image_2_209 <= io_pixelVal_in_2_1;
      end else if (10'hd1 == _T_15[9:0]) begin
        image_2_209 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_210 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd2 == _T_37[9:0]) begin
        image_2_210 <= io_pixelVal_in_2_7;
      end else if (10'hd2 == _T_34[9:0]) begin
        image_2_210 <= io_pixelVal_in_2_6;
      end else if (10'hd2 == _T_31[9:0]) begin
        image_2_210 <= io_pixelVal_in_2_5;
      end else if (10'hd2 == _T_28[9:0]) begin
        image_2_210 <= io_pixelVal_in_2_4;
      end else if (10'hd2 == _T_25[9:0]) begin
        image_2_210 <= io_pixelVal_in_2_3;
      end else if (10'hd2 == _T_22[9:0]) begin
        image_2_210 <= io_pixelVal_in_2_2;
      end else if (10'hd2 == _T_19[9:0]) begin
        image_2_210 <= io_pixelVal_in_2_1;
      end else if (10'hd2 == _T_15[9:0]) begin
        image_2_210 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_211 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd3 == _T_37[9:0]) begin
        image_2_211 <= io_pixelVal_in_2_7;
      end else if (10'hd3 == _T_34[9:0]) begin
        image_2_211 <= io_pixelVal_in_2_6;
      end else if (10'hd3 == _T_31[9:0]) begin
        image_2_211 <= io_pixelVal_in_2_5;
      end else if (10'hd3 == _T_28[9:0]) begin
        image_2_211 <= io_pixelVal_in_2_4;
      end else if (10'hd3 == _T_25[9:0]) begin
        image_2_211 <= io_pixelVal_in_2_3;
      end else if (10'hd3 == _T_22[9:0]) begin
        image_2_211 <= io_pixelVal_in_2_2;
      end else if (10'hd3 == _T_19[9:0]) begin
        image_2_211 <= io_pixelVal_in_2_1;
      end else if (10'hd3 == _T_15[9:0]) begin
        image_2_211 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_212 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd4 == _T_37[9:0]) begin
        image_2_212 <= io_pixelVal_in_2_7;
      end else if (10'hd4 == _T_34[9:0]) begin
        image_2_212 <= io_pixelVal_in_2_6;
      end else if (10'hd4 == _T_31[9:0]) begin
        image_2_212 <= io_pixelVal_in_2_5;
      end else if (10'hd4 == _T_28[9:0]) begin
        image_2_212 <= io_pixelVal_in_2_4;
      end else if (10'hd4 == _T_25[9:0]) begin
        image_2_212 <= io_pixelVal_in_2_3;
      end else if (10'hd4 == _T_22[9:0]) begin
        image_2_212 <= io_pixelVal_in_2_2;
      end else if (10'hd4 == _T_19[9:0]) begin
        image_2_212 <= io_pixelVal_in_2_1;
      end else if (10'hd4 == _T_15[9:0]) begin
        image_2_212 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_213 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd5 == _T_37[9:0]) begin
        image_2_213 <= io_pixelVal_in_2_7;
      end else if (10'hd5 == _T_34[9:0]) begin
        image_2_213 <= io_pixelVal_in_2_6;
      end else if (10'hd5 == _T_31[9:0]) begin
        image_2_213 <= io_pixelVal_in_2_5;
      end else if (10'hd5 == _T_28[9:0]) begin
        image_2_213 <= io_pixelVal_in_2_4;
      end else if (10'hd5 == _T_25[9:0]) begin
        image_2_213 <= io_pixelVal_in_2_3;
      end else if (10'hd5 == _T_22[9:0]) begin
        image_2_213 <= io_pixelVal_in_2_2;
      end else if (10'hd5 == _T_19[9:0]) begin
        image_2_213 <= io_pixelVal_in_2_1;
      end else if (10'hd5 == _T_15[9:0]) begin
        image_2_213 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_214 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd6 == _T_37[9:0]) begin
        image_2_214 <= io_pixelVal_in_2_7;
      end else if (10'hd6 == _T_34[9:0]) begin
        image_2_214 <= io_pixelVal_in_2_6;
      end else if (10'hd6 == _T_31[9:0]) begin
        image_2_214 <= io_pixelVal_in_2_5;
      end else if (10'hd6 == _T_28[9:0]) begin
        image_2_214 <= io_pixelVal_in_2_4;
      end else if (10'hd6 == _T_25[9:0]) begin
        image_2_214 <= io_pixelVal_in_2_3;
      end else if (10'hd6 == _T_22[9:0]) begin
        image_2_214 <= io_pixelVal_in_2_2;
      end else if (10'hd6 == _T_19[9:0]) begin
        image_2_214 <= io_pixelVal_in_2_1;
      end else if (10'hd6 == _T_15[9:0]) begin
        image_2_214 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_215 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd7 == _T_37[9:0]) begin
        image_2_215 <= io_pixelVal_in_2_7;
      end else if (10'hd7 == _T_34[9:0]) begin
        image_2_215 <= io_pixelVal_in_2_6;
      end else if (10'hd7 == _T_31[9:0]) begin
        image_2_215 <= io_pixelVal_in_2_5;
      end else if (10'hd7 == _T_28[9:0]) begin
        image_2_215 <= io_pixelVal_in_2_4;
      end else if (10'hd7 == _T_25[9:0]) begin
        image_2_215 <= io_pixelVal_in_2_3;
      end else if (10'hd7 == _T_22[9:0]) begin
        image_2_215 <= io_pixelVal_in_2_2;
      end else if (10'hd7 == _T_19[9:0]) begin
        image_2_215 <= io_pixelVal_in_2_1;
      end else if (10'hd7 == _T_15[9:0]) begin
        image_2_215 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_216 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd8 == _T_37[9:0]) begin
        image_2_216 <= io_pixelVal_in_2_7;
      end else if (10'hd8 == _T_34[9:0]) begin
        image_2_216 <= io_pixelVal_in_2_6;
      end else if (10'hd8 == _T_31[9:0]) begin
        image_2_216 <= io_pixelVal_in_2_5;
      end else if (10'hd8 == _T_28[9:0]) begin
        image_2_216 <= io_pixelVal_in_2_4;
      end else if (10'hd8 == _T_25[9:0]) begin
        image_2_216 <= io_pixelVal_in_2_3;
      end else if (10'hd8 == _T_22[9:0]) begin
        image_2_216 <= io_pixelVal_in_2_2;
      end else if (10'hd8 == _T_19[9:0]) begin
        image_2_216 <= io_pixelVal_in_2_1;
      end else if (10'hd8 == _T_15[9:0]) begin
        image_2_216 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_217 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hd9 == _T_37[9:0]) begin
        image_2_217 <= io_pixelVal_in_2_7;
      end else if (10'hd9 == _T_34[9:0]) begin
        image_2_217 <= io_pixelVal_in_2_6;
      end else if (10'hd9 == _T_31[9:0]) begin
        image_2_217 <= io_pixelVal_in_2_5;
      end else if (10'hd9 == _T_28[9:0]) begin
        image_2_217 <= io_pixelVal_in_2_4;
      end else if (10'hd9 == _T_25[9:0]) begin
        image_2_217 <= io_pixelVal_in_2_3;
      end else if (10'hd9 == _T_22[9:0]) begin
        image_2_217 <= io_pixelVal_in_2_2;
      end else if (10'hd9 == _T_19[9:0]) begin
        image_2_217 <= io_pixelVal_in_2_1;
      end else if (10'hd9 == _T_15[9:0]) begin
        image_2_217 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_218 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hda == _T_37[9:0]) begin
        image_2_218 <= io_pixelVal_in_2_7;
      end else if (10'hda == _T_34[9:0]) begin
        image_2_218 <= io_pixelVal_in_2_6;
      end else if (10'hda == _T_31[9:0]) begin
        image_2_218 <= io_pixelVal_in_2_5;
      end else if (10'hda == _T_28[9:0]) begin
        image_2_218 <= io_pixelVal_in_2_4;
      end else if (10'hda == _T_25[9:0]) begin
        image_2_218 <= io_pixelVal_in_2_3;
      end else if (10'hda == _T_22[9:0]) begin
        image_2_218 <= io_pixelVal_in_2_2;
      end else if (10'hda == _T_19[9:0]) begin
        image_2_218 <= io_pixelVal_in_2_1;
      end else if (10'hda == _T_15[9:0]) begin
        image_2_218 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_219 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hdb == _T_37[9:0]) begin
        image_2_219 <= io_pixelVal_in_2_7;
      end else if (10'hdb == _T_34[9:0]) begin
        image_2_219 <= io_pixelVal_in_2_6;
      end else if (10'hdb == _T_31[9:0]) begin
        image_2_219 <= io_pixelVal_in_2_5;
      end else if (10'hdb == _T_28[9:0]) begin
        image_2_219 <= io_pixelVal_in_2_4;
      end else if (10'hdb == _T_25[9:0]) begin
        image_2_219 <= io_pixelVal_in_2_3;
      end else if (10'hdb == _T_22[9:0]) begin
        image_2_219 <= io_pixelVal_in_2_2;
      end else if (10'hdb == _T_19[9:0]) begin
        image_2_219 <= io_pixelVal_in_2_1;
      end else if (10'hdb == _T_15[9:0]) begin
        image_2_219 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_220 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hdc == _T_37[9:0]) begin
        image_2_220 <= io_pixelVal_in_2_7;
      end else if (10'hdc == _T_34[9:0]) begin
        image_2_220 <= io_pixelVal_in_2_6;
      end else if (10'hdc == _T_31[9:0]) begin
        image_2_220 <= io_pixelVal_in_2_5;
      end else if (10'hdc == _T_28[9:0]) begin
        image_2_220 <= io_pixelVal_in_2_4;
      end else if (10'hdc == _T_25[9:0]) begin
        image_2_220 <= io_pixelVal_in_2_3;
      end else if (10'hdc == _T_22[9:0]) begin
        image_2_220 <= io_pixelVal_in_2_2;
      end else if (10'hdc == _T_19[9:0]) begin
        image_2_220 <= io_pixelVal_in_2_1;
      end else if (10'hdc == _T_15[9:0]) begin
        image_2_220 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_221 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hdd == _T_37[9:0]) begin
        image_2_221 <= io_pixelVal_in_2_7;
      end else if (10'hdd == _T_34[9:0]) begin
        image_2_221 <= io_pixelVal_in_2_6;
      end else if (10'hdd == _T_31[9:0]) begin
        image_2_221 <= io_pixelVal_in_2_5;
      end else if (10'hdd == _T_28[9:0]) begin
        image_2_221 <= io_pixelVal_in_2_4;
      end else if (10'hdd == _T_25[9:0]) begin
        image_2_221 <= io_pixelVal_in_2_3;
      end else if (10'hdd == _T_22[9:0]) begin
        image_2_221 <= io_pixelVal_in_2_2;
      end else if (10'hdd == _T_19[9:0]) begin
        image_2_221 <= io_pixelVal_in_2_1;
      end else if (10'hdd == _T_15[9:0]) begin
        image_2_221 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_222 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hde == _T_37[9:0]) begin
        image_2_222 <= io_pixelVal_in_2_7;
      end else if (10'hde == _T_34[9:0]) begin
        image_2_222 <= io_pixelVal_in_2_6;
      end else if (10'hde == _T_31[9:0]) begin
        image_2_222 <= io_pixelVal_in_2_5;
      end else if (10'hde == _T_28[9:0]) begin
        image_2_222 <= io_pixelVal_in_2_4;
      end else if (10'hde == _T_25[9:0]) begin
        image_2_222 <= io_pixelVal_in_2_3;
      end else if (10'hde == _T_22[9:0]) begin
        image_2_222 <= io_pixelVal_in_2_2;
      end else if (10'hde == _T_19[9:0]) begin
        image_2_222 <= io_pixelVal_in_2_1;
      end else if (10'hde == _T_15[9:0]) begin
        image_2_222 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_223 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hdf == _T_37[9:0]) begin
        image_2_223 <= io_pixelVal_in_2_7;
      end else if (10'hdf == _T_34[9:0]) begin
        image_2_223 <= io_pixelVal_in_2_6;
      end else if (10'hdf == _T_31[9:0]) begin
        image_2_223 <= io_pixelVal_in_2_5;
      end else if (10'hdf == _T_28[9:0]) begin
        image_2_223 <= io_pixelVal_in_2_4;
      end else if (10'hdf == _T_25[9:0]) begin
        image_2_223 <= io_pixelVal_in_2_3;
      end else if (10'hdf == _T_22[9:0]) begin
        image_2_223 <= io_pixelVal_in_2_2;
      end else if (10'hdf == _T_19[9:0]) begin
        image_2_223 <= io_pixelVal_in_2_1;
      end else if (10'hdf == _T_15[9:0]) begin
        image_2_223 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_224 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he0 == _T_37[9:0]) begin
        image_2_224 <= io_pixelVal_in_2_7;
      end else if (10'he0 == _T_34[9:0]) begin
        image_2_224 <= io_pixelVal_in_2_6;
      end else if (10'he0 == _T_31[9:0]) begin
        image_2_224 <= io_pixelVal_in_2_5;
      end else if (10'he0 == _T_28[9:0]) begin
        image_2_224 <= io_pixelVal_in_2_4;
      end else if (10'he0 == _T_25[9:0]) begin
        image_2_224 <= io_pixelVal_in_2_3;
      end else if (10'he0 == _T_22[9:0]) begin
        image_2_224 <= io_pixelVal_in_2_2;
      end else if (10'he0 == _T_19[9:0]) begin
        image_2_224 <= io_pixelVal_in_2_1;
      end else if (10'he0 == _T_15[9:0]) begin
        image_2_224 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_225 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he1 == _T_37[9:0]) begin
        image_2_225 <= io_pixelVal_in_2_7;
      end else if (10'he1 == _T_34[9:0]) begin
        image_2_225 <= io_pixelVal_in_2_6;
      end else if (10'he1 == _T_31[9:0]) begin
        image_2_225 <= io_pixelVal_in_2_5;
      end else if (10'he1 == _T_28[9:0]) begin
        image_2_225 <= io_pixelVal_in_2_4;
      end else if (10'he1 == _T_25[9:0]) begin
        image_2_225 <= io_pixelVal_in_2_3;
      end else if (10'he1 == _T_22[9:0]) begin
        image_2_225 <= io_pixelVal_in_2_2;
      end else if (10'he1 == _T_19[9:0]) begin
        image_2_225 <= io_pixelVal_in_2_1;
      end else if (10'he1 == _T_15[9:0]) begin
        image_2_225 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_226 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he2 == _T_37[9:0]) begin
        image_2_226 <= io_pixelVal_in_2_7;
      end else if (10'he2 == _T_34[9:0]) begin
        image_2_226 <= io_pixelVal_in_2_6;
      end else if (10'he2 == _T_31[9:0]) begin
        image_2_226 <= io_pixelVal_in_2_5;
      end else if (10'he2 == _T_28[9:0]) begin
        image_2_226 <= io_pixelVal_in_2_4;
      end else if (10'he2 == _T_25[9:0]) begin
        image_2_226 <= io_pixelVal_in_2_3;
      end else if (10'he2 == _T_22[9:0]) begin
        image_2_226 <= io_pixelVal_in_2_2;
      end else if (10'he2 == _T_19[9:0]) begin
        image_2_226 <= io_pixelVal_in_2_1;
      end else if (10'he2 == _T_15[9:0]) begin
        image_2_226 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_227 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he3 == _T_37[9:0]) begin
        image_2_227 <= io_pixelVal_in_2_7;
      end else if (10'he3 == _T_34[9:0]) begin
        image_2_227 <= io_pixelVal_in_2_6;
      end else if (10'he3 == _T_31[9:0]) begin
        image_2_227 <= io_pixelVal_in_2_5;
      end else if (10'he3 == _T_28[9:0]) begin
        image_2_227 <= io_pixelVal_in_2_4;
      end else if (10'he3 == _T_25[9:0]) begin
        image_2_227 <= io_pixelVal_in_2_3;
      end else if (10'he3 == _T_22[9:0]) begin
        image_2_227 <= io_pixelVal_in_2_2;
      end else if (10'he3 == _T_19[9:0]) begin
        image_2_227 <= io_pixelVal_in_2_1;
      end else if (10'he3 == _T_15[9:0]) begin
        image_2_227 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_228 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he4 == _T_37[9:0]) begin
        image_2_228 <= io_pixelVal_in_2_7;
      end else if (10'he4 == _T_34[9:0]) begin
        image_2_228 <= io_pixelVal_in_2_6;
      end else if (10'he4 == _T_31[9:0]) begin
        image_2_228 <= io_pixelVal_in_2_5;
      end else if (10'he4 == _T_28[9:0]) begin
        image_2_228 <= io_pixelVal_in_2_4;
      end else if (10'he4 == _T_25[9:0]) begin
        image_2_228 <= io_pixelVal_in_2_3;
      end else if (10'he4 == _T_22[9:0]) begin
        image_2_228 <= io_pixelVal_in_2_2;
      end else if (10'he4 == _T_19[9:0]) begin
        image_2_228 <= io_pixelVal_in_2_1;
      end else if (10'he4 == _T_15[9:0]) begin
        image_2_228 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_229 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he5 == _T_37[9:0]) begin
        image_2_229 <= io_pixelVal_in_2_7;
      end else if (10'he5 == _T_34[9:0]) begin
        image_2_229 <= io_pixelVal_in_2_6;
      end else if (10'he5 == _T_31[9:0]) begin
        image_2_229 <= io_pixelVal_in_2_5;
      end else if (10'he5 == _T_28[9:0]) begin
        image_2_229 <= io_pixelVal_in_2_4;
      end else if (10'he5 == _T_25[9:0]) begin
        image_2_229 <= io_pixelVal_in_2_3;
      end else if (10'he5 == _T_22[9:0]) begin
        image_2_229 <= io_pixelVal_in_2_2;
      end else if (10'he5 == _T_19[9:0]) begin
        image_2_229 <= io_pixelVal_in_2_1;
      end else if (10'he5 == _T_15[9:0]) begin
        image_2_229 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_230 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he6 == _T_37[9:0]) begin
        image_2_230 <= io_pixelVal_in_2_7;
      end else if (10'he6 == _T_34[9:0]) begin
        image_2_230 <= io_pixelVal_in_2_6;
      end else if (10'he6 == _T_31[9:0]) begin
        image_2_230 <= io_pixelVal_in_2_5;
      end else if (10'he6 == _T_28[9:0]) begin
        image_2_230 <= io_pixelVal_in_2_4;
      end else if (10'he6 == _T_25[9:0]) begin
        image_2_230 <= io_pixelVal_in_2_3;
      end else if (10'he6 == _T_22[9:0]) begin
        image_2_230 <= io_pixelVal_in_2_2;
      end else if (10'he6 == _T_19[9:0]) begin
        image_2_230 <= io_pixelVal_in_2_1;
      end else if (10'he6 == _T_15[9:0]) begin
        image_2_230 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_231 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he7 == _T_37[9:0]) begin
        image_2_231 <= io_pixelVal_in_2_7;
      end else if (10'he7 == _T_34[9:0]) begin
        image_2_231 <= io_pixelVal_in_2_6;
      end else if (10'he7 == _T_31[9:0]) begin
        image_2_231 <= io_pixelVal_in_2_5;
      end else if (10'he7 == _T_28[9:0]) begin
        image_2_231 <= io_pixelVal_in_2_4;
      end else if (10'he7 == _T_25[9:0]) begin
        image_2_231 <= io_pixelVal_in_2_3;
      end else if (10'he7 == _T_22[9:0]) begin
        image_2_231 <= io_pixelVal_in_2_2;
      end else if (10'he7 == _T_19[9:0]) begin
        image_2_231 <= io_pixelVal_in_2_1;
      end else if (10'he7 == _T_15[9:0]) begin
        image_2_231 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_232 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he8 == _T_37[9:0]) begin
        image_2_232 <= io_pixelVal_in_2_7;
      end else if (10'he8 == _T_34[9:0]) begin
        image_2_232 <= io_pixelVal_in_2_6;
      end else if (10'he8 == _T_31[9:0]) begin
        image_2_232 <= io_pixelVal_in_2_5;
      end else if (10'he8 == _T_28[9:0]) begin
        image_2_232 <= io_pixelVal_in_2_4;
      end else if (10'he8 == _T_25[9:0]) begin
        image_2_232 <= io_pixelVal_in_2_3;
      end else if (10'he8 == _T_22[9:0]) begin
        image_2_232 <= io_pixelVal_in_2_2;
      end else if (10'he8 == _T_19[9:0]) begin
        image_2_232 <= io_pixelVal_in_2_1;
      end else if (10'he8 == _T_15[9:0]) begin
        image_2_232 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_233 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'he9 == _T_37[9:0]) begin
        image_2_233 <= io_pixelVal_in_2_7;
      end else if (10'he9 == _T_34[9:0]) begin
        image_2_233 <= io_pixelVal_in_2_6;
      end else if (10'he9 == _T_31[9:0]) begin
        image_2_233 <= io_pixelVal_in_2_5;
      end else if (10'he9 == _T_28[9:0]) begin
        image_2_233 <= io_pixelVal_in_2_4;
      end else if (10'he9 == _T_25[9:0]) begin
        image_2_233 <= io_pixelVal_in_2_3;
      end else if (10'he9 == _T_22[9:0]) begin
        image_2_233 <= io_pixelVal_in_2_2;
      end else if (10'he9 == _T_19[9:0]) begin
        image_2_233 <= io_pixelVal_in_2_1;
      end else if (10'he9 == _T_15[9:0]) begin
        image_2_233 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_234 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hea == _T_37[9:0]) begin
        image_2_234 <= io_pixelVal_in_2_7;
      end else if (10'hea == _T_34[9:0]) begin
        image_2_234 <= io_pixelVal_in_2_6;
      end else if (10'hea == _T_31[9:0]) begin
        image_2_234 <= io_pixelVal_in_2_5;
      end else if (10'hea == _T_28[9:0]) begin
        image_2_234 <= io_pixelVal_in_2_4;
      end else if (10'hea == _T_25[9:0]) begin
        image_2_234 <= io_pixelVal_in_2_3;
      end else if (10'hea == _T_22[9:0]) begin
        image_2_234 <= io_pixelVal_in_2_2;
      end else if (10'hea == _T_19[9:0]) begin
        image_2_234 <= io_pixelVal_in_2_1;
      end else if (10'hea == _T_15[9:0]) begin
        image_2_234 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_235 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'heb == _T_37[9:0]) begin
        image_2_235 <= io_pixelVal_in_2_7;
      end else if (10'heb == _T_34[9:0]) begin
        image_2_235 <= io_pixelVal_in_2_6;
      end else if (10'heb == _T_31[9:0]) begin
        image_2_235 <= io_pixelVal_in_2_5;
      end else if (10'heb == _T_28[9:0]) begin
        image_2_235 <= io_pixelVal_in_2_4;
      end else if (10'heb == _T_25[9:0]) begin
        image_2_235 <= io_pixelVal_in_2_3;
      end else if (10'heb == _T_22[9:0]) begin
        image_2_235 <= io_pixelVal_in_2_2;
      end else if (10'heb == _T_19[9:0]) begin
        image_2_235 <= io_pixelVal_in_2_1;
      end else if (10'heb == _T_15[9:0]) begin
        image_2_235 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_236 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hec == _T_37[9:0]) begin
        image_2_236 <= io_pixelVal_in_2_7;
      end else if (10'hec == _T_34[9:0]) begin
        image_2_236 <= io_pixelVal_in_2_6;
      end else if (10'hec == _T_31[9:0]) begin
        image_2_236 <= io_pixelVal_in_2_5;
      end else if (10'hec == _T_28[9:0]) begin
        image_2_236 <= io_pixelVal_in_2_4;
      end else if (10'hec == _T_25[9:0]) begin
        image_2_236 <= io_pixelVal_in_2_3;
      end else if (10'hec == _T_22[9:0]) begin
        image_2_236 <= io_pixelVal_in_2_2;
      end else if (10'hec == _T_19[9:0]) begin
        image_2_236 <= io_pixelVal_in_2_1;
      end else if (10'hec == _T_15[9:0]) begin
        image_2_236 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_237 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hed == _T_37[9:0]) begin
        image_2_237 <= io_pixelVal_in_2_7;
      end else if (10'hed == _T_34[9:0]) begin
        image_2_237 <= io_pixelVal_in_2_6;
      end else if (10'hed == _T_31[9:0]) begin
        image_2_237 <= io_pixelVal_in_2_5;
      end else if (10'hed == _T_28[9:0]) begin
        image_2_237 <= io_pixelVal_in_2_4;
      end else if (10'hed == _T_25[9:0]) begin
        image_2_237 <= io_pixelVal_in_2_3;
      end else if (10'hed == _T_22[9:0]) begin
        image_2_237 <= io_pixelVal_in_2_2;
      end else if (10'hed == _T_19[9:0]) begin
        image_2_237 <= io_pixelVal_in_2_1;
      end else if (10'hed == _T_15[9:0]) begin
        image_2_237 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_238 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hee == _T_37[9:0]) begin
        image_2_238 <= io_pixelVal_in_2_7;
      end else if (10'hee == _T_34[9:0]) begin
        image_2_238 <= io_pixelVal_in_2_6;
      end else if (10'hee == _T_31[9:0]) begin
        image_2_238 <= io_pixelVal_in_2_5;
      end else if (10'hee == _T_28[9:0]) begin
        image_2_238 <= io_pixelVal_in_2_4;
      end else if (10'hee == _T_25[9:0]) begin
        image_2_238 <= io_pixelVal_in_2_3;
      end else if (10'hee == _T_22[9:0]) begin
        image_2_238 <= io_pixelVal_in_2_2;
      end else if (10'hee == _T_19[9:0]) begin
        image_2_238 <= io_pixelVal_in_2_1;
      end else if (10'hee == _T_15[9:0]) begin
        image_2_238 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_239 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hef == _T_37[9:0]) begin
        image_2_239 <= io_pixelVal_in_2_7;
      end else if (10'hef == _T_34[9:0]) begin
        image_2_239 <= io_pixelVal_in_2_6;
      end else if (10'hef == _T_31[9:0]) begin
        image_2_239 <= io_pixelVal_in_2_5;
      end else if (10'hef == _T_28[9:0]) begin
        image_2_239 <= io_pixelVal_in_2_4;
      end else if (10'hef == _T_25[9:0]) begin
        image_2_239 <= io_pixelVal_in_2_3;
      end else if (10'hef == _T_22[9:0]) begin
        image_2_239 <= io_pixelVal_in_2_2;
      end else if (10'hef == _T_19[9:0]) begin
        image_2_239 <= io_pixelVal_in_2_1;
      end else if (10'hef == _T_15[9:0]) begin
        image_2_239 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_240 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf0 == _T_37[9:0]) begin
        image_2_240 <= io_pixelVal_in_2_7;
      end else if (10'hf0 == _T_34[9:0]) begin
        image_2_240 <= io_pixelVal_in_2_6;
      end else if (10'hf0 == _T_31[9:0]) begin
        image_2_240 <= io_pixelVal_in_2_5;
      end else if (10'hf0 == _T_28[9:0]) begin
        image_2_240 <= io_pixelVal_in_2_4;
      end else if (10'hf0 == _T_25[9:0]) begin
        image_2_240 <= io_pixelVal_in_2_3;
      end else if (10'hf0 == _T_22[9:0]) begin
        image_2_240 <= io_pixelVal_in_2_2;
      end else if (10'hf0 == _T_19[9:0]) begin
        image_2_240 <= io_pixelVal_in_2_1;
      end else if (10'hf0 == _T_15[9:0]) begin
        image_2_240 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_241 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf1 == _T_37[9:0]) begin
        image_2_241 <= io_pixelVal_in_2_7;
      end else if (10'hf1 == _T_34[9:0]) begin
        image_2_241 <= io_pixelVal_in_2_6;
      end else if (10'hf1 == _T_31[9:0]) begin
        image_2_241 <= io_pixelVal_in_2_5;
      end else if (10'hf1 == _T_28[9:0]) begin
        image_2_241 <= io_pixelVal_in_2_4;
      end else if (10'hf1 == _T_25[9:0]) begin
        image_2_241 <= io_pixelVal_in_2_3;
      end else if (10'hf1 == _T_22[9:0]) begin
        image_2_241 <= io_pixelVal_in_2_2;
      end else if (10'hf1 == _T_19[9:0]) begin
        image_2_241 <= io_pixelVal_in_2_1;
      end else if (10'hf1 == _T_15[9:0]) begin
        image_2_241 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_242 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf2 == _T_37[9:0]) begin
        image_2_242 <= io_pixelVal_in_2_7;
      end else if (10'hf2 == _T_34[9:0]) begin
        image_2_242 <= io_pixelVal_in_2_6;
      end else if (10'hf2 == _T_31[9:0]) begin
        image_2_242 <= io_pixelVal_in_2_5;
      end else if (10'hf2 == _T_28[9:0]) begin
        image_2_242 <= io_pixelVal_in_2_4;
      end else if (10'hf2 == _T_25[9:0]) begin
        image_2_242 <= io_pixelVal_in_2_3;
      end else if (10'hf2 == _T_22[9:0]) begin
        image_2_242 <= io_pixelVal_in_2_2;
      end else if (10'hf2 == _T_19[9:0]) begin
        image_2_242 <= io_pixelVal_in_2_1;
      end else if (10'hf2 == _T_15[9:0]) begin
        image_2_242 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_243 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf3 == _T_37[9:0]) begin
        image_2_243 <= io_pixelVal_in_2_7;
      end else if (10'hf3 == _T_34[9:0]) begin
        image_2_243 <= io_pixelVal_in_2_6;
      end else if (10'hf3 == _T_31[9:0]) begin
        image_2_243 <= io_pixelVal_in_2_5;
      end else if (10'hf3 == _T_28[9:0]) begin
        image_2_243 <= io_pixelVal_in_2_4;
      end else if (10'hf3 == _T_25[9:0]) begin
        image_2_243 <= io_pixelVal_in_2_3;
      end else if (10'hf3 == _T_22[9:0]) begin
        image_2_243 <= io_pixelVal_in_2_2;
      end else if (10'hf3 == _T_19[9:0]) begin
        image_2_243 <= io_pixelVal_in_2_1;
      end else if (10'hf3 == _T_15[9:0]) begin
        image_2_243 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_244 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf4 == _T_37[9:0]) begin
        image_2_244 <= io_pixelVal_in_2_7;
      end else if (10'hf4 == _T_34[9:0]) begin
        image_2_244 <= io_pixelVal_in_2_6;
      end else if (10'hf4 == _T_31[9:0]) begin
        image_2_244 <= io_pixelVal_in_2_5;
      end else if (10'hf4 == _T_28[9:0]) begin
        image_2_244 <= io_pixelVal_in_2_4;
      end else if (10'hf4 == _T_25[9:0]) begin
        image_2_244 <= io_pixelVal_in_2_3;
      end else if (10'hf4 == _T_22[9:0]) begin
        image_2_244 <= io_pixelVal_in_2_2;
      end else if (10'hf4 == _T_19[9:0]) begin
        image_2_244 <= io_pixelVal_in_2_1;
      end else if (10'hf4 == _T_15[9:0]) begin
        image_2_244 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_245 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf5 == _T_37[9:0]) begin
        image_2_245 <= io_pixelVal_in_2_7;
      end else if (10'hf5 == _T_34[9:0]) begin
        image_2_245 <= io_pixelVal_in_2_6;
      end else if (10'hf5 == _T_31[9:0]) begin
        image_2_245 <= io_pixelVal_in_2_5;
      end else if (10'hf5 == _T_28[9:0]) begin
        image_2_245 <= io_pixelVal_in_2_4;
      end else if (10'hf5 == _T_25[9:0]) begin
        image_2_245 <= io_pixelVal_in_2_3;
      end else if (10'hf5 == _T_22[9:0]) begin
        image_2_245 <= io_pixelVal_in_2_2;
      end else if (10'hf5 == _T_19[9:0]) begin
        image_2_245 <= io_pixelVal_in_2_1;
      end else if (10'hf5 == _T_15[9:0]) begin
        image_2_245 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_246 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf6 == _T_37[9:0]) begin
        image_2_246 <= io_pixelVal_in_2_7;
      end else if (10'hf6 == _T_34[9:0]) begin
        image_2_246 <= io_pixelVal_in_2_6;
      end else if (10'hf6 == _T_31[9:0]) begin
        image_2_246 <= io_pixelVal_in_2_5;
      end else if (10'hf6 == _T_28[9:0]) begin
        image_2_246 <= io_pixelVal_in_2_4;
      end else if (10'hf6 == _T_25[9:0]) begin
        image_2_246 <= io_pixelVal_in_2_3;
      end else if (10'hf6 == _T_22[9:0]) begin
        image_2_246 <= io_pixelVal_in_2_2;
      end else if (10'hf6 == _T_19[9:0]) begin
        image_2_246 <= io_pixelVal_in_2_1;
      end else if (10'hf6 == _T_15[9:0]) begin
        image_2_246 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_247 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf7 == _T_37[9:0]) begin
        image_2_247 <= io_pixelVal_in_2_7;
      end else if (10'hf7 == _T_34[9:0]) begin
        image_2_247 <= io_pixelVal_in_2_6;
      end else if (10'hf7 == _T_31[9:0]) begin
        image_2_247 <= io_pixelVal_in_2_5;
      end else if (10'hf7 == _T_28[9:0]) begin
        image_2_247 <= io_pixelVal_in_2_4;
      end else if (10'hf7 == _T_25[9:0]) begin
        image_2_247 <= io_pixelVal_in_2_3;
      end else if (10'hf7 == _T_22[9:0]) begin
        image_2_247 <= io_pixelVal_in_2_2;
      end else if (10'hf7 == _T_19[9:0]) begin
        image_2_247 <= io_pixelVal_in_2_1;
      end else if (10'hf7 == _T_15[9:0]) begin
        image_2_247 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_248 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf8 == _T_37[9:0]) begin
        image_2_248 <= io_pixelVal_in_2_7;
      end else if (10'hf8 == _T_34[9:0]) begin
        image_2_248 <= io_pixelVal_in_2_6;
      end else if (10'hf8 == _T_31[9:0]) begin
        image_2_248 <= io_pixelVal_in_2_5;
      end else if (10'hf8 == _T_28[9:0]) begin
        image_2_248 <= io_pixelVal_in_2_4;
      end else if (10'hf8 == _T_25[9:0]) begin
        image_2_248 <= io_pixelVal_in_2_3;
      end else if (10'hf8 == _T_22[9:0]) begin
        image_2_248 <= io_pixelVal_in_2_2;
      end else if (10'hf8 == _T_19[9:0]) begin
        image_2_248 <= io_pixelVal_in_2_1;
      end else if (10'hf8 == _T_15[9:0]) begin
        image_2_248 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_249 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hf9 == _T_37[9:0]) begin
        image_2_249 <= io_pixelVal_in_2_7;
      end else if (10'hf9 == _T_34[9:0]) begin
        image_2_249 <= io_pixelVal_in_2_6;
      end else if (10'hf9 == _T_31[9:0]) begin
        image_2_249 <= io_pixelVal_in_2_5;
      end else if (10'hf9 == _T_28[9:0]) begin
        image_2_249 <= io_pixelVal_in_2_4;
      end else if (10'hf9 == _T_25[9:0]) begin
        image_2_249 <= io_pixelVal_in_2_3;
      end else if (10'hf9 == _T_22[9:0]) begin
        image_2_249 <= io_pixelVal_in_2_2;
      end else if (10'hf9 == _T_19[9:0]) begin
        image_2_249 <= io_pixelVal_in_2_1;
      end else if (10'hf9 == _T_15[9:0]) begin
        image_2_249 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_250 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hfa == _T_37[9:0]) begin
        image_2_250 <= io_pixelVal_in_2_7;
      end else if (10'hfa == _T_34[9:0]) begin
        image_2_250 <= io_pixelVal_in_2_6;
      end else if (10'hfa == _T_31[9:0]) begin
        image_2_250 <= io_pixelVal_in_2_5;
      end else if (10'hfa == _T_28[9:0]) begin
        image_2_250 <= io_pixelVal_in_2_4;
      end else if (10'hfa == _T_25[9:0]) begin
        image_2_250 <= io_pixelVal_in_2_3;
      end else if (10'hfa == _T_22[9:0]) begin
        image_2_250 <= io_pixelVal_in_2_2;
      end else if (10'hfa == _T_19[9:0]) begin
        image_2_250 <= io_pixelVal_in_2_1;
      end else if (10'hfa == _T_15[9:0]) begin
        image_2_250 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_251 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hfb == _T_37[9:0]) begin
        image_2_251 <= io_pixelVal_in_2_7;
      end else if (10'hfb == _T_34[9:0]) begin
        image_2_251 <= io_pixelVal_in_2_6;
      end else if (10'hfb == _T_31[9:0]) begin
        image_2_251 <= io_pixelVal_in_2_5;
      end else if (10'hfb == _T_28[9:0]) begin
        image_2_251 <= io_pixelVal_in_2_4;
      end else if (10'hfb == _T_25[9:0]) begin
        image_2_251 <= io_pixelVal_in_2_3;
      end else if (10'hfb == _T_22[9:0]) begin
        image_2_251 <= io_pixelVal_in_2_2;
      end else if (10'hfb == _T_19[9:0]) begin
        image_2_251 <= io_pixelVal_in_2_1;
      end else if (10'hfb == _T_15[9:0]) begin
        image_2_251 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_252 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hfc == _T_37[9:0]) begin
        image_2_252 <= io_pixelVal_in_2_7;
      end else if (10'hfc == _T_34[9:0]) begin
        image_2_252 <= io_pixelVal_in_2_6;
      end else if (10'hfc == _T_31[9:0]) begin
        image_2_252 <= io_pixelVal_in_2_5;
      end else if (10'hfc == _T_28[9:0]) begin
        image_2_252 <= io_pixelVal_in_2_4;
      end else if (10'hfc == _T_25[9:0]) begin
        image_2_252 <= io_pixelVal_in_2_3;
      end else if (10'hfc == _T_22[9:0]) begin
        image_2_252 <= io_pixelVal_in_2_2;
      end else if (10'hfc == _T_19[9:0]) begin
        image_2_252 <= io_pixelVal_in_2_1;
      end else if (10'hfc == _T_15[9:0]) begin
        image_2_252 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_253 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hfd == _T_37[9:0]) begin
        image_2_253 <= io_pixelVal_in_2_7;
      end else if (10'hfd == _T_34[9:0]) begin
        image_2_253 <= io_pixelVal_in_2_6;
      end else if (10'hfd == _T_31[9:0]) begin
        image_2_253 <= io_pixelVal_in_2_5;
      end else if (10'hfd == _T_28[9:0]) begin
        image_2_253 <= io_pixelVal_in_2_4;
      end else if (10'hfd == _T_25[9:0]) begin
        image_2_253 <= io_pixelVal_in_2_3;
      end else if (10'hfd == _T_22[9:0]) begin
        image_2_253 <= io_pixelVal_in_2_2;
      end else if (10'hfd == _T_19[9:0]) begin
        image_2_253 <= io_pixelVal_in_2_1;
      end else if (10'hfd == _T_15[9:0]) begin
        image_2_253 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_254 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hfe == _T_37[9:0]) begin
        image_2_254 <= io_pixelVal_in_2_7;
      end else if (10'hfe == _T_34[9:0]) begin
        image_2_254 <= io_pixelVal_in_2_6;
      end else if (10'hfe == _T_31[9:0]) begin
        image_2_254 <= io_pixelVal_in_2_5;
      end else if (10'hfe == _T_28[9:0]) begin
        image_2_254 <= io_pixelVal_in_2_4;
      end else if (10'hfe == _T_25[9:0]) begin
        image_2_254 <= io_pixelVal_in_2_3;
      end else if (10'hfe == _T_22[9:0]) begin
        image_2_254 <= io_pixelVal_in_2_2;
      end else if (10'hfe == _T_19[9:0]) begin
        image_2_254 <= io_pixelVal_in_2_1;
      end else if (10'hfe == _T_15[9:0]) begin
        image_2_254 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_255 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'hff == _T_37[9:0]) begin
        image_2_255 <= io_pixelVal_in_2_7;
      end else if (10'hff == _T_34[9:0]) begin
        image_2_255 <= io_pixelVal_in_2_6;
      end else if (10'hff == _T_31[9:0]) begin
        image_2_255 <= io_pixelVal_in_2_5;
      end else if (10'hff == _T_28[9:0]) begin
        image_2_255 <= io_pixelVal_in_2_4;
      end else if (10'hff == _T_25[9:0]) begin
        image_2_255 <= io_pixelVal_in_2_3;
      end else if (10'hff == _T_22[9:0]) begin
        image_2_255 <= io_pixelVal_in_2_2;
      end else if (10'hff == _T_19[9:0]) begin
        image_2_255 <= io_pixelVal_in_2_1;
      end else if (10'hff == _T_15[9:0]) begin
        image_2_255 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_256 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h100 == _T_37[9:0]) begin
        image_2_256 <= io_pixelVal_in_2_7;
      end else if (10'h100 == _T_34[9:0]) begin
        image_2_256 <= io_pixelVal_in_2_6;
      end else if (10'h100 == _T_31[9:0]) begin
        image_2_256 <= io_pixelVal_in_2_5;
      end else if (10'h100 == _T_28[9:0]) begin
        image_2_256 <= io_pixelVal_in_2_4;
      end else if (10'h100 == _T_25[9:0]) begin
        image_2_256 <= io_pixelVal_in_2_3;
      end else if (10'h100 == _T_22[9:0]) begin
        image_2_256 <= io_pixelVal_in_2_2;
      end else if (10'h100 == _T_19[9:0]) begin
        image_2_256 <= io_pixelVal_in_2_1;
      end else if (10'h100 == _T_15[9:0]) begin
        image_2_256 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_257 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h101 == _T_37[9:0]) begin
        image_2_257 <= io_pixelVal_in_2_7;
      end else if (10'h101 == _T_34[9:0]) begin
        image_2_257 <= io_pixelVal_in_2_6;
      end else if (10'h101 == _T_31[9:0]) begin
        image_2_257 <= io_pixelVal_in_2_5;
      end else if (10'h101 == _T_28[9:0]) begin
        image_2_257 <= io_pixelVal_in_2_4;
      end else if (10'h101 == _T_25[9:0]) begin
        image_2_257 <= io_pixelVal_in_2_3;
      end else if (10'h101 == _T_22[9:0]) begin
        image_2_257 <= io_pixelVal_in_2_2;
      end else if (10'h101 == _T_19[9:0]) begin
        image_2_257 <= io_pixelVal_in_2_1;
      end else if (10'h101 == _T_15[9:0]) begin
        image_2_257 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_258 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h102 == _T_37[9:0]) begin
        image_2_258 <= io_pixelVal_in_2_7;
      end else if (10'h102 == _T_34[9:0]) begin
        image_2_258 <= io_pixelVal_in_2_6;
      end else if (10'h102 == _T_31[9:0]) begin
        image_2_258 <= io_pixelVal_in_2_5;
      end else if (10'h102 == _T_28[9:0]) begin
        image_2_258 <= io_pixelVal_in_2_4;
      end else if (10'h102 == _T_25[9:0]) begin
        image_2_258 <= io_pixelVal_in_2_3;
      end else if (10'h102 == _T_22[9:0]) begin
        image_2_258 <= io_pixelVal_in_2_2;
      end else if (10'h102 == _T_19[9:0]) begin
        image_2_258 <= io_pixelVal_in_2_1;
      end else if (10'h102 == _T_15[9:0]) begin
        image_2_258 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_259 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h103 == _T_37[9:0]) begin
        image_2_259 <= io_pixelVal_in_2_7;
      end else if (10'h103 == _T_34[9:0]) begin
        image_2_259 <= io_pixelVal_in_2_6;
      end else if (10'h103 == _T_31[9:0]) begin
        image_2_259 <= io_pixelVal_in_2_5;
      end else if (10'h103 == _T_28[9:0]) begin
        image_2_259 <= io_pixelVal_in_2_4;
      end else if (10'h103 == _T_25[9:0]) begin
        image_2_259 <= io_pixelVal_in_2_3;
      end else if (10'h103 == _T_22[9:0]) begin
        image_2_259 <= io_pixelVal_in_2_2;
      end else if (10'h103 == _T_19[9:0]) begin
        image_2_259 <= io_pixelVal_in_2_1;
      end else if (10'h103 == _T_15[9:0]) begin
        image_2_259 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_260 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h104 == _T_37[9:0]) begin
        image_2_260 <= io_pixelVal_in_2_7;
      end else if (10'h104 == _T_34[9:0]) begin
        image_2_260 <= io_pixelVal_in_2_6;
      end else if (10'h104 == _T_31[9:0]) begin
        image_2_260 <= io_pixelVal_in_2_5;
      end else if (10'h104 == _T_28[9:0]) begin
        image_2_260 <= io_pixelVal_in_2_4;
      end else if (10'h104 == _T_25[9:0]) begin
        image_2_260 <= io_pixelVal_in_2_3;
      end else if (10'h104 == _T_22[9:0]) begin
        image_2_260 <= io_pixelVal_in_2_2;
      end else if (10'h104 == _T_19[9:0]) begin
        image_2_260 <= io_pixelVal_in_2_1;
      end else if (10'h104 == _T_15[9:0]) begin
        image_2_260 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_261 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h105 == _T_37[9:0]) begin
        image_2_261 <= io_pixelVal_in_2_7;
      end else if (10'h105 == _T_34[9:0]) begin
        image_2_261 <= io_pixelVal_in_2_6;
      end else if (10'h105 == _T_31[9:0]) begin
        image_2_261 <= io_pixelVal_in_2_5;
      end else if (10'h105 == _T_28[9:0]) begin
        image_2_261 <= io_pixelVal_in_2_4;
      end else if (10'h105 == _T_25[9:0]) begin
        image_2_261 <= io_pixelVal_in_2_3;
      end else if (10'h105 == _T_22[9:0]) begin
        image_2_261 <= io_pixelVal_in_2_2;
      end else if (10'h105 == _T_19[9:0]) begin
        image_2_261 <= io_pixelVal_in_2_1;
      end else if (10'h105 == _T_15[9:0]) begin
        image_2_261 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_262 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h106 == _T_37[9:0]) begin
        image_2_262 <= io_pixelVal_in_2_7;
      end else if (10'h106 == _T_34[9:0]) begin
        image_2_262 <= io_pixelVal_in_2_6;
      end else if (10'h106 == _T_31[9:0]) begin
        image_2_262 <= io_pixelVal_in_2_5;
      end else if (10'h106 == _T_28[9:0]) begin
        image_2_262 <= io_pixelVal_in_2_4;
      end else if (10'h106 == _T_25[9:0]) begin
        image_2_262 <= io_pixelVal_in_2_3;
      end else if (10'h106 == _T_22[9:0]) begin
        image_2_262 <= io_pixelVal_in_2_2;
      end else if (10'h106 == _T_19[9:0]) begin
        image_2_262 <= io_pixelVal_in_2_1;
      end else if (10'h106 == _T_15[9:0]) begin
        image_2_262 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_263 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h107 == _T_37[9:0]) begin
        image_2_263 <= io_pixelVal_in_2_7;
      end else if (10'h107 == _T_34[9:0]) begin
        image_2_263 <= io_pixelVal_in_2_6;
      end else if (10'h107 == _T_31[9:0]) begin
        image_2_263 <= io_pixelVal_in_2_5;
      end else if (10'h107 == _T_28[9:0]) begin
        image_2_263 <= io_pixelVal_in_2_4;
      end else if (10'h107 == _T_25[9:0]) begin
        image_2_263 <= io_pixelVal_in_2_3;
      end else if (10'h107 == _T_22[9:0]) begin
        image_2_263 <= io_pixelVal_in_2_2;
      end else if (10'h107 == _T_19[9:0]) begin
        image_2_263 <= io_pixelVal_in_2_1;
      end else if (10'h107 == _T_15[9:0]) begin
        image_2_263 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_264 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h108 == _T_37[9:0]) begin
        image_2_264 <= io_pixelVal_in_2_7;
      end else if (10'h108 == _T_34[9:0]) begin
        image_2_264 <= io_pixelVal_in_2_6;
      end else if (10'h108 == _T_31[9:0]) begin
        image_2_264 <= io_pixelVal_in_2_5;
      end else if (10'h108 == _T_28[9:0]) begin
        image_2_264 <= io_pixelVal_in_2_4;
      end else if (10'h108 == _T_25[9:0]) begin
        image_2_264 <= io_pixelVal_in_2_3;
      end else if (10'h108 == _T_22[9:0]) begin
        image_2_264 <= io_pixelVal_in_2_2;
      end else if (10'h108 == _T_19[9:0]) begin
        image_2_264 <= io_pixelVal_in_2_1;
      end else if (10'h108 == _T_15[9:0]) begin
        image_2_264 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_265 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h109 == _T_37[9:0]) begin
        image_2_265 <= io_pixelVal_in_2_7;
      end else if (10'h109 == _T_34[9:0]) begin
        image_2_265 <= io_pixelVal_in_2_6;
      end else if (10'h109 == _T_31[9:0]) begin
        image_2_265 <= io_pixelVal_in_2_5;
      end else if (10'h109 == _T_28[9:0]) begin
        image_2_265 <= io_pixelVal_in_2_4;
      end else if (10'h109 == _T_25[9:0]) begin
        image_2_265 <= io_pixelVal_in_2_3;
      end else if (10'h109 == _T_22[9:0]) begin
        image_2_265 <= io_pixelVal_in_2_2;
      end else if (10'h109 == _T_19[9:0]) begin
        image_2_265 <= io_pixelVal_in_2_1;
      end else if (10'h109 == _T_15[9:0]) begin
        image_2_265 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_266 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h10a == _T_37[9:0]) begin
        image_2_266 <= io_pixelVal_in_2_7;
      end else if (10'h10a == _T_34[9:0]) begin
        image_2_266 <= io_pixelVal_in_2_6;
      end else if (10'h10a == _T_31[9:0]) begin
        image_2_266 <= io_pixelVal_in_2_5;
      end else if (10'h10a == _T_28[9:0]) begin
        image_2_266 <= io_pixelVal_in_2_4;
      end else if (10'h10a == _T_25[9:0]) begin
        image_2_266 <= io_pixelVal_in_2_3;
      end else if (10'h10a == _T_22[9:0]) begin
        image_2_266 <= io_pixelVal_in_2_2;
      end else if (10'h10a == _T_19[9:0]) begin
        image_2_266 <= io_pixelVal_in_2_1;
      end else if (10'h10a == _T_15[9:0]) begin
        image_2_266 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_267 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h10b == _T_37[9:0]) begin
        image_2_267 <= io_pixelVal_in_2_7;
      end else if (10'h10b == _T_34[9:0]) begin
        image_2_267 <= io_pixelVal_in_2_6;
      end else if (10'h10b == _T_31[9:0]) begin
        image_2_267 <= io_pixelVal_in_2_5;
      end else if (10'h10b == _T_28[9:0]) begin
        image_2_267 <= io_pixelVal_in_2_4;
      end else if (10'h10b == _T_25[9:0]) begin
        image_2_267 <= io_pixelVal_in_2_3;
      end else if (10'h10b == _T_22[9:0]) begin
        image_2_267 <= io_pixelVal_in_2_2;
      end else if (10'h10b == _T_19[9:0]) begin
        image_2_267 <= io_pixelVal_in_2_1;
      end else if (10'h10b == _T_15[9:0]) begin
        image_2_267 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_268 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h10c == _T_37[9:0]) begin
        image_2_268 <= io_pixelVal_in_2_7;
      end else if (10'h10c == _T_34[9:0]) begin
        image_2_268 <= io_pixelVal_in_2_6;
      end else if (10'h10c == _T_31[9:0]) begin
        image_2_268 <= io_pixelVal_in_2_5;
      end else if (10'h10c == _T_28[9:0]) begin
        image_2_268 <= io_pixelVal_in_2_4;
      end else if (10'h10c == _T_25[9:0]) begin
        image_2_268 <= io_pixelVal_in_2_3;
      end else if (10'h10c == _T_22[9:0]) begin
        image_2_268 <= io_pixelVal_in_2_2;
      end else if (10'h10c == _T_19[9:0]) begin
        image_2_268 <= io_pixelVal_in_2_1;
      end else if (10'h10c == _T_15[9:0]) begin
        image_2_268 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_269 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h10d == _T_37[9:0]) begin
        image_2_269 <= io_pixelVal_in_2_7;
      end else if (10'h10d == _T_34[9:0]) begin
        image_2_269 <= io_pixelVal_in_2_6;
      end else if (10'h10d == _T_31[9:0]) begin
        image_2_269 <= io_pixelVal_in_2_5;
      end else if (10'h10d == _T_28[9:0]) begin
        image_2_269 <= io_pixelVal_in_2_4;
      end else if (10'h10d == _T_25[9:0]) begin
        image_2_269 <= io_pixelVal_in_2_3;
      end else if (10'h10d == _T_22[9:0]) begin
        image_2_269 <= io_pixelVal_in_2_2;
      end else if (10'h10d == _T_19[9:0]) begin
        image_2_269 <= io_pixelVal_in_2_1;
      end else if (10'h10d == _T_15[9:0]) begin
        image_2_269 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_270 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h10e == _T_37[9:0]) begin
        image_2_270 <= io_pixelVal_in_2_7;
      end else if (10'h10e == _T_34[9:0]) begin
        image_2_270 <= io_pixelVal_in_2_6;
      end else if (10'h10e == _T_31[9:0]) begin
        image_2_270 <= io_pixelVal_in_2_5;
      end else if (10'h10e == _T_28[9:0]) begin
        image_2_270 <= io_pixelVal_in_2_4;
      end else if (10'h10e == _T_25[9:0]) begin
        image_2_270 <= io_pixelVal_in_2_3;
      end else if (10'h10e == _T_22[9:0]) begin
        image_2_270 <= io_pixelVal_in_2_2;
      end else if (10'h10e == _T_19[9:0]) begin
        image_2_270 <= io_pixelVal_in_2_1;
      end else if (10'h10e == _T_15[9:0]) begin
        image_2_270 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_271 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h10f == _T_37[9:0]) begin
        image_2_271 <= io_pixelVal_in_2_7;
      end else if (10'h10f == _T_34[9:0]) begin
        image_2_271 <= io_pixelVal_in_2_6;
      end else if (10'h10f == _T_31[9:0]) begin
        image_2_271 <= io_pixelVal_in_2_5;
      end else if (10'h10f == _T_28[9:0]) begin
        image_2_271 <= io_pixelVal_in_2_4;
      end else if (10'h10f == _T_25[9:0]) begin
        image_2_271 <= io_pixelVal_in_2_3;
      end else if (10'h10f == _T_22[9:0]) begin
        image_2_271 <= io_pixelVal_in_2_2;
      end else if (10'h10f == _T_19[9:0]) begin
        image_2_271 <= io_pixelVal_in_2_1;
      end else if (10'h10f == _T_15[9:0]) begin
        image_2_271 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_272 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h110 == _T_37[9:0]) begin
        image_2_272 <= io_pixelVal_in_2_7;
      end else if (10'h110 == _T_34[9:0]) begin
        image_2_272 <= io_pixelVal_in_2_6;
      end else if (10'h110 == _T_31[9:0]) begin
        image_2_272 <= io_pixelVal_in_2_5;
      end else if (10'h110 == _T_28[9:0]) begin
        image_2_272 <= io_pixelVal_in_2_4;
      end else if (10'h110 == _T_25[9:0]) begin
        image_2_272 <= io_pixelVal_in_2_3;
      end else if (10'h110 == _T_22[9:0]) begin
        image_2_272 <= io_pixelVal_in_2_2;
      end else if (10'h110 == _T_19[9:0]) begin
        image_2_272 <= io_pixelVal_in_2_1;
      end else if (10'h110 == _T_15[9:0]) begin
        image_2_272 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_273 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h111 == _T_37[9:0]) begin
        image_2_273 <= io_pixelVal_in_2_7;
      end else if (10'h111 == _T_34[9:0]) begin
        image_2_273 <= io_pixelVal_in_2_6;
      end else if (10'h111 == _T_31[9:0]) begin
        image_2_273 <= io_pixelVal_in_2_5;
      end else if (10'h111 == _T_28[9:0]) begin
        image_2_273 <= io_pixelVal_in_2_4;
      end else if (10'h111 == _T_25[9:0]) begin
        image_2_273 <= io_pixelVal_in_2_3;
      end else if (10'h111 == _T_22[9:0]) begin
        image_2_273 <= io_pixelVal_in_2_2;
      end else if (10'h111 == _T_19[9:0]) begin
        image_2_273 <= io_pixelVal_in_2_1;
      end else if (10'h111 == _T_15[9:0]) begin
        image_2_273 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_274 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h112 == _T_37[9:0]) begin
        image_2_274 <= io_pixelVal_in_2_7;
      end else if (10'h112 == _T_34[9:0]) begin
        image_2_274 <= io_pixelVal_in_2_6;
      end else if (10'h112 == _T_31[9:0]) begin
        image_2_274 <= io_pixelVal_in_2_5;
      end else if (10'h112 == _T_28[9:0]) begin
        image_2_274 <= io_pixelVal_in_2_4;
      end else if (10'h112 == _T_25[9:0]) begin
        image_2_274 <= io_pixelVal_in_2_3;
      end else if (10'h112 == _T_22[9:0]) begin
        image_2_274 <= io_pixelVal_in_2_2;
      end else if (10'h112 == _T_19[9:0]) begin
        image_2_274 <= io_pixelVal_in_2_1;
      end else if (10'h112 == _T_15[9:0]) begin
        image_2_274 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_275 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h113 == _T_37[9:0]) begin
        image_2_275 <= io_pixelVal_in_2_7;
      end else if (10'h113 == _T_34[9:0]) begin
        image_2_275 <= io_pixelVal_in_2_6;
      end else if (10'h113 == _T_31[9:0]) begin
        image_2_275 <= io_pixelVal_in_2_5;
      end else if (10'h113 == _T_28[9:0]) begin
        image_2_275 <= io_pixelVal_in_2_4;
      end else if (10'h113 == _T_25[9:0]) begin
        image_2_275 <= io_pixelVal_in_2_3;
      end else if (10'h113 == _T_22[9:0]) begin
        image_2_275 <= io_pixelVal_in_2_2;
      end else if (10'h113 == _T_19[9:0]) begin
        image_2_275 <= io_pixelVal_in_2_1;
      end else if (10'h113 == _T_15[9:0]) begin
        image_2_275 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_276 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h114 == _T_37[9:0]) begin
        image_2_276 <= io_pixelVal_in_2_7;
      end else if (10'h114 == _T_34[9:0]) begin
        image_2_276 <= io_pixelVal_in_2_6;
      end else if (10'h114 == _T_31[9:0]) begin
        image_2_276 <= io_pixelVal_in_2_5;
      end else if (10'h114 == _T_28[9:0]) begin
        image_2_276 <= io_pixelVal_in_2_4;
      end else if (10'h114 == _T_25[9:0]) begin
        image_2_276 <= io_pixelVal_in_2_3;
      end else if (10'h114 == _T_22[9:0]) begin
        image_2_276 <= io_pixelVal_in_2_2;
      end else if (10'h114 == _T_19[9:0]) begin
        image_2_276 <= io_pixelVal_in_2_1;
      end else if (10'h114 == _T_15[9:0]) begin
        image_2_276 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_277 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h115 == _T_37[9:0]) begin
        image_2_277 <= io_pixelVal_in_2_7;
      end else if (10'h115 == _T_34[9:0]) begin
        image_2_277 <= io_pixelVal_in_2_6;
      end else if (10'h115 == _T_31[9:0]) begin
        image_2_277 <= io_pixelVal_in_2_5;
      end else if (10'h115 == _T_28[9:0]) begin
        image_2_277 <= io_pixelVal_in_2_4;
      end else if (10'h115 == _T_25[9:0]) begin
        image_2_277 <= io_pixelVal_in_2_3;
      end else if (10'h115 == _T_22[9:0]) begin
        image_2_277 <= io_pixelVal_in_2_2;
      end else if (10'h115 == _T_19[9:0]) begin
        image_2_277 <= io_pixelVal_in_2_1;
      end else if (10'h115 == _T_15[9:0]) begin
        image_2_277 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_278 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h116 == _T_37[9:0]) begin
        image_2_278 <= io_pixelVal_in_2_7;
      end else if (10'h116 == _T_34[9:0]) begin
        image_2_278 <= io_pixelVal_in_2_6;
      end else if (10'h116 == _T_31[9:0]) begin
        image_2_278 <= io_pixelVal_in_2_5;
      end else if (10'h116 == _T_28[9:0]) begin
        image_2_278 <= io_pixelVal_in_2_4;
      end else if (10'h116 == _T_25[9:0]) begin
        image_2_278 <= io_pixelVal_in_2_3;
      end else if (10'h116 == _T_22[9:0]) begin
        image_2_278 <= io_pixelVal_in_2_2;
      end else if (10'h116 == _T_19[9:0]) begin
        image_2_278 <= io_pixelVal_in_2_1;
      end else if (10'h116 == _T_15[9:0]) begin
        image_2_278 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_279 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h117 == _T_37[9:0]) begin
        image_2_279 <= io_pixelVal_in_2_7;
      end else if (10'h117 == _T_34[9:0]) begin
        image_2_279 <= io_pixelVal_in_2_6;
      end else if (10'h117 == _T_31[9:0]) begin
        image_2_279 <= io_pixelVal_in_2_5;
      end else if (10'h117 == _T_28[9:0]) begin
        image_2_279 <= io_pixelVal_in_2_4;
      end else if (10'h117 == _T_25[9:0]) begin
        image_2_279 <= io_pixelVal_in_2_3;
      end else if (10'h117 == _T_22[9:0]) begin
        image_2_279 <= io_pixelVal_in_2_2;
      end else if (10'h117 == _T_19[9:0]) begin
        image_2_279 <= io_pixelVal_in_2_1;
      end else if (10'h117 == _T_15[9:0]) begin
        image_2_279 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_280 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h118 == _T_37[9:0]) begin
        image_2_280 <= io_pixelVal_in_2_7;
      end else if (10'h118 == _T_34[9:0]) begin
        image_2_280 <= io_pixelVal_in_2_6;
      end else if (10'h118 == _T_31[9:0]) begin
        image_2_280 <= io_pixelVal_in_2_5;
      end else if (10'h118 == _T_28[9:0]) begin
        image_2_280 <= io_pixelVal_in_2_4;
      end else if (10'h118 == _T_25[9:0]) begin
        image_2_280 <= io_pixelVal_in_2_3;
      end else if (10'h118 == _T_22[9:0]) begin
        image_2_280 <= io_pixelVal_in_2_2;
      end else if (10'h118 == _T_19[9:0]) begin
        image_2_280 <= io_pixelVal_in_2_1;
      end else if (10'h118 == _T_15[9:0]) begin
        image_2_280 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_281 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h119 == _T_37[9:0]) begin
        image_2_281 <= io_pixelVal_in_2_7;
      end else if (10'h119 == _T_34[9:0]) begin
        image_2_281 <= io_pixelVal_in_2_6;
      end else if (10'h119 == _T_31[9:0]) begin
        image_2_281 <= io_pixelVal_in_2_5;
      end else if (10'h119 == _T_28[9:0]) begin
        image_2_281 <= io_pixelVal_in_2_4;
      end else if (10'h119 == _T_25[9:0]) begin
        image_2_281 <= io_pixelVal_in_2_3;
      end else if (10'h119 == _T_22[9:0]) begin
        image_2_281 <= io_pixelVal_in_2_2;
      end else if (10'h119 == _T_19[9:0]) begin
        image_2_281 <= io_pixelVal_in_2_1;
      end else if (10'h119 == _T_15[9:0]) begin
        image_2_281 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_282 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h11a == _T_37[9:0]) begin
        image_2_282 <= io_pixelVal_in_2_7;
      end else if (10'h11a == _T_34[9:0]) begin
        image_2_282 <= io_pixelVal_in_2_6;
      end else if (10'h11a == _T_31[9:0]) begin
        image_2_282 <= io_pixelVal_in_2_5;
      end else if (10'h11a == _T_28[9:0]) begin
        image_2_282 <= io_pixelVal_in_2_4;
      end else if (10'h11a == _T_25[9:0]) begin
        image_2_282 <= io_pixelVal_in_2_3;
      end else if (10'h11a == _T_22[9:0]) begin
        image_2_282 <= io_pixelVal_in_2_2;
      end else if (10'h11a == _T_19[9:0]) begin
        image_2_282 <= io_pixelVal_in_2_1;
      end else if (10'h11a == _T_15[9:0]) begin
        image_2_282 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_283 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h11b == _T_37[9:0]) begin
        image_2_283 <= io_pixelVal_in_2_7;
      end else if (10'h11b == _T_34[9:0]) begin
        image_2_283 <= io_pixelVal_in_2_6;
      end else if (10'h11b == _T_31[9:0]) begin
        image_2_283 <= io_pixelVal_in_2_5;
      end else if (10'h11b == _T_28[9:0]) begin
        image_2_283 <= io_pixelVal_in_2_4;
      end else if (10'h11b == _T_25[9:0]) begin
        image_2_283 <= io_pixelVal_in_2_3;
      end else if (10'h11b == _T_22[9:0]) begin
        image_2_283 <= io_pixelVal_in_2_2;
      end else if (10'h11b == _T_19[9:0]) begin
        image_2_283 <= io_pixelVal_in_2_1;
      end else if (10'h11b == _T_15[9:0]) begin
        image_2_283 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_284 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h11c == _T_37[9:0]) begin
        image_2_284 <= io_pixelVal_in_2_7;
      end else if (10'h11c == _T_34[9:0]) begin
        image_2_284 <= io_pixelVal_in_2_6;
      end else if (10'h11c == _T_31[9:0]) begin
        image_2_284 <= io_pixelVal_in_2_5;
      end else if (10'h11c == _T_28[9:0]) begin
        image_2_284 <= io_pixelVal_in_2_4;
      end else if (10'h11c == _T_25[9:0]) begin
        image_2_284 <= io_pixelVal_in_2_3;
      end else if (10'h11c == _T_22[9:0]) begin
        image_2_284 <= io_pixelVal_in_2_2;
      end else if (10'h11c == _T_19[9:0]) begin
        image_2_284 <= io_pixelVal_in_2_1;
      end else if (10'h11c == _T_15[9:0]) begin
        image_2_284 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_285 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h11d == _T_37[9:0]) begin
        image_2_285 <= io_pixelVal_in_2_7;
      end else if (10'h11d == _T_34[9:0]) begin
        image_2_285 <= io_pixelVal_in_2_6;
      end else if (10'h11d == _T_31[9:0]) begin
        image_2_285 <= io_pixelVal_in_2_5;
      end else if (10'h11d == _T_28[9:0]) begin
        image_2_285 <= io_pixelVal_in_2_4;
      end else if (10'h11d == _T_25[9:0]) begin
        image_2_285 <= io_pixelVal_in_2_3;
      end else if (10'h11d == _T_22[9:0]) begin
        image_2_285 <= io_pixelVal_in_2_2;
      end else if (10'h11d == _T_19[9:0]) begin
        image_2_285 <= io_pixelVal_in_2_1;
      end else if (10'h11d == _T_15[9:0]) begin
        image_2_285 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_286 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h11e == _T_37[9:0]) begin
        image_2_286 <= io_pixelVal_in_2_7;
      end else if (10'h11e == _T_34[9:0]) begin
        image_2_286 <= io_pixelVal_in_2_6;
      end else if (10'h11e == _T_31[9:0]) begin
        image_2_286 <= io_pixelVal_in_2_5;
      end else if (10'h11e == _T_28[9:0]) begin
        image_2_286 <= io_pixelVal_in_2_4;
      end else if (10'h11e == _T_25[9:0]) begin
        image_2_286 <= io_pixelVal_in_2_3;
      end else if (10'h11e == _T_22[9:0]) begin
        image_2_286 <= io_pixelVal_in_2_2;
      end else if (10'h11e == _T_19[9:0]) begin
        image_2_286 <= io_pixelVal_in_2_1;
      end else if (10'h11e == _T_15[9:0]) begin
        image_2_286 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_287 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h11f == _T_37[9:0]) begin
        image_2_287 <= io_pixelVal_in_2_7;
      end else if (10'h11f == _T_34[9:0]) begin
        image_2_287 <= io_pixelVal_in_2_6;
      end else if (10'h11f == _T_31[9:0]) begin
        image_2_287 <= io_pixelVal_in_2_5;
      end else if (10'h11f == _T_28[9:0]) begin
        image_2_287 <= io_pixelVal_in_2_4;
      end else if (10'h11f == _T_25[9:0]) begin
        image_2_287 <= io_pixelVal_in_2_3;
      end else if (10'h11f == _T_22[9:0]) begin
        image_2_287 <= io_pixelVal_in_2_2;
      end else if (10'h11f == _T_19[9:0]) begin
        image_2_287 <= io_pixelVal_in_2_1;
      end else if (10'h11f == _T_15[9:0]) begin
        image_2_287 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_288 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h120 == _T_37[9:0]) begin
        image_2_288 <= io_pixelVal_in_2_7;
      end else if (10'h120 == _T_34[9:0]) begin
        image_2_288 <= io_pixelVal_in_2_6;
      end else if (10'h120 == _T_31[9:0]) begin
        image_2_288 <= io_pixelVal_in_2_5;
      end else if (10'h120 == _T_28[9:0]) begin
        image_2_288 <= io_pixelVal_in_2_4;
      end else if (10'h120 == _T_25[9:0]) begin
        image_2_288 <= io_pixelVal_in_2_3;
      end else if (10'h120 == _T_22[9:0]) begin
        image_2_288 <= io_pixelVal_in_2_2;
      end else if (10'h120 == _T_19[9:0]) begin
        image_2_288 <= io_pixelVal_in_2_1;
      end else if (10'h120 == _T_15[9:0]) begin
        image_2_288 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_289 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h121 == _T_37[9:0]) begin
        image_2_289 <= io_pixelVal_in_2_7;
      end else if (10'h121 == _T_34[9:0]) begin
        image_2_289 <= io_pixelVal_in_2_6;
      end else if (10'h121 == _T_31[9:0]) begin
        image_2_289 <= io_pixelVal_in_2_5;
      end else if (10'h121 == _T_28[9:0]) begin
        image_2_289 <= io_pixelVal_in_2_4;
      end else if (10'h121 == _T_25[9:0]) begin
        image_2_289 <= io_pixelVal_in_2_3;
      end else if (10'h121 == _T_22[9:0]) begin
        image_2_289 <= io_pixelVal_in_2_2;
      end else if (10'h121 == _T_19[9:0]) begin
        image_2_289 <= io_pixelVal_in_2_1;
      end else if (10'h121 == _T_15[9:0]) begin
        image_2_289 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_290 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h122 == _T_37[9:0]) begin
        image_2_290 <= io_pixelVal_in_2_7;
      end else if (10'h122 == _T_34[9:0]) begin
        image_2_290 <= io_pixelVal_in_2_6;
      end else if (10'h122 == _T_31[9:0]) begin
        image_2_290 <= io_pixelVal_in_2_5;
      end else if (10'h122 == _T_28[9:0]) begin
        image_2_290 <= io_pixelVal_in_2_4;
      end else if (10'h122 == _T_25[9:0]) begin
        image_2_290 <= io_pixelVal_in_2_3;
      end else if (10'h122 == _T_22[9:0]) begin
        image_2_290 <= io_pixelVal_in_2_2;
      end else if (10'h122 == _T_19[9:0]) begin
        image_2_290 <= io_pixelVal_in_2_1;
      end else if (10'h122 == _T_15[9:0]) begin
        image_2_290 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_291 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h123 == _T_37[9:0]) begin
        image_2_291 <= io_pixelVal_in_2_7;
      end else if (10'h123 == _T_34[9:0]) begin
        image_2_291 <= io_pixelVal_in_2_6;
      end else if (10'h123 == _T_31[9:0]) begin
        image_2_291 <= io_pixelVal_in_2_5;
      end else if (10'h123 == _T_28[9:0]) begin
        image_2_291 <= io_pixelVal_in_2_4;
      end else if (10'h123 == _T_25[9:0]) begin
        image_2_291 <= io_pixelVal_in_2_3;
      end else if (10'h123 == _T_22[9:0]) begin
        image_2_291 <= io_pixelVal_in_2_2;
      end else if (10'h123 == _T_19[9:0]) begin
        image_2_291 <= io_pixelVal_in_2_1;
      end else if (10'h123 == _T_15[9:0]) begin
        image_2_291 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_292 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h124 == _T_37[9:0]) begin
        image_2_292 <= io_pixelVal_in_2_7;
      end else if (10'h124 == _T_34[9:0]) begin
        image_2_292 <= io_pixelVal_in_2_6;
      end else if (10'h124 == _T_31[9:0]) begin
        image_2_292 <= io_pixelVal_in_2_5;
      end else if (10'h124 == _T_28[9:0]) begin
        image_2_292 <= io_pixelVal_in_2_4;
      end else if (10'h124 == _T_25[9:0]) begin
        image_2_292 <= io_pixelVal_in_2_3;
      end else if (10'h124 == _T_22[9:0]) begin
        image_2_292 <= io_pixelVal_in_2_2;
      end else if (10'h124 == _T_19[9:0]) begin
        image_2_292 <= io_pixelVal_in_2_1;
      end else if (10'h124 == _T_15[9:0]) begin
        image_2_292 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_293 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h125 == _T_37[9:0]) begin
        image_2_293 <= io_pixelVal_in_2_7;
      end else if (10'h125 == _T_34[9:0]) begin
        image_2_293 <= io_pixelVal_in_2_6;
      end else if (10'h125 == _T_31[9:0]) begin
        image_2_293 <= io_pixelVal_in_2_5;
      end else if (10'h125 == _T_28[9:0]) begin
        image_2_293 <= io_pixelVal_in_2_4;
      end else if (10'h125 == _T_25[9:0]) begin
        image_2_293 <= io_pixelVal_in_2_3;
      end else if (10'h125 == _T_22[9:0]) begin
        image_2_293 <= io_pixelVal_in_2_2;
      end else if (10'h125 == _T_19[9:0]) begin
        image_2_293 <= io_pixelVal_in_2_1;
      end else if (10'h125 == _T_15[9:0]) begin
        image_2_293 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_294 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h126 == _T_37[9:0]) begin
        image_2_294 <= io_pixelVal_in_2_7;
      end else if (10'h126 == _T_34[9:0]) begin
        image_2_294 <= io_pixelVal_in_2_6;
      end else if (10'h126 == _T_31[9:0]) begin
        image_2_294 <= io_pixelVal_in_2_5;
      end else if (10'h126 == _T_28[9:0]) begin
        image_2_294 <= io_pixelVal_in_2_4;
      end else if (10'h126 == _T_25[9:0]) begin
        image_2_294 <= io_pixelVal_in_2_3;
      end else if (10'h126 == _T_22[9:0]) begin
        image_2_294 <= io_pixelVal_in_2_2;
      end else if (10'h126 == _T_19[9:0]) begin
        image_2_294 <= io_pixelVal_in_2_1;
      end else if (10'h126 == _T_15[9:0]) begin
        image_2_294 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_295 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h127 == _T_37[9:0]) begin
        image_2_295 <= io_pixelVal_in_2_7;
      end else if (10'h127 == _T_34[9:0]) begin
        image_2_295 <= io_pixelVal_in_2_6;
      end else if (10'h127 == _T_31[9:0]) begin
        image_2_295 <= io_pixelVal_in_2_5;
      end else if (10'h127 == _T_28[9:0]) begin
        image_2_295 <= io_pixelVal_in_2_4;
      end else if (10'h127 == _T_25[9:0]) begin
        image_2_295 <= io_pixelVal_in_2_3;
      end else if (10'h127 == _T_22[9:0]) begin
        image_2_295 <= io_pixelVal_in_2_2;
      end else if (10'h127 == _T_19[9:0]) begin
        image_2_295 <= io_pixelVal_in_2_1;
      end else if (10'h127 == _T_15[9:0]) begin
        image_2_295 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_296 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h128 == _T_37[9:0]) begin
        image_2_296 <= io_pixelVal_in_2_7;
      end else if (10'h128 == _T_34[9:0]) begin
        image_2_296 <= io_pixelVal_in_2_6;
      end else if (10'h128 == _T_31[9:0]) begin
        image_2_296 <= io_pixelVal_in_2_5;
      end else if (10'h128 == _T_28[9:0]) begin
        image_2_296 <= io_pixelVal_in_2_4;
      end else if (10'h128 == _T_25[9:0]) begin
        image_2_296 <= io_pixelVal_in_2_3;
      end else if (10'h128 == _T_22[9:0]) begin
        image_2_296 <= io_pixelVal_in_2_2;
      end else if (10'h128 == _T_19[9:0]) begin
        image_2_296 <= io_pixelVal_in_2_1;
      end else if (10'h128 == _T_15[9:0]) begin
        image_2_296 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_297 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h129 == _T_37[9:0]) begin
        image_2_297 <= io_pixelVal_in_2_7;
      end else if (10'h129 == _T_34[9:0]) begin
        image_2_297 <= io_pixelVal_in_2_6;
      end else if (10'h129 == _T_31[9:0]) begin
        image_2_297 <= io_pixelVal_in_2_5;
      end else if (10'h129 == _T_28[9:0]) begin
        image_2_297 <= io_pixelVal_in_2_4;
      end else if (10'h129 == _T_25[9:0]) begin
        image_2_297 <= io_pixelVal_in_2_3;
      end else if (10'h129 == _T_22[9:0]) begin
        image_2_297 <= io_pixelVal_in_2_2;
      end else if (10'h129 == _T_19[9:0]) begin
        image_2_297 <= io_pixelVal_in_2_1;
      end else if (10'h129 == _T_15[9:0]) begin
        image_2_297 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_298 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h12a == _T_37[9:0]) begin
        image_2_298 <= io_pixelVal_in_2_7;
      end else if (10'h12a == _T_34[9:0]) begin
        image_2_298 <= io_pixelVal_in_2_6;
      end else if (10'h12a == _T_31[9:0]) begin
        image_2_298 <= io_pixelVal_in_2_5;
      end else if (10'h12a == _T_28[9:0]) begin
        image_2_298 <= io_pixelVal_in_2_4;
      end else if (10'h12a == _T_25[9:0]) begin
        image_2_298 <= io_pixelVal_in_2_3;
      end else if (10'h12a == _T_22[9:0]) begin
        image_2_298 <= io_pixelVal_in_2_2;
      end else if (10'h12a == _T_19[9:0]) begin
        image_2_298 <= io_pixelVal_in_2_1;
      end else if (10'h12a == _T_15[9:0]) begin
        image_2_298 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_299 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h12b == _T_37[9:0]) begin
        image_2_299 <= io_pixelVal_in_2_7;
      end else if (10'h12b == _T_34[9:0]) begin
        image_2_299 <= io_pixelVal_in_2_6;
      end else if (10'h12b == _T_31[9:0]) begin
        image_2_299 <= io_pixelVal_in_2_5;
      end else if (10'h12b == _T_28[9:0]) begin
        image_2_299 <= io_pixelVal_in_2_4;
      end else if (10'h12b == _T_25[9:0]) begin
        image_2_299 <= io_pixelVal_in_2_3;
      end else if (10'h12b == _T_22[9:0]) begin
        image_2_299 <= io_pixelVal_in_2_2;
      end else if (10'h12b == _T_19[9:0]) begin
        image_2_299 <= io_pixelVal_in_2_1;
      end else if (10'h12b == _T_15[9:0]) begin
        image_2_299 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_300 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h12c == _T_37[9:0]) begin
        image_2_300 <= io_pixelVal_in_2_7;
      end else if (10'h12c == _T_34[9:0]) begin
        image_2_300 <= io_pixelVal_in_2_6;
      end else if (10'h12c == _T_31[9:0]) begin
        image_2_300 <= io_pixelVal_in_2_5;
      end else if (10'h12c == _T_28[9:0]) begin
        image_2_300 <= io_pixelVal_in_2_4;
      end else if (10'h12c == _T_25[9:0]) begin
        image_2_300 <= io_pixelVal_in_2_3;
      end else if (10'h12c == _T_22[9:0]) begin
        image_2_300 <= io_pixelVal_in_2_2;
      end else if (10'h12c == _T_19[9:0]) begin
        image_2_300 <= io_pixelVal_in_2_1;
      end else if (10'h12c == _T_15[9:0]) begin
        image_2_300 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_301 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h12d == _T_37[9:0]) begin
        image_2_301 <= io_pixelVal_in_2_7;
      end else if (10'h12d == _T_34[9:0]) begin
        image_2_301 <= io_pixelVal_in_2_6;
      end else if (10'h12d == _T_31[9:0]) begin
        image_2_301 <= io_pixelVal_in_2_5;
      end else if (10'h12d == _T_28[9:0]) begin
        image_2_301 <= io_pixelVal_in_2_4;
      end else if (10'h12d == _T_25[9:0]) begin
        image_2_301 <= io_pixelVal_in_2_3;
      end else if (10'h12d == _T_22[9:0]) begin
        image_2_301 <= io_pixelVal_in_2_2;
      end else if (10'h12d == _T_19[9:0]) begin
        image_2_301 <= io_pixelVal_in_2_1;
      end else if (10'h12d == _T_15[9:0]) begin
        image_2_301 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_302 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h12e == _T_37[9:0]) begin
        image_2_302 <= io_pixelVal_in_2_7;
      end else if (10'h12e == _T_34[9:0]) begin
        image_2_302 <= io_pixelVal_in_2_6;
      end else if (10'h12e == _T_31[9:0]) begin
        image_2_302 <= io_pixelVal_in_2_5;
      end else if (10'h12e == _T_28[9:0]) begin
        image_2_302 <= io_pixelVal_in_2_4;
      end else if (10'h12e == _T_25[9:0]) begin
        image_2_302 <= io_pixelVal_in_2_3;
      end else if (10'h12e == _T_22[9:0]) begin
        image_2_302 <= io_pixelVal_in_2_2;
      end else if (10'h12e == _T_19[9:0]) begin
        image_2_302 <= io_pixelVal_in_2_1;
      end else if (10'h12e == _T_15[9:0]) begin
        image_2_302 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_303 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h12f == _T_37[9:0]) begin
        image_2_303 <= io_pixelVal_in_2_7;
      end else if (10'h12f == _T_34[9:0]) begin
        image_2_303 <= io_pixelVal_in_2_6;
      end else if (10'h12f == _T_31[9:0]) begin
        image_2_303 <= io_pixelVal_in_2_5;
      end else if (10'h12f == _T_28[9:0]) begin
        image_2_303 <= io_pixelVal_in_2_4;
      end else if (10'h12f == _T_25[9:0]) begin
        image_2_303 <= io_pixelVal_in_2_3;
      end else if (10'h12f == _T_22[9:0]) begin
        image_2_303 <= io_pixelVal_in_2_2;
      end else if (10'h12f == _T_19[9:0]) begin
        image_2_303 <= io_pixelVal_in_2_1;
      end else if (10'h12f == _T_15[9:0]) begin
        image_2_303 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_304 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h130 == _T_37[9:0]) begin
        image_2_304 <= io_pixelVal_in_2_7;
      end else if (10'h130 == _T_34[9:0]) begin
        image_2_304 <= io_pixelVal_in_2_6;
      end else if (10'h130 == _T_31[9:0]) begin
        image_2_304 <= io_pixelVal_in_2_5;
      end else if (10'h130 == _T_28[9:0]) begin
        image_2_304 <= io_pixelVal_in_2_4;
      end else if (10'h130 == _T_25[9:0]) begin
        image_2_304 <= io_pixelVal_in_2_3;
      end else if (10'h130 == _T_22[9:0]) begin
        image_2_304 <= io_pixelVal_in_2_2;
      end else if (10'h130 == _T_19[9:0]) begin
        image_2_304 <= io_pixelVal_in_2_1;
      end else if (10'h130 == _T_15[9:0]) begin
        image_2_304 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_305 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h131 == _T_37[9:0]) begin
        image_2_305 <= io_pixelVal_in_2_7;
      end else if (10'h131 == _T_34[9:0]) begin
        image_2_305 <= io_pixelVal_in_2_6;
      end else if (10'h131 == _T_31[9:0]) begin
        image_2_305 <= io_pixelVal_in_2_5;
      end else if (10'h131 == _T_28[9:0]) begin
        image_2_305 <= io_pixelVal_in_2_4;
      end else if (10'h131 == _T_25[9:0]) begin
        image_2_305 <= io_pixelVal_in_2_3;
      end else if (10'h131 == _T_22[9:0]) begin
        image_2_305 <= io_pixelVal_in_2_2;
      end else if (10'h131 == _T_19[9:0]) begin
        image_2_305 <= io_pixelVal_in_2_1;
      end else if (10'h131 == _T_15[9:0]) begin
        image_2_305 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_306 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h132 == _T_37[9:0]) begin
        image_2_306 <= io_pixelVal_in_2_7;
      end else if (10'h132 == _T_34[9:0]) begin
        image_2_306 <= io_pixelVal_in_2_6;
      end else if (10'h132 == _T_31[9:0]) begin
        image_2_306 <= io_pixelVal_in_2_5;
      end else if (10'h132 == _T_28[9:0]) begin
        image_2_306 <= io_pixelVal_in_2_4;
      end else if (10'h132 == _T_25[9:0]) begin
        image_2_306 <= io_pixelVal_in_2_3;
      end else if (10'h132 == _T_22[9:0]) begin
        image_2_306 <= io_pixelVal_in_2_2;
      end else if (10'h132 == _T_19[9:0]) begin
        image_2_306 <= io_pixelVal_in_2_1;
      end else if (10'h132 == _T_15[9:0]) begin
        image_2_306 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_307 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h133 == _T_37[9:0]) begin
        image_2_307 <= io_pixelVal_in_2_7;
      end else if (10'h133 == _T_34[9:0]) begin
        image_2_307 <= io_pixelVal_in_2_6;
      end else if (10'h133 == _T_31[9:0]) begin
        image_2_307 <= io_pixelVal_in_2_5;
      end else if (10'h133 == _T_28[9:0]) begin
        image_2_307 <= io_pixelVal_in_2_4;
      end else if (10'h133 == _T_25[9:0]) begin
        image_2_307 <= io_pixelVal_in_2_3;
      end else if (10'h133 == _T_22[9:0]) begin
        image_2_307 <= io_pixelVal_in_2_2;
      end else if (10'h133 == _T_19[9:0]) begin
        image_2_307 <= io_pixelVal_in_2_1;
      end else if (10'h133 == _T_15[9:0]) begin
        image_2_307 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_308 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h134 == _T_37[9:0]) begin
        image_2_308 <= io_pixelVal_in_2_7;
      end else if (10'h134 == _T_34[9:0]) begin
        image_2_308 <= io_pixelVal_in_2_6;
      end else if (10'h134 == _T_31[9:0]) begin
        image_2_308 <= io_pixelVal_in_2_5;
      end else if (10'h134 == _T_28[9:0]) begin
        image_2_308 <= io_pixelVal_in_2_4;
      end else if (10'h134 == _T_25[9:0]) begin
        image_2_308 <= io_pixelVal_in_2_3;
      end else if (10'h134 == _T_22[9:0]) begin
        image_2_308 <= io_pixelVal_in_2_2;
      end else if (10'h134 == _T_19[9:0]) begin
        image_2_308 <= io_pixelVal_in_2_1;
      end else if (10'h134 == _T_15[9:0]) begin
        image_2_308 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_309 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h135 == _T_37[9:0]) begin
        image_2_309 <= io_pixelVal_in_2_7;
      end else if (10'h135 == _T_34[9:0]) begin
        image_2_309 <= io_pixelVal_in_2_6;
      end else if (10'h135 == _T_31[9:0]) begin
        image_2_309 <= io_pixelVal_in_2_5;
      end else if (10'h135 == _T_28[9:0]) begin
        image_2_309 <= io_pixelVal_in_2_4;
      end else if (10'h135 == _T_25[9:0]) begin
        image_2_309 <= io_pixelVal_in_2_3;
      end else if (10'h135 == _T_22[9:0]) begin
        image_2_309 <= io_pixelVal_in_2_2;
      end else if (10'h135 == _T_19[9:0]) begin
        image_2_309 <= io_pixelVal_in_2_1;
      end else if (10'h135 == _T_15[9:0]) begin
        image_2_309 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_310 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h136 == _T_37[9:0]) begin
        image_2_310 <= io_pixelVal_in_2_7;
      end else if (10'h136 == _T_34[9:0]) begin
        image_2_310 <= io_pixelVal_in_2_6;
      end else if (10'h136 == _T_31[9:0]) begin
        image_2_310 <= io_pixelVal_in_2_5;
      end else if (10'h136 == _T_28[9:0]) begin
        image_2_310 <= io_pixelVal_in_2_4;
      end else if (10'h136 == _T_25[9:0]) begin
        image_2_310 <= io_pixelVal_in_2_3;
      end else if (10'h136 == _T_22[9:0]) begin
        image_2_310 <= io_pixelVal_in_2_2;
      end else if (10'h136 == _T_19[9:0]) begin
        image_2_310 <= io_pixelVal_in_2_1;
      end else if (10'h136 == _T_15[9:0]) begin
        image_2_310 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_311 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h137 == _T_37[9:0]) begin
        image_2_311 <= io_pixelVal_in_2_7;
      end else if (10'h137 == _T_34[9:0]) begin
        image_2_311 <= io_pixelVal_in_2_6;
      end else if (10'h137 == _T_31[9:0]) begin
        image_2_311 <= io_pixelVal_in_2_5;
      end else if (10'h137 == _T_28[9:0]) begin
        image_2_311 <= io_pixelVal_in_2_4;
      end else if (10'h137 == _T_25[9:0]) begin
        image_2_311 <= io_pixelVal_in_2_3;
      end else if (10'h137 == _T_22[9:0]) begin
        image_2_311 <= io_pixelVal_in_2_2;
      end else if (10'h137 == _T_19[9:0]) begin
        image_2_311 <= io_pixelVal_in_2_1;
      end else if (10'h137 == _T_15[9:0]) begin
        image_2_311 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_312 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h138 == _T_37[9:0]) begin
        image_2_312 <= io_pixelVal_in_2_7;
      end else if (10'h138 == _T_34[9:0]) begin
        image_2_312 <= io_pixelVal_in_2_6;
      end else if (10'h138 == _T_31[9:0]) begin
        image_2_312 <= io_pixelVal_in_2_5;
      end else if (10'h138 == _T_28[9:0]) begin
        image_2_312 <= io_pixelVal_in_2_4;
      end else if (10'h138 == _T_25[9:0]) begin
        image_2_312 <= io_pixelVal_in_2_3;
      end else if (10'h138 == _T_22[9:0]) begin
        image_2_312 <= io_pixelVal_in_2_2;
      end else if (10'h138 == _T_19[9:0]) begin
        image_2_312 <= io_pixelVal_in_2_1;
      end else if (10'h138 == _T_15[9:0]) begin
        image_2_312 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_313 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h139 == _T_37[9:0]) begin
        image_2_313 <= io_pixelVal_in_2_7;
      end else if (10'h139 == _T_34[9:0]) begin
        image_2_313 <= io_pixelVal_in_2_6;
      end else if (10'h139 == _T_31[9:0]) begin
        image_2_313 <= io_pixelVal_in_2_5;
      end else if (10'h139 == _T_28[9:0]) begin
        image_2_313 <= io_pixelVal_in_2_4;
      end else if (10'h139 == _T_25[9:0]) begin
        image_2_313 <= io_pixelVal_in_2_3;
      end else if (10'h139 == _T_22[9:0]) begin
        image_2_313 <= io_pixelVal_in_2_2;
      end else if (10'h139 == _T_19[9:0]) begin
        image_2_313 <= io_pixelVal_in_2_1;
      end else if (10'h139 == _T_15[9:0]) begin
        image_2_313 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_314 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h13a == _T_37[9:0]) begin
        image_2_314 <= io_pixelVal_in_2_7;
      end else if (10'h13a == _T_34[9:0]) begin
        image_2_314 <= io_pixelVal_in_2_6;
      end else if (10'h13a == _T_31[9:0]) begin
        image_2_314 <= io_pixelVal_in_2_5;
      end else if (10'h13a == _T_28[9:0]) begin
        image_2_314 <= io_pixelVal_in_2_4;
      end else if (10'h13a == _T_25[9:0]) begin
        image_2_314 <= io_pixelVal_in_2_3;
      end else if (10'h13a == _T_22[9:0]) begin
        image_2_314 <= io_pixelVal_in_2_2;
      end else if (10'h13a == _T_19[9:0]) begin
        image_2_314 <= io_pixelVal_in_2_1;
      end else if (10'h13a == _T_15[9:0]) begin
        image_2_314 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_315 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h13b == _T_37[9:0]) begin
        image_2_315 <= io_pixelVal_in_2_7;
      end else if (10'h13b == _T_34[9:0]) begin
        image_2_315 <= io_pixelVal_in_2_6;
      end else if (10'h13b == _T_31[9:0]) begin
        image_2_315 <= io_pixelVal_in_2_5;
      end else if (10'h13b == _T_28[9:0]) begin
        image_2_315 <= io_pixelVal_in_2_4;
      end else if (10'h13b == _T_25[9:0]) begin
        image_2_315 <= io_pixelVal_in_2_3;
      end else if (10'h13b == _T_22[9:0]) begin
        image_2_315 <= io_pixelVal_in_2_2;
      end else if (10'h13b == _T_19[9:0]) begin
        image_2_315 <= io_pixelVal_in_2_1;
      end else if (10'h13b == _T_15[9:0]) begin
        image_2_315 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_316 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h13c == _T_37[9:0]) begin
        image_2_316 <= io_pixelVal_in_2_7;
      end else if (10'h13c == _T_34[9:0]) begin
        image_2_316 <= io_pixelVal_in_2_6;
      end else if (10'h13c == _T_31[9:0]) begin
        image_2_316 <= io_pixelVal_in_2_5;
      end else if (10'h13c == _T_28[9:0]) begin
        image_2_316 <= io_pixelVal_in_2_4;
      end else if (10'h13c == _T_25[9:0]) begin
        image_2_316 <= io_pixelVal_in_2_3;
      end else if (10'h13c == _T_22[9:0]) begin
        image_2_316 <= io_pixelVal_in_2_2;
      end else if (10'h13c == _T_19[9:0]) begin
        image_2_316 <= io_pixelVal_in_2_1;
      end else if (10'h13c == _T_15[9:0]) begin
        image_2_316 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_317 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h13d == _T_37[9:0]) begin
        image_2_317 <= io_pixelVal_in_2_7;
      end else if (10'h13d == _T_34[9:0]) begin
        image_2_317 <= io_pixelVal_in_2_6;
      end else if (10'h13d == _T_31[9:0]) begin
        image_2_317 <= io_pixelVal_in_2_5;
      end else if (10'h13d == _T_28[9:0]) begin
        image_2_317 <= io_pixelVal_in_2_4;
      end else if (10'h13d == _T_25[9:0]) begin
        image_2_317 <= io_pixelVal_in_2_3;
      end else if (10'h13d == _T_22[9:0]) begin
        image_2_317 <= io_pixelVal_in_2_2;
      end else if (10'h13d == _T_19[9:0]) begin
        image_2_317 <= io_pixelVal_in_2_1;
      end else if (10'h13d == _T_15[9:0]) begin
        image_2_317 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_318 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h13e == _T_37[9:0]) begin
        image_2_318 <= io_pixelVal_in_2_7;
      end else if (10'h13e == _T_34[9:0]) begin
        image_2_318 <= io_pixelVal_in_2_6;
      end else if (10'h13e == _T_31[9:0]) begin
        image_2_318 <= io_pixelVal_in_2_5;
      end else if (10'h13e == _T_28[9:0]) begin
        image_2_318 <= io_pixelVal_in_2_4;
      end else if (10'h13e == _T_25[9:0]) begin
        image_2_318 <= io_pixelVal_in_2_3;
      end else if (10'h13e == _T_22[9:0]) begin
        image_2_318 <= io_pixelVal_in_2_2;
      end else if (10'h13e == _T_19[9:0]) begin
        image_2_318 <= io_pixelVal_in_2_1;
      end else if (10'h13e == _T_15[9:0]) begin
        image_2_318 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_319 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h13f == _T_37[9:0]) begin
        image_2_319 <= io_pixelVal_in_2_7;
      end else if (10'h13f == _T_34[9:0]) begin
        image_2_319 <= io_pixelVal_in_2_6;
      end else if (10'h13f == _T_31[9:0]) begin
        image_2_319 <= io_pixelVal_in_2_5;
      end else if (10'h13f == _T_28[9:0]) begin
        image_2_319 <= io_pixelVal_in_2_4;
      end else if (10'h13f == _T_25[9:0]) begin
        image_2_319 <= io_pixelVal_in_2_3;
      end else if (10'h13f == _T_22[9:0]) begin
        image_2_319 <= io_pixelVal_in_2_2;
      end else if (10'h13f == _T_19[9:0]) begin
        image_2_319 <= io_pixelVal_in_2_1;
      end else if (10'h13f == _T_15[9:0]) begin
        image_2_319 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_320 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h140 == _T_37[9:0]) begin
        image_2_320 <= io_pixelVal_in_2_7;
      end else if (10'h140 == _T_34[9:0]) begin
        image_2_320 <= io_pixelVal_in_2_6;
      end else if (10'h140 == _T_31[9:0]) begin
        image_2_320 <= io_pixelVal_in_2_5;
      end else if (10'h140 == _T_28[9:0]) begin
        image_2_320 <= io_pixelVal_in_2_4;
      end else if (10'h140 == _T_25[9:0]) begin
        image_2_320 <= io_pixelVal_in_2_3;
      end else if (10'h140 == _T_22[9:0]) begin
        image_2_320 <= io_pixelVal_in_2_2;
      end else if (10'h140 == _T_19[9:0]) begin
        image_2_320 <= io_pixelVal_in_2_1;
      end else if (10'h140 == _T_15[9:0]) begin
        image_2_320 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_321 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h141 == _T_37[9:0]) begin
        image_2_321 <= io_pixelVal_in_2_7;
      end else if (10'h141 == _T_34[9:0]) begin
        image_2_321 <= io_pixelVal_in_2_6;
      end else if (10'h141 == _T_31[9:0]) begin
        image_2_321 <= io_pixelVal_in_2_5;
      end else if (10'h141 == _T_28[9:0]) begin
        image_2_321 <= io_pixelVal_in_2_4;
      end else if (10'h141 == _T_25[9:0]) begin
        image_2_321 <= io_pixelVal_in_2_3;
      end else if (10'h141 == _T_22[9:0]) begin
        image_2_321 <= io_pixelVal_in_2_2;
      end else if (10'h141 == _T_19[9:0]) begin
        image_2_321 <= io_pixelVal_in_2_1;
      end else if (10'h141 == _T_15[9:0]) begin
        image_2_321 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_322 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h142 == _T_37[9:0]) begin
        image_2_322 <= io_pixelVal_in_2_7;
      end else if (10'h142 == _T_34[9:0]) begin
        image_2_322 <= io_pixelVal_in_2_6;
      end else if (10'h142 == _T_31[9:0]) begin
        image_2_322 <= io_pixelVal_in_2_5;
      end else if (10'h142 == _T_28[9:0]) begin
        image_2_322 <= io_pixelVal_in_2_4;
      end else if (10'h142 == _T_25[9:0]) begin
        image_2_322 <= io_pixelVal_in_2_3;
      end else if (10'h142 == _T_22[9:0]) begin
        image_2_322 <= io_pixelVal_in_2_2;
      end else if (10'h142 == _T_19[9:0]) begin
        image_2_322 <= io_pixelVal_in_2_1;
      end else if (10'h142 == _T_15[9:0]) begin
        image_2_322 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_323 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h143 == _T_37[9:0]) begin
        image_2_323 <= io_pixelVal_in_2_7;
      end else if (10'h143 == _T_34[9:0]) begin
        image_2_323 <= io_pixelVal_in_2_6;
      end else if (10'h143 == _T_31[9:0]) begin
        image_2_323 <= io_pixelVal_in_2_5;
      end else if (10'h143 == _T_28[9:0]) begin
        image_2_323 <= io_pixelVal_in_2_4;
      end else if (10'h143 == _T_25[9:0]) begin
        image_2_323 <= io_pixelVal_in_2_3;
      end else if (10'h143 == _T_22[9:0]) begin
        image_2_323 <= io_pixelVal_in_2_2;
      end else if (10'h143 == _T_19[9:0]) begin
        image_2_323 <= io_pixelVal_in_2_1;
      end else if (10'h143 == _T_15[9:0]) begin
        image_2_323 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_324 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h144 == _T_37[9:0]) begin
        image_2_324 <= io_pixelVal_in_2_7;
      end else if (10'h144 == _T_34[9:0]) begin
        image_2_324 <= io_pixelVal_in_2_6;
      end else if (10'h144 == _T_31[9:0]) begin
        image_2_324 <= io_pixelVal_in_2_5;
      end else if (10'h144 == _T_28[9:0]) begin
        image_2_324 <= io_pixelVal_in_2_4;
      end else if (10'h144 == _T_25[9:0]) begin
        image_2_324 <= io_pixelVal_in_2_3;
      end else if (10'h144 == _T_22[9:0]) begin
        image_2_324 <= io_pixelVal_in_2_2;
      end else if (10'h144 == _T_19[9:0]) begin
        image_2_324 <= io_pixelVal_in_2_1;
      end else if (10'h144 == _T_15[9:0]) begin
        image_2_324 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_325 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h145 == _T_37[9:0]) begin
        image_2_325 <= io_pixelVal_in_2_7;
      end else if (10'h145 == _T_34[9:0]) begin
        image_2_325 <= io_pixelVal_in_2_6;
      end else if (10'h145 == _T_31[9:0]) begin
        image_2_325 <= io_pixelVal_in_2_5;
      end else if (10'h145 == _T_28[9:0]) begin
        image_2_325 <= io_pixelVal_in_2_4;
      end else if (10'h145 == _T_25[9:0]) begin
        image_2_325 <= io_pixelVal_in_2_3;
      end else if (10'h145 == _T_22[9:0]) begin
        image_2_325 <= io_pixelVal_in_2_2;
      end else if (10'h145 == _T_19[9:0]) begin
        image_2_325 <= io_pixelVal_in_2_1;
      end else if (10'h145 == _T_15[9:0]) begin
        image_2_325 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_326 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h146 == _T_37[9:0]) begin
        image_2_326 <= io_pixelVal_in_2_7;
      end else if (10'h146 == _T_34[9:0]) begin
        image_2_326 <= io_pixelVal_in_2_6;
      end else if (10'h146 == _T_31[9:0]) begin
        image_2_326 <= io_pixelVal_in_2_5;
      end else if (10'h146 == _T_28[9:0]) begin
        image_2_326 <= io_pixelVal_in_2_4;
      end else if (10'h146 == _T_25[9:0]) begin
        image_2_326 <= io_pixelVal_in_2_3;
      end else if (10'h146 == _T_22[9:0]) begin
        image_2_326 <= io_pixelVal_in_2_2;
      end else if (10'h146 == _T_19[9:0]) begin
        image_2_326 <= io_pixelVal_in_2_1;
      end else if (10'h146 == _T_15[9:0]) begin
        image_2_326 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_327 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h147 == _T_37[9:0]) begin
        image_2_327 <= io_pixelVal_in_2_7;
      end else if (10'h147 == _T_34[9:0]) begin
        image_2_327 <= io_pixelVal_in_2_6;
      end else if (10'h147 == _T_31[9:0]) begin
        image_2_327 <= io_pixelVal_in_2_5;
      end else if (10'h147 == _T_28[9:0]) begin
        image_2_327 <= io_pixelVal_in_2_4;
      end else if (10'h147 == _T_25[9:0]) begin
        image_2_327 <= io_pixelVal_in_2_3;
      end else if (10'h147 == _T_22[9:0]) begin
        image_2_327 <= io_pixelVal_in_2_2;
      end else if (10'h147 == _T_19[9:0]) begin
        image_2_327 <= io_pixelVal_in_2_1;
      end else if (10'h147 == _T_15[9:0]) begin
        image_2_327 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_328 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h148 == _T_37[9:0]) begin
        image_2_328 <= io_pixelVal_in_2_7;
      end else if (10'h148 == _T_34[9:0]) begin
        image_2_328 <= io_pixelVal_in_2_6;
      end else if (10'h148 == _T_31[9:0]) begin
        image_2_328 <= io_pixelVal_in_2_5;
      end else if (10'h148 == _T_28[9:0]) begin
        image_2_328 <= io_pixelVal_in_2_4;
      end else if (10'h148 == _T_25[9:0]) begin
        image_2_328 <= io_pixelVal_in_2_3;
      end else if (10'h148 == _T_22[9:0]) begin
        image_2_328 <= io_pixelVal_in_2_2;
      end else if (10'h148 == _T_19[9:0]) begin
        image_2_328 <= io_pixelVal_in_2_1;
      end else if (10'h148 == _T_15[9:0]) begin
        image_2_328 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_329 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h149 == _T_37[9:0]) begin
        image_2_329 <= io_pixelVal_in_2_7;
      end else if (10'h149 == _T_34[9:0]) begin
        image_2_329 <= io_pixelVal_in_2_6;
      end else if (10'h149 == _T_31[9:0]) begin
        image_2_329 <= io_pixelVal_in_2_5;
      end else if (10'h149 == _T_28[9:0]) begin
        image_2_329 <= io_pixelVal_in_2_4;
      end else if (10'h149 == _T_25[9:0]) begin
        image_2_329 <= io_pixelVal_in_2_3;
      end else if (10'h149 == _T_22[9:0]) begin
        image_2_329 <= io_pixelVal_in_2_2;
      end else if (10'h149 == _T_19[9:0]) begin
        image_2_329 <= io_pixelVal_in_2_1;
      end else if (10'h149 == _T_15[9:0]) begin
        image_2_329 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_330 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h14a == _T_37[9:0]) begin
        image_2_330 <= io_pixelVal_in_2_7;
      end else if (10'h14a == _T_34[9:0]) begin
        image_2_330 <= io_pixelVal_in_2_6;
      end else if (10'h14a == _T_31[9:0]) begin
        image_2_330 <= io_pixelVal_in_2_5;
      end else if (10'h14a == _T_28[9:0]) begin
        image_2_330 <= io_pixelVal_in_2_4;
      end else if (10'h14a == _T_25[9:0]) begin
        image_2_330 <= io_pixelVal_in_2_3;
      end else if (10'h14a == _T_22[9:0]) begin
        image_2_330 <= io_pixelVal_in_2_2;
      end else if (10'h14a == _T_19[9:0]) begin
        image_2_330 <= io_pixelVal_in_2_1;
      end else if (10'h14a == _T_15[9:0]) begin
        image_2_330 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_331 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h14b == _T_37[9:0]) begin
        image_2_331 <= io_pixelVal_in_2_7;
      end else if (10'h14b == _T_34[9:0]) begin
        image_2_331 <= io_pixelVal_in_2_6;
      end else if (10'h14b == _T_31[9:0]) begin
        image_2_331 <= io_pixelVal_in_2_5;
      end else if (10'h14b == _T_28[9:0]) begin
        image_2_331 <= io_pixelVal_in_2_4;
      end else if (10'h14b == _T_25[9:0]) begin
        image_2_331 <= io_pixelVal_in_2_3;
      end else if (10'h14b == _T_22[9:0]) begin
        image_2_331 <= io_pixelVal_in_2_2;
      end else if (10'h14b == _T_19[9:0]) begin
        image_2_331 <= io_pixelVal_in_2_1;
      end else if (10'h14b == _T_15[9:0]) begin
        image_2_331 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_332 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h14c == _T_37[9:0]) begin
        image_2_332 <= io_pixelVal_in_2_7;
      end else if (10'h14c == _T_34[9:0]) begin
        image_2_332 <= io_pixelVal_in_2_6;
      end else if (10'h14c == _T_31[9:0]) begin
        image_2_332 <= io_pixelVal_in_2_5;
      end else if (10'h14c == _T_28[9:0]) begin
        image_2_332 <= io_pixelVal_in_2_4;
      end else if (10'h14c == _T_25[9:0]) begin
        image_2_332 <= io_pixelVal_in_2_3;
      end else if (10'h14c == _T_22[9:0]) begin
        image_2_332 <= io_pixelVal_in_2_2;
      end else if (10'h14c == _T_19[9:0]) begin
        image_2_332 <= io_pixelVal_in_2_1;
      end else if (10'h14c == _T_15[9:0]) begin
        image_2_332 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_333 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h14d == _T_37[9:0]) begin
        image_2_333 <= io_pixelVal_in_2_7;
      end else if (10'h14d == _T_34[9:0]) begin
        image_2_333 <= io_pixelVal_in_2_6;
      end else if (10'h14d == _T_31[9:0]) begin
        image_2_333 <= io_pixelVal_in_2_5;
      end else if (10'h14d == _T_28[9:0]) begin
        image_2_333 <= io_pixelVal_in_2_4;
      end else if (10'h14d == _T_25[9:0]) begin
        image_2_333 <= io_pixelVal_in_2_3;
      end else if (10'h14d == _T_22[9:0]) begin
        image_2_333 <= io_pixelVal_in_2_2;
      end else if (10'h14d == _T_19[9:0]) begin
        image_2_333 <= io_pixelVal_in_2_1;
      end else if (10'h14d == _T_15[9:0]) begin
        image_2_333 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_334 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h14e == _T_37[9:0]) begin
        image_2_334 <= io_pixelVal_in_2_7;
      end else if (10'h14e == _T_34[9:0]) begin
        image_2_334 <= io_pixelVal_in_2_6;
      end else if (10'h14e == _T_31[9:0]) begin
        image_2_334 <= io_pixelVal_in_2_5;
      end else if (10'h14e == _T_28[9:0]) begin
        image_2_334 <= io_pixelVal_in_2_4;
      end else if (10'h14e == _T_25[9:0]) begin
        image_2_334 <= io_pixelVal_in_2_3;
      end else if (10'h14e == _T_22[9:0]) begin
        image_2_334 <= io_pixelVal_in_2_2;
      end else if (10'h14e == _T_19[9:0]) begin
        image_2_334 <= io_pixelVal_in_2_1;
      end else if (10'h14e == _T_15[9:0]) begin
        image_2_334 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_335 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h14f == _T_37[9:0]) begin
        image_2_335 <= io_pixelVal_in_2_7;
      end else if (10'h14f == _T_34[9:0]) begin
        image_2_335 <= io_pixelVal_in_2_6;
      end else if (10'h14f == _T_31[9:0]) begin
        image_2_335 <= io_pixelVal_in_2_5;
      end else if (10'h14f == _T_28[9:0]) begin
        image_2_335 <= io_pixelVal_in_2_4;
      end else if (10'h14f == _T_25[9:0]) begin
        image_2_335 <= io_pixelVal_in_2_3;
      end else if (10'h14f == _T_22[9:0]) begin
        image_2_335 <= io_pixelVal_in_2_2;
      end else if (10'h14f == _T_19[9:0]) begin
        image_2_335 <= io_pixelVal_in_2_1;
      end else if (10'h14f == _T_15[9:0]) begin
        image_2_335 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_336 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h150 == _T_37[9:0]) begin
        image_2_336 <= io_pixelVal_in_2_7;
      end else if (10'h150 == _T_34[9:0]) begin
        image_2_336 <= io_pixelVal_in_2_6;
      end else if (10'h150 == _T_31[9:0]) begin
        image_2_336 <= io_pixelVal_in_2_5;
      end else if (10'h150 == _T_28[9:0]) begin
        image_2_336 <= io_pixelVal_in_2_4;
      end else if (10'h150 == _T_25[9:0]) begin
        image_2_336 <= io_pixelVal_in_2_3;
      end else if (10'h150 == _T_22[9:0]) begin
        image_2_336 <= io_pixelVal_in_2_2;
      end else if (10'h150 == _T_19[9:0]) begin
        image_2_336 <= io_pixelVal_in_2_1;
      end else if (10'h150 == _T_15[9:0]) begin
        image_2_336 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_337 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h151 == _T_37[9:0]) begin
        image_2_337 <= io_pixelVal_in_2_7;
      end else if (10'h151 == _T_34[9:0]) begin
        image_2_337 <= io_pixelVal_in_2_6;
      end else if (10'h151 == _T_31[9:0]) begin
        image_2_337 <= io_pixelVal_in_2_5;
      end else if (10'h151 == _T_28[9:0]) begin
        image_2_337 <= io_pixelVal_in_2_4;
      end else if (10'h151 == _T_25[9:0]) begin
        image_2_337 <= io_pixelVal_in_2_3;
      end else if (10'h151 == _T_22[9:0]) begin
        image_2_337 <= io_pixelVal_in_2_2;
      end else if (10'h151 == _T_19[9:0]) begin
        image_2_337 <= io_pixelVal_in_2_1;
      end else if (10'h151 == _T_15[9:0]) begin
        image_2_337 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_338 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h152 == _T_37[9:0]) begin
        image_2_338 <= io_pixelVal_in_2_7;
      end else if (10'h152 == _T_34[9:0]) begin
        image_2_338 <= io_pixelVal_in_2_6;
      end else if (10'h152 == _T_31[9:0]) begin
        image_2_338 <= io_pixelVal_in_2_5;
      end else if (10'h152 == _T_28[9:0]) begin
        image_2_338 <= io_pixelVal_in_2_4;
      end else if (10'h152 == _T_25[9:0]) begin
        image_2_338 <= io_pixelVal_in_2_3;
      end else if (10'h152 == _T_22[9:0]) begin
        image_2_338 <= io_pixelVal_in_2_2;
      end else if (10'h152 == _T_19[9:0]) begin
        image_2_338 <= io_pixelVal_in_2_1;
      end else if (10'h152 == _T_15[9:0]) begin
        image_2_338 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_339 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h153 == _T_37[9:0]) begin
        image_2_339 <= io_pixelVal_in_2_7;
      end else if (10'h153 == _T_34[9:0]) begin
        image_2_339 <= io_pixelVal_in_2_6;
      end else if (10'h153 == _T_31[9:0]) begin
        image_2_339 <= io_pixelVal_in_2_5;
      end else if (10'h153 == _T_28[9:0]) begin
        image_2_339 <= io_pixelVal_in_2_4;
      end else if (10'h153 == _T_25[9:0]) begin
        image_2_339 <= io_pixelVal_in_2_3;
      end else if (10'h153 == _T_22[9:0]) begin
        image_2_339 <= io_pixelVal_in_2_2;
      end else if (10'h153 == _T_19[9:0]) begin
        image_2_339 <= io_pixelVal_in_2_1;
      end else if (10'h153 == _T_15[9:0]) begin
        image_2_339 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_340 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h154 == _T_37[9:0]) begin
        image_2_340 <= io_pixelVal_in_2_7;
      end else if (10'h154 == _T_34[9:0]) begin
        image_2_340 <= io_pixelVal_in_2_6;
      end else if (10'h154 == _T_31[9:0]) begin
        image_2_340 <= io_pixelVal_in_2_5;
      end else if (10'h154 == _T_28[9:0]) begin
        image_2_340 <= io_pixelVal_in_2_4;
      end else if (10'h154 == _T_25[9:0]) begin
        image_2_340 <= io_pixelVal_in_2_3;
      end else if (10'h154 == _T_22[9:0]) begin
        image_2_340 <= io_pixelVal_in_2_2;
      end else if (10'h154 == _T_19[9:0]) begin
        image_2_340 <= io_pixelVal_in_2_1;
      end else if (10'h154 == _T_15[9:0]) begin
        image_2_340 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_341 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h155 == _T_37[9:0]) begin
        image_2_341 <= io_pixelVal_in_2_7;
      end else if (10'h155 == _T_34[9:0]) begin
        image_2_341 <= io_pixelVal_in_2_6;
      end else if (10'h155 == _T_31[9:0]) begin
        image_2_341 <= io_pixelVal_in_2_5;
      end else if (10'h155 == _T_28[9:0]) begin
        image_2_341 <= io_pixelVal_in_2_4;
      end else if (10'h155 == _T_25[9:0]) begin
        image_2_341 <= io_pixelVal_in_2_3;
      end else if (10'h155 == _T_22[9:0]) begin
        image_2_341 <= io_pixelVal_in_2_2;
      end else if (10'h155 == _T_19[9:0]) begin
        image_2_341 <= io_pixelVal_in_2_1;
      end else if (10'h155 == _T_15[9:0]) begin
        image_2_341 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_342 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h156 == _T_37[9:0]) begin
        image_2_342 <= io_pixelVal_in_2_7;
      end else if (10'h156 == _T_34[9:0]) begin
        image_2_342 <= io_pixelVal_in_2_6;
      end else if (10'h156 == _T_31[9:0]) begin
        image_2_342 <= io_pixelVal_in_2_5;
      end else if (10'h156 == _T_28[9:0]) begin
        image_2_342 <= io_pixelVal_in_2_4;
      end else if (10'h156 == _T_25[9:0]) begin
        image_2_342 <= io_pixelVal_in_2_3;
      end else if (10'h156 == _T_22[9:0]) begin
        image_2_342 <= io_pixelVal_in_2_2;
      end else if (10'h156 == _T_19[9:0]) begin
        image_2_342 <= io_pixelVal_in_2_1;
      end else if (10'h156 == _T_15[9:0]) begin
        image_2_342 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_343 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h157 == _T_37[9:0]) begin
        image_2_343 <= io_pixelVal_in_2_7;
      end else if (10'h157 == _T_34[9:0]) begin
        image_2_343 <= io_pixelVal_in_2_6;
      end else if (10'h157 == _T_31[9:0]) begin
        image_2_343 <= io_pixelVal_in_2_5;
      end else if (10'h157 == _T_28[9:0]) begin
        image_2_343 <= io_pixelVal_in_2_4;
      end else if (10'h157 == _T_25[9:0]) begin
        image_2_343 <= io_pixelVal_in_2_3;
      end else if (10'h157 == _T_22[9:0]) begin
        image_2_343 <= io_pixelVal_in_2_2;
      end else if (10'h157 == _T_19[9:0]) begin
        image_2_343 <= io_pixelVal_in_2_1;
      end else if (10'h157 == _T_15[9:0]) begin
        image_2_343 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_344 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h158 == _T_37[9:0]) begin
        image_2_344 <= io_pixelVal_in_2_7;
      end else if (10'h158 == _T_34[9:0]) begin
        image_2_344 <= io_pixelVal_in_2_6;
      end else if (10'h158 == _T_31[9:0]) begin
        image_2_344 <= io_pixelVal_in_2_5;
      end else if (10'h158 == _T_28[9:0]) begin
        image_2_344 <= io_pixelVal_in_2_4;
      end else if (10'h158 == _T_25[9:0]) begin
        image_2_344 <= io_pixelVal_in_2_3;
      end else if (10'h158 == _T_22[9:0]) begin
        image_2_344 <= io_pixelVal_in_2_2;
      end else if (10'h158 == _T_19[9:0]) begin
        image_2_344 <= io_pixelVal_in_2_1;
      end else if (10'h158 == _T_15[9:0]) begin
        image_2_344 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_345 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h159 == _T_37[9:0]) begin
        image_2_345 <= io_pixelVal_in_2_7;
      end else if (10'h159 == _T_34[9:0]) begin
        image_2_345 <= io_pixelVal_in_2_6;
      end else if (10'h159 == _T_31[9:0]) begin
        image_2_345 <= io_pixelVal_in_2_5;
      end else if (10'h159 == _T_28[9:0]) begin
        image_2_345 <= io_pixelVal_in_2_4;
      end else if (10'h159 == _T_25[9:0]) begin
        image_2_345 <= io_pixelVal_in_2_3;
      end else if (10'h159 == _T_22[9:0]) begin
        image_2_345 <= io_pixelVal_in_2_2;
      end else if (10'h159 == _T_19[9:0]) begin
        image_2_345 <= io_pixelVal_in_2_1;
      end else if (10'h159 == _T_15[9:0]) begin
        image_2_345 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_346 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h15a == _T_37[9:0]) begin
        image_2_346 <= io_pixelVal_in_2_7;
      end else if (10'h15a == _T_34[9:0]) begin
        image_2_346 <= io_pixelVal_in_2_6;
      end else if (10'h15a == _T_31[9:0]) begin
        image_2_346 <= io_pixelVal_in_2_5;
      end else if (10'h15a == _T_28[9:0]) begin
        image_2_346 <= io_pixelVal_in_2_4;
      end else if (10'h15a == _T_25[9:0]) begin
        image_2_346 <= io_pixelVal_in_2_3;
      end else if (10'h15a == _T_22[9:0]) begin
        image_2_346 <= io_pixelVal_in_2_2;
      end else if (10'h15a == _T_19[9:0]) begin
        image_2_346 <= io_pixelVal_in_2_1;
      end else if (10'h15a == _T_15[9:0]) begin
        image_2_346 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_347 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h15b == _T_37[9:0]) begin
        image_2_347 <= io_pixelVal_in_2_7;
      end else if (10'h15b == _T_34[9:0]) begin
        image_2_347 <= io_pixelVal_in_2_6;
      end else if (10'h15b == _T_31[9:0]) begin
        image_2_347 <= io_pixelVal_in_2_5;
      end else if (10'h15b == _T_28[9:0]) begin
        image_2_347 <= io_pixelVal_in_2_4;
      end else if (10'h15b == _T_25[9:0]) begin
        image_2_347 <= io_pixelVal_in_2_3;
      end else if (10'h15b == _T_22[9:0]) begin
        image_2_347 <= io_pixelVal_in_2_2;
      end else if (10'h15b == _T_19[9:0]) begin
        image_2_347 <= io_pixelVal_in_2_1;
      end else if (10'h15b == _T_15[9:0]) begin
        image_2_347 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_348 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h15c == _T_37[9:0]) begin
        image_2_348 <= io_pixelVal_in_2_7;
      end else if (10'h15c == _T_34[9:0]) begin
        image_2_348 <= io_pixelVal_in_2_6;
      end else if (10'h15c == _T_31[9:0]) begin
        image_2_348 <= io_pixelVal_in_2_5;
      end else if (10'h15c == _T_28[9:0]) begin
        image_2_348 <= io_pixelVal_in_2_4;
      end else if (10'h15c == _T_25[9:0]) begin
        image_2_348 <= io_pixelVal_in_2_3;
      end else if (10'h15c == _T_22[9:0]) begin
        image_2_348 <= io_pixelVal_in_2_2;
      end else if (10'h15c == _T_19[9:0]) begin
        image_2_348 <= io_pixelVal_in_2_1;
      end else if (10'h15c == _T_15[9:0]) begin
        image_2_348 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_349 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h15d == _T_37[9:0]) begin
        image_2_349 <= io_pixelVal_in_2_7;
      end else if (10'h15d == _T_34[9:0]) begin
        image_2_349 <= io_pixelVal_in_2_6;
      end else if (10'h15d == _T_31[9:0]) begin
        image_2_349 <= io_pixelVal_in_2_5;
      end else if (10'h15d == _T_28[9:0]) begin
        image_2_349 <= io_pixelVal_in_2_4;
      end else if (10'h15d == _T_25[9:0]) begin
        image_2_349 <= io_pixelVal_in_2_3;
      end else if (10'h15d == _T_22[9:0]) begin
        image_2_349 <= io_pixelVal_in_2_2;
      end else if (10'h15d == _T_19[9:0]) begin
        image_2_349 <= io_pixelVal_in_2_1;
      end else if (10'h15d == _T_15[9:0]) begin
        image_2_349 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_350 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h15e == _T_37[9:0]) begin
        image_2_350 <= io_pixelVal_in_2_7;
      end else if (10'h15e == _T_34[9:0]) begin
        image_2_350 <= io_pixelVal_in_2_6;
      end else if (10'h15e == _T_31[9:0]) begin
        image_2_350 <= io_pixelVal_in_2_5;
      end else if (10'h15e == _T_28[9:0]) begin
        image_2_350 <= io_pixelVal_in_2_4;
      end else if (10'h15e == _T_25[9:0]) begin
        image_2_350 <= io_pixelVal_in_2_3;
      end else if (10'h15e == _T_22[9:0]) begin
        image_2_350 <= io_pixelVal_in_2_2;
      end else if (10'h15e == _T_19[9:0]) begin
        image_2_350 <= io_pixelVal_in_2_1;
      end else if (10'h15e == _T_15[9:0]) begin
        image_2_350 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_351 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h15f == _T_37[9:0]) begin
        image_2_351 <= io_pixelVal_in_2_7;
      end else if (10'h15f == _T_34[9:0]) begin
        image_2_351 <= io_pixelVal_in_2_6;
      end else if (10'h15f == _T_31[9:0]) begin
        image_2_351 <= io_pixelVal_in_2_5;
      end else if (10'h15f == _T_28[9:0]) begin
        image_2_351 <= io_pixelVal_in_2_4;
      end else if (10'h15f == _T_25[9:0]) begin
        image_2_351 <= io_pixelVal_in_2_3;
      end else if (10'h15f == _T_22[9:0]) begin
        image_2_351 <= io_pixelVal_in_2_2;
      end else if (10'h15f == _T_19[9:0]) begin
        image_2_351 <= io_pixelVal_in_2_1;
      end else if (10'h15f == _T_15[9:0]) begin
        image_2_351 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_352 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h160 == _T_37[9:0]) begin
        image_2_352 <= io_pixelVal_in_2_7;
      end else if (10'h160 == _T_34[9:0]) begin
        image_2_352 <= io_pixelVal_in_2_6;
      end else if (10'h160 == _T_31[9:0]) begin
        image_2_352 <= io_pixelVal_in_2_5;
      end else if (10'h160 == _T_28[9:0]) begin
        image_2_352 <= io_pixelVal_in_2_4;
      end else if (10'h160 == _T_25[9:0]) begin
        image_2_352 <= io_pixelVal_in_2_3;
      end else if (10'h160 == _T_22[9:0]) begin
        image_2_352 <= io_pixelVal_in_2_2;
      end else if (10'h160 == _T_19[9:0]) begin
        image_2_352 <= io_pixelVal_in_2_1;
      end else if (10'h160 == _T_15[9:0]) begin
        image_2_352 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_353 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h161 == _T_37[9:0]) begin
        image_2_353 <= io_pixelVal_in_2_7;
      end else if (10'h161 == _T_34[9:0]) begin
        image_2_353 <= io_pixelVal_in_2_6;
      end else if (10'h161 == _T_31[9:0]) begin
        image_2_353 <= io_pixelVal_in_2_5;
      end else if (10'h161 == _T_28[9:0]) begin
        image_2_353 <= io_pixelVal_in_2_4;
      end else if (10'h161 == _T_25[9:0]) begin
        image_2_353 <= io_pixelVal_in_2_3;
      end else if (10'h161 == _T_22[9:0]) begin
        image_2_353 <= io_pixelVal_in_2_2;
      end else if (10'h161 == _T_19[9:0]) begin
        image_2_353 <= io_pixelVal_in_2_1;
      end else if (10'h161 == _T_15[9:0]) begin
        image_2_353 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_354 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h162 == _T_37[9:0]) begin
        image_2_354 <= io_pixelVal_in_2_7;
      end else if (10'h162 == _T_34[9:0]) begin
        image_2_354 <= io_pixelVal_in_2_6;
      end else if (10'h162 == _T_31[9:0]) begin
        image_2_354 <= io_pixelVal_in_2_5;
      end else if (10'h162 == _T_28[9:0]) begin
        image_2_354 <= io_pixelVal_in_2_4;
      end else if (10'h162 == _T_25[9:0]) begin
        image_2_354 <= io_pixelVal_in_2_3;
      end else if (10'h162 == _T_22[9:0]) begin
        image_2_354 <= io_pixelVal_in_2_2;
      end else if (10'h162 == _T_19[9:0]) begin
        image_2_354 <= io_pixelVal_in_2_1;
      end else if (10'h162 == _T_15[9:0]) begin
        image_2_354 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_355 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h163 == _T_37[9:0]) begin
        image_2_355 <= io_pixelVal_in_2_7;
      end else if (10'h163 == _T_34[9:0]) begin
        image_2_355 <= io_pixelVal_in_2_6;
      end else if (10'h163 == _T_31[9:0]) begin
        image_2_355 <= io_pixelVal_in_2_5;
      end else if (10'h163 == _T_28[9:0]) begin
        image_2_355 <= io_pixelVal_in_2_4;
      end else if (10'h163 == _T_25[9:0]) begin
        image_2_355 <= io_pixelVal_in_2_3;
      end else if (10'h163 == _T_22[9:0]) begin
        image_2_355 <= io_pixelVal_in_2_2;
      end else if (10'h163 == _T_19[9:0]) begin
        image_2_355 <= io_pixelVal_in_2_1;
      end else if (10'h163 == _T_15[9:0]) begin
        image_2_355 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_356 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h164 == _T_37[9:0]) begin
        image_2_356 <= io_pixelVal_in_2_7;
      end else if (10'h164 == _T_34[9:0]) begin
        image_2_356 <= io_pixelVal_in_2_6;
      end else if (10'h164 == _T_31[9:0]) begin
        image_2_356 <= io_pixelVal_in_2_5;
      end else if (10'h164 == _T_28[9:0]) begin
        image_2_356 <= io_pixelVal_in_2_4;
      end else if (10'h164 == _T_25[9:0]) begin
        image_2_356 <= io_pixelVal_in_2_3;
      end else if (10'h164 == _T_22[9:0]) begin
        image_2_356 <= io_pixelVal_in_2_2;
      end else if (10'h164 == _T_19[9:0]) begin
        image_2_356 <= io_pixelVal_in_2_1;
      end else if (10'h164 == _T_15[9:0]) begin
        image_2_356 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_357 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h165 == _T_37[9:0]) begin
        image_2_357 <= io_pixelVal_in_2_7;
      end else if (10'h165 == _T_34[9:0]) begin
        image_2_357 <= io_pixelVal_in_2_6;
      end else if (10'h165 == _T_31[9:0]) begin
        image_2_357 <= io_pixelVal_in_2_5;
      end else if (10'h165 == _T_28[9:0]) begin
        image_2_357 <= io_pixelVal_in_2_4;
      end else if (10'h165 == _T_25[9:0]) begin
        image_2_357 <= io_pixelVal_in_2_3;
      end else if (10'h165 == _T_22[9:0]) begin
        image_2_357 <= io_pixelVal_in_2_2;
      end else if (10'h165 == _T_19[9:0]) begin
        image_2_357 <= io_pixelVal_in_2_1;
      end else if (10'h165 == _T_15[9:0]) begin
        image_2_357 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_358 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h166 == _T_37[9:0]) begin
        image_2_358 <= io_pixelVal_in_2_7;
      end else if (10'h166 == _T_34[9:0]) begin
        image_2_358 <= io_pixelVal_in_2_6;
      end else if (10'h166 == _T_31[9:0]) begin
        image_2_358 <= io_pixelVal_in_2_5;
      end else if (10'h166 == _T_28[9:0]) begin
        image_2_358 <= io_pixelVal_in_2_4;
      end else if (10'h166 == _T_25[9:0]) begin
        image_2_358 <= io_pixelVal_in_2_3;
      end else if (10'h166 == _T_22[9:0]) begin
        image_2_358 <= io_pixelVal_in_2_2;
      end else if (10'h166 == _T_19[9:0]) begin
        image_2_358 <= io_pixelVal_in_2_1;
      end else if (10'h166 == _T_15[9:0]) begin
        image_2_358 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_359 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h167 == _T_37[9:0]) begin
        image_2_359 <= io_pixelVal_in_2_7;
      end else if (10'h167 == _T_34[9:0]) begin
        image_2_359 <= io_pixelVal_in_2_6;
      end else if (10'h167 == _T_31[9:0]) begin
        image_2_359 <= io_pixelVal_in_2_5;
      end else if (10'h167 == _T_28[9:0]) begin
        image_2_359 <= io_pixelVal_in_2_4;
      end else if (10'h167 == _T_25[9:0]) begin
        image_2_359 <= io_pixelVal_in_2_3;
      end else if (10'h167 == _T_22[9:0]) begin
        image_2_359 <= io_pixelVal_in_2_2;
      end else if (10'h167 == _T_19[9:0]) begin
        image_2_359 <= io_pixelVal_in_2_1;
      end else if (10'h167 == _T_15[9:0]) begin
        image_2_359 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_360 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h168 == _T_37[9:0]) begin
        image_2_360 <= io_pixelVal_in_2_7;
      end else if (10'h168 == _T_34[9:0]) begin
        image_2_360 <= io_pixelVal_in_2_6;
      end else if (10'h168 == _T_31[9:0]) begin
        image_2_360 <= io_pixelVal_in_2_5;
      end else if (10'h168 == _T_28[9:0]) begin
        image_2_360 <= io_pixelVal_in_2_4;
      end else if (10'h168 == _T_25[9:0]) begin
        image_2_360 <= io_pixelVal_in_2_3;
      end else if (10'h168 == _T_22[9:0]) begin
        image_2_360 <= io_pixelVal_in_2_2;
      end else if (10'h168 == _T_19[9:0]) begin
        image_2_360 <= io_pixelVal_in_2_1;
      end else if (10'h168 == _T_15[9:0]) begin
        image_2_360 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_361 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h169 == _T_37[9:0]) begin
        image_2_361 <= io_pixelVal_in_2_7;
      end else if (10'h169 == _T_34[9:0]) begin
        image_2_361 <= io_pixelVal_in_2_6;
      end else if (10'h169 == _T_31[9:0]) begin
        image_2_361 <= io_pixelVal_in_2_5;
      end else if (10'h169 == _T_28[9:0]) begin
        image_2_361 <= io_pixelVal_in_2_4;
      end else if (10'h169 == _T_25[9:0]) begin
        image_2_361 <= io_pixelVal_in_2_3;
      end else if (10'h169 == _T_22[9:0]) begin
        image_2_361 <= io_pixelVal_in_2_2;
      end else if (10'h169 == _T_19[9:0]) begin
        image_2_361 <= io_pixelVal_in_2_1;
      end else if (10'h169 == _T_15[9:0]) begin
        image_2_361 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_362 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h16a == _T_37[9:0]) begin
        image_2_362 <= io_pixelVal_in_2_7;
      end else if (10'h16a == _T_34[9:0]) begin
        image_2_362 <= io_pixelVal_in_2_6;
      end else if (10'h16a == _T_31[9:0]) begin
        image_2_362 <= io_pixelVal_in_2_5;
      end else if (10'h16a == _T_28[9:0]) begin
        image_2_362 <= io_pixelVal_in_2_4;
      end else if (10'h16a == _T_25[9:0]) begin
        image_2_362 <= io_pixelVal_in_2_3;
      end else if (10'h16a == _T_22[9:0]) begin
        image_2_362 <= io_pixelVal_in_2_2;
      end else if (10'h16a == _T_19[9:0]) begin
        image_2_362 <= io_pixelVal_in_2_1;
      end else if (10'h16a == _T_15[9:0]) begin
        image_2_362 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_363 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h16b == _T_37[9:0]) begin
        image_2_363 <= io_pixelVal_in_2_7;
      end else if (10'h16b == _T_34[9:0]) begin
        image_2_363 <= io_pixelVal_in_2_6;
      end else if (10'h16b == _T_31[9:0]) begin
        image_2_363 <= io_pixelVal_in_2_5;
      end else if (10'h16b == _T_28[9:0]) begin
        image_2_363 <= io_pixelVal_in_2_4;
      end else if (10'h16b == _T_25[9:0]) begin
        image_2_363 <= io_pixelVal_in_2_3;
      end else if (10'h16b == _T_22[9:0]) begin
        image_2_363 <= io_pixelVal_in_2_2;
      end else if (10'h16b == _T_19[9:0]) begin
        image_2_363 <= io_pixelVal_in_2_1;
      end else if (10'h16b == _T_15[9:0]) begin
        image_2_363 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_364 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h16c == _T_37[9:0]) begin
        image_2_364 <= io_pixelVal_in_2_7;
      end else if (10'h16c == _T_34[9:0]) begin
        image_2_364 <= io_pixelVal_in_2_6;
      end else if (10'h16c == _T_31[9:0]) begin
        image_2_364 <= io_pixelVal_in_2_5;
      end else if (10'h16c == _T_28[9:0]) begin
        image_2_364 <= io_pixelVal_in_2_4;
      end else if (10'h16c == _T_25[9:0]) begin
        image_2_364 <= io_pixelVal_in_2_3;
      end else if (10'h16c == _T_22[9:0]) begin
        image_2_364 <= io_pixelVal_in_2_2;
      end else if (10'h16c == _T_19[9:0]) begin
        image_2_364 <= io_pixelVal_in_2_1;
      end else if (10'h16c == _T_15[9:0]) begin
        image_2_364 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_365 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h16d == _T_37[9:0]) begin
        image_2_365 <= io_pixelVal_in_2_7;
      end else if (10'h16d == _T_34[9:0]) begin
        image_2_365 <= io_pixelVal_in_2_6;
      end else if (10'h16d == _T_31[9:0]) begin
        image_2_365 <= io_pixelVal_in_2_5;
      end else if (10'h16d == _T_28[9:0]) begin
        image_2_365 <= io_pixelVal_in_2_4;
      end else if (10'h16d == _T_25[9:0]) begin
        image_2_365 <= io_pixelVal_in_2_3;
      end else if (10'h16d == _T_22[9:0]) begin
        image_2_365 <= io_pixelVal_in_2_2;
      end else if (10'h16d == _T_19[9:0]) begin
        image_2_365 <= io_pixelVal_in_2_1;
      end else if (10'h16d == _T_15[9:0]) begin
        image_2_365 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_366 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h16e == _T_37[9:0]) begin
        image_2_366 <= io_pixelVal_in_2_7;
      end else if (10'h16e == _T_34[9:0]) begin
        image_2_366 <= io_pixelVal_in_2_6;
      end else if (10'h16e == _T_31[9:0]) begin
        image_2_366 <= io_pixelVal_in_2_5;
      end else if (10'h16e == _T_28[9:0]) begin
        image_2_366 <= io_pixelVal_in_2_4;
      end else if (10'h16e == _T_25[9:0]) begin
        image_2_366 <= io_pixelVal_in_2_3;
      end else if (10'h16e == _T_22[9:0]) begin
        image_2_366 <= io_pixelVal_in_2_2;
      end else if (10'h16e == _T_19[9:0]) begin
        image_2_366 <= io_pixelVal_in_2_1;
      end else if (10'h16e == _T_15[9:0]) begin
        image_2_366 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_367 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h16f == _T_37[9:0]) begin
        image_2_367 <= io_pixelVal_in_2_7;
      end else if (10'h16f == _T_34[9:0]) begin
        image_2_367 <= io_pixelVal_in_2_6;
      end else if (10'h16f == _T_31[9:0]) begin
        image_2_367 <= io_pixelVal_in_2_5;
      end else if (10'h16f == _T_28[9:0]) begin
        image_2_367 <= io_pixelVal_in_2_4;
      end else if (10'h16f == _T_25[9:0]) begin
        image_2_367 <= io_pixelVal_in_2_3;
      end else if (10'h16f == _T_22[9:0]) begin
        image_2_367 <= io_pixelVal_in_2_2;
      end else if (10'h16f == _T_19[9:0]) begin
        image_2_367 <= io_pixelVal_in_2_1;
      end else if (10'h16f == _T_15[9:0]) begin
        image_2_367 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_368 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h170 == _T_37[9:0]) begin
        image_2_368 <= io_pixelVal_in_2_7;
      end else if (10'h170 == _T_34[9:0]) begin
        image_2_368 <= io_pixelVal_in_2_6;
      end else if (10'h170 == _T_31[9:0]) begin
        image_2_368 <= io_pixelVal_in_2_5;
      end else if (10'h170 == _T_28[9:0]) begin
        image_2_368 <= io_pixelVal_in_2_4;
      end else if (10'h170 == _T_25[9:0]) begin
        image_2_368 <= io_pixelVal_in_2_3;
      end else if (10'h170 == _T_22[9:0]) begin
        image_2_368 <= io_pixelVal_in_2_2;
      end else if (10'h170 == _T_19[9:0]) begin
        image_2_368 <= io_pixelVal_in_2_1;
      end else if (10'h170 == _T_15[9:0]) begin
        image_2_368 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_369 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h171 == _T_37[9:0]) begin
        image_2_369 <= io_pixelVal_in_2_7;
      end else if (10'h171 == _T_34[9:0]) begin
        image_2_369 <= io_pixelVal_in_2_6;
      end else if (10'h171 == _T_31[9:0]) begin
        image_2_369 <= io_pixelVal_in_2_5;
      end else if (10'h171 == _T_28[9:0]) begin
        image_2_369 <= io_pixelVal_in_2_4;
      end else if (10'h171 == _T_25[9:0]) begin
        image_2_369 <= io_pixelVal_in_2_3;
      end else if (10'h171 == _T_22[9:0]) begin
        image_2_369 <= io_pixelVal_in_2_2;
      end else if (10'h171 == _T_19[9:0]) begin
        image_2_369 <= io_pixelVal_in_2_1;
      end else if (10'h171 == _T_15[9:0]) begin
        image_2_369 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_370 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h172 == _T_37[9:0]) begin
        image_2_370 <= io_pixelVal_in_2_7;
      end else if (10'h172 == _T_34[9:0]) begin
        image_2_370 <= io_pixelVal_in_2_6;
      end else if (10'h172 == _T_31[9:0]) begin
        image_2_370 <= io_pixelVal_in_2_5;
      end else if (10'h172 == _T_28[9:0]) begin
        image_2_370 <= io_pixelVal_in_2_4;
      end else if (10'h172 == _T_25[9:0]) begin
        image_2_370 <= io_pixelVal_in_2_3;
      end else if (10'h172 == _T_22[9:0]) begin
        image_2_370 <= io_pixelVal_in_2_2;
      end else if (10'h172 == _T_19[9:0]) begin
        image_2_370 <= io_pixelVal_in_2_1;
      end else if (10'h172 == _T_15[9:0]) begin
        image_2_370 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_371 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h173 == _T_37[9:0]) begin
        image_2_371 <= io_pixelVal_in_2_7;
      end else if (10'h173 == _T_34[9:0]) begin
        image_2_371 <= io_pixelVal_in_2_6;
      end else if (10'h173 == _T_31[9:0]) begin
        image_2_371 <= io_pixelVal_in_2_5;
      end else if (10'h173 == _T_28[9:0]) begin
        image_2_371 <= io_pixelVal_in_2_4;
      end else if (10'h173 == _T_25[9:0]) begin
        image_2_371 <= io_pixelVal_in_2_3;
      end else if (10'h173 == _T_22[9:0]) begin
        image_2_371 <= io_pixelVal_in_2_2;
      end else if (10'h173 == _T_19[9:0]) begin
        image_2_371 <= io_pixelVal_in_2_1;
      end else if (10'h173 == _T_15[9:0]) begin
        image_2_371 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_372 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h174 == _T_37[9:0]) begin
        image_2_372 <= io_pixelVal_in_2_7;
      end else if (10'h174 == _T_34[9:0]) begin
        image_2_372 <= io_pixelVal_in_2_6;
      end else if (10'h174 == _T_31[9:0]) begin
        image_2_372 <= io_pixelVal_in_2_5;
      end else if (10'h174 == _T_28[9:0]) begin
        image_2_372 <= io_pixelVal_in_2_4;
      end else if (10'h174 == _T_25[9:0]) begin
        image_2_372 <= io_pixelVal_in_2_3;
      end else if (10'h174 == _T_22[9:0]) begin
        image_2_372 <= io_pixelVal_in_2_2;
      end else if (10'h174 == _T_19[9:0]) begin
        image_2_372 <= io_pixelVal_in_2_1;
      end else if (10'h174 == _T_15[9:0]) begin
        image_2_372 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_373 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h175 == _T_37[9:0]) begin
        image_2_373 <= io_pixelVal_in_2_7;
      end else if (10'h175 == _T_34[9:0]) begin
        image_2_373 <= io_pixelVal_in_2_6;
      end else if (10'h175 == _T_31[9:0]) begin
        image_2_373 <= io_pixelVal_in_2_5;
      end else if (10'h175 == _T_28[9:0]) begin
        image_2_373 <= io_pixelVal_in_2_4;
      end else if (10'h175 == _T_25[9:0]) begin
        image_2_373 <= io_pixelVal_in_2_3;
      end else if (10'h175 == _T_22[9:0]) begin
        image_2_373 <= io_pixelVal_in_2_2;
      end else if (10'h175 == _T_19[9:0]) begin
        image_2_373 <= io_pixelVal_in_2_1;
      end else if (10'h175 == _T_15[9:0]) begin
        image_2_373 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_374 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h176 == _T_37[9:0]) begin
        image_2_374 <= io_pixelVal_in_2_7;
      end else if (10'h176 == _T_34[9:0]) begin
        image_2_374 <= io_pixelVal_in_2_6;
      end else if (10'h176 == _T_31[9:0]) begin
        image_2_374 <= io_pixelVal_in_2_5;
      end else if (10'h176 == _T_28[9:0]) begin
        image_2_374 <= io_pixelVal_in_2_4;
      end else if (10'h176 == _T_25[9:0]) begin
        image_2_374 <= io_pixelVal_in_2_3;
      end else if (10'h176 == _T_22[9:0]) begin
        image_2_374 <= io_pixelVal_in_2_2;
      end else if (10'h176 == _T_19[9:0]) begin
        image_2_374 <= io_pixelVal_in_2_1;
      end else if (10'h176 == _T_15[9:0]) begin
        image_2_374 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_375 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h177 == _T_37[9:0]) begin
        image_2_375 <= io_pixelVal_in_2_7;
      end else if (10'h177 == _T_34[9:0]) begin
        image_2_375 <= io_pixelVal_in_2_6;
      end else if (10'h177 == _T_31[9:0]) begin
        image_2_375 <= io_pixelVal_in_2_5;
      end else if (10'h177 == _T_28[9:0]) begin
        image_2_375 <= io_pixelVal_in_2_4;
      end else if (10'h177 == _T_25[9:0]) begin
        image_2_375 <= io_pixelVal_in_2_3;
      end else if (10'h177 == _T_22[9:0]) begin
        image_2_375 <= io_pixelVal_in_2_2;
      end else if (10'h177 == _T_19[9:0]) begin
        image_2_375 <= io_pixelVal_in_2_1;
      end else if (10'h177 == _T_15[9:0]) begin
        image_2_375 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_376 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h178 == _T_37[9:0]) begin
        image_2_376 <= io_pixelVal_in_2_7;
      end else if (10'h178 == _T_34[9:0]) begin
        image_2_376 <= io_pixelVal_in_2_6;
      end else if (10'h178 == _T_31[9:0]) begin
        image_2_376 <= io_pixelVal_in_2_5;
      end else if (10'h178 == _T_28[9:0]) begin
        image_2_376 <= io_pixelVal_in_2_4;
      end else if (10'h178 == _T_25[9:0]) begin
        image_2_376 <= io_pixelVal_in_2_3;
      end else if (10'h178 == _T_22[9:0]) begin
        image_2_376 <= io_pixelVal_in_2_2;
      end else if (10'h178 == _T_19[9:0]) begin
        image_2_376 <= io_pixelVal_in_2_1;
      end else if (10'h178 == _T_15[9:0]) begin
        image_2_376 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_377 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h179 == _T_37[9:0]) begin
        image_2_377 <= io_pixelVal_in_2_7;
      end else if (10'h179 == _T_34[9:0]) begin
        image_2_377 <= io_pixelVal_in_2_6;
      end else if (10'h179 == _T_31[9:0]) begin
        image_2_377 <= io_pixelVal_in_2_5;
      end else if (10'h179 == _T_28[9:0]) begin
        image_2_377 <= io_pixelVal_in_2_4;
      end else if (10'h179 == _T_25[9:0]) begin
        image_2_377 <= io_pixelVal_in_2_3;
      end else if (10'h179 == _T_22[9:0]) begin
        image_2_377 <= io_pixelVal_in_2_2;
      end else if (10'h179 == _T_19[9:0]) begin
        image_2_377 <= io_pixelVal_in_2_1;
      end else if (10'h179 == _T_15[9:0]) begin
        image_2_377 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_378 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h17a == _T_37[9:0]) begin
        image_2_378 <= io_pixelVal_in_2_7;
      end else if (10'h17a == _T_34[9:0]) begin
        image_2_378 <= io_pixelVal_in_2_6;
      end else if (10'h17a == _T_31[9:0]) begin
        image_2_378 <= io_pixelVal_in_2_5;
      end else if (10'h17a == _T_28[9:0]) begin
        image_2_378 <= io_pixelVal_in_2_4;
      end else if (10'h17a == _T_25[9:0]) begin
        image_2_378 <= io_pixelVal_in_2_3;
      end else if (10'h17a == _T_22[9:0]) begin
        image_2_378 <= io_pixelVal_in_2_2;
      end else if (10'h17a == _T_19[9:0]) begin
        image_2_378 <= io_pixelVal_in_2_1;
      end else if (10'h17a == _T_15[9:0]) begin
        image_2_378 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_379 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h17b == _T_37[9:0]) begin
        image_2_379 <= io_pixelVal_in_2_7;
      end else if (10'h17b == _T_34[9:0]) begin
        image_2_379 <= io_pixelVal_in_2_6;
      end else if (10'h17b == _T_31[9:0]) begin
        image_2_379 <= io_pixelVal_in_2_5;
      end else if (10'h17b == _T_28[9:0]) begin
        image_2_379 <= io_pixelVal_in_2_4;
      end else if (10'h17b == _T_25[9:0]) begin
        image_2_379 <= io_pixelVal_in_2_3;
      end else if (10'h17b == _T_22[9:0]) begin
        image_2_379 <= io_pixelVal_in_2_2;
      end else if (10'h17b == _T_19[9:0]) begin
        image_2_379 <= io_pixelVal_in_2_1;
      end else if (10'h17b == _T_15[9:0]) begin
        image_2_379 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_380 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h17c == _T_37[9:0]) begin
        image_2_380 <= io_pixelVal_in_2_7;
      end else if (10'h17c == _T_34[9:0]) begin
        image_2_380 <= io_pixelVal_in_2_6;
      end else if (10'h17c == _T_31[9:0]) begin
        image_2_380 <= io_pixelVal_in_2_5;
      end else if (10'h17c == _T_28[9:0]) begin
        image_2_380 <= io_pixelVal_in_2_4;
      end else if (10'h17c == _T_25[9:0]) begin
        image_2_380 <= io_pixelVal_in_2_3;
      end else if (10'h17c == _T_22[9:0]) begin
        image_2_380 <= io_pixelVal_in_2_2;
      end else if (10'h17c == _T_19[9:0]) begin
        image_2_380 <= io_pixelVal_in_2_1;
      end else if (10'h17c == _T_15[9:0]) begin
        image_2_380 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_381 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h17d == _T_37[9:0]) begin
        image_2_381 <= io_pixelVal_in_2_7;
      end else if (10'h17d == _T_34[9:0]) begin
        image_2_381 <= io_pixelVal_in_2_6;
      end else if (10'h17d == _T_31[9:0]) begin
        image_2_381 <= io_pixelVal_in_2_5;
      end else if (10'h17d == _T_28[9:0]) begin
        image_2_381 <= io_pixelVal_in_2_4;
      end else if (10'h17d == _T_25[9:0]) begin
        image_2_381 <= io_pixelVal_in_2_3;
      end else if (10'h17d == _T_22[9:0]) begin
        image_2_381 <= io_pixelVal_in_2_2;
      end else if (10'h17d == _T_19[9:0]) begin
        image_2_381 <= io_pixelVal_in_2_1;
      end else if (10'h17d == _T_15[9:0]) begin
        image_2_381 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_382 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h17e == _T_37[9:0]) begin
        image_2_382 <= io_pixelVal_in_2_7;
      end else if (10'h17e == _T_34[9:0]) begin
        image_2_382 <= io_pixelVal_in_2_6;
      end else if (10'h17e == _T_31[9:0]) begin
        image_2_382 <= io_pixelVal_in_2_5;
      end else if (10'h17e == _T_28[9:0]) begin
        image_2_382 <= io_pixelVal_in_2_4;
      end else if (10'h17e == _T_25[9:0]) begin
        image_2_382 <= io_pixelVal_in_2_3;
      end else if (10'h17e == _T_22[9:0]) begin
        image_2_382 <= io_pixelVal_in_2_2;
      end else if (10'h17e == _T_19[9:0]) begin
        image_2_382 <= io_pixelVal_in_2_1;
      end else if (10'h17e == _T_15[9:0]) begin
        image_2_382 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_383 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h17f == _T_37[9:0]) begin
        image_2_383 <= io_pixelVal_in_2_7;
      end else if (10'h17f == _T_34[9:0]) begin
        image_2_383 <= io_pixelVal_in_2_6;
      end else if (10'h17f == _T_31[9:0]) begin
        image_2_383 <= io_pixelVal_in_2_5;
      end else if (10'h17f == _T_28[9:0]) begin
        image_2_383 <= io_pixelVal_in_2_4;
      end else if (10'h17f == _T_25[9:0]) begin
        image_2_383 <= io_pixelVal_in_2_3;
      end else if (10'h17f == _T_22[9:0]) begin
        image_2_383 <= io_pixelVal_in_2_2;
      end else if (10'h17f == _T_19[9:0]) begin
        image_2_383 <= io_pixelVal_in_2_1;
      end else if (10'h17f == _T_15[9:0]) begin
        image_2_383 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_384 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h180 == _T_37[9:0]) begin
        image_2_384 <= io_pixelVal_in_2_7;
      end else if (10'h180 == _T_34[9:0]) begin
        image_2_384 <= io_pixelVal_in_2_6;
      end else if (10'h180 == _T_31[9:0]) begin
        image_2_384 <= io_pixelVal_in_2_5;
      end else if (10'h180 == _T_28[9:0]) begin
        image_2_384 <= io_pixelVal_in_2_4;
      end else if (10'h180 == _T_25[9:0]) begin
        image_2_384 <= io_pixelVal_in_2_3;
      end else if (10'h180 == _T_22[9:0]) begin
        image_2_384 <= io_pixelVal_in_2_2;
      end else if (10'h180 == _T_19[9:0]) begin
        image_2_384 <= io_pixelVal_in_2_1;
      end else if (10'h180 == _T_15[9:0]) begin
        image_2_384 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_385 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h181 == _T_37[9:0]) begin
        image_2_385 <= io_pixelVal_in_2_7;
      end else if (10'h181 == _T_34[9:0]) begin
        image_2_385 <= io_pixelVal_in_2_6;
      end else if (10'h181 == _T_31[9:0]) begin
        image_2_385 <= io_pixelVal_in_2_5;
      end else if (10'h181 == _T_28[9:0]) begin
        image_2_385 <= io_pixelVal_in_2_4;
      end else if (10'h181 == _T_25[9:0]) begin
        image_2_385 <= io_pixelVal_in_2_3;
      end else if (10'h181 == _T_22[9:0]) begin
        image_2_385 <= io_pixelVal_in_2_2;
      end else if (10'h181 == _T_19[9:0]) begin
        image_2_385 <= io_pixelVal_in_2_1;
      end else if (10'h181 == _T_15[9:0]) begin
        image_2_385 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_386 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h182 == _T_37[9:0]) begin
        image_2_386 <= io_pixelVal_in_2_7;
      end else if (10'h182 == _T_34[9:0]) begin
        image_2_386 <= io_pixelVal_in_2_6;
      end else if (10'h182 == _T_31[9:0]) begin
        image_2_386 <= io_pixelVal_in_2_5;
      end else if (10'h182 == _T_28[9:0]) begin
        image_2_386 <= io_pixelVal_in_2_4;
      end else if (10'h182 == _T_25[9:0]) begin
        image_2_386 <= io_pixelVal_in_2_3;
      end else if (10'h182 == _T_22[9:0]) begin
        image_2_386 <= io_pixelVal_in_2_2;
      end else if (10'h182 == _T_19[9:0]) begin
        image_2_386 <= io_pixelVal_in_2_1;
      end else if (10'h182 == _T_15[9:0]) begin
        image_2_386 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_387 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h183 == _T_37[9:0]) begin
        image_2_387 <= io_pixelVal_in_2_7;
      end else if (10'h183 == _T_34[9:0]) begin
        image_2_387 <= io_pixelVal_in_2_6;
      end else if (10'h183 == _T_31[9:0]) begin
        image_2_387 <= io_pixelVal_in_2_5;
      end else if (10'h183 == _T_28[9:0]) begin
        image_2_387 <= io_pixelVal_in_2_4;
      end else if (10'h183 == _T_25[9:0]) begin
        image_2_387 <= io_pixelVal_in_2_3;
      end else if (10'h183 == _T_22[9:0]) begin
        image_2_387 <= io_pixelVal_in_2_2;
      end else if (10'h183 == _T_19[9:0]) begin
        image_2_387 <= io_pixelVal_in_2_1;
      end else if (10'h183 == _T_15[9:0]) begin
        image_2_387 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_388 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h184 == _T_37[9:0]) begin
        image_2_388 <= io_pixelVal_in_2_7;
      end else if (10'h184 == _T_34[9:0]) begin
        image_2_388 <= io_pixelVal_in_2_6;
      end else if (10'h184 == _T_31[9:0]) begin
        image_2_388 <= io_pixelVal_in_2_5;
      end else if (10'h184 == _T_28[9:0]) begin
        image_2_388 <= io_pixelVal_in_2_4;
      end else if (10'h184 == _T_25[9:0]) begin
        image_2_388 <= io_pixelVal_in_2_3;
      end else if (10'h184 == _T_22[9:0]) begin
        image_2_388 <= io_pixelVal_in_2_2;
      end else if (10'h184 == _T_19[9:0]) begin
        image_2_388 <= io_pixelVal_in_2_1;
      end else if (10'h184 == _T_15[9:0]) begin
        image_2_388 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_389 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h185 == _T_37[9:0]) begin
        image_2_389 <= io_pixelVal_in_2_7;
      end else if (10'h185 == _T_34[9:0]) begin
        image_2_389 <= io_pixelVal_in_2_6;
      end else if (10'h185 == _T_31[9:0]) begin
        image_2_389 <= io_pixelVal_in_2_5;
      end else if (10'h185 == _T_28[9:0]) begin
        image_2_389 <= io_pixelVal_in_2_4;
      end else if (10'h185 == _T_25[9:0]) begin
        image_2_389 <= io_pixelVal_in_2_3;
      end else if (10'h185 == _T_22[9:0]) begin
        image_2_389 <= io_pixelVal_in_2_2;
      end else if (10'h185 == _T_19[9:0]) begin
        image_2_389 <= io_pixelVal_in_2_1;
      end else if (10'h185 == _T_15[9:0]) begin
        image_2_389 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_390 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h186 == _T_37[9:0]) begin
        image_2_390 <= io_pixelVal_in_2_7;
      end else if (10'h186 == _T_34[9:0]) begin
        image_2_390 <= io_pixelVal_in_2_6;
      end else if (10'h186 == _T_31[9:0]) begin
        image_2_390 <= io_pixelVal_in_2_5;
      end else if (10'h186 == _T_28[9:0]) begin
        image_2_390 <= io_pixelVal_in_2_4;
      end else if (10'h186 == _T_25[9:0]) begin
        image_2_390 <= io_pixelVal_in_2_3;
      end else if (10'h186 == _T_22[9:0]) begin
        image_2_390 <= io_pixelVal_in_2_2;
      end else if (10'h186 == _T_19[9:0]) begin
        image_2_390 <= io_pixelVal_in_2_1;
      end else if (10'h186 == _T_15[9:0]) begin
        image_2_390 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_391 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h187 == _T_37[9:0]) begin
        image_2_391 <= io_pixelVal_in_2_7;
      end else if (10'h187 == _T_34[9:0]) begin
        image_2_391 <= io_pixelVal_in_2_6;
      end else if (10'h187 == _T_31[9:0]) begin
        image_2_391 <= io_pixelVal_in_2_5;
      end else if (10'h187 == _T_28[9:0]) begin
        image_2_391 <= io_pixelVal_in_2_4;
      end else if (10'h187 == _T_25[9:0]) begin
        image_2_391 <= io_pixelVal_in_2_3;
      end else if (10'h187 == _T_22[9:0]) begin
        image_2_391 <= io_pixelVal_in_2_2;
      end else if (10'h187 == _T_19[9:0]) begin
        image_2_391 <= io_pixelVal_in_2_1;
      end else if (10'h187 == _T_15[9:0]) begin
        image_2_391 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_392 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h188 == _T_37[9:0]) begin
        image_2_392 <= io_pixelVal_in_2_7;
      end else if (10'h188 == _T_34[9:0]) begin
        image_2_392 <= io_pixelVal_in_2_6;
      end else if (10'h188 == _T_31[9:0]) begin
        image_2_392 <= io_pixelVal_in_2_5;
      end else if (10'h188 == _T_28[9:0]) begin
        image_2_392 <= io_pixelVal_in_2_4;
      end else if (10'h188 == _T_25[9:0]) begin
        image_2_392 <= io_pixelVal_in_2_3;
      end else if (10'h188 == _T_22[9:0]) begin
        image_2_392 <= io_pixelVal_in_2_2;
      end else if (10'h188 == _T_19[9:0]) begin
        image_2_392 <= io_pixelVal_in_2_1;
      end else if (10'h188 == _T_15[9:0]) begin
        image_2_392 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_393 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h189 == _T_37[9:0]) begin
        image_2_393 <= io_pixelVal_in_2_7;
      end else if (10'h189 == _T_34[9:0]) begin
        image_2_393 <= io_pixelVal_in_2_6;
      end else if (10'h189 == _T_31[9:0]) begin
        image_2_393 <= io_pixelVal_in_2_5;
      end else if (10'h189 == _T_28[9:0]) begin
        image_2_393 <= io_pixelVal_in_2_4;
      end else if (10'h189 == _T_25[9:0]) begin
        image_2_393 <= io_pixelVal_in_2_3;
      end else if (10'h189 == _T_22[9:0]) begin
        image_2_393 <= io_pixelVal_in_2_2;
      end else if (10'h189 == _T_19[9:0]) begin
        image_2_393 <= io_pixelVal_in_2_1;
      end else if (10'h189 == _T_15[9:0]) begin
        image_2_393 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_394 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h18a == _T_37[9:0]) begin
        image_2_394 <= io_pixelVal_in_2_7;
      end else if (10'h18a == _T_34[9:0]) begin
        image_2_394 <= io_pixelVal_in_2_6;
      end else if (10'h18a == _T_31[9:0]) begin
        image_2_394 <= io_pixelVal_in_2_5;
      end else if (10'h18a == _T_28[9:0]) begin
        image_2_394 <= io_pixelVal_in_2_4;
      end else if (10'h18a == _T_25[9:0]) begin
        image_2_394 <= io_pixelVal_in_2_3;
      end else if (10'h18a == _T_22[9:0]) begin
        image_2_394 <= io_pixelVal_in_2_2;
      end else if (10'h18a == _T_19[9:0]) begin
        image_2_394 <= io_pixelVal_in_2_1;
      end else if (10'h18a == _T_15[9:0]) begin
        image_2_394 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_395 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h18b == _T_37[9:0]) begin
        image_2_395 <= io_pixelVal_in_2_7;
      end else if (10'h18b == _T_34[9:0]) begin
        image_2_395 <= io_pixelVal_in_2_6;
      end else if (10'h18b == _T_31[9:0]) begin
        image_2_395 <= io_pixelVal_in_2_5;
      end else if (10'h18b == _T_28[9:0]) begin
        image_2_395 <= io_pixelVal_in_2_4;
      end else if (10'h18b == _T_25[9:0]) begin
        image_2_395 <= io_pixelVal_in_2_3;
      end else if (10'h18b == _T_22[9:0]) begin
        image_2_395 <= io_pixelVal_in_2_2;
      end else if (10'h18b == _T_19[9:0]) begin
        image_2_395 <= io_pixelVal_in_2_1;
      end else if (10'h18b == _T_15[9:0]) begin
        image_2_395 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_396 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h18c == _T_37[9:0]) begin
        image_2_396 <= io_pixelVal_in_2_7;
      end else if (10'h18c == _T_34[9:0]) begin
        image_2_396 <= io_pixelVal_in_2_6;
      end else if (10'h18c == _T_31[9:0]) begin
        image_2_396 <= io_pixelVal_in_2_5;
      end else if (10'h18c == _T_28[9:0]) begin
        image_2_396 <= io_pixelVal_in_2_4;
      end else if (10'h18c == _T_25[9:0]) begin
        image_2_396 <= io_pixelVal_in_2_3;
      end else if (10'h18c == _T_22[9:0]) begin
        image_2_396 <= io_pixelVal_in_2_2;
      end else if (10'h18c == _T_19[9:0]) begin
        image_2_396 <= io_pixelVal_in_2_1;
      end else if (10'h18c == _T_15[9:0]) begin
        image_2_396 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_397 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h18d == _T_37[9:0]) begin
        image_2_397 <= io_pixelVal_in_2_7;
      end else if (10'h18d == _T_34[9:0]) begin
        image_2_397 <= io_pixelVal_in_2_6;
      end else if (10'h18d == _T_31[9:0]) begin
        image_2_397 <= io_pixelVal_in_2_5;
      end else if (10'h18d == _T_28[9:0]) begin
        image_2_397 <= io_pixelVal_in_2_4;
      end else if (10'h18d == _T_25[9:0]) begin
        image_2_397 <= io_pixelVal_in_2_3;
      end else if (10'h18d == _T_22[9:0]) begin
        image_2_397 <= io_pixelVal_in_2_2;
      end else if (10'h18d == _T_19[9:0]) begin
        image_2_397 <= io_pixelVal_in_2_1;
      end else if (10'h18d == _T_15[9:0]) begin
        image_2_397 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_398 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h18e == _T_37[9:0]) begin
        image_2_398 <= io_pixelVal_in_2_7;
      end else if (10'h18e == _T_34[9:0]) begin
        image_2_398 <= io_pixelVal_in_2_6;
      end else if (10'h18e == _T_31[9:0]) begin
        image_2_398 <= io_pixelVal_in_2_5;
      end else if (10'h18e == _T_28[9:0]) begin
        image_2_398 <= io_pixelVal_in_2_4;
      end else if (10'h18e == _T_25[9:0]) begin
        image_2_398 <= io_pixelVal_in_2_3;
      end else if (10'h18e == _T_22[9:0]) begin
        image_2_398 <= io_pixelVal_in_2_2;
      end else if (10'h18e == _T_19[9:0]) begin
        image_2_398 <= io_pixelVal_in_2_1;
      end else if (10'h18e == _T_15[9:0]) begin
        image_2_398 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_399 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h18f == _T_37[9:0]) begin
        image_2_399 <= io_pixelVal_in_2_7;
      end else if (10'h18f == _T_34[9:0]) begin
        image_2_399 <= io_pixelVal_in_2_6;
      end else if (10'h18f == _T_31[9:0]) begin
        image_2_399 <= io_pixelVal_in_2_5;
      end else if (10'h18f == _T_28[9:0]) begin
        image_2_399 <= io_pixelVal_in_2_4;
      end else if (10'h18f == _T_25[9:0]) begin
        image_2_399 <= io_pixelVal_in_2_3;
      end else if (10'h18f == _T_22[9:0]) begin
        image_2_399 <= io_pixelVal_in_2_2;
      end else if (10'h18f == _T_19[9:0]) begin
        image_2_399 <= io_pixelVal_in_2_1;
      end else if (10'h18f == _T_15[9:0]) begin
        image_2_399 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_400 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h190 == _T_37[9:0]) begin
        image_2_400 <= io_pixelVal_in_2_7;
      end else if (10'h190 == _T_34[9:0]) begin
        image_2_400 <= io_pixelVal_in_2_6;
      end else if (10'h190 == _T_31[9:0]) begin
        image_2_400 <= io_pixelVal_in_2_5;
      end else if (10'h190 == _T_28[9:0]) begin
        image_2_400 <= io_pixelVal_in_2_4;
      end else if (10'h190 == _T_25[9:0]) begin
        image_2_400 <= io_pixelVal_in_2_3;
      end else if (10'h190 == _T_22[9:0]) begin
        image_2_400 <= io_pixelVal_in_2_2;
      end else if (10'h190 == _T_19[9:0]) begin
        image_2_400 <= io_pixelVal_in_2_1;
      end else if (10'h190 == _T_15[9:0]) begin
        image_2_400 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_401 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h191 == _T_37[9:0]) begin
        image_2_401 <= io_pixelVal_in_2_7;
      end else if (10'h191 == _T_34[9:0]) begin
        image_2_401 <= io_pixelVal_in_2_6;
      end else if (10'h191 == _T_31[9:0]) begin
        image_2_401 <= io_pixelVal_in_2_5;
      end else if (10'h191 == _T_28[9:0]) begin
        image_2_401 <= io_pixelVal_in_2_4;
      end else if (10'h191 == _T_25[9:0]) begin
        image_2_401 <= io_pixelVal_in_2_3;
      end else if (10'h191 == _T_22[9:0]) begin
        image_2_401 <= io_pixelVal_in_2_2;
      end else if (10'h191 == _T_19[9:0]) begin
        image_2_401 <= io_pixelVal_in_2_1;
      end else if (10'h191 == _T_15[9:0]) begin
        image_2_401 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_402 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h192 == _T_37[9:0]) begin
        image_2_402 <= io_pixelVal_in_2_7;
      end else if (10'h192 == _T_34[9:0]) begin
        image_2_402 <= io_pixelVal_in_2_6;
      end else if (10'h192 == _T_31[9:0]) begin
        image_2_402 <= io_pixelVal_in_2_5;
      end else if (10'h192 == _T_28[9:0]) begin
        image_2_402 <= io_pixelVal_in_2_4;
      end else if (10'h192 == _T_25[9:0]) begin
        image_2_402 <= io_pixelVal_in_2_3;
      end else if (10'h192 == _T_22[9:0]) begin
        image_2_402 <= io_pixelVal_in_2_2;
      end else if (10'h192 == _T_19[9:0]) begin
        image_2_402 <= io_pixelVal_in_2_1;
      end else if (10'h192 == _T_15[9:0]) begin
        image_2_402 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_403 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h193 == _T_37[9:0]) begin
        image_2_403 <= io_pixelVal_in_2_7;
      end else if (10'h193 == _T_34[9:0]) begin
        image_2_403 <= io_pixelVal_in_2_6;
      end else if (10'h193 == _T_31[9:0]) begin
        image_2_403 <= io_pixelVal_in_2_5;
      end else if (10'h193 == _T_28[9:0]) begin
        image_2_403 <= io_pixelVal_in_2_4;
      end else if (10'h193 == _T_25[9:0]) begin
        image_2_403 <= io_pixelVal_in_2_3;
      end else if (10'h193 == _T_22[9:0]) begin
        image_2_403 <= io_pixelVal_in_2_2;
      end else if (10'h193 == _T_19[9:0]) begin
        image_2_403 <= io_pixelVal_in_2_1;
      end else if (10'h193 == _T_15[9:0]) begin
        image_2_403 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_404 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h194 == _T_37[9:0]) begin
        image_2_404 <= io_pixelVal_in_2_7;
      end else if (10'h194 == _T_34[9:0]) begin
        image_2_404 <= io_pixelVal_in_2_6;
      end else if (10'h194 == _T_31[9:0]) begin
        image_2_404 <= io_pixelVal_in_2_5;
      end else if (10'h194 == _T_28[9:0]) begin
        image_2_404 <= io_pixelVal_in_2_4;
      end else if (10'h194 == _T_25[9:0]) begin
        image_2_404 <= io_pixelVal_in_2_3;
      end else if (10'h194 == _T_22[9:0]) begin
        image_2_404 <= io_pixelVal_in_2_2;
      end else if (10'h194 == _T_19[9:0]) begin
        image_2_404 <= io_pixelVal_in_2_1;
      end else if (10'h194 == _T_15[9:0]) begin
        image_2_404 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_405 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h195 == _T_37[9:0]) begin
        image_2_405 <= io_pixelVal_in_2_7;
      end else if (10'h195 == _T_34[9:0]) begin
        image_2_405 <= io_pixelVal_in_2_6;
      end else if (10'h195 == _T_31[9:0]) begin
        image_2_405 <= io_pixelVal_in_2_5;
      end else if (10'h195 == _T_28[9:0]) begin
        image_2_405 <= io_pixelVal_in_2_4;
      end else if (10'h195 == _T_25[9:0]) begin
        image_2_405 <= io_pixelVal_in_2_3;
      end else if (10'h195 == _T_22[9:0]) begin
        image_2_405 <= io_pixelVal_in_2_2;
      end else if (10'h195 == _T_19[9:0]) begin
        image_2_405 <= io_pixelVal_in_2_1;
      end else if (10'h195 == _T_15[9:0]) begin
        image_2_405 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_406 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h196 == _T_37[9:0]) begin
        image_2_406 <= io_pixelVal_in_2_7;
      end else if (10'h196 == _T_34[9:0]) begin
        image_2_406 <= io_pixelVal_in_2_6;
      end else if (10'h196 == _T_31[9:0]) begin
        image_2_406 <= io_pixelVal_in_2_5;
      end else if (10'h196 == _T_28[9:0]) begin
        image_2_406 <= io_pixelVal_in_2_4;
      end else if (10'h196 == _T_25[9:0]) begin
        image_2_406 <= io_pixelVal_in_2_3;
      end else if (10'h196 == _T_22[9:0]) begin
        image_2_406 <= io_pixelVal_in_2_2;
      end else if (10'h196 == _T_19[9:0]) begin
        image_2_406 <= io_pixelVal_in_2_1;
      end else if (10'h196 == _T_15[9:0]) begin
        image_2_406 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_407 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h197 == _T_37[9:0]) begin
        image_2_407 <= io_pixelVal_in_2_7;
      end else if (10'h197 == _T_34[9:0]) begin
        image_2_407 <= io_pixelVal_in_2_6;
      end else if (10'h197 == _T_31[9:0]) begin
        image_2_407 <= io_pixelVal_in_2_5;
      end else if (10'h197 == _T_28[9:0]) begin
        image_2_407 <= io_pixelVal_in_2_4;
      end else if (10'h197 == _T_25[9:0]) begin
        image_2_407 <= io_pixelVal_in_2_3;
      end else if (10'h197 == _T_22[9:0]) begin
        image_2_407 <= io_pixelVal_in_2_2;
      end else if (10'h197 == _T_19[9:0]) begin
        image_2_407 <= io_pixelVal_in_2_1;
      end else if (10'h197 == _T_15[9:0]) begin
        image_2_407 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_408 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h198 == _T_37[9:0]) begin
        image_2_408 <= io_pixelVal_in_2_7;
      end else if (10'h198 == _T_34[9:0]) begin
        image_2_408 <= io_pixelVal_in_2_6;
      end else if (10'h198 == _T_31[9:0]) begin
        image_2_408 <= io_pixelVal_in_2_5;
      end else if (10'h198 == _T_28[9:0]) begin
        image_2_408 <= io_pixelVal_in_2_4;
      end else if (10'h198 == _T_25[9:0]) begin
        image_2_408 <= io_pixelVal_in_2_3;
      end else if (10'h198 == _T_22[9:0]) begin
        image_2_408 <= io_pixelVal_in_2_2;
      end else if (10'h198 == _T_19[9:0]) begin
        image_2_408 <= io_pixelVal_in_2_1;
      end else if (10'h198 == _T_15[9:0]) begin
        image_2_408 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_409 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h199 == _T_37[9:0]) begin
        image_2_409 <= io_pixelVal_in_2_7;
      end else if (10'h199 == _T_34[9:0]) begin
        image_2_409 <= io_pixelVal_in_2_6;
      end else if (10'h199 == _T_31[9:0]) begin
        image_2_409 <= io_pixelVal_in_2_5;
      end else if (10'h199 == _T_28[9:0]) begin
        image_2_409 <= io_pixelVal_in_2_4;
      end else if (10'h199 == _T_25[9:0]) begin
        image_2_409 <= io_pixelVal_in_2_3;
      end else if (10'h199 == _T_22[9:0]) begin
        image_2_409 <= io_pixelVal_in_2_2;
      end else if (10'h199 == _T_19[9:0]) begin
        image_2_409 <= io_pixelVal_in_2_1;
      end else if (10'h199 == _T_15[9:0]) begin
        image_2_409 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_410 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h19a == _T_37[9:0]) begin
        image_2_410 <= io_pixelVal_in_2_7;
      end else if (10'h19a == _T_34[9:0]) begin
        image_2_410 <= io_pixelVal_in_2_6;
      end else if (10'h19a == _T_31[9:0]) begin
        image_2_410 <= io_pixelVal_in_2_5;
      end else if (10'h19a == _T_28[9:0]) begin
        image_2_410 <= io_pixelVal_in_2_4;
      end else if (10'h19a == _T_25[9:0]) begin
        image_2_410 <= io_pixelVal_in_2_3;
      end else if (10'h19a == _T_22[9:0]) begin
        image_2_410 <= io_pixelVal_in_2_2;
      end else if (10'h19a == _T_19[9:0]) begin
        image_2_410 <= io_pixelVal_in_2_1;
      end else if (10'h19a == _T_15[9:0]) begin
        image_2_410 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_411 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h19b == _T_37[9:0]) begin
        image_2_411 <= io_pixelVal_in_2_7;
      end else if (10'h19b == _T_34[9:0]) begin
        image_2_411 <= io_pixelVal_in_2_6;
      end else if (10'h19b == _T_31[9:0]) begin
        image_2_411 <= io_pixelVal_in_2_5;
      end else if (10'h19b == _T_28[9:0]) begin
        image_2_411 <= io_pixelVal_in_2_4;
      end else if (10'h19b == _T_25[9:0]) begin
        image_2_411 <= io_pixelVal_in_2_3;
      end else if (10'h19b == _T_22[9:0]) begin
        image_2_411 <= io_pixelVal_in_2_2;
      end else if (10'h19b == _T_19[9:0]) begin
        image_2_411 <= io_pixelVal_in_2_1;
      end else if (10'h19b == _T_15[9:0]) begin
        image_2_411 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_412 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h19c == _T_37[9:0]) begin
        image_2_412 <= io_pixelVal_in_2_7;
      end else if (10'h19c == _T_34[9:0]) begin
        image_2_412 <= io_pixelVal_in_2_6;
      end else if (10'h19c == _T_31[9:0]) begin
        image_2_412 <= io_pixelVal_in_2_5;
      end else if (10'h19c == _T_28[9:0]) begin
        image_2_412 <= io_pixelVal_in_2_4;
      end else if (10'h19c == _T_25[9:0]) begin
        image_2_412 <= io_pixelVal_in_2_3;
      end else if (10'h19c == _T_22[9:0]) begin
        image_2_412 <= io_pixelVal_in_2_2;
      end else if (10'h19c == _T_19[9:0]) begin
        image_2_412 <= io_pixelVal_in_2_1;
      end else if (10'h19c == _T_15[9:0]) begin
        image_2_412 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_413 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h19d == _T_37[9:0]) begin
        image_2_413 <= io_pixelVal_in_2_7;
      end else if (10'h19d == _T_34[9:0]) begin
        image_2_413 <= io_pixelVal_in_2_6;
      end else if (10'h19d == _T_31[9:0]) begin
        image_2_413 <= io_pixelVal_in_2_5;
      end else if (10'h19d == _T_28[9:0]) begin
        image_2_413 <= io_pixelVal_in_2_4;
      end else if (10'h19d == _T_25[9:0]) begin
        image_2_413 <= io_pixelVal_in_2_3;
      end else if (10'h19d == _T_22[9:0]) begin
        image_2_413 <= io_pixelVal_in_2_2;
      end else if (10'h19d == _T_19[9:0]) begin
        image_2_413 <= io_pixelVal_in_2_1;
      end else if (10'h19d == _T_15[9:0]) begin
        image_2_413 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_414 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h19e == _T_37[9:0]) begin
        image_2_414 <= io_pixelVal_in_2_7;
      end else if (10'h19e == _T_34[9:0]) begin
        image_2_414 <= io_pixelVal_in_2_6;
      end else if (10'h19e == _T_31[9:0]) begin
        image_2_414 <= io_pixelVal_in_2_5;
      end else if (10'h19e == _T_28[9:0]) begin
        image_2_414 <= io_pixelVal_in_2_4;
      end else if (10'h19e == _T_25[9:0]) begin
        image_2_414 <= io_pixelVal_in_2_3;
      end else if (10'h19e == _T_22[9:0]) begin
        image_2_414 <= io_pixelVal_in_2_2;
      end else if (10'h19e == _T_19[9:0]) begin
        image_2_414 <= io_pixelVal_in_2_1;
      end else if (10'h19e == _T_15[9:0]) begin
        image_2_414 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_415 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h19f == _T_37[9:0]) begin
        image_2_415 <= io_pixelVal_in_2_7;
      end else if (10'h19f == _T_34[9:0]) begin
        image_2_415 <= io_pixelVal_in_2_6;
      end else if (10'h19f == _T_31[9:0]) begin
        image_2_415 <= io_pixelVal_in_2_5;
      end else if (10'h19f == _T_28[9:0]) begin
        image_2_415 <= io_pixelVal_in_2_4;
      end else if (10'h19f == _T_25[9:0]) begin
        image_2_415 <= io_pixelVal_in_2_3;
      end else if (10'h19f == _T_22[9:0]) begin
        image_2_415 <= io_pixelVal_in_2_2;
      end else if (10'h19f == _T_19[9:0]) begin
        image_2_415 <= io_pixelVal_in_2_1;
      end else if (10'h19f == _T_15[9:0]) begin
        image_2_415 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_416 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a0 == _T_37[9:0]) begin
        image_2_416 <= io_pixelVal_in_2_7;
      end else if (10'h1a0 == _T_34[9:0]) begin
        image_2_416 <= io_pixelVal_in_2_6;
      end else if (10'h1a0 == _T_31[9:0]) begin
        image_2_416 <= io_pixelVal_in_2_5;
      end else if (10'h1a0 == _T_28[9:0]) begin
        image_2_416 <= io_pixelVal_in_2_4;
      end else if (10'h1a0 == _T_25[9:0]) begin
        image_2_416 <= io_pixelVal_in_2_3;
      end else if (10'h1a0 == _T_22[9:0]) begin
        image_2_416 <= io_pixelVal_in_2_2;
      end else if (10'h1a0 == _T_19[9:0]) begin
        image_2_416 <= io_pixelVal_in_2_1;
      end else if (10'h1a0 == _T_15[9:0]) begin
        image_2_416 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_417 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a1 == _T_37[9:0]) begin
        image_2_417 <= io_pixelVal_in_2_7;
      end else if (10'h1a1 == _T_34[9:0]) begin
        image_2_417 <= io_pixelVal_in_2_6;
      end else if (10'h1a1 == _T_31[9:0]) begin
        image_2_417 <= io_pixelVal_in_2_5;
      end else if (10'h1a1 == _T_28[9:0]) begin
        image_2_417 <= io_pixelVal_in_2_4;
      end else if (10'h1a1 == _T_25[9:0]) begin
        image_2_417 <= io_pixelVal_in_2_3;
      end else if (10'h1a1 == _T_22[9:0]) begin
        image_2_417 <= io_pixelVal_in_2_2;
      end else if (10'h1a1 == _T_19[9:0]) begin
        image_2_417 <= io_pixelVal_in_2_1;
      end else if (10'h1a1 == _T_15[9:0]) begin
        image_2_417 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_418 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a2 == _T_37[9:0]) begin
        image_2_418 <= io_pixelVal_in_2_7;
      end else if (10'h1a2 == _T_34[9:0]) begin
        image_2_418 <= io_pixelVal_in_2_6;
      end else if (10'h1a2 == _T_31[9:0]) begin
        image_2_418 <= io_pixelVal_in_2_5;
      end else if (10'h1a2 == _T_28[9:0]) begin
        image_2_418 <= io_pixelVal_in_2_4;
      end else if (10'h1a2 == _T_25[9:0]) begin
        image_2_418 <= io_pixelVal_in_2_3;
      end else if (10'h1a2 == _T_22[9:0]) begin
        image_2_418 <= io_pixelVal_in_2_2;
      end else if (10'h1a2 == _T_19[9:0]) begin
        image_2_418 <= io_pixelVal_in_2_1;
      end else if (10'h1a2 == _T_15[9:0]) begin
        image_2_418 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_419 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a3 == _T_37[9:0]) begin
        image_2_419 <= io_pixelVal_in_2_7;
      end else if (10'h1a3 == _T_34[9:0]) begin
        image_2_419 <= io_pixelVal_in_2_6;
      end else if (10'h1a3 == _T_31[9:0]) begin
        image_2_419 <= io_pixelVal_in_2_5;
      end else if (10'h1a3 == _T_28[9:0]) begin
        image_2_419 <= io_pixelVal_in_2_4;
      end else if (10'h1a3 == _T_25[9:0]) begin
        image_2_419 <= io_pixelVal_in_2_3;
      end else if (10'h1a3 == _T_22[9:0]) begin
        image_2_419 <= io_pixelVal_in_2_2;
      end else if (10'h1a3 == _T_19[9:0]) begin
        image_2_419 <= io_pixelVal_in_2_1;
      end else if (10'h1a3 == _T_15[9:0]) begin
        image_2_419 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_420 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a4 == _T_37[9:0]) begin
        image_2_420 <= io_pixelVal_in_2_7;
      end else if (10'h1a4 == _T_34[9:0]) begin
        image_2_420 <= io_pixelVal_in_2_6;
      end else if (10'h1a4 == _T_31[9:0]) begin
        image_2_420 <= io_pixelVal_in_2_5;
      end else if (10'h1a4 == _T_28[9:0]) begin
        image_2_420 <= io_pixelVal_in_2_4;
      end else if (10'h1a4 == _T_25[9:0]) begin
        image_2_420 <= io_pixelVal_in_2_3;
      end else if (10'h1a4 == _T_22[9:0]) begin
        image_2_420 <= io_pixelVal_in_2_2;
      end else if (10'h1a4 == _T_19[9:0]) begin
        image_2_420 <= io_pixelVal_in_2_1;
      end else if (10'h1a4 == _T_15[9:0]) begin
        image_2_420 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_421 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a5 == _T_37[9:0]) begin
        image_2_421 <= io_pixelVal_in_2_7;
      end else if (10'h1a5 == _T_34[9:0]) begin
        image_2_421 <= io_pixelVal_in_2_6;
      end else if (10'h1a5 == _T_31[9:0]) begin
        image_2_421 <= io_pixelVal_in_2_5;
      end else if (10'h1a5 == _T_28[9:0]) begin
        image_2_421 <= io_pixelVal_in_2_4;
      end else if (10'h1a5 == _T_25[9:0]) begin
        image_2_421 <= io_pixelVal_in_2_3;
      end else if (10'h1a5 == _T_22[9:0]) begin
        image_2_421 <= io_pixelVal_in_2_2;
      end else if (10'h1a5 == _T_19[9:0]) begin
        image_2_421 <= io_pixelVal_in_2_1;
      end else if (10'h1a5 == _T_15[9:0]) begin
        image_2_421 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_422 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a6 == _T_37[9:0]) begin
        image_2_422 <= io_pixelVal_in_2_7;
      end else if (10'h1a6 == _T_34[9:0]) begin
        image_2_422 <= io_pixelVal_in_2_6;
      end else if (10'h1a6 == _T_31[9:0]) begin
        image_2_422 <= io_pixelVal_in_2_5;
      end else if (10'h1a6 == _T_28[9:0]) begin
        image_2_422 <= io_pixelVal_in_2_4;
      end else if (10'h1a6 == _T_25[9:0]) begin
        image_2_422 <= io_pixelVal_in_2_3;
      end else if (10'h1a6 == _T_22[9:0]) begin
        image_2_422 <= io_pixelVal_in_2_2;
      end else if (10'h1a6 == _T_19[9:0]) begin
        image_2_422 <= io_pixelVal_in_2_1;
      end else if (10'h1a6 == _T_15[9:0]) begin
        image_2_422 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_423 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a7 == _T_37[9:0]) begin
        image_2_423 <= io_pixelVal_in_2_7;
      end else if (10'h1a7 == _T_34[9:0]) begin
        image_2_423 <= io_pixelVal_in_2_6;
      end else if (10'h1a7 == _T_31[9:0]) begin
        image_2_423 <= io_pixelVal_in_2_5;
      end else if (10'h1a7 == _T_28[9:0]) begin
        image_2_423 <= io_pixelVal_in_2_4;
      end else if (10'h1a7 == _T_25[9:0]) begin
        image_2_423 <= io_pixelVal_in_2_3;
      end else if (10'h1a7 == _T_22[9:0]) begin
        image_2_423 <= io_pixelVal_in_2_2;
      end else if (10'h1a7 == _T_19[9:0]) begin
        image_2_423 <= io_pixelVal_in_2_1;
      end else if (10'h1a7 == _T_15[9:0]) begin
        image_2_423 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_424 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a8 == _T_37[9:0]) begin
        image_2_424 <= io_pixelVal_in_2_7;
      end else if (10'h1a8 == _T_34[9:0]) begin
        image_2_424 <= io_pixelVal_in_2_6;
      end else if (10'h1a8 == _T_31[9:0]) begin
        image_2_424 <= io_pixelVal_in_2_5;
      end else if (10'h1a8 == _T_28[9:0]) begin
        image_2_424 <= io_pixelVal_in_2_4;
      end else if (10'h1a8 == _T_25[9:0]) begin
        image_2_424 <= io_pixelVal_in_2_3;
      end else if (10'h1a8 == _T_22[9:0]) begin
        image_2_424 <= io_pixelVal_in_2_2;
      end else if (10'h1a8 == _T_19[9:0]) begin
        image_2_424 <= io_pixelVal_in_2_1;
      end else if (10'h1a8 == _T_15[9:0]) begin
        image_2_424 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_425 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1a9 == _T_37[9:0]) begin
        image_2_425 <= io_pixelVal_in_2_7;
      end else if (10'h1a9 == _T_34[9:0]) begin
        image_2_425 <= io_pixelVal_in_2_6;
      end else if (10'h1a9 == _T_31[9:0]) begin
        image_2_425 <= io_pixelVal_in_2_5;
      end else if (10'h1a9 == _T_28[9:0]) begin
        image_2_425 <= io_pixelVal_in_2_4;
      end else if (10'h1a9 == _T_25[9:0]) begin
        image_2_425 <= io_pixelVal_in_2_3;
      end else if (10'h1a9 == _T_22[9:0]) begin
        image_2_425 <= io_pixelVal_in_2_2;
      end else if (10'h1a9 == _T_19[9:0]) begin
        image_2_425 <= io_pixelVal_in_2_1;
      end else if (10'h1a9 == _T_15[9:0]) begin
        image_2_425 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_426 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1aa == _T_37[9:0]) begin
        image_2_426 <= io_pixelVal_in_2_7;
      end else if (10'h1aa == _T_34[9:0]) begin
        image_2_426 <= io_pixelVal_in_2_6;
      end else if (10'h1aa == _T_31[9:0]) begin
        image_2_426 <= io_pixelVal_in_2_5;
      end else if (10'h1aa == _T_28[9:0]) begin
        image_2_426 <= io_pixelVal_in_2_4;
      end else if (10'h1aa == _T_25[9:0]) begin
        image_2_426 <= io_pixelVal_in_2_3;
      end else if (10'h1aa == _T_22[9:0]) begin
        image_2_426 <= io_pixelVal_in_2_2;
      end else if (10'h1aa == _T_19[9:0]) begin
        image_2_426 <= io_pixelVal_in_2_1;
      end else if (10'h1aa == _T_15[9:0]) begin
        image_2_426 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_427 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ab == _T_37[9:0]) begin
        image_2_427 <= io_pixelVal_in_2_7;
      end else if (10'h1ab == _T_34[9:0]) begin
        image_2_427 <= io_pixelVal_in_2_6;
      end else if (10'h1ab == _T_31[9:0]) begin
        image_2_427 <= io_pixelVal_in_2_5;
      end else if (10'h1ab == _T_28[9:0]) begin
        image_2_427 <= io_pixelVal_in_2_4;
      end else if (10'h1ab == _T_25[9:0]) begin
        image_2_427 <= io_pixelVal_in_2_3;
      end else if (10'h1ab == _T_22[9:0]) begin
        image_2_427 <= io_pixelVal_in_2_2;
      end else if (10'h1ab == _T_19[9:0]) begin
        image_2_427 <= io_pixelVal_in_2_1;
      end else if (10'h1ab == _T_15[9:0]) begin
        image_2_427 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_428 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ac == _T_37[9:0]) begin
        image_2_428 <= io_pixelVal_in_2_7;
      end else if (10'h1ac == _T_34[9:0]) begin
        image_2_428 <= io_pixelVal_in_2_6;
      end else if (10'h1ac == _T_31[9:0]) begin
        image_2_428 <= io_pixelVal_in_2_5;
      end else if (10'h1ac == _T_28[9:0]) begin
        image_2_428 <= io_pixelVal_in_2_4;
      end else if (10'h1ac == _T_25[9:0]) begin
        image_2_428 <= io_pixelVal_in_2_3;
      end else if (10'h1ac == _T_22[9:0]) begin
        image_2_428 <= io_pixelVal_in_2_2;
      end else if (10'h1ac == _T_19[9:0]) begin
        image_2_428 <= io_pixelVal_in_2_1;
      end else if (10'h1ac == _T_15[9:0]) begin
        image_2_428 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_429 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ad == _T_37[9:0]) begin
        image_2_429 <= io_pixelVal_in_2_7;
      end else if (10'h1ad == _T_34[9:0]) begin
        image_2_429 <= io_pixelVal_in_2_6;
      end else if (10'h1ad == _T_31[9:0]) begin
        image_2_429 <= io_pixelVal_in_2_5;
      end else if (10'h1ad == _T_28[9:0]) begin
        image_2_429 <= io_pixelVal_in_2_4;
      end else if (10'h1ad == _T_25[9:0]) begin
        image_2_429 <= io_pixelVal_in_2_3;
      end else if (10'h1ad == _T_22[9:0]) begin
        image_2_429 <= io_pixelVal_in_2_2;
      end else if (10'h1ad == _T_19[9:0]) begin
        image_2_429 <= io_pixelVal_in_2_1;
      end else if (10'h1ad == _T_15[9:0]) begin
        image_2_429 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_430 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ae == _T_37[9:0]) begin
        image_2_430 <= io_pixelVal_in_2_7;
      end else if (10'h1ae == _T_34[9:0]) begin
        image_2_430 <= io_pixelVal_in_2_6;
      end else if (10'h1ae == _T_31[9:0]) begin
        image_2_430 <= io_pixelVal_in_2_5;
      end else if (10'h1ae == _T_28[9:0]) begin
        image_2_430 <= io_pixelVal_in_2_4;
      end else if (10'h1ae == _T_25[9:0]) begin
        image_2_430 <= io_pixelVal_in_2_3;
      end else if (10'h1ae == _T_22[9:0]) begin
        image_2_430 <= io_pixelVal_in_2_2;
      end else if (10'h1ae == _T_19[9:0]) begin
        image_2_430 <= io_pixelVal_in_2_1;
      end else if (10'h1ae == _T_15[9:0]) begin
        image_2_430 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_431 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1af == _T_37[9:0]) begin
        image_2_431 <= io_pixelVal_in_2_7;
      end else if (10'h1af == _T_34[9:0]) begin
        image_2_431 <= io_pixelVal_in_2_6;
      end else if (10'h1af == _T_31[9:0]) begin
        image_2_431 <= io_pixelVal_in_2_5;
      end else if (10'h1af == _T_28[9:0]) begin
        image_2_431 <= io_pixelVal_in_2_4;
      end else if (10'h1af == _T_25[9:0]) begin
        image_2_431 <= io_pixelVal_in_2_3;
      end else if (10'h1af == _T_22[9:0]) begin
        image_2_431 <= io_pixelVal_in_2_2;
      end else if (10'h1af == _T_19[9:0]) begin
        image_2_431 <= io_pixelVal_in_2_1;
      end else if (10'h1af == _T_15[9:0]) begin
        image_2_431 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_432 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b0 == _T_37[9:0]) begin
        image_2_432 <= io_pixelVal_in_2_7;
      end else if (10'h1b0 == _T_34[9:0]) begin
        image_2_432 <= io_pixelVal_in_2_6;
      end else if (10'h1b0 == _T_31[9:0]) begin
        image_2_432 <= io_pixelVal_in_2_5;
      end else if (10'h1b0 == _T_28[9:0]) begin
        image_2_432 <= io_pixelVal_in_2_4;
      end else if (10'h1b0 == _T_25[9:0]) begin
        image_2_432 <= io_pixelVal_in_2_3;
      end else if (10'h1b0 == _T_22[9:0]) begin
        image_2_432 <= io_pixelVal_in_2_2;
      end else if (10'h1b0 == _T_19[9:0]) begin
        image_2_432 <= io_pixelVal_in_2_1;
      end else if (10'h1b0 == _T_15[9:0]) begin
        image_2_432 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_433 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b1 == _T_37[9:0]) begin
        image_2_433 <= io_pixelVal_in_2_7;
      end else if (10'h1b1 == _T_34[9:0]) begin
        image_2_433 <= io_pixelVal_in_2_6;
      end else if (10'h1b1 == _T_31[9:0]) begin
        image_2_433 <= io_pixelVal_in_2_5;
      end else if (10'h1b1 == _T_28[9:0]) begin
        image_2_433 <= io_pixelVal_in_2_4;
      end else if (10'h1b1 == _T_25[9:0]) begin
        image_2_433 <= io_pixelVal_in_2_3;
      end else if (10'h1b1 == _T_22[9:0]) begin
        image_2_433 <= io_pixelVal_in_2_2;
      end else if (10'h1b1 == _T_19[9:0]) begin
        image_2_433 <= io_pixelVal_in_2_1;
      end else if (10'h1b1 == _T_15[9:0]) begin
        image_2_433 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_434 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b2 == _T_37[9:0]) begin
        image_2_434 <= io_pixelVal_in_2_7;
      end else if (10'h1b2 == _T_34[9:0]) begin
        image_2_434 <= io_pixelVal_in_2_6;
      end else if (10'h1b2 == _T_31[9:0]) begin
        image_2_434 <= io_pixelVal_in_2_5;
      end else if (10'h1b2 == _T_28[9:0]) begin
        image_2_434 <= io_pixelVal_in_2_4;
      end else if (10'h1b2 == _T_25[9:0]) begin
        image_2_434 <= io_pixelVal_in_2_3;
      end else if (10'h1b2 == _T_22[9:0]) begin
        image_2_434 <= io_pixelVal_in_2_2;
      end else if (10'h1b2 == _T_19[9:0]) begin
        image_2_434 <= io_pixelVal_in_2_1;
      end else if (10'h1b2 == _T_15[9:0]) begin
        image_2_434 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_435 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b3 == _T_37[9:0]) begin
        image_2_435 <= io_pixelVal_in_2_7;
      end else if (10'h1b3 == _T_34[9:0]) begin
        image_2_435 <= io_pixelVal_in_2_6;
      end else if (10'h1b3 == _T_31[9:0]) begin
        image_2_435 <= io_pixelVal_in_2_5;
      end else if (10'h1b3 == _T_28[9:0]) begin
        image_2_435 <= io_pixelVal_in_2_4;
      end else if (10'h1b3 == _T_25[9:0]) begin
        image_2_435 <= io_pixelVal_in_2_3;
      end else if (10'h1b3 == _T_22[9:0]) begin
        image_2_435 <= io_pixelVal_in_2_2;
      end else if (10'h1b3 == _T_19[9:0]) begin
        image_2_435 <= io_pixelVal_in_2_1;
      end else if (10'h1b3 == _T_15[9:0]) begin
        image_2_435 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_436 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b4 == _T_37[9:0]) begin
        image_2_436 <= io_pixelVal_in_2_7;
      end else if (10'h1b4 == _T_34[9:0]) begin
        image_2_436 <= io_pixelVal_in_2_6;
      end else if (10'h1b4 == _T_31[9:0]) begin
        image_2_436 <= io_pixelVal_in_2_5;
      end else if (10'h1b4 == _T_28[9:0]) begin
        image_2_436 <= io_pixelVal_in_2_4;
      end else if (10'h1b4 == _T_25[9:0]) begin
        image_2_436 <= io_pixelVal_in_2_3;
      end else if (10'h1b4 == _T_22[9:0]) begin
        image_2_436 <= io_pixelVal_in_2_2;
      end else if (10'h1b4 == _T_19[9:0]) begin
        image_2_436 <= io_pixelVal_in_2_1;
      end else if (10'h1b4 == _T_15[9:0]) begin
        image_2_436 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_437 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b5 == _T_37[9:0]) begin
        image_2_437 <= io_pixelVal_in_2_7;
      end else if (10'h1b5 == _T_34[9:0]) begin
        image_2_437 <= io_pixelVal_in_2_6;
      end else if (10'h1b5 == _T_31[9:0]) begin
        image_2_437 <= io_pixelVal_in_2_5;
      end else if (10'h1b5 == _T_28[9:0]) begin
        image_2_437 <= io_pixelVal_in_2_4;
      end else if (10'h1b5 == _T_25[9:0]) begin
        image_2_437 <= io_pixelVal_in_2_3;
      end else if (10'h1b5 == _T_22[9:0]) begin
        image_2_437 <= io_pixelVal_in_2_2;
      end else if (10'h1b5 == _T_19[9:0]) begin
        image_2_437 <= io_pixelVal_in_2_1;
      end else if (10'h1b5 == _T_15[9:0]) begin
        image_2_437 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_438 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b6 == _T_37[9:0]) begin
        image_2_438 <= io_pixelVal_in_2_7;
      end else if (10'h1b6 == _T_34[9:0]) begin
        image_2_438 <= io_pixelVal_in_2_6;
      end else if (10'h1b6 == _T_31[9:0]) begin
        image_2_438 <= io_pixelVal_in_2_5;
      end else if (10'h1b6 == _T_28[9:0]) begin
        image_2_438 <= io_pixelVal_in_2_4;
      end else if (10'h1b6 == _T_25[9:0]) begin
        image_2_438 <= io_pixelVal_in_2_3;
      end else if (10'h1b6 == _T_22[9:0]) begin
        image_2_438 <= io_pixelVal_in_2_2;
      end else if (10'h1b6 == _T_19[9:0]) begin
        image_2_438 <= io_pixelVal_in_2_1;
      end else if (10'h1b6 == _T_15[9:0]) begin
        image_2_438 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_439 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b7 == _T_37[9:0]) begin
        image_2_439 <= io_pixelVal_in_2_7;
      end else if (10'h1b7 == _T_34[9:0]) begin
        image_2_439 <= io_pixelVal_in_2_6;
      end else if (10'h1b7 == _T_31[9:0]) begin
        image_2_439 <= io_pixelVal_in_2_5;
      end else if (10'h1b7 == _T_28[9:0]) begin
        image_2_439 <= io_pixelVal_in_2_4;
      end else if (10'h1b7 == _T_25[9:0]) begin
        image_2_439 <= io_pixelVal_in_2_3;
      end else if (10'h1b7 == _T_22[9:0]) begin
        image_2_439 <= io_pixelVal_in_2_2;
      end else if (10'h1b7 == _T_19[9:0]) begin
        image_2_439 <= io_pixelVal_in_2_1;
      end else if (10'h1b7 == _T_15[9:0]) begin
        image_2_439 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_440 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b8 == _T_37[9:0]) begin
        image_2_440 <= io_pixelVal_in_2_7;
      end else if (10'h1b8 == _T_34[9:0]) begin
        image_2_440 <= io_pixelVal_in_2_6;
      end else if (10'h1b8 == _T_31[9:0]) begin
        image_2_440 <= io_pixelVal_in_2_5;
      end else if (10'h1b8 == _T_28[9:0]) begin
        image_2_440 <= io_pixelVal_in_2_4;
      end else if (10'h1b8 == _T_25[9:0]) begin
        image_2_440 <= io_pixelVal_in_2_3;
      end else if (10'h1b8 == _T_22[9:0]) begin
        image_2_440 <= io_pixelVal_in_2_2;
      end else if (10'h1b8 == _T_19[9:0]) begin
        image_2_440 <= io_pixelVal_in_2_1;
      end else if (10'h1b8 == _T_15[9:0]) begin
        image_2_440 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_441 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1b9 == _T_37[9:0]) begin
        image_2_441 <= io_pixelVal_in_2_7;
      end else if (10'h1b9 == _T_34[9:0]) begin
        image_2_441 <= io_pixelVal_in_2_6;
      end else if (10'h1b9 == _T_31[9:0]) begin
        image_2_441 <= io_pixelVal_in_2_5;
      end else if (10'h1b9 == _T_28[9:0]) begin
        image_2_441 <= io_pixelVal_in_2_4;
      end else if (10'h1b9 == _T_25[9:0]) begin
        image_2_441 <= io_pixelVal_in_2_3;
      end else if (10'h1b9 == _T_22[9:0]) begin
        image_2_441 <= io_pixelVal_in_2_2;
      end else if (10'h1b9 == _T_19[9:0]) begin
        image_2_441 <= io_pixelVal_in_2_1;
      end else if (10'h1b9 == _T_15[9:0]) begin
        image_2_441 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_442 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ba == _T_37[9:0]) begin
        image_2_442 <= io_pixelVal_in_2_7;
      end else if (10'h1ba == _T_34[9:0]) begin
        image_2_442 <= io_pixelVal_in_2_6;
      end else if (10'h1ba == _T_31[9:0]) begin
        image_2_442 <= io_pixelVal_in_2_5;
      end else if (10'h1ba == _T_28[9:0]) begin
        image_2_442 <= io_pixelVal_in_2_4;
      end else if (10'h1ba == _T_25[9:0]) begin
        image_2_442 <= io_pixelVal_in_2_3;
      end else if (10'h1ba == _T_22[9:0]) begin
        image_2_442 <= io_pixelVal_in_2_2;
      end else if (10'h1ba == _T_19[9:0]) begin
        image_2_442 <= io_pixelVal_in_2_1;
      end else if (10'h1ba == _T_15[9:0]) begin
        image_2_442 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_443 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1bb == _T_37[9:0]) begin
        image_2_443 <= io_pixelVal_in_2_7;
      end else if (10'h1bb == _T_34[9:0]) begin
        image_2_443 <= io_pixelVal_in_2_6;
      end else if (10'h1bb == _T_31[9:0]) begin
        image_2_443 <= io_pixelVal_in_2_5;
      end else if (10'h1bb == _T_28[9:0]) begin
        image_2_443 <= io_pixelVal_in_2_4;
      end else if (10'h1bb == _T_25[9:0]) begin
        image_2_443 <= io_pixelVal_in_2_3;
      end else if (10'h1bb == _T_22[9:0]) begin
        image_2_443 <= io_pixelVal_in_2_2;
      end else if (10'h1bb == _T_19[9:0]) begin
        image_2_443 <= io_pixelVal_in_2_1;
      end else if (10'h1bb == _T_15[9:0]) begin
        image_2_443 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_444 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1bc == _T_37[9:0]) begin
        image_2_444 <= io_pixelVal_in_2_7;
      end else if (10'h1bc == _T_34[9:0]) begin
        image_2_444 <= io_pixelVal_in_2_6;
      end else if (10'h1bc == _T_31[9:0]) begin
        image_2_444 <= io_pixelVal_in_2_5;
      end else if (10'h1bc == _T_28[9:0]) begin
        image_2_444 <= io_pixelVal_in_2_4;
      end else if (10'h1bc == _T_25[9:0]) begin
        image_2_444 <= io_pixelVal_in_2_3;
      end else if (10'h1bc == _T_22[9:0]) begin
        image_2_444 <= io_pixelVal_in_2_2;
      end else if (10'h1bc == _T_19[9:0]) begin
        image_2_444 <= io_pixelVal_in_2_1;
      end else if (10'h1bc == _T_15[9:0]) begin
        image_2_444 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_445 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1bd == _T_37[9:0]) begin
        image_2_445 <= io_pixelVal_in_2_7;
      end else if (10'h1bd == _T_34[9:0]) begin
        image_2_445 <= io_pixelVal_in_2_6;
      end else if (10'h1bd == _T_31[9:0]) begin
        image_2_445 <= io_pixelVal_in_2_5;
      end else if (10'h1bd == _T_28[9:0]) begin
        image_2_445 <= io_pixelVal_in_2_4;
      end else if (10'h1bd == _T_25[9:0]) begin
        image_2_445 <= io_pixelVal_in_2_3;
      end else if (10'h1bd == _T_22[9:0]) begin
        image_2_445 <= io_pixelVal_in_2_2;
      end else if (10'h1bd == _T_19[9:0]) begin
        image_2_445 <= io_pixelVal_in_2_1;
      end else if (10'h1bd == _T_15[9:0]) begin
        image_2_445 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_446 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1be == _T_37[9:0]) begin
        image_2_446 <= io_pixelVal_in_2_7;
      end else if (10'h1be == _T_34[9:0]) begin
        image_2_446 <= io_pixelVal_in_2_6;
      end else if (10'h1be == _T_31[9:0]) begin
        image_2_446 <= io_pixelVal_in_2_5;
      end else if (10'h1be == _T_28[9:0]) begin
        image_2_446 <= io_pixelVal_in_2_4;
      end else if (10'h1be == _T_25[9:0]) begin
        image_2_446 <= io_pixelVal_in_2_3;
      end else if (10'h1be == _T_22[9:0]) begin
        image_2_446 <= io_pixelVal_in_2_2;
      end else if (10'h1be == _T_19[9:0]) begin
        image_2_446 <= io_pixelVal_in_2_1;
      end else if (10'h1be == _T_15[9:0]) begin
        image_2_446 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_447 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1bf == _T_37[9:0]) begin
        image_2_447 <= io_pixelVal_in_2_7;
      end else if (10'h1bf == _T_34[9:0]) begin
        image_2_447 <= io_pixelVal_in_2_6;
      end else if (10'h1bf == _T_31[9:0]) begin
        image_2_447 <= io_pixelVal_in_2_5;
      end else if (10'h1bf == _T_28[9:0]) begin
        image_2_447 <= io_pixelVal_in_2_4;
      end else if (10'h1bf == _T_25[9:0]) begin
        image_2_447 <= io_pixelVal_in_2_3;
      end else if (10'h1bf == _T_22[9:0]) begin
        image_2_447 <= io_pixelVal_in_2_2;
      end else if (10'h1bf == _T_19[9:0]) begin
        image_2_447 <= io_pixelVal_in_2_1;
      end else if (10'h1bf == _T_15[9:0]) begin
        image_2_447 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_448 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c0 == _T_37[9:0]) begin
        image_2_448 <= io_pixelVal_in_2_7;
      end else if (10'h1c0 == _T_34[9:0]) begin
        image_2_448 <= io_pixelVal_in_2_6;
      end else if (10'h1c0 == _T_31[9:0]) begin
        image_2_448 <= io_pixelVal_in_2_5;
      end else if (10'h1c0 == _T_28[9:0]) begin
        image_2_448 <= io_pixelVal_in_2_4;
      end else if (10'h1c0 == _T_25[9:0]) begin
        image_2_448 <= io_pixelVal_in_2_3;
      end else if (10'h1c0 == _T_22[9:0]) begin
        image_2_448 <= io_pixelVal_in_2_2;
      end else if (10'h1c0 == _T_19[9:0]) begin
        image_2_448 <= io_pixelVal_in_2_1;
      end else if (10'h1c0 == _T_15[9:0]) begin
        image_2_448 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_449 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c1 == _T_37[9:0]) begin
        image_2_449 <= io_pixelVal_in_2_7;
      end else if (10'h1c1 == _T_34[9:0]) begin
        image_2_449 <= io_pixelVal_in_2_6;
      end else if (10'h1c1 == _T_31[9:0]) begin
        image_2_449 <= io_pixelVal_in_2_5;
      end else if (10'h1c1 == _T_28[9:0]) begin
        image_2_449 <= io_pixelVal_in_2_4;
      end else if (10'h1c1 == _T_25[9:0]) begin
        image_2_449 <= io_pixelVal_in_2_3;
      end else if (10'h1c1 == _T_22[9:0]) begin
        image_2_449 <= io_pixelVal_in_2_2;
      end else if (10'h1c1 == _T_19[9:0]) begin
        image_2_449 <= io_pixelVal_in_2_1;
      end else if (10'h1c1 == _T_15[9:0]) begin
        image_2_449 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_450 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c2 == _T_37[9:0]) begin
        image_2_450 <= io_pixelVal_in_2_7;
      end else if (10'h1c2 == _T_34[9:0]) begin
        image_2_450 <= io_pixelVal_in_2_6;
      end else if (10'h1c2 == _T_31[9:0]) begin
        image_2_450 <= io_pixelVal_in_2_5;
      end else if (10'h1c2 == _T_28[9:0]) begin
        image_2_450 <= io_pixelVal_in_2_4;
      end else if (10'h1c2 == _T_25[9:0]) begin
        image_2_450 <= io_pixelVal_in_2_3;
      end else if (10'h1c2 == _T_22[9:0]) begin
        image_2_450 <= io_pixelVal_in_2_2;
      end else if (10'h1c2 == _T_19[9:0]) begin
        image_2_450 <= io_pixelVal_in_2_1;
      end else if (10'h1c2 == _T_15[9:0]) begin
        image_2_450 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_451 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c3 == _T_37[9:0]) begin
        image_2_451 <= io_pixelVal_in_2_7;
      end else if (10'h1c3 == _T_34[9:0]) begin
        image_2_451 <= io_pixelVal_in_2_6;
      end else if (10'h1c3 == _T_31[9:0]) begin
        image_2_451 <= io_pixelVal_in_2_5;
      end else if (10'h1c3 == _T_28[9:0]) begin
        image_2_451 <= io_pixelVal_in_2_4;
      end else if (10'h1c3 == _T_25[9:0]) begin
        image_2_451 <= io_pixelVal_in_2_3;
      end else if (10'h1c3 == _T_22[9:0]) begin
        image_2_451 <= io_pixelVal_in_2_2;
      end else if (10'h1c3 == _T_19[9:0]) begin
        image_2_451 <= io_pixelVal_in_2_1;
      end else if (10'h1c3 == _T_15[9:0]) begin
        image_2_451 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_452 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c4 == _T_37[9:0]) begin
        image_2_452 <= io_pixelVal_in_2_7;
      end else if (10'h1c4 == _T_34[9:0]) begin
        image_2_452 <= io_pixelVal_in_2_6;
      end else if (10'h1c4 == _T_31[9:0]) begin
        image_2_452 <= io_pixelVal_in_2_5;
      end else if (10'h1c4 == _T_28[9:0]) begin
        image_2_452 <= io_pixelVal_in_2_4;
      end else if (10'h1c4 == _T_25[9:0]) begin
        image_2_452 <= io_pixelVal_in_2_3;
      end else if (10'h1c4 == _T_22[9:0]) begin
        image_2_452 <= io_pixelVal_in_2_2;
      end else if (10'h1c4 == _T_19[9:0]) begin
        image_2_452 <= io_pixelVal_in_2_1;
      end else if (10'h1c4 == _T_15[9:0]) begin
        image_2_452 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_453 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c5 == _T_37[9:0]) begin
        image_2_453 <= io_pixelVal_in_2_7;
      end else if (10'h1c5 == _T_34[9:0]) begin
        image_2_453 <= io_pixelVal_in_2_6;
      end else if (10'h1c5 == _T_31[9:0]) begin
        image_2_453 <= io_pixelVal_in_2_5;
      end else if (10'h1c5 == _T_28[9:0]) begin
        image_2_453 <= io_pixelVal_in_2_4;
      end else if (10'h1c5 == _T_25[9:0]) begin
        image_2_453 <= io_pixelVal_in_2_3;
      end else if (10'h1c5 == _T_22[9:0]) begin
        image_2_453 <= io_pixelVal_in_2_2;
      end else if (10'h1c5 == _T_19[9:0]) begin
        image_2_453 <= io_pixelVal_in_2_1;
      end else if (10'h1c5 == _T_15[9:0]) begin
        image_2_453 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_454 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c6 == _T_37[9:0]) begin
        image_2_454 <= io_pixelVal_in_2_7;
      end else if (10'h1c6 == _T_34[9:0]) begin
        image_2_454 <= io_pixelVal_in_2_6;
      end else if (10'h1c6 == _T_31[9:0]) begin
        image_2_454 <= io_pixelVal_in_2_5;
      end else if (10'h1c6 == _T_28[9:0]) begin
        image_2_454 <= io_pixelVal_in_2_4;
      end else if (10'h1c6 == _T_25[9:0]) begin
        image_2_454 <= io_pixelVal_in_2_3;
      end else if (10'h1c6 == _T_22[9:0]) begin
        image_2_454 <= io_pixelVal_in_2_2;
      end else if (10'h1c6 == _T_19[9:0]) begin
        image_2_454 <= io_pixelVal_in_2_1;
      end else if (10'h1c6 == _T_15[9:0]) begin
        image_2_454 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_455 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c7 == _T_37[9:0]) begin
        image_2_455 <= io_pixelVal_in_2_7;
      end else if (10'h1c7 == _T_34[9:0]) begin
        image_2_455 <= io_pixelVal_in_2_6;
      end else if (10'h1c7 == _T_31[9:0]) begin
        image_2_455 <= io_pixelVal_in_2_5;
      end else if (10'h1c7 == _T_28[9:0]) begin
        image_2_455 <= io_pixelVal_in_2_4;
      end else if (10'h1c7 == _T_25[9:0]) begin
        image_2_455 <= io_pixelVal_in_2_3;
      end else if (10'h1c7 == _T_22[9:0]) begin
        image_2_455 <= io_pixelVal_in_2_2;
      end else if (10'h1c7 == _T_19[9:0]) begin
        image_2_455 <= io_pixelVal_in_2_1;
      end else if (10'h1c7 == _T_15[9:0]) begin
        image_2_455 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_456 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c8 == _T_37[9:0]) begin
        image_2_456 <= io_pixelVal_in_2_7;
      end else if (10'h1c8 == _T_34[9:0]) begin
        image_2_456 <= io_pixelVal_in_2_6;
      end else if (10'h1c8 == _T_31[9:0]) begin
        image_2_456 <= io_pixelVal_in_2_5;
      end else if (10'h1c8 == _T_28[9:0]) begin
        image_2_456 <= io_pixelVal_in_2_4;
      end else if (10'h1c8 == _T_25[9:0]) begin
        image_2_456 <= io_pixelVal_in_2_3;
      end else if (10'h1c8 == _T_22[9:0]) begin
        image_2_456 <= io_pixelVal_in_2_2;
      end else if (10'h1c8 == _T_19[9:0]) begin
        image_2_456 <= io_pixelVal_in_2_1;
      end else if (10'h1c8 == _T_15[9:0]) begin
        image_2_456 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_457 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1c9 == _T_37[9:0]) begin
        image_2_457 <= io_pixelVal_in_2_7;
      end else if (10'h1c9 == _T_34[9:0]) begin
        image_2_457 <= io_pixelVal_in_2_6;
      end else if (10'h1c9 == _T_31[9:0]) begin
        image_2_457 <= io_pixelVal_in_2_5;
      end else if (10'h1c9 == _T_28[9:0]) begin
        image_2_457 <= io_pixelVal_in_2_4;
      end else if (10'h1c9 == _T_25[9:0]) begin
        image_2_457 <= io_pixelVal_in_2_3;
      end else if (10'h1c9 == _T_22[9:0]) begin
        image_2_457 <= io_pixelVal_in_2_2;
      end else if (10'h1c9 == _T_19[9:0]) begin
        image_2_457 <= io_pixelVal_in_2_1;
      end else if (10'h1c9 == _T_15[9:0]) begin
        image_2_457 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_458 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ca == _T_37[9:0]) begin
        image_2_458 <= io_pixelVal_in_2_7;
      end else if (10'h1ca == _T_34[9:0]) begin
        image_2_458 <= io_pixelVal_in_2_6;
      end else if (10'h1ca == _T_31[9:0]) begin
        image_2_458 <= io_pixelVal_in_2_5;
      end else if (10'h1ca == _T_28[9:0]) begin
        image_2_458 <= io_pixelVal_in_2_4;
      end else if (10'h1ca == _T_25[9:0]) begin
        image_2_458 <= io_pixelVal_in_2_3;
      end else if (10'h1ca == _T_22[9:0]) begin
        image_2_458 <= io_pixelVal_in_2_2;
      end else if (10'h1ca == _T_19[9:0]) begin
        image_2_458 <= io_pixelVal_in_2_1;
      end else if (10'h1ca == _T_15[9:0]) begin
        image_2_458 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_459 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1cb == _T_37[9:0]) begin
        image_2_459 <= io_pixelVal_in_2_7;
      end else if (10'h1cb == _T_34[9:0]) begin
        image_2_459 <= io_pixelVal_in_2_6;
      end else if (10'h1cb == _T_31[9:0]) begin
        image_2_459 <= io_pixelVal_in_2_5;
      end else if (10'h1cb == _T_28[9:0]) begin
        image_2_459 <= io_pixelVal_in_2_4;
      end else if (10'h1cb == _T_25[9:0]) begin
        image_2_459 <= io_pixelVal_in_2_3;
      end else if (10'h1cb == _T_22[9:0]) begin
        image_2_459 <= io_pixelVal_in_2_2;
      end else if (10'h1cb == _T_19[9:0]) begin
        image_2_459 <= io_pixelVal_in_2_1;
      end else if (10'h1cb == _T_15[9:0]) begin
        image_2_459 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_460 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1cc == _T_37[9:0]) begin
        image_2_460 <= io_pixelVal_in_2_7;
      end else if (10'h1cc == _T_34[9:0]) begin
        image_2_460 <= io_pixelVal_in_2_6;
      end else if (10'h1cc == _T_31[9:0]) begin
        image_2_460 <= io_pixelVal_in_2_5;
      end else if (10'h1cc == _T_28[9:0]) begin
        image_2_460 <= io_pixelVal_in_2_4;
      end else if (10'h1cc == _T_25[9:0]) begin
        image_2_460 <= io_pixelVal_in_2_3;
      end else if (10'h1cc == _T_22[9:0]) begin
        image_2_460 <= io_pixelVal_in_2_2;
      end else if (10'h1cc == _T_19[9:0]) begin
        image_2_460 <= io_pixelVal_in_2_1;
      end else if (10'h1cc == _T_15[9:0]) begin
        image_2_460 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_461 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1cd == _T_37[9:0]) begin
        image_2_461 <= io_pixelVal_in_2_7;
      end else if (10'h1cd == _T_34[9:0]) begin
        image_2_461 <= io_pixelVal_in_2_6;
      end else if (10'h1cd == _T_31[9:0]) begin
        image_2_461 <= io_pixelVal_in_2_5;
      end else if (10'h1cd == _T_28[9:0]) begin
        image_2_461 <= io_pixelVal_in_2_4;
      end else if (10'h1cd == _T_25[9:0]) begin
        image_2_461 <= io_pixelVal_in_2_3;
      end else if (10'h1cd == _T_22[9:0]) begin
        image_2_461 <= io_pixelVal_in_2_2;
      end else if (10'h1cd == _T_19[9:0]) begin
        image_2_461 <= io_pixelVal_in_2_1;
      end else if (10'h1cd == _T_15[9:0]) begin
        image_2_461 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_462 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ce == _T_37[9:0]) begin
        image_2_462 <= io_pixelVal_in_2_7;
      end else if (10'h1ce == _T_34[9:0]) begin
        image_2_462 <= io_pixelVal_in_2_6;
      end else if (10'h1ce == _T_31[9:0]) begin
        image_2_462 <= io_pixelVal_in_2_5;
      end else if (10'h1ce == _T_28[9:0]) begin
        image_2_462 <= io_pixelVal_in_2_4;
      end else if (10'h1ce == _T_25[9:0]) begin
        image_2_462 <= io_pixelVal_in_2_3;
      end else if (10'h1ce == _T_22[9:0]) begin
        image_2_462 <= io_pixelVal_in_2_2;
      end else if (10'h1ce == _T_19[9:0]) begin
        image_2_462 <= io_pixelVal_in_2_1;
      end else if (10'h1ce == _T_15[9:0]) begin
        image_2_462 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_463 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1cf == _T_37[9:0]) begin
        image_2_463 <= io_pixelVal_in_2_7;
      end else if (10'h1cf == _T_34[9:0]) begin
        image_2_463 <= io_pixelVal_in_2_6;
      end else if (10'h1cf == _T_31[9:0]) begin
        image_2_463 <= io_pixelVal_in_2_5;
      end else if (10'h1cf == _T_28[9:0]) begin
        image_2_463 <= io_pixelVal_in_2_4;
      end else if (10'h1cf == _T_25[9:0]) begin
        image_2_463 <= io_pixelVal_in_2_3;
      end else if (10'h1cf == _T_22[9:0]) begin
        image_2_463 <= io_pixelVal_in_2_2;
      end else if (10'h1cf == _T_19[9:0]) begin
        image_2_463 <= io_pixelVal_in_2_1;
      end else if (10'h1cf == _T_15[9:0]) begin
        image_2_463 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_464 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d0 == _T_37[9:0]) begin
        image_2_464 <= io_pixelVal_in_2_7;
      end else if (10'h1d0 == _T_34[9:0]) begin
        image_2_464 <= io_pixelVal_in_2_6;
      end else if (10'h1d0 == _T_31[9:0]) begin
        image_2_464 <= io_pixelVal_in_2_5;
      end else if (10'h1d0 == _T_28[9:0]) begin
        image_2_464 <= io_pixelVal_in_2_4;
      end else if (10'h1d0 == _T_25[9:0]) begin
        image_2_464 <= io_pixelVal_in_2_3;
      end else if (10'h1d0 == _T_22[9:0]) begin
        image_2_464 <= io_pixelVal_in_2_2;
      end else if (10'h1d0 == _T_19[9:0]) begin
        image_2_464 <= io_pixelVal_in_2_1;
      end else if (10'h1d0 == _T_15[9:0]) begin
        image_2_464 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_465 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d1 == _T_37[9:0]) begin
        image_2_465 <= io_pixelVal_in_2_7;
      end else if (10'h1d1 == _T_34[9:0]) begin
        image_2_465 <= io_pixelVal_in_2_6;
      end else if (10'h1d1 == _T_31[9:0]) begin
        image_2_465 <= io_pixelVal_in_2_5;
      end else if (10'h1d1 == _T_28[9:0]) begin
        image_2_465 <= io_pixelVal_in_2_4;
      end else if (10'h1d1 == _T_25[9:0]) begin
        image_2_465 <= io_pixelVal_in_2_3;
      end else if (10'h1d1 == _T_22[9:0]) begin
        image_2_465 <= io_pixelVal_in_2_2;
      end else if (10'h1d1 == _T_19[9:0]) begin
        image_2_465 <= io_pixelVal_in_2_1;
      end else if (10'h1d1 == _T_15[9:0]) begin
        image_2_465 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_466 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d2 == _T_37[9:0]) begin
        image_2_466 <= io_pixelVal_in_2_7;
      end else if (10'h1d2 == _T_34[9:0]) begin
        image_2_466 <= io_pixelVal_in_2_6;
      end else if (10'h1d2 == _T_31[9:0]) begin
        image_2_466 <= io_pixelVal_in_2_5;
      end else if (10'h1d2 == _T_28[9:0]) begin
        image_2_466 <= io_pixelVal_in_2_4;
      end else if (10'h1d2 == _T_25[9:0]) begin
        image_2_466 <= io_pixelVal_in_2_3;
      end else if (10'h1d2 == _T_22[9:0]) begin
        image_2_466 <= io_pixelVal_in_2_2;
      end else if (10'h1d2 == _T_19[9:0]) begin
        image_2_466 <= io_pixelVal_in_2_1;
      end else if (10'h1d2 == _T_15[9:0]) begin
        image_2_466 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_467 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d3 == _T_37[9:0]) begin
        image_2_467 <= io_pixelVal_in_2_7;
      end else if (10'h1d3 == _T_34[9:0]) begin
        image_2_467 <= io_pixelVal_in_2_6;
      end else if (10'h1d3 == _T_31[9:0]) begin
        image_2_467 <= io_pixelVal_in_2_5;
      end else if (10'h1d3 == _T_28[9:0]) begin
        image_2_467 <= io_pixelVal_in_2_4;
      end else if (10'h1d3 == _T_25[9:0]) begin
        image_2_467 <= io_pixelVal_in_2_3;
      end else if (10'h1d3 == _T_22[9:0]) begin
        image_2_467 <= io_pixelVal_in_2_2;
      end else if (10'h1d3 == _T_19[9:0]) begin
        image_2_467 <= io_pixelVal_in_2_1;
      end else if (10'h1d3 == _T_15[9:0]) begin
        image_2_467 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_468 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d4 == _T_37[9:0]) begin
        image_2_468 <= io_pixelVal_in_2_7;
      end else if (10'h1d4 == _T_34[9:0]) begin
        image_2_468 <= io_pixelVal_in_2_6;
      end else if (10'h1d4 == _T_31[9:0]) begin
        image_2_468 <= io_pixelVal_in_2_5;
      end else if (10'h1d4 == _T_28[9:0]) begin
        image_2_468 <= io_pixelVal_in_2_4;
      end else if (10'h1d4 == _T_25[9:0]) begin
        image_2_468 <= io_pixelVal_in_2_3;
      end else if (10'h1d4 == _T_22[9:0]) begin
        image_2_468 <= io_pixelVal_in_2_2;
      end else if (10'h1d4 == _T_19[9:0]) begin
        image_2_468 <= io_pixelVal_in_2_1;
      end else if (10'h1d4 == _T_15[9:0]) begin
        image_2_468 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_469 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d5 == _T_37[9:0]) begin
        image_2_469 <= io_pixelVal_in_2_7;
      end else if (10'h1d5 == _T_34[9:0]) begin
        image_2_469 <= io_pixelVal_in_2_6;
      end else if (10'h1d5 == _T_31[9:0]) begin
        image_2_469 <= io_pixelVal_in_2_5;
      end else if (10'h1d5 == _T_28[9:0]) begin
        image_2_469 <= io_pixelVal_in_2_4;
      end else if (10'h1d5 == _T_25[9:0]) begin
        image_2_469 <= io_pixelVal_in_2_3;
      end else if (10'h1d5 == _T_22[9:0]) begin
        image_2_469 <= io_pixelVal_in_2_2;
      end else if (10'h1d5 == _T_19[9:0]) begin
        image_2_469 <= io_pixelVal_in_2_1;
      end else if (10'h1d5 == _T_15[9:0]) begin
        image_2_469 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_470 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d6 == _T_37[9:0]) begin
        image_2_470 <= io_pixelVal_in_2_7;
      end else if (10'h1d6 == _T_34[9:0]) begin
        image_2_470 <= io_pixelVal_in_2_6;
      end else if (10'h1d6 == _T_31[9:0]) begin
        image_2_470 <= io_pixelVal_in_2_5;
      end else if (10'h1d6 == _T_28[9:0]) begin
        image_2_470 <= io_pixelVal_in_2_4;
      end else if (10'h1d6 == _T_25[9:0]) begin
        image_2_470 <= io_pixelVal_in_2_3;
      end else if (10'h1d6 == _T_22[9:0]) begin
        image_2_470 <= io_pixelVal_in_2_2;
      end else if (10'h1d6 == _T_19[9:0]) begin
        image_2_470 <= io_pixelVal_in_2_1;
      end else if (10'h1d6 == _T_15[9:0]) begin
        image_2_470 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_471 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d7 == _T_37[9:0]) begin
        image_2_471 <= io_pixelVal_in_2_7;
      end else if (10'h1d7 == _T_34[9:0]) begin
        image_2_471 <= io_pixelVal_in_2_6;
      end else if (10'h1d7 == _T_31[9:0]) begin
        image_2_471 <= io_pixelVal_in_2_5;
      end else if (10'h1d7 == _T_28[9:0]) begin
        image_2_471 <= io_pixelVal_in_2_4;
      end else if (10'h1d7 == _T_25[9:0]) begin
        image_2_471 <= io_pixelVal_in_2_3;
      end else if (10'h1d7 == _T_22[9:0]) begin
        image_2_471 <= io_pixelVal_in_2_2;
      end else if (10'h1d7 == _T_19[9:0]) begin
        image_2_471 <= io_pixelVal_in_2_1;
      end else if (10'h1d7 == _T_15[9:0]) begin
        image_2_471 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_472 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d8 == _T_37[9:0]) begin
        image_2_472 <= io_pixelVal_in_2_7;
      end else if (10'h1d8 == _T_34[9:0]) begin
        image_2_472 <= io_pixelVal_in_2_6;
      end else if (10'h1d8 == _T_31[9:0]) begin
        image_2_472 <= io_pixelVal_in_2_5;
      end else if (10'h1d8 == _T_28[9:0]) begin
        image_2_472 <= io_pixelVal_in_2_4;
      end else if (10'h1d8 == _T_25[9:0]) begin
        image_2_472 <= io_pixelVal_in_2_3;
      end else if (10'h1d8 == _T_22[9:0]) begin
        image_2_472 <= io_pixelVal_in_2_2;
      end else if (10'h1d8 == _T_19[9:0]) begin
        image_2_472 <= io_pixelVal_in_2_1;
      end else if (10'h1d8 == _T_15[9:0]) begin
        image_2_472 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_473 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1d9 == _T_37[9:0]) begin
        image_2_473 <= io_pixelVal_in_2_7;
      end else if (10'h1d9 == _T_34[9:0]) begin
        image_2_473 <= io_pixelVal_in_2_6;
      end else if (10'h1d9 == _T_31[9:0]) begin
        image_2_473 <= io_pixelVal_in_2_5;
      end else if (10'h1d9 == _T_28[9:0]) begin
        image_2_473 <= io_pixelVal_in_2_4;
      end else if (10'h1d9 == _T_25[9:0]) begin
        image_2_473 <= io_pixelVal_in_2_3;
      end else if (10'h1d9 == _T_22[9:0]) begin
        image_2_473 <= io_pixelVal_in_2_2;
      end else if (10'h1d9 == _T_19[9:0]) begin
        image_2_473 <= io_pixelVal_in_2_1;
      end else if (10'h1d9 == _T_15[9:0]) begin
        image_2_473 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_474 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1da == _T_37[9:0]) begin
        image_2_474 <= io_pixelVal_in_2_7;
      end else if (10'h1da == _T_34[9:0]) begin
        image_2_474 <= io_pixelVal_in_2_6;
      end else if (10'h1da == _T_31[9:0]) begin
        image_2_474 <= io_pixelVal_in_2_5;
      end else if (10'h1da == _T_28[9:0]) begin
        image_2_474 <= io_pixelVal_in_2_4;
      end else if (10'h1da == _T_25[9:0]) begin
        image_2_474 <= io_pixelVal_in_2_3;
      end else if (10'h1da == _T_22[9:0]) begin
        image_2_474 <= io_pixelVal_in_2_2;
      end else if (10'h1da == _T_19[9:0]) begin
        image_2_474 <= io_pixelVal_in_2_1;
      end else if (10'h1da == _T_15[9:0]) begin
        image_2_474 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_475 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1db == _T_37[9:0]) begin
        image_2_475 <= io_pixelVal_in_2_7;
      end else if (10'h1db == _T_34[9:0]) begin
        image_2_475 <= io_pixelVal_in_2_6;
      end else if (10'h1db == _T_31[9:0]) begin
        image_2_475 <= io_pixelVal_in_2_5;
      end else if (10'h1db == _T_28[9:0]) begin
        image_2_475 <= io_pixelVal_in_2_4;
      end else if (10'h1db == _T_25[9:0]) begin
        image_2_475 <= io_pixelVal_in_2_3;
      end else if (10'h1db == _T_22[9:0]) begin
        image_2_475 <= io_pixelVal_in_2_2;
      end else if (10'h1db == _T_19[9:0]) begin
        image_2_475 <= io_pixelVal_in_2_1;
      end else if (10'h1db == _T_15[9:0]) begin
        image_2_475 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_476 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1dc == _T_37[9:0]) begin
        image_2_476 <= io_pixelVal_in_2_7;
      end else if (10'h1dc == _T_34[9:0]) begin
        image_2_476 <= io_pixelVal_in_2_6;
      end else if (10'h1dc == _T_31[9:0]) begin
        image_2_476 <= io_pixelVal_in_2_5;
      end else if (10'h1dc == _T_28[9:0]) begin
        image_2_476 <= io_pixelVal_in_2_4;
      end else if (10'h1dc == _T_25[9:0]) begin
        image_2_476 <= io_pixelVal_in_2_3;
      end else if (10'h1dc == _T_22[9:0]) begin
        image_2_476 <= io_pixelVal_in_2_2;
      end else if (10'h1dc == _T_19[9:0]) begin
        image_2_476 <= io_pixelVal_in_2_1;
      end else if (10'h1dc == _T_15[9:0]) begin
        image_2_476 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_477 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1dd == _T_37[9:0]) begin
        image_2_477 <= io_pixelVal_in_2_7;
      end else if (10'h1dd == _T_34[9:0]) begin
        image_2_477 <= io_pixelVal_in_2_6;
      end else if (10'h1dd == _T_31[9:0]) begin
        image_2_477 <= io_pixelVal_in_2_5;
      end else if (10'h1dd == _T_28[9:0]) begin
        image_2_477 <= io_pixelVal_in_2_4;
      end else if (10'h1dd == _T_25[9:0]) begin
        image_2_477 <= io_pixelVal_in_2_3;
      end else if (10'h1dd == _T_22[9:0]) begin
        image_2_477 <= io_pixelVal_in_2_2;
      end else if (10'h1dd == _T_19[9:0]) begin
        image_2_477 <= io_pixelVal_in_2_1;
      end else if (10'h1dd == _T_15[9:0]) begin
        image_2_477 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_478 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1de == _T_37[9:0]) begin
        image_2_478 <= io_pixelVal_in_2_7;
      end else if (10'h1de == _T_34[9:0]) begin
        image_2_478 <= io_pixelVal_in_2_6;
      end else if (10'h1de == _T_31[9:0]) begin
        image_2_478 <= io_pixelVal_in_2_5;
      end else if (10'h1de == _T_28[9:0]) begin
        image_2_478 <= io_pixelVal_in_2_4;
      end else if (10'h1de == _T_25[9:0]) begin
        image_2_478 <= io_pixelVal_in_2_3;
      end else if (10'h1de == _T_22[9:0]) begin
        image_2_478 <= io_pixelVal_in_2_2;
      end else if (10'h1de == _T_19[9:0]) begin
        image_2_478 <= io_pixelVal_in_2_1;
      end else if (10'h1de == _T_15[9:0]) begin
        image_2_478 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_479 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1df == _T_37[9:0]) begin
        image_2_479 <= io_pixelVal_in_2_7;
      end else if (10'h1df == _T_34[9:0]) begin
        image_2_479 <= io_pixelVal_in_2_6;
      end else if (10'h1df == _T_31[9:0]) begin
        image_2_479 <= io_pixelVal_in_2_5;
      end else if (10'h1df == _T_28[9:0]) begin
        image_2_479 <= io_pixelVal_in_2_4;
      end else if (10'h1df == _T_25[9:0]) begin
        image_2_479 <= io_pixelVal_in_2_3;
      end else if (10'h1df == _T_22[9:0]) begin
        image_2_479 <= io_pixelVal_in_2_2;
      end else if (10'h1df == _T_19[9:0]) begin
        image_2_479 <= io_pixelVal_in_2_1;
      end else if (10'h1df == _T_15[9:0]) begin
        image_2_479 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_480 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e0 == _T_37[9:0]) begin
        image_2_480 <= io_pixelVal_in_2_7;
      end else if (10'h1e0 == _T_34[9:0]) begin
        image_2_480 <= io_pixelVal_in_2_6;
      end else if (10'h1e0 == _T_31[9:0]) begin
        image_2_480 <= io_pixelVal_in_2_5;
      end else if (10'h1e0 == _T_28[9:0]) begin
        image_2_480 <= io_pixelVal_in_2_4;
      end else if (10'h1e0 == _T_25[9:0]) begin
        image_2_480 <= io_pixelVal_in_2_3;
      end else if (10'h1e0 == _T_22[9:0]) begin
        image_2_480 <= io_pixelVal_in_2_2;
      end else if (10'h1e0 == _T_19[9:0]) begin
        image_2_480 <= io_pixelVal_in_2_1;
      end else if (10'h1e0 == _T_15[9:0]) begin
        image_2_480 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_481 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e1 == _T_37[9:0]) begin
        image_2_481 <= io_pixelVal_in_2_7;
      end else if (10'h1e1 == _T_34[9:0]) begin
        image_2_481 <= io_pixelVal_in_2_6;
      end else if (10'h1e1 == _T_31[9:0]) begin
        image_2_481 <= io_pixelVal_in_2_5;
      end else if (10'h1e1 == _T_28[9:0]) begin
        image_2_481 <= io_pixelVal_in_2_4;
      end else if (10'h1e1 == _T_25[9:0]) begin
        image_2_481 <= io_pixelVal_in_2_3;
      end else if (10'h1e1 == _T_22[9:0]) begin
        image_2_481 <= io_pixelVal_in_2_2;
      end else if (10'h1e1 == _T_19[9:0]) begin
        image_2_481 <= io_pixelVal_in_2_1;
      end else if (10'h1e1 == _T_15[9:0]) begin
        image_2_481 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_482 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e2 == _T_37[9:0]) begin
        image_2_482 <= io_pixelVal_in_2_7;
      end else if (10'h1e2 == _T_34[9:0]) begin
        image_2_482 <= io_pixelVal_in_2_6;
      end else if (10'h1e2 == _T_31[9:0]) begin
        image_2_482 <= io_pixelVal_in_2_5;
      end else if (10'h1e2 == _T_28[9:0]) begin
        image_2_482 <= io_pixelVal_in_2_4;
      end else if (10'h1e2 == _T_25[9:0]) begin
        image_2_482 <= io_pixelVal_in_2_3;
      end else if (10'h1e2 == _T_22[9:0]) begin
        image_2_482 <= io_pixelVal_in_2_2;
      end else if (10'h1e2 == _T_19[9:0]) begin
        image_2_482 <= io_pixelVal_in_2_1;
      end else if (10'h1e2 == _T_15[9:0]) begin
        image_2_482 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_483 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e3 == _T_37[9:0]) begin
        image_2_483 <= io_pixelVal_in_2_7;
      end else if (10'h1e3 == _T_34[9:0]) begin
        image_2_483 <= io_pixelVal_in_2_6;
      end else if (10'h1e3 == _T_31[9:0]) begin
        image_2_483 <= io_pixelVal_in_2_5;
      end else if (10'h1e3 == _T_28[9:0]) begin
        image_2_483 <= io_pixelVal_in_2_4;
      end else if (10'h1e3 == _T_25[9:0]) begin
        image_2_483 <= io_pixelVal_in_2_3;
      end else if (10'h1e3 == _T_22[9:0]) begin
        image_2_483 <= io_pixelVal_in_2_2;
      end else if (10'h1e3 == _T_19[9:0]) begin
        image_2_483 <= io_pixelVal_in_2_1;
      end else if (10'h1e3 == _T_15[9:0]) begin
        image_2_483 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_484 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e4 == _T_37[9:0]) begin
        image_2_484 <= io_pixelVal_in_2_7;
      end else if (10'h1e4 == _T_34[9:0]) begin
        image_2_484 <= io_pixelVal_in_2_6;
      end else if (10'h1e4 == _T_31[9:0]) begin
        image_2_484 <= io_pixelVal_in_2_5;
      end else if (10'h1e4 == _T_28[9:0]) begin
        image_2_484 <= io_pixelVal_in_2_4;
      end else if (10'h1e4 == _T_25[9:0]) begin
        image_2_484 <= io_pixelVal_in_2_3;
      end else if (10'h1e4 == _T_22[9:0]) begin
        image_2_484 <= io_pixelVal_in_2_2;
      end else if (10'h1e4 == _T_19[9:0]) begin
        image_2_484 <= io_pixelVal_in_2_1;
      end else if (10'h1e4 == _T_15[9:0]) begin
        image_2_484 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_485 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e5 == _T_37[9:0]) begin
        image_2_485 <= io_pixelVal_in_2_7;
      end else if (10'h1e5 == _T_34[9:0]) begin
        image_2_485 <= io_pixelVal_in_2_6;
      end else if (10'h1e5 == _T_31[9:0]) begin
        image_2_485 <= io_pixelVal_in_2_5;
      end else if (10'h1e5 == _T_28[9:0]) begin
        image_2_485 <= io_pixelVal_in_2_4;
      end else if (10'h1e5 == _T_25[9:0]) begin
        image_2_485 <= io_pixelVal_in_2_3;
      end else if (10'h1e5 == _T_22[9:0]) begin
        image_2_485 <= io_pixelVal_in_2_2;
      end else if (10'h1e5 == _T_19[9:0]) begin
        image_2_485 <= io_pixelVal_in_2_1;
      end else if (10'h1e5 == _T_15[9:0]) begin
        image_2_485 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_486 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e6 == _T_37[9:0]) begin
        image_2_486 <= io_pixelVal_in_2_7;
      end else if (10'h1e6 == _T_34[9:0]) begin
        image_2_486 <= io_pixelVal_in_2_6;
      end else if (10'h1e6 == _T_31[9:0]) begin
        image_2_486 <= io_pixelVal_in_2_5;
      end else if (10'h1e6 == _T_28[9:0]) begin
        image_2_486 <= io_pixelVal_in_2_4;
      end else if (10'h1e6 == _T_25[9:0]) begin
        image_2_486 <= io_pixelVal_in_2_3;
      end else if (10'h1e6 == _T_22[9:0]) begin
        image_2_486 <= io_pixelVal_in_2_2;
      end else if (10'h1e6 == _T_19[9:0]) begin
        image_2_486 <= io_pixelVal_in_2_1;
      end else if (10'h1e6 == _T_15[9:0]) begin
        image_2_486 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_487 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e7 == _T_37[9:0]) begin
        image_2_487 <= io_pixelVal_in_2_7;
      end else if (10'h1e7 == _T_34[9:0]) begin
        image_2_487 <= io_pixelVal_in_2_6;
      end else if (10'h1e7 == _T_31[9:0]) begin
        image_2_487 <= io_pixelVal_in_2_5;
      end else if (10'h1e7 == _T_28[9:0]) begin
        image_2_487 <= io_pixelVal_in_2_4;
      end else if (10'h1e7 == _T_25[9:0]) begin
        image_2_487 <= io_pixelVal_in_2_3;
      end else if (10'h1e7 == _T_22[9:0]) begin
        image_2_487 <= io_pixelVal_in_2_2;
      end else if (10'h1e7 == _T_19[9:0]) begin
        image_2_487 <= io_pixelVal_in_2_1;
      end else if (10'h1e7 == _T_15[9:0]) begin
        image_2_487 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_488 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e8 == _T_37[9:0]) begin
        image_2_488 <= io_pixelVal_in_2_7;
      end else if (10'h1e8 == _T_34[9:0]) begin
        image_2_488 <= io_pixelVal_in_2_6;
      end else if (10'h1e8 == _T_31[9:0]) begin
        image_2_488 <= io_pixelVal_in_2_5;
      end else if (10'h1e8 == _T_28[9:0]) begin
        image_2_488 <= io_pixelVal_in_2_4;
      end else if (10'h1e8 == _T_25[9:0]) begin
        image_2_488 <= io_pixelVal_in_2_3;
      end else if (10'h1e8 == _T_22[9:0]) begin
        image_2_488 <= io_pixelVal_in_2_2;
      end else if (10'h1e8 == _T_19[9:0]) begin
        image_2_488 <= io_pixelVal_in_2_1;
      end else if (10'h1e8 == _T_15[9:0]) begin
        image_2_488 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_489 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1e9 == _T_37[9:0]) begin
        image_2_489 <= io_pixelVal_in_2_7;
      end else if (10'h1e9 == _T_34[9:0]) begin
        image_2_489 <= io_pixelVal_in_2_6;
      end else if (10'h1e9 == _T_31[9:0]) begin
        image_2_489 <= io_pixelVal_in_2_5;
      end else if (10'h1e9 == _T_28[9:0]) begin
        image_2_489 <= io_pixelVal_in_2_4;
      end else if (10'h1e9 == _T_25[9:0]) begin
        image_2_489 <= io_pixelVal_in_2_3;
      end else if (10'h1e9 == _T_22[9:0]) begin
        image_2_489 <= io_pixelVal_in_2_2;
      end else if (10'h1e9 == _T_19[9:0]) begin
        image_2_489 <= io_pixelVal_in_2_1;
      end else if (10'h1e9 == _T_15[9:0]) begin
        image_2_489 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_490 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ea == _T_37[9:0]) begin
        image_2_490 <= io_pixelVal_in_2_7;
      end else if (10'h1ea == _T_34[9:0]) begin
        image_2_490 <= io_pixelVal_in_2_6;
      end else if (10'h1ea == _T_31[9:0]) begin
        image_2_490 <= io_pixelVal_in_2_5;
      end else if (10'h1ea == _T_28[9:0]) begin
        image_2_490 <= io_pixelVal_in_2_4;
      end else if (10'h1ea == _T_25[9:0]) begin
        image_2_490 <= io_pixelVal_in_2_3;
      end else if (10'h1ea == _T_22[9:0]) begin
        image_2_490 <= io_pixelVal_in_2_2;
      end else if (10'h1ea == _T_19[9:0]) begin
        image_2_490 <= io_pixelVal_in_2_1;
      end else if (10'h1ea == _T_15[9:0]) begin
        image_2_490 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_491 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1eb == _T_37[9:0]) begin
        image_2_491 <= io_pixelVal_in_2_7;
      end else if (10'h1eb == _T_34[9:0]) begin
        image_2_491 <= io_pixelVal_in_2_6;
      end else if (10'h1eb == _T_31[9:0]) begin
        image_2_491 <= io_pixelVal_in_2_5;
      end else if (10'h1eb == _T_28[9:0]) begin
        image_2_491 <= io_pixelVal_in_2_4;
      end else if (10'h1eb == _T_25[9:0]) begin
        image_2_491 <= io_pixelVal_in_2_3;
      end else if (10'h1eb == _T_22[9:0]) begin
        image_2_491 <= io_pixelVal_in_2_2;
      end else if (10'h1eb == _T_19[9:0]) begin
        image_2_491 <= io_pixelVal_in_2_1;
      end else if (10'h1eb == _T_15[9:0]) begin
        image_2_491 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_492 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ec == _T_37[9:0]) begin
        image_2_492 <= io_pixelVal_in_2_7;
      end else if (10'h1ec == _T_34[9:0]) begin
        image_2_492 <= io_pixelVal_in_2_6;
      end else if (10'h1ec == _T_31[9:0]) begin
        image_2_492 <= io_pixelVal_in_2_5;
      end else if (10'h1ec == _T_28[9:0]) begin
        image_2_492 <= io_pixelVal_in_2_4;
      end else if (10'h1ec == _T_25[9:0]) begin
        image_2_492 <= io_pixelVal_in_2_3;
      end else if (10'h1ec == _T_22[9:0]) begin
        image_2_492 <= io_pixelVal_in_2_2;
      end else if (10'h1ec == _T_19[9:0]) begin
        image_2_492 <= io_pixelVal_in_2_1;
      end else if (10'h1ec == _T_15[9:0]) begin
        image_2_492 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_493 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ed == _T_37[9:0]) begin
        image_2_493 <= io_pixelVal_in_2_7;
      end else if (10'h1ed == _T_34[9:0]) begin
        image_2_493 <= io_pixelVal_in_2_6;
      end else if (10'h1ed == _T_31[9:0]) begin
        image_2_493 <= io_pixelVal_in_2_5;
      end else if (10'h1ed == _T_28[9:0]) begin
        image_2_493 <= io_pixelVal_in_2_4;
      end else if (10'h1ed == _T_25[9:0]) begin
        image_2_493 <= io_pixelVal_in_2_3;
      end else if (10'h1ed == _T_22[9:0]) begin
        image_2_493 <= io_pixelVal_in_2_2;
      end else if (10'h1ed == _T_19[9:0]) begin
        image_2_493 <= io_pixelVal_in_2_1;
      end else if (10'h1ed == _T_15[9:0]) begin
        image_2_493 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_494 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ee == _T_37[9:0]) begin
        image_2_494 <= io_pixelVal_in_2_7;
      end else if (10'h1ee == _T_34[9:0]) begin
        image_2_494 <= io_pixelVal_in_2_6;
      end else if (10'h1ee == _T_31[9:0]) begin
        image_2_494 <= io_pixelVal_in_2_5;
      end else if (10'h1ee == _T_28[9:0]) begin
        image_2_494 <= io_pixelVal_in_2_4;
      end else if (10'h1ee == _T_25[9:0]) begin
        image_2_494 <= io_pixelVal_in_2_3;
      end else if (10'h1ee == _T_22[9:0]) begin
        image_2_494 <= io_pixelVal_in_2_2;
      end else if (10'h1ee == _T_19[9:0]) begin
        image_2_494 <= io_pixelVal_in_2_1;
      end else if (10'h1ee == _T_15[9:0]) begin
        image_2_494 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_495 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ef == _T_37[9:0]) begin
        image_2_495 <= io_pixelVal_in_2_7;
      end else if (10'h1ef == _T_34[9:0]) begin
        image_2_495 <= io_pixelVal_in_2_6;
      end else if (10'h1ef == _T_31[9:0]) begin
        image_2_495 <= io_pixelVal_in_2_5;
      end else if (10'h1ef == _T_28[9:0]) begin
        image_2_495 <= io_pixelVal_in_2_4;
      end else if (10'h1ef == _T_25[9:0]) begin
        image_2_495 <= io_pixelVal_in_2_3;
      end else if (10'h1ef == _T_22[9:0]) begin
        image_2_495 <= io_pixelVal_in_2_2;
      end else if (10'h1ef == _T_19[9:0]) begin
        image_2_495 <= io_pixelVal_in_2_1;
      end else if (10'h1ef == _T_15[9:0]) begin
        image_2_495 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_496 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f0 == _T_37[9:0]) begin
        image_2_496 <= io_pixelVal_in_2_7;
      end else if (10'h1f0 == _T_34[9:0]) begin
        image_2_496 <= io_pixelVal_in_2_6;
      end else if (10'h1f0 == _T_31[9:0]) begin
        image_2_496 <= io_pixelVal_in_2_5;
      end else if (10'h1f0 == _T_28[9:0]) begin
        image_2_496 <= io_pixelVal_in_2_4;
      end else if (10'h1f0 == _T_25[9:0]) begin
        image_2_496 <= io_pixelVal_in_2_3;
      end else if (10'h1f0 == _T_22[9:0]) begin
        image_2_496 <= io_pixelVal_in_2_2;
      end else if (10'h1f0 == _T_19[9:0]) begin
        image_2_496 <= io_pixelVal_in_2_1;
      end else if (10'h1f0 == _T_15[9:0]) begin
        image_2_496 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_497 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f1 == _T_37[9:0]) begin
        image_2_497 <= io_pixelVal_in_2_7;
      end else if (10'h1f1 == _T_34[9:0]) begin
        image_2_497 <= io_pixelVal_in_2_6;
      end else if (10'h1f1 == _T_31[9:0]) begin
        image_2_497 <= io_pixelVal_in_2_5;
      end else if (10'h1f1 == _T_28[9:0]) begin
        image_2_497 <= io_pixelVal_in_2_4;
      end else if (10'h1f1 == _T_25[9:0]) begin
        image_2_497 <= io_pixelVal_in_2_3;
      end else if (10'h1f1 == _T_22[9:0]) begin
        image_2_497 <= io_pixelVal_in_2_2;
      end else if (10'h1f1 == _T_19[9:0]) begin
        image_2_497 <= io_pixelVal_in_2_1;
      end else if (10'h1f1 == _T_15[9:0]) begin
        image_2_497 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_498 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f2 == _T_37[9:0]) begin
        image_2_498 <= io_pixelVal_in_2_7;
      end else if (10'h1f2 == _T_34[9:0]) begin
        image_2_498 <= io_pixelVal_in_2_6;
      end else if (10'h1f2 == _T_31[9:0]) begin
        image_2_498 <= io_pixelVal_in_2_5;
      end else if (10'h1f2 == _T_28[9:0]) begin
        image_2_498 <= io_pixelVal_in_2_4;
      end else if (10'h1f2 == _T_25[9:0]) begin
        image_2_498 <= io_pixelVal_in_2_3;
      end else if (10'h1f2 == _T_22[9:0]) begin
        image_2_498 <= io_pixelVal_in_2_2;
      end else if (10'h1f2 == _T_19[9:0]) begin
        image_2_498 <= io_pixelVal_in_2_1;
      end else if (10'h1f2 == _T_15[9:0]) begin
        image_2_498 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_499 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f3 == _T_37[9:0]) begin
        image_2_499 <= io_pixelVal_in_2_7;
      end else if (10'h1f3 == _T_34[9:0]) begin
        image_2_499 <= io_pixelVal_in_2_6;
      end else if (10'h1f3 == _T_31[9:0]) begin
        image_2_499 <= io_pixelVal_in_2_5;
      end else if (10'h1f3 == _T_28[9:0]) begin
        image_2_499 <= io_pixelVal_in_2_4;
      end else if (10'h1f3 == _T_25[9:0]) begin
        image_2_499 <= io_pixelVal_in_2_3;
      end else if (10'h1f3 == _T_22[9:0]) begin
        image_2_499 <= io_pixelVal_in_2_2;
      end else if (10'h1f3 == _T_19[9:0]) begin
        image_2_499 <= io_pixelVal_in_2_1;
      end else if (10'h1f3 == _T_15[9:0]) begin
        image_2_499 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_500 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f4 == _T_37[9:0]) begin
        image_2_500 <= io_pixelVal_in_2_7;
      end else if (10'h1f4 == _T_34[9:0]) begin
        image_2_500 <= io_pixelVal_in_2_6;
      end else if (10'h1f4 == _T_31[9:0]) begin
        image_2_500 <= io_pixelVal_in_2_5;
      end else if (10'h1f4 == _T_28[9:0]) begin
        image_2_500 <= io_pixelVal_in_2_4;
      end else if (10'h1f4 == _T_25[9:0]) begin
        image_2_500 <= io_pixelVal_in_2_3;
      end else if (10'h1f4 == _T_22[9:0]) begin
        image_2_500 <= io_pixelVal_in_2_2;
      end else if (10'h1f4 == _T_19[9:0]) begin
        image_2_500 <= io_pixelVal_in_2_1;
      end else if (10'h1f4 == _T_15[9:0]) begin
        image_2_500 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_501 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f5 == _T_37[9:0]) begin
        image_2_501 <= io_pixelVal_in_2_7;
      end else if (10'h1f5 == _T_34[9:0]) begin
        image_2_501 <= io_pixelVal_in_2_6;
      end else if (10'h1f5 == _T_31[9:0]) begin
        image_2_501 <= io_pixelVal_in_2_5;
      end else if (10'h1f5 == _T_28[9:0]) begin
        image_2_501 <= io_pixelVal_in_2_4;
      end else if (10'h1f5 == _T_25[9:0]) begin
        image_2_501 <= io_pixelVal_in_2_3;
      end else if (10'h1f5 == _T_22[9:0]) begin
        image_2_501 <= io_pixelVal_in_2_2;
      end else if (10'h1f5 == _T_19[9:0]) begin
        image_2_501 <= io_pixelVal_in_2_1;
      end else if (10'h1f5 == _T_15[9:0]) begin
        image_2_501 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_502 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f6 == _T_37[9:0]) begin
        image_2_502 <= io_pixelVal_in_2_7;
      end else if (10'h1f6 == _T_34[9:0]) begin
        image_2_502 <= io_pixelVal_in_2_6;
      end else if (10'h1f6 == _T_31[9:0]) begin
        image_2_502 <= io_pixelVal_in_2_5;
      end else if (10'h1f6 == _T_28[9:0]) begin
        image_2_502 <= io_pixelVal_in_2_4;
      end else if (10'h1f6 == _T_25[9:0]) begin
        image_2_502 <= io_pixelVal_in_2_3;
      end else if (10'h1f6 == _T_22[9:0]) begin
        image_2_502 <= io_pixelVal_in_2_2;
      end else if (10'h1f6 == _T_19[9:0]) begin
        image_2_502 <= io_pixelVal_in_2_1;
      end else if (10'h1f6 == _T_15[9:0]) begin
        image_2_502 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_503 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f7 == _T_37[9:0]) begin
        image_2_503 <= io_pixelVal_in_2_7;
      end else if (10'h1f7 == _T_34[9:0]) begin
        image_2_503 <= io_pixelVal_in_2_6;
      end else if (10'h1f7 == _T_31[9:0]) begin
        image_2_503 <= io_pixelVal_in_2_5;
      end else if (10'h1f7 == _T_28[9:0]) begin
        image_2_503 <= io_pixelVal_in_2_4;
      end else if (10'h1f7 == _T_25[9:0]) begin
        image_2_503 <= io_pixelVal_in_2_3;
      end else if (10'h1f7 == _T_22[9:0]) begin
        image_2_503 <= io_pixelVal_in_2_2;
      end else if (10'h1f7 == _T_19[9:0]) begin
        image_2_503 <= io_pixelVal_in_2_1;
      end else if (10'h1f7 == _T_15[9:0]) begin
        image_2_503 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_504 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f8 == _T_37[9:0]) begin
        image_2_504 <= io_pixelVal_in_2_7;
      end else if (10'h1f8 == _T_34[9:0]) begin
        image_2_504 <= io_pixelVal_in_2_6;
      end else if (10'h1f8 == _T_31[9:0]) begin
        image_2_504 <= io_pixelVal_in_2_5;
      end else if (10'h1f8 == _T_28[9:0]) begin
        image_2_504 <= io_pixelVal_in_2_4;
      end else if (10'h1f8 == _T_25[9:0]) begin
        image_2_504 <= io_pixelVal_in_2_3;
      end else if (10'h1f8 == _T_22[9:0]) begin
        image_2_504 <= io_pixelVal_in_2_2;
      end else if (10'h1f8 == _T_19[9:0]) begin
        image_2_504 <= io_pixelVal_in_2_1;
      end else if (10'h1f8 == _T_15[9:0]) begin
        image_2_504 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_505 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1f9 == _T_37[9:0]) begin
        image_2_505 <= io_pixelVal_in_2_7;
      end else if (10'h1f9 == _T_34[9:0]) begin
        image_2_505 <= io_pixelVal_in_2_6;
      end else if (10'h1f9 == _T_31[9:0]) begin
        image_2_505 <= io_pixelVal_in_2_5;
      end else if (10'h1f9 == _T_28[9:0]) begin
        image_2_505 <= io_pixelVal_in_2_4;
      end else if (10'h1f9 == _T_25[9:0]) begin
        image_2_505 <= io_pixelVal_in_2_3;
      end else if (10'h1f9 == _T_22[9:0]) begin
        image_2_505 <= io_pixelVal_in_2_2;
      end else if (10'h1f9 == _T_19[9:0]) begin
        image_2_505 <= io_pixelVal_in_2_1;
      end else if (10'h1f9 == _T_15[9:0]) begin
        image_2_505 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_506 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1fa == _T_37[9:0]) begin
        image_2_506 <= io_pixelVal_in_2_7;
      end else if (10'h1fa == _T_34[9:0]) begin
        image_2_506 <= io_pixelVal_in_2_6;
      end else if (10'h1fa == _T_31[9:0]) begin
        image_2_506 <= io_pixelVal_in_2_5;
      end else if (10'h1fa == _T_28[9:0]) begin
        image_2_506 <= io_pixelVal_in_2_4;
      end else if (10'h1fa == _T_25[9:0]) begin
        image_2_506 <= io_pixelVal_in_2_3;
      end else if (10'h1fa == _T_22[9:0]) begin
        image_2_506 <= io_pixelVal_in_2_2;
      end else if (10'h1fa == _T_19[9:0]) begin
        image_2_506 <= io_pixelVal_in_2_1;
      end else if (10'h1fa == _T_15[9:0]) begin
        image_2_506 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_507 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1fb == _T_37[9:0]) begin
        image_2_507 <= io_pixelVal_in_2_7;
      end else if (10'h1fb == _T_34[9:0]) begin
        image_2_507 <= io_pixelVal_in_2_6;
      end else if (10'h1fb == _T_31[9:0]) begin
        image_2_507 <= io_pixelVal_in_2_5;
      end else if (10'h1fb == _T_28[9:0]) begin
        image_2_507 <= io_pixelVal_in_2_4;
      end else if (10'h1fb == _T_25[9:0]) begin
        image_2_507 <= io_pixelVal_in_2_3;
      end else if (10'h1fb == _T_22[9:0]) begin
        image_2_507 <= io_pixelVal_in_2_2;
      end else if (10'h1fb == _T_19[9:0]) begin
        image_2_507 <= io_pixelVal_in_2_1;
      end else if (10'h1fb == _T_15[9:0]) begin
        image_2_507 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_508 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1fc == _T_37[9:0]) begin
        image_2_508 <= io_pixelVal_in_2_7;
      end else if (10'h1fc == _T_34[9:0]) begin
        image_2_508 <= io_pixelVal_in_2_6;
      end else if (10'h1fc == _T_31[9:0]) begin
        image_2_508 <= io_pixelVal_in_2_5;
      end else if (10'h1fc == _T_28[9:0]) begin
        image_2_508 <= io_pixelVal_in_2_4;
      end else if (10'h1fc == _T_25[9:0]) begin
        image_2_508 <= io_pixelVal_in_2_3;
      end else if (10'h1fc == _T_22[9:0]) begin
        image_2_508 <= io_pixelVal_in_2_2;
      end else if (10'h1fc == _T_19[9:0]) begin
        image_2_508 <= io_pixelVal_in_2_1;
      end else if (10'h1fc == _T_15[9:0]) begin
        image_2_508 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_509 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1fd == _T_37[9:0]) begin
        image_2_509 <= io_pixelVal_in_2_7;
      end else if (10'h1fd == _T_34[9:0]) begin
        image_2_509 <= io_pixelVal_in_2_6;
      end else if (10'h1fd == _T_31[9:0]) begin
        image_2_509 <= io_pixelVal_in_2_5;
      end else if (10'h1fd == _T_28[9:0]) begin
        image_2_509 <= io_pixelVal_in_2_4;
      end else if (10'h1fd == _T_25[9:0]) begin
        image_2_509 <= io_pixelVal_in_2_3;
      end else if (10'h1fd == _T_22[9:0]) begin
        image_2_509 <= io_pixelVal_in_2_2;
      end else if (10'h1fd == _T_19[9:0]) begin
        image_2_509 <= io_pixelVal_in_2_1;
      end else if (10'h1fd == _T_15[9:0]) begin
        image_2_509 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_510 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1fe == _T_37[9:0]) begin
        image_2_510 <= io_pixelVal_in_2_7;
      end else if (10'h1fe == _T_34[9:0]) begin
        image_2_510 <= io_pixelVal_in_2_6;
      end else if (10'h1fe == _T_31[9:0]) begin
        image_2_510 <= io_pixelVal_in_2_5;
      end else if (10'h1fe == _T_28[9:0]) begin
        image_2_510 <= io_pixelVal_in_2_4;
      end else if (10'h1fe == _T_25[9:0]) begin
        image_2_510 <= io_pixelVal_in_2_3;
      end else if (10'h1fe == _T_22[9:0]) begin
        image_2_510 <= io_pixelVal_in_2_2;
      end else if (10'h1fe == _T_19[9:0]) begin
        image_2_510 <= io_pixelVal_in_2_1;
      end else if (10'h1fe == _T_15[9:0]) begin
        image_2_510 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_511 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h1ff == _T_37[9:0]) begin
        image_2_511 <= io_pixelVal_in_2_7;
      end else if (10'h1ff == _T_34[9:0]) begin
        image_2_511 <= io_pixelVal_in_2_6;
      end else if (10'h1ff == _T_31[9:0]) begin
        image_2_511 <= io_pixelVal_in_2_5;
      end else if (10'h1ff == _T_28[9:0]) begin
        image_2_511 <= io_pixelVal_in_2_4;
      end else if (10'h1ff == _T_25[9:0]) begin
        image_2_511 <= io_pixelVal_in_2_3;
      end else if (10'h1ff == _T_22[9:0]) begin
        image_2_511 <= io_pixelVal_in_2_2;
      end else if (10'h1ff == _T_19[9:0]) begin
        image_2_511 <= io_pixelVal_in_2_1;
      end else if (10'h1ff == _T_15[9:0]) begin
        image_2_511 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_512 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h200 == _T_37[9:0]) begin
        image_2_512 <= io_pixelVal_in_2_7;
      end else if (10'h200 == _T_34[9:0]) begin
        image_2_512 <= io_pixelVal_in_2_6;
      end else if (10'h200 == _T_31[9:0]) begin
        image_2_512 <= io_pixelVal_in_2_5;
      end else if (10'h200 == _T_28[9:0]) begin
        image_2_512 <= io_pixelVal_in_2_4;
      end else if (10'h200 == _T_25[9:0]) begin
        image_2_512 <= io_pixelVal_in_2_3;
      end else if (10'h200 == _T_22[9:0]) begin
        image_2_512 <= io_pixelVal_in_2_2;
      end else if (10'h200 == _T_19[9:0]) begin
        image_2_512 <= io_pixelVal_in_2_1;
      end else if (10'h200 == _T_15[9:0]) begin
        image_2_512 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_513 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h201 == _T_37[9:0]) begin
        image_2_513 <= io_pixelVal_in_2_7;
      end else if (10'h201 == _T_34[9:0]) begin
        image_2_513 <= io_pixelVal_in_2_6;
      end else if (10'h201 == _T_31[9:0]) begin
        image_2_513 <= io_pixelVal_in_2_5;
      end else if (10'h201 == _T_28[9:0]) begin
        image_2_513 <= io_pixelVal_in_2_4;
      end else if (10'h201 == _T_25[9:0]) begin
        image_2_513 <= io_pixelVal_in_2_3;
      end else if (10'h201 == _T_22[9:0]) begin
        image_2_513 <= io_pixelVal_in_2_2;
      end else if (10'h201 == _T_19[9:0]) begin
        image_2_513 <= io_pixelVal_in_2_1;
      end else if (10'h201 == _T_15[9:0]) begin
        image_2_513 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_514 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h202 == _T_37[9:0]) begin
        image_2_514 <= io_pixelVal_in_2_7;
      end else if (10'h202 == _T_34[9:0]) begin
        image_2_514 <= io_pixelVal_in_2_6;
      end else if (10'h202 == _T_31[9:0]) begin
        image_2_514 <= io_pixelVal_in_2_5;
      end else if (10'h202 == _T_28[9:0]) begin
        image_2_514 <= io_pixelVal_in_2_4;
      end else if (10'h202 == _T_25[9:0]) begin
        image_2_514 <= io_pixelVal_in_2_3;
      end else if (10'h202 == _T_22[9:0]) begin
        image_2_514 <= io_pixelVal_in_2_2;
      end else if (10'h202 == _T_19[9:0]) begin
        image_2_514 <= io_pixelVal_in_2_1;
      end else if (10'h202 == _T_15[9:0]) begin
        image_2_514 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_515 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h203 == _T_37[9:0]) begin
        image_2_515 <= io_pixelVal_in_2_7;
      end else if (10'h203 == _T_34[9:0]) begin
        image_2_515 <= io_pixelVal_in_2_6;
      end else if (10'h203 == _T_31[9:0]) begin
        image_2_515 <= io_pixelVal_in_2_5;
      end else if (10'h203 == _T_28[9:0]) begin
        image_2_515 <= io_pixelVal_in_2_4;
      end else if (10'h203 == _T_25[9:0]) begin
        image_2_515 <= io_pixelVal_in_2_3;
      end else if (10'h203 == _T_22[9:0]) begin
        image_2_515 <= io_pixelVal_in_2_2;
      end else if (10'h203 == _T_19[9:0]) begin
        image_2_515 <= io_pixelVal_in_2_1;
      end else if (10'h203 == _T_15[9:0]) begin
        image_2_515 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_516 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h204 == _T_37[9:0]) begin
        image_2_516 <= io_pixelVal_in_2_7;
      end else if (10'h204 == _T_34[9:0]) begin
        image_2_516 <= io_pixelVal_in_2_6;
      end else if (10'h204 == _T_31[9:0]) begin
        image_2_516 <= io_pixelVal_in_2_5;
      end else if (10'h204 == _T_28[9:0]) begin
        image_2_516 <= io_pixelVal_in_2_4;
      end else if (10'h204 == _T_25[9:0]) begin
        image_2_516 <= io_pixelVal_in_2_3;
      end else if (10'h204 == _T_22[9:0]) begin
        image_2_516 <= io_pixelVal_in_2_2;
      end else if (10'h204 == _T_19[9:0]) begin
        image_2_516 <= io_pixelVal_in_2_1;
      end else if (10'h204 == _T_15[9:0]) begin
        image_2_516 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_517 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h205 == _T_37[9:0]) begin
        image_2_517 <= io_pixelVal_in_2_7;
      end else if (10'h205 == _T_34[9:0]) begin
        image_2_517 <= io_pixelVal_in_2_6;
      end else if (10'h205 == _T_31[9:0]) begin
        image_2_517 <= io_pixelVal_in_2_5;
      end else if (10'h205 == _T_28[9:0]) begin
        image_2_517 <= io_pixelVal_in_2_4;
      end else if (10'h205 == _T_25[9:0]) begin
        image_2_517 <= io_pixelVal_in_2_3;
      end else if (10'h205 == _T_22[9:0]) begin
        image_2_517 <= io_pixelVal_in_2_2;
      end else if (10'h205 == _T_19[9:0]) begin
        image_2_517 <= io_pixelVal_in_2_1;
      end else if (10'h205 == _T_15[9:0]) begin
        image_2_517 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_518 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h206 == _T_37[9:0]) begin
        image_2_518 <= io_pixelVal_in_2_7;
      end else if (10'h206 == _T_34[9:0]) begin
        image_2_518 <= io_pixelVal_in_2_6;
      end else if (10'h206 == _T_31[9:0]) begin
        image_2_518 <= io_pixelVal_in_2_5;
      end else if (10'h206 == _T_28[9:0]) begin
        image_2_518 <= io_pixelVal_in_2_4;
      end else if (10'h206 == _T_25[9:0]) begin
        image_2_518 <= io_pixelVal_in_2_3;
      end else if (10'h206 == _T_22[9:0]) begin
        image_2_518 <= io_pixelVal_in_2_2;
      end else if (10'h206 == _T_19[9:0]) begin
        image_2_518 <= io_pixelVal_in_2_1;
      end else if (10'h206 == _T_15[9:0]) begin
        image_2_518 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_519 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h207 == _T_37[9:0]) begin
        image_2_519 <= io_pixelVal_in_2_7;
      end else if (10'h207 == _T_34[9:0]) begin
        image_2_519 <= io_pixelVal_in_2_6;
      end else if (10'h207 == _T_31[9:0]) begin
        image_2_519 <= io_pixelVal_in_2_5;
      end else if (10'h207 == _T_28[9:0]) begin
        image_2_519 <= io_pixelVal_in_2_4;
      end else if (10'h207 == _T_25[9:0]) begin
        image_2_519 <= io_pixelVal_in_2_3;
      end else if (10'h207 == _T_22[9:0]) begin
        image_2_519 <= io_pixelVal_in_2_2;
      end else if (10'h207 == _T_19[9:0]) begin
        image_2_519 <= io_pixelVal_in_2_1;
      end else if (10'h207 == _T_15[9:0]) begin
        image_2_519 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_520 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h208 == _T_37[9:0]) begin
        image_2_520 <= io_pixelVal_in_2_7;
      end else if (10'h208 == _T_34[9:0]) begin
        image_2_520 <= io_pixelVal_in_2_6;
      end else if (10'h208 == _T_31[9:0]) begin
        image_2_520 <= io_pixelVal_in_2_5;
      end else if (10'h208 == _T_28[9:0]) begin
        image_2_520 <= io_pixelVal_in_2_4;
      end else if (10'h208 == _T_25[9:0]) begin
        image_2_520 <= io_pixelVal_in_2_3;
      end else if (10'h208 == _T_22[9:0]) begin
        image_2_520 <= io_pixelVal_in_2_2;
      end else if (10'h208 == _T_19[9:0]) begin
        image_2_520 <= io_pixelVal_in_2_1;
      end else if (10'h208 == _T_15[9:0]) begin
        image_2_520 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_521 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h209 == _T_37[9:0]) begin
        image_2_521 <= io_pixelVal_in_2_7;
      end else if (10'h209 == _T_34[9:0]) begin
        image_2_521 <= io_pixelVal_in_2_6;
      end else if (10'h209 == _T_31[9:0]) begin
        image_2_521 <= io_pixelVal_in_2_5;
      end else if (10'h209 == _T_28[9:0]) begin
        image_2_521 <= io_pixelVal_in_2_4;
      end else if (10'h209 == _T_25[9:0]) begin
        image_2_521 <= io_pixelVal_in_2_3;
      end else if (10'h209 == _T_22[9:0]) begin
        image_2_521 <= io_pixelVal_in_2_2;
      end else if (10'h209 == _T_19[9:0]) begin
        image_2_521 <= io_pixelVal_in_2_1;
      end else if (10'h209 == _T_15[9:0]) begin
        image_2_521 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_522 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h20a == _T_37[9:0]) begin
        image_2_522 <= io_pixelVal_in_2_7;
      end else if (10'h20a == _T_34[9:0]) begin
        image_2_522 <= io_pixelVal_in_2_6;
      end else if (10'h20a == _T_31[9:0]) begin
        image_2_522 <= io_pixelVal_in_2_5;
      end else if (10'h20a == _T_28[9:0]) begin
        image_2_522 <= io_pixelVal_in_2_4;
      end else if (10'h20a == _T_25[9:0]) begin
        image_2_522 <= io_pixelVal_in_2_3;
      end else if (10'h20a == _T_22[9:0]) begin
        image_2_522 <= io_pixelVal_in_2_2;
      end else if (10'h20a == _T_19[9:0]) begin
        image_2_522 <= io_pixelVal_in_2_1;
      end else if (10'h20a == _T_15[9:0]) begin
        image_2_522 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_523 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h20b == _T_37[9:0]) begin
        image_2_523 <= io_pixelVal_in_2_7;
      end else if (10'h20b == _T_34[9:0]) begin
        image_2_523 <= io_pixelVal_in_2_6;
      end else if (10'h20b == _T_31[9:0]) begin
        image_2_523 <= io_pixelVal_in_2_5;
      end else if (10'h20b == _T_28[9:0]) begin
        image_2_523 <= io_pixelVal_in_2_4;
      end else if (10'h20b == _T_25[9:0]) begin
        image_2_523 <= io_pixelVal_in_2_3;
      end else if (10'h20b == _T_22[9:0]) begin
        image_2_523 <= io_pixelVal_in_2_2;
      end else if (10'h20b == _T_19[9:0]) begin
        image_2_523 <= io_pixelVal_in_2_1;
      end else if (10'h20b == _T_15[9:0]) begin
        image_2_523 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_524 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h20c == _T_37[9:0]) begin
        image_2_524 <= io_pixelVal_in_2_7;
      end else if (10'h20c == _T_34[9:0]) begin
        image_2_524 <= io_pixelVal_in_2_6;
      end else if (10'h20c == _T_31[9:0]) begin
        image_2_524 <= io_pixelVal_in_2_5;
      end else if (10'h20c == _T_28[9:0]) begin
        image_2_524 <= io_pixelVal_in_2_4;
      end else if (10'h20c == _T_25[9:0]) begin
        image_2_524 <= io_pixelVal_in_2_3;
      end else if (10'h20c == _T_22[9:0]) begin
        image_2_524 <= io_pixelVal_in_2_2;
      end else if (10'h20c == _T_19[9:0]) begin
        image_2_524 <= io_pixelVal_in_2_1;
      end else if (10'h20c == _T_15[9:0]) begin
        image_2_524 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_525 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h20d == _T_37[9:0]) begin
        image_2_525 <= io_pixelVal_in_2_7;
      end else if (10'h20d == _T_34[9:0]) begin
        image_2_525 <= io_pixelVal_in_2_6;
      end else if (10'h20d == _T_31[9:0]) begin
        image_2_525 <= io_pixelVal_in_2_5;
      end else if (10'h20d == _T_28[9:0]) begin
        image_2_525 <= io_pixelVal_in_2_4;
      end else if (10'h20d == _T_25[9:0]) begin
        image_2_525 <= io_pixelVal_in_2_3;
      end else if (10'h20d == _T_22[9:0]) begin
        image_2_525 <= io_pixelVal_in_2_2;
      end else if (10'h20d == _T_19[9:0]) begin
        image_2_525 <= io_pixelVal_in_2_1;
      end else if (10'h20d == _T_15[9:0]) begin
        image_2_525 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_526 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h20e == _T_37[9:0]) begin
        image_2_526 <= io_pixelVal_in_2_7;
      end else if (10'h20e == _T_34[9:0]) begin
        image_2_526 <= io_pixelVal_in_2_6;
      end else if (10'h20e == _T_31[9:0]) begin
        image_2_526 <= io_pixelVal_in_2_5;
      end else if (10'h20e == _T_28[9:0]) begin
        image_2_526 <= io_pixelVal_in_2_4;
      end else if (10'h20e == _T_25[9:0]) begin
        image_2_526 <= io_pixelVal_in_2_3;
      end else if (10'h20e == _T_22[9:0]) begin
        image_2_526 <= io_pixelVal_in_2_2;
      end else if (10'h20e == _T_19[9:0]) begin
        image_2_526 <= io_pixelVal_in_2_1;
      end else if (10'h20e == _T_15[9:0]) begin
        image_2_526 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_527 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h20f == _T_37[9:0]) begin
        image_2_527 <= io_pixelVal_in_2_7;
      end else if (10'h20f == _T_34[9:0]) begin
        image_2_527 <= io_pixelVal_in_2_6;
      end else if (10'h20f == _T_31[9:0]) begin
        image_2_527 <= io_pixelVal_in_2_5;
      end else if (10'h20f == _T_28[9:0]) begin
        image_2_527 <= io_pixelVal_in_2_4;
      end else if (10'h20f == _T_25[9:0]) begin
        image_2_527 <= io_pixelVal_in_2_3;
      end else if (10'h20f == _T_22[9:0]) begin
        image_2_527 <= io_pixelVal_in_2_2;
      end else if (10'h20f == _T_19[9:0]) begin
        image_2_527 <= io_pixelVal_in_2_1;
      end else if (10'h20f == _T_15[9:0]) begin
        image_2_527 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_528 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h210 == _T_37[9:0]) begin
        image_2_528 <= io_pixelVal_in_2_7;
      end else if (10'h210 == _T_34[9:0]) begin
        image_2_528 <= io_pixelVal_in_2_6;
      end else if (10'h210 == _T_31[9:0]) begin
        image_2_528 <= io_pixelVal_in_2_5;
      end else if (10'h210 == _T_28[9:0]) begin
        image_2_528 <= io_pixelVal_in_2_4;
      end else if (10'h210 == _T_25[9:0]) begin
        image_2_528 <= io_pixelVal_in_2_3;
      end else if (10'h210 == _T_22[9:0]) begin
        image_2_528 <= io_pixelVal_in_2_2;
      end else if (10'h210 == _T_19[9:0]) begin
        image_2_528 <= io_pixelVal_in_2_1;
      end else if (10'h210 == _T_15[9:0]) begin
        image_2_528 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_529 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h211 == _T_37[9:0]) begin
        image_2_529 <= io_pixelVal_in_2_7;
      end else if (10'h211 == _T_34[9:0]) begin
        image_2_529 <= io_pixelVal_in_2_6;
      end else if (10'h211 == _T_31[9:0]) begin
        image_2_529 <= io_pixelVal_in_2_5;
      end else if (10'h211 == _T_28[9:0]) begin
        image_2_529 <= io_pixelVal_in_2_4;
      end else if (10'h211 == _T_25[9:0]) begin
        image_2_529 <= io_pixelVal_in_2_3;
      end else if (10'h211 == _T_22[9:0]) begin
        image_2_529 <= io_pixelVal_in_2_2;
      end else if (10'h211 == _T_19[9:0]) begin
        image_2_529 <= io_pixelVal_in_2_1;
      end else if (10'h211 == _T_15[9:0]) begin
        image_2_529 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_530 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h212 == _T_37[9:0]) begin
        image_2_530 <= io_pixelVal_in_2_7;
      end else if (10'h212 == _T_34[9:0]) begin
        image_2_530 <= io_pixelVal_in_2_6;
      end else if (10'h212 == _T_31[9:0]) begin
        image_2_530 <= io_pixelVal_in_2_5;
      end else if (10'h212 == _T_28[9:0]) begin
        image_2_530 <= io_pixelVal_in_2_4;
      end else if (10'h212 == _T_25[9:0]) begin
        image_2_530 <= io_pixelVal_in_2_3;
      end else if (10'h212 == _T_22[9:0]) begin
        image_2_530 <= io_pixelVal_in_2_2;
      end else if (10'h212 == _T_19[9:0]) begin
        image_2_530 <= io_pixelVal_in_2_1;
      end else if (10'h212 == _T_15[9:0]) begin
        image_2_530 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_531 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h213 == _T_37[9:0]) begin
        image_2_531 <= io_pixelVal_in_2_7;
      end else if (10'h213 == _T_34[9:0]) begin
        image_2_531 <= io_pixelVal_in_2_6;
      end else if (10'h213 == _T_31[9:0]) begin
        image_2_531 <= io_pixelVal_in_2_5;
      end else if (10'h213 == _T_28[9:0]) begin
        image_2_531 <= io_pixelVal_in_2_4;
      end else if (10'h213 == _T_25[9:0]) begin
        image_2_531 <= io_pixelVal_in_2_3;
      end else if (10'h213 == _T_22[9:0]) begin
        image_2_531 <= io_pixelVal_in_2_2;
      end else if (10'h213 == _T_19[9:0]) begin
        image_2_531 <= io_pixelVal_in_2_1;
      end else if (10'h213 == _T_15[9:0]) begin
        image_2_531 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_532 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h214 == _T_37[9:0]) begin
        image_2_532 <= io_pixelVal_in_2_7;
      end else if (10'h214 == _T_34[9:0]) begin
        image_2_532 <= io_pixelVal_in_2_6;
      end else if (10'h214 == _T_31[9:0]) begin
        image_2_532 <= io_pixelVal_in_2_5;
      end else if (10'h214 == _T_28[9:0]) begin
        image_2_532 <= io_pixelVal_in_2_4;
      end else if (10'h214 == _T_25[9:0]) begin
        image_2_532 <= io_pixelVal_in_2_3;
      end else if (10'h214 == _T_22[9:0]) begin
        image_2_532 <= io_pixelVal_in_2_2;
      end else if (10'h214 == _T_19[9:0]) begin
        image_2_532 <= io_pixelVal_in_2_1;
      end else if (10'h214 == _T_15[9:0]) begin
        image_2_532 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_533 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h215 == _T_37[9:0]) begin
        image_2_533 <= io_pixelVal_in_2_7;
      end else if (10'h215 == _T_34[9:0]) begin
        image_2_533 <= io_pixelVal_in_2_6;
      end else if (10'h215 == _T_31[9:0]) begin
        image_2_533 <= io_pixelVal_in_2_5;
      end else if (10'h215 == _T_28[9:0]) begin
        image_2_533 <= io_pixelVal_in_2_4;
      end else if (10'h215 == _T_25[9:0]) begin
        image_2_533 <= io_pixelVal_in_2_3;
      end else if (10'h215 == _T_22[9:0]) begin
        image_2_533 <= io_pixelVal_in_2_2;
      end else if (10'h215 == _T_19[9:0]) begin
        image_2_533 <= io_pixelVal_in_2_1;
      end else if (10'h215 == _T_15[9:0]) begin
        image_2_533 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_534 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h216 == _T_37[9:0]) begin
        image_2_534 <= io_pixelVal_in_2_7;
      end else if (10'h216 == _T_34[9:0]) begin
        image_2_534 <= io_pixelVal_in_2_6;
      end else if (10'h216 == _T_31[9:0]) begin
        image_2_534 <= io_pixelVal_in_2_5;
      end else if (10'h216 == _T_28[9:0]) begin
        image_2_534 <= io_pixelVal_in_2_4;
      end else if (10'h216 == _T_25[9:0]) begin
        image_2_534 <= io_pixelVal_in_2_3;
      end else if (10'h216 == _T_22[9:0]) begin
        image_2_534 <= io_pixelVal_in_2_2;
      end else if (10'h216 == _T_19[9:0]) begin
        image_2_534 <= io_pixelVal_in_2_1;
      end else if (10'h216 == _T_15[9:0]) begin
        image_2_534 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_535 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h217 == _T_37[9:0]) begin
        image_2_535 <= io_pixelVal_in_2_7;
      end else if (10'h217 == _T_34[9:0]) begin
        image_2_535 <= io_pixelVal_in_2_6;
      end else if (10'h217 == _T_31[9:0]) begin
        image_2_535 <= io_pixelVal_in_2_5;
      end else if (10'h217 == _T_28[9:0]) begin
        image_2_535 <= io_pixelVal_in_2_4;
      end else if (10'h217 == _T_25[9:0]) begin
        image_2_535 <= io_pixelVal_in_2_3;
      end else if (10'h217 == _T_22[9:0]) begin
        image_2_535 <= io_pixelVal_in_2_2;
      end else if (10'h217 == _T_19[9:0]) begin
        image_2_535 <= io_pixelVal_in_2_1;
      end else if (10'h217 == _T_15[9:0]) begin
        image_2_535 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_536 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h218 == _T_37[9:0]) begin
        image_2_536 <= io_pixelVal_in_2_7;
      end else if (10'h218 == _T_34[9:0]) begin
        image_2_536 <= io_pixelVal_in_2_6;
      end else if (10'h218 == _T_31[9:0]) begin
        image_2_536 <= io_pixelVal_in_2_5;
      end else if (10'h218 == _T_28[9:0]) begin
        image_2_536 <= io_pixelVal_in_2_4;
      end else if (10'h218 == _T_25[9:0]) begin
        image_2_536 <= io_pixelVal_in_2_3;
      end else if (10'h218 == _T_22[9:0]) begin
        image_2_536 <= io_pixelVal_in_2_2;
      end else if (10'h218 == _T_19[9:0]) begin
        image_2_536 <= io_pixelVal_in_2_1;
      end else if (10'h218 == _T_15[9:0]) begin
        image_2_536 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_537 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h219 == _T_37[9:0]) begin
        image_2_537 <= io_pixelVal_in_2_7;
      end else if (10'h219 == _T_34[9:0]) begin
        image_2_537 <= io_pixelVal_in_2_6;
      end else if (10'h219 == _T_31[9:0]) begin
        image_2_537 <= io_pixelVal_in_2_5;
      end else if (10'h219 == _T_28[9:0]) begin
        image_2_537 <= io_pixelVal_in_2_4;
      end else if (10'h219 == _T_25[9:0]) begin
        image_2_537 <= io_pixelVal_in_2_3;
      end else if (10'h219 == _T_22[9:0]) begin
        image_2_537 <= io_pixelVal_in_2_2;
      end else if (10'h219 == _T_19[9:0]) begin
        image_2_537 <= io_pixelVal_in_2_1;
      end else if (10'h219 == _T_15[9:0]) begin
        image_2_537 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_538 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h21a == _T_37[9:0]) begin
        image_2_538 <= io_pixelVal_in_2_7;
      end else if (10'h21a == _T_34[9:0]) begin
        image_2_538 <= io_pixelVal_in_2_6;
      end else if (10'h21a == _T_31[9:0]) begin
        image_2_538 <= io_pixelVal_in_2_5;
      end else if (10'h21a == _T_28[9:0]) begin
        image_2_538 <= io_pixelVal_in_2_4;
      end else if (10'h21a == _T_25[9:0]) begin
        image_2_538 <= io_pixelVal_in_2_3;
      end else if (10'h21a == _T_22[9:0]) begin
        image_2_538 <= io_pixelVal_in_2_2;
      end else if (10'h21a == _T_19[9:0]) begin
        image_2_538 <= io_pixelVal_in_2_1;
      end else if (10'h21a == _T_15[9:0]) begin
        image_2_538 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_539 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h21b == _T_37[9:0]) begin
        image_2_539 <= io_pixelVal_in_2_7;
      end else if (10'h21b == _T_34[9:0]) begin
        image_2_539 <= io_pixelVal_in_2_6;
      end else if (10'h21b == _T_31[9:0]) begin
        image_2_539 <= io_pixelVal_in_2_5;
      end else if (10'h21b == _T_28[9:0]) begin
        image_2_539 <= io_pixelVal_in_2_4;
      end else if (10'h21b == _T_25[9:0]) begin
        image_2_539 <= io_pixelVal_in_2_3;
      end else if (10'h21b == _T_22[9:0]) begin
        image_2_539 <= io_pixelVal_in_2_2;
      end else if (10'h21b == _T_19[9:0]) begin
        image_2_539 <= io_pixelVal_in_2_1;
      end else if (10'h21b == _T_15[9:0]) begin
        image_2_539 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_540 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h21c == _T_37[9:0]) begin
        image_2_540 <= io_pixelVal_in_2_7;
      end else if (10'h21c == _T_34[9:0]) begin
        image_2_540 <= io_pixelVal_in_2_6;
      end else if (10'h21c == _T_31[9:0]) begin
        image_2_540 <= io_pixelVal_in_2_5;
      end else if (10'h21c == _T_28[9:0]) begin
        image_2_540 <= io_pixelVal_in_2_4;
      end else if (10'h21c == _T_25[9:0]) begin
        image_2_540 <= io_pixelVal_in_2_3;
      end else if (10'h21c == _T_22[9:0]) begin
        image_2_540 <= io_pixelVal_in_2_2;
      end else if (10'h21c == _T_19[9:0]) begin
        image_2_540 <= io_pixelVal_in_2_1;
      end else if (10'h21c == _T_15[9:0]) begin
        image_2_540 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_541 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h21d == _T_37[9:0]) begin
        image_2_541 <= io_pixelVal_in_2_7;
      end else if (10'h21d == _T_34[9:0]) begin
        image_2_541 <= io_pixelVal_in_2_6;
      end else if (10'h21d == _T_31[9:0]) begin
        image_2_541 <= io_pixelVal_in_2_5;
      end else if (10'h21d == _T_28[9:0]) begin
        image_2_541 <= io_pixelVal_in_2_4;
      end else if (10'h21d == _T_25[9:0]) begin
        image_2_541 <= io_pixelVal_in_2_3;
      end else if (10'h21d == _T_22[9:0]) begin
        image_2_541 <= io_pixelVal_in_2_2;
      end else if (10'h21d == _T_19[9:0]) begin
        image_2_541 <= io_pixelVal_in_2_1;
      end else if (10'h21d == _T_15[9:0]) begin
        image_2_541 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_542 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h21e == _T_37[9:0]) begin
        image_2_542 <= io_pixelVal_in_2_7;
      end else if (10'h21e == _T_34[9:0]) begin
        image_2_542 <= io_pixelVal_in_2_6;
      end else if (10'h21e == _T_31[9:0]) begin
        image_2_542 <= io_pixelVal_in_2_5;
      end else if (10'h21e == _T_28[9:0]) begin
        image_2_542 <= io_pixelVal_in_2_4;
      end else if (10'h21e == _T_25[9:0]) begin
        image_2_542 <= io_pixelVal_in_2_3;
      end else if (10'h21e == _T_22[9:0]) begin
        image_2_542 <= io_pixelVal_in_2_2;
      end else if (10'h21e == _T_19[9:0]) begin
        image_2_542 <= io_pixelVal_in_2_1;
      end else if (10'h21e == _T_15[9:0]) begin
        image_2_542 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_543 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h21f == _T_37[9:0]) begin
        image_2_543 <= io_pixelVal_in_2_7;
      end else if (10'h21f == _T_34[9:0]) begin
        image_2_543 <= io_pixelVal_in_2_6;
      end else if (10'h21f == _T_31[9:0]) begin
        image_2_543 <= io_pixelVal_in_2_5;
      end else if (10'h21f == _T_28[9:0]) begin
        image_2_543 <= io_pixelVal_in_2_4;
      end else if (10'h21f == _T_25[9:0]) begin
        image_2_543 <= io_pixelVal_in_2_3;
      end else if (10'h21f == _T_22[9:0]) begin
        image_2_543 <= io_pixelVal_in_2_2;
      end else if (10'h21f == _T_19[9:0]) begin
        image_2_543 <= io_pixelVal_in_2_1;
      end else if (10'h21f == _T_15[9:0]) begin
        image_2_543 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_544 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h220 == _T_37[9:0]) begin
        image_2_544 <= io_pixelVal_in_2_7;
      end else if (10'h220 == _T_34[9:0]) begin
        image_2_544 <= io_pixelVal_in_2_6;
      end else if (10'h220 == _T_31[9:0]) begin
        image_2_544 <= io_pixelVal_in_2_5;
      end else if (10'h220 == _T_28[9:0]) begin
        image_2_544 <= io_pixelVal_in_2_4;
      end else if (10'h220 == _T_25[9:0]) begin
        image_2_544 <= io_pixelVal_in_2_3;
      end else if (10'h220 == _T_22[9:0]) begin
        image_2_544 <= io_pixelVal_in_2_2;
      end else if (10'h220 == _T_19[9:0]) begin
        image_2_544 <= io_pixelVal_in_2_1;
      end else if (10'h220 == _T_15[9:0]) begin
        image_2_544 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_545 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h221 == _T_37[9:0]) begin
        image_2_545 <= io_pixelVal_in_2_7;
      end else if (10'h221 == _T_34[9:0]) begin
        image_2_545 <= io_pixelVal_in_2_6;
      end else if (10'h221 == _T_31[9:0]) begin
        image_2_545 <= io_pixelVal_in_2_5;
      end else if (10'h221 == _T_28[9:0]) begin
        image_2_545 <= io_pixelVal_in_2_4;
      end else if (10'h221 == _T_25[9:0]) begin
        image_2_545 <= io_pixelVal_in_2_3;
      end else if (10'h221 == _T_22[9:0]) begin
        image_2_545 <= io_pixelVal_in_2_2;
      end else if (10'h221 == _T_19[9:0]) begin
        image_2_545 <= io_pixelVal_in_2_1;
      end else if (10'h221 == _T_15[9:0]) begin
        image_2_545 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_546 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h222 == _T_37[9:0]) begin
        image_2_546 <= io_pixelVal_in_2_7;
      end else if (10'h222 == _T_34[9:0]) begin
        image_2_546 <= io_pixelVal_in_2_6;
      end else if (10'h222 == _T_31[9:0]) begin
        image_2_546 <= io_pixelVal_in_2_5;
      end else if (10'h222 == _T_28[9:0]) begin
        image_2_546 <= io_pixelVal_in_2_4;
      end else if (10'h222 == _T_25[9:0]) begin
        image_2_546 <= io_pixelVal_in_2_3;
      end else if (10'h222 == _T_22[9:0]) begin
        image_2_546 <= io_pixelVal_in_2_2;
      end else if (10'h222 == _T_19[9:0]) begin
        image_2_546 <= io_pixelVal_in_2_1;
      end else if (10'h222 == _T_15[9:0]) begin
        image_2_546 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_547 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h223 == _T_37[9:0]) begin
        image_2_547 <= io_pixelVal_in_2_7;
      end else if (10'h223 == _T_34[9:0]) begin
        image_2_547 <= io_pixelVal_in_2_6;
      end else if (10'h223 == _T_31[9:0]) begin
        image_2_547 <= io_pixelVal_in_2_5;
      end else if (10'h223 == _T_28[9:0]) begin
        image_2_547 <= io_pixelVal_in_2_4;
      end else if (10'h223 == _T_25[9:0]) begin
        image_2_547 <= io_pixelVal_in_2_3;
      end else if (10'h223 == _T_22[9:0]) begin
        image_2_547 <= io_pixelVal_in_2_2;
      end else if (10'h223 == _T_19[9:0]) begin
        image_2_547 <= io_pixelVal_in_2_1;
      end else if (10'h223 == _T_15[9:0]) begin
        image_2_547 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_548 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h224 == _T_37[9:0]) begin
        image_2_548 <= io_pixelVal_in_2_7;
      end else if (10'h224 == _T_34[9:0]) begin
        image_2_548 <= io_pixelVal_in_2_6;
      end else if (10'h224 == _T_31[9:0]) begin
        image_2_548 <= io_pixelVal_in_2_5;
      end else if (10'h224 == _T_28[9:0]) begin
        image_2_548 <= io_pixelVal_in_2_4;
      end else if (10'h224 == _T_25[9:0]) begin
        image_2_548 <= io_pixelVal_in_2_3;
      end else if (10'h224 == _T_22[9:0]) begin
        image_2_548 <= io_pixelVal_in_2_2;
      end else if (10'h224 == _T_19[9:0]) begin
        image_2_548 <= io_pixelVal_in_2_1;
      end else if (10'h224 == _T_15[9:0]) begin
        image_2_548 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_549 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h225 == _T_37[9:0]) begin
        image_2_549 <= io_pixelVal_in_2_7;
      end else if (10'h225 == _T_34[9:0]) begin
        image_2_549 <= io_pixelVal_in_2_6;
      end else if (10'h225 == _T_31[9:0]) begin
        image_2_549 <= io_pixelVal_in_2_5;
      end else if (10'h225 == _T_28[9:0]) begin
        image_2_549 <= io_pixelVal_in_2_4;
      end else if (10'h225 == _T_25[9:0]) begin
        image_2_549 <= io_pixelVal_in_2_3;
      end else if (10'h225 == _T_22[9:0]) begin
        image_2_549 <= io_pixelVal_in_2_2;
      end else if (10'h225 == _T_19[9:0]) begin
        image_2_549 <= io_pixelVal_in_2_1;
      end else if (10'h225 == _T_15[9:0]) begin
        image_2_549 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_550 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h226 == _T_37[9:0]) begin
        image_2_550 <= io_pixelVal_in_2_7;
      end else if (10'h226 == _T_34[9:0]) begin
        image_2_550 <= io_pixelVal_in_2_6;
      end else if (10'h226 == _T_31[9:0]) begin
        image_2_550 <= io_pixelVal_in_2_5;
      end else if (10'h226 == _T_28[9:0]) begin
        image_2_550 <= io_pixelVal_in_2_4;
      end else if (10'h226 == _T_25[9:0]) begin
        image_2_550 <= io_pixelVal_in_2_3;
      end else if (10'h226 == _T_22[9:0]) begin
        image_2_550 <= io_pixelVal_in_2_2;
      end else if (10'h226 == _T_19[9:0]) begin
        image_2_550 <= io_pixelVal_in_2_1;
      end else if (10'h226 == _T_15[9:0]) begin
        image_2_550 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_551 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h227 == _T_37[9:0]) begin
        image_2_551 <= io_pixelVal_in_2_7;
      end else if (10'h227 == _T_34[9:0]) begin
        image_2_551 <= io_pixelVal_in_2_6;
      end else if (10'h227 == _T_31[9:0]) begin
        image_2_551 <= io_pixelVal_in_2_5;
      end else if (10'h227 == _T_28[9:0]) begin
        image_2_551 <= io_pixelVal_in_2_4;
      end else if (10'h227 == _T_25[9:0]) begin
        image_2_551 <= io_pixelVal_in_2_3;
      end else if (10'h227 == _T_22[9:0]) begin
        image_2_551 <= io_pixelVal_in_2_2;
      end else if (10'h227 == _T_19[9:0]) begin
        image_2_551 <= io_pixelVal_in_2_1;
      end else if (10'h227 == _T_15[9:0]) begin
        image_2_551 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_552 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h228 == _T_37[9:0]) begin
        image_2_552 <= io_pixelVal_in_2_7;
      end else if (10'h228 == _T_34[9:0]) begin
        image_2_552 <= io_pixelVal_in_2_6;
      end else if (10'h228 == _T_31[9:0]) begin
        image_2_552 <= io_pixelVal_in_2_5;
      end else if (10'h228 == _T_28[9:0]) begin
        image_2_552 <= io_pixelVal_in_2_4;
      end else if (10'h228 == _T_25[9:0]) begin
        image_2_552 <= io_pixelVal_in_2_3;
      end else if (10'h228 == _T_22[9:0]) begin
        image_2_552 <= io_pixelVal_in_2_2;
      end else if (10'h228 == _T_19[9:0]) begin
        image_2_552 <= io_pixelVal_in_2_1;
      end else if (10'h228 == _T_15[9:0]) begin
        image_2_552 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_553 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h229 == _T_37[9:0]) begin
        image_2_553 <= io_pixelVal_in_2_7;
      end else if (10'h229 == _T_34[9:0]) begin
        image_2_553 <= io_pixelVal_in_2_6;
      end else if (10'h229 == _T_31[9:0]) begin
        image_2_553 <= io_pixelVal_in_2_5;
      end else if (10'h229 == _T_28[9:0]) begin
        image_2_553 <= io_pixelVal_in_2_4;
      end else if (10'h229 == _T_25[9:0]) begin
        image_2_553 <= io_pixelVal_in_2_3;
      end else if (10'h229 == _T_22[9:0]) begin
        image_2_553 <= io_pixelVal_in_2_2;
      end else if (10'h229 == _T_19[9:0]) begin
        image_2_553 <= io_pixelVal_in_2_1;
      end else if (10'h229 == _T_15[9:0]) begin
        image_2_553 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_554 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h22a == _T_37[9:0]) begin
        image_2_554 <= io_pixelVal_in_2_7;
      end else if (10'h22a == _T_34[9:0]) begin
        image_2_554 <= io_pixelVal_in_2_6;
      end else if (10'h22a == _T_31[9:0]) begin
        image_2_554 <= io_pixelVal_in_2_5;
      end else if (10'h22a == _T_28[9:0]) begin
        image_2_554 <= io_pixelVal_in_2_4;
      end else if (10'h22a == _T_25[9:0]) begin
        image_2_554 <= io_pixelVal_in_2_3;
      end else if (10'h22a == _T_22[9:0]) begin
        image_2_554 <= io_pixelVal_in_2_2;
      end else if (10'h22a == _T_19[9:0]) begin
        image_2_554 <= io_pixelVal_in_2_1;
      end else if (10'h22a == _T_15[9:0]) begin
        image_2_554 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_555 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h22b == _T_37[9:0]) begin
        image_2_555 <= io_pixelVal_in_2_7;
      end else if (10'h22b == _T_34[9:0]) begin
        image_2_555 <= io_pixelVal_in_2_6;
      end else if (10'h22b == _T_31[9:0]) begin
        image_2_555 <= io_pixelVal_in_2_5;
      end else if (10'h22b == _T_28[9:0]) begin
        image_2_555 <= io_pixelVal_in_2_4;
      end else if (10'h22b == _T_25[9:0]) begin
        image_2_555 <= io_pixelVal_in_2_3;
      end else if (10'h22b == _T_22[9:0]) begin
        image_2_555 <= io_pixelVal_in_2_2;
      end else if (10'h22b == _T_19[9:0]) begin
        image_2_555 <= io_pixelVal_in_2_1;
      end else if (10'h22b == _T_15[9:0]) begin
        image_2_555 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_556 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h22c == _T_37[9:0]) begin
        image_2_556 <= io_pixelVal_in_2_7;
      end else if (10'h22c == _T_34[9:0]) begin
        image_2_556 <= io_pixelVal_in_2_6;
      end else if (10'h22c == _T_31[9:0]) begin
        image_2_556 <= io_pixelVal_in_2_5;
      end else if (10'h22c == _T_28[9:0]) begin
        image_2_556 <= io_pixelVal_in_2_4;
      end else if (10'h22c == _T_25[9:0]) begin
        image_2_556 <= io_pixelVal_in_2_3;
      end else if (10'h22c == _T_22[9:0]) begin
        image_2_556 <= io_pixelVal_in_2_2;
      end else if (10'h22c == _T_19[9:0]) begin
        image_2_556 <= io_pixelVal_in_2_1;
      end else if (10'h22c == _T_15[9:0]) begin
        image_2_556 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_557 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h22d == _T_37[9:0]) begin
        image_2_557 <= io_pixelVal_in_2_7;
      end else if (10'h22d == _T_34[9:0]) begin
        image_2_557 <= io_pixelVal_in_2_6;
      end else if (10'h22d == _T_31[9:0]) begin
        image_2_557 <= io_pixelVal_in_2_5;
      end else if (10'h22d == _T_28[9:0]) begin
        image_2_557 <= io_pixelVal_in_2_4;
      end else if (10'h22d == _T_25[9:0]) begin
        image_2_557 <= io_pixelVal_in_2_3;
      end else if (10'h22d == _T_22[9:0]) begin
        image_2_557 <= io_pixelVal_in_2_2;
      end else if (10'h22d == _T_19[9:0]) begin
        image_2_557 <= io_pixelVal_in_2_1;
      end else if (10'h22d == _T_15[9:0]) begin
        image_2_557 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_558 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h22e == _T_37[9:0]) begin
        image_2_558 <= io_pixelVal_in_2_7;
      end else if (10'h22e == _T_34[9:0]) begin
        image_2_558 <= io_pixelVal_in_2_6;
      end else if (10'h22e == _T_31[9:0]) begin
        image_2_558 <= io_pixelVal_in_2_5;
      end else if (10'h22e == _T_28[9:0]) begin
        image_2_558 <= io_pixelVal_in_2_4;
      end else if (10'h22e == _T_25[9:0]) begin
        image_2_558 <= io_pixelVal_in_2_3;
      end else if (10'h22e == _T_22[9:0]) begin
        image_2_558 <= io_pixelVal_in_2_2;
      end else if (10'h22e == _T_19[9:0]) begin
        image_2_558 <= io_pixelVal_in_2_1;
      end else if (10'h22e == _T_15[9:0]) begin
        image_2_558 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_559 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h22f == _T_37[9:0]) begin
        image_2_559 <= io_pixelVal_in_2_7;
      end else if (10'h22f == _T_34[9:0]) begin
        image_2_559 <= io_pixelVal_in_2_6;
      end else if (10'h22f == _T_31[9:0]) begin
        image_2_559 <= io_pixelVal_in_2_5;
      end else if (10'h22f == _T_28[9:0]) begin
        image_2_559 <= io_pixelVal_in_2_4;
      end else if (10'h22f == _T_25[9:0]) begin
        image_2_559 <= io_pixelVal_in_2_3;
      end else if (10'h22f == _T_22[9:0]) begin
        image_2_559 <= io_pixelVal_in_2_2;
      end else if (10'h22f == _T_19[9:0]) begin
        image_2_559 <= io_pixelVal_in_2_1;
      end else if (10'h22f == _T_15[9:0]) begin
        image_2_559 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_560 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h230 == _T_37[9:0]) begin
        image_2_560 <= io_pixelVal_in_2_7;
      end else if (10'h230 == _T_34[9:0]) begin
        image_2_560 <= io_pixelVal_in_2_6;
      end else if (10'h230 == _T_31[9:0]) begin
        image_2_560 <= io_pixelVal_in_2_5;
      end else if (10'h230 == _T_28[9:0]) begin
        image_2_560 <= io_pixelVal_in_2_4;
      end else if (10'h230 == _T_25[9:0]) begin
        image_2_560 <= io_pixelVal_in_2_3;
      end else if (10'h230 == _T_22[9:0]) begin
        image_2_560 <= io_pixelVal_in_2_2;
      end else if (10'h230 == _T_19[9:0]) begin
        image_2_560 <= io_pixelVal_in_2_1;
      end else if (10'h230 == _T_15[9:0]) begin
        image_2_560 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_561 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h231 == _T_37[9:0]) begin
        image_2_561 <= io_pixelVal_in_2_7;
      end else if (10'h231 == _T_34[9:0]) begin
        image_2_561 <= io_pixelVal_in_2_6;
      end else if (10'h231 == _T_31[9:0]) begin
        image_2_561 <= io_pixelVal_in_2_5;
      end else if (10'h231 == _T_28[9:0]) begin
        image_2_561 <= io_pixelVal_in_2_4;
      end else if (10'h231 == _T_25[9:0]) begin
        image_2_561 <= io_pixelVal_in_2_3;
      end else if (10'h231 == _T_22[9:0]) begin
        image_2_561 <= io_pixelVal_in_2_2;
      end else if (10'h231 == _T_19[9:0]) begin
        image_2_561 <= io_pixelVal_in_2_1;
      end else if (10'h231 == _T_15[9:0]) begin
        image_2_561 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_562 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h232 == _T_37[9:0]) begin
        image_2_562 <= io_pixelVal_in_2_7;
      end else if (10'h232 == _T_34[9:0]) begin
        image_2_562 <= io_pixelVal_in_2_6;
      end else if (10'h232 == _T_31[9:0]) begin
        image_2_562 <= io_pixelVal_in_2_5;
      end else if (10'h232 == _T_28[9:0]) begin
        image_2_562 <= io_pixelVal_in_2_4;
      end else if (10'h232 == _T_25[9:0]) begin
        image_2_562 <= io_pixelVal_in_2_3;
      end else if (10'h232 == _T_22[9:0]) begin
        image_2_562 <= io_pixelVal_in_2_2;
      end else if (10'h232 == _T_19[9:0]) begin
        image_2_562 <= io_pixelVal_in_2_1;
      end else if (10'h232 == _T_15[9:0]) begin
        image_2_562 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_563 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h233 == _T_37[9:0]) begin
        image_2_563 <= io_pixelVal_in_2_7;
      end else if (10'h233 == _T_34[9:0]) begin
        image_2_563 <= io_pixelVal_in_2_6;
      end else if (10'h233 == _T_31[9:0]) begin
        image_2_563 <= io_pixelVal_in_2_5;
      end else if (10'h233 == _T_28[9:0]) begin
        image_2_563 <= io_pixelVal_in_2_4;
      end else if (10'h233 == _T_25[9:0]) begin
        image_2_563 <= io_pixelVal_in_2_3;
      end else if (10'h233 == _T_22[9:0]) begin
        image_2_563 <= io_pixelVal_in_2_2;
      end else if (10'h233 == _T_19[9:0]) begin
        image_2_563 <= io_pixelVal_in_2_1;
      end else if (10'h233 == _T_15[9:0]) begin
        image_2_563 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_564 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h234 == _T_37[9:0]) begin
        image_2_564 <= io_pixelVal_in_2_7;
      end else if (10'h234 == _T_34[9:0]) begin
        image_2_564 <= io_pixelVal_in_2_6;
      end else if (10'h234 == _T_31[9:0]) begin
        image_2_564 <= io_pixelVal_in_2_5;
      end else if (10'h234 == _T_28[9:0]) begin
        image_2_564 <= io_pixelVal_in_2_4;
      end else if (10'h234 == _T_25[9:0]) begin
        image_2_564 <= io_pixelVal_in_2_3;
      end else if (10'h234 == _T_22[9:0]) begin
        image_2_564 <= io_pixelVal_in_2_2;
      end else if (10'h234 == _T_19[9:0]) begin
        image_2_564 <= io_pixelVal_in_2_1;
      end else if (10'h234 == _T_15[9:0]) begin
        image_2_564 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_565 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h235 == _T_37[9:0]) begin
        image_2_565 <= io_pixelVal_in_2_7;
      end else if (10'h235 == _T_34[9:0]) begin
        image_2_565 <= io_pixelVal_in_2_6;
      end else if (10'h235 == _T_31[9:0]) begin
        image_2_565 <= io_pixelVal_in_2_5;
      end else if (10'h235 == _T_28[9:0]) begin
        image_2_565 <= io_pixelVal_in_2_4;
      end else if (10'h235 == _T_25[9:0]) begin
        image_2_565 <= io_pixelVal_in_2_3;
      end else if (10'h235 == _T_22[9:0]) begin
        image_2_565 <= io_pixelVal_in_2_2;
      end else if (10'h235 == _T_19[9:0]) begin
        image_2_565 <= io_pixelVal_in_2_1;
      end else if (10'h235 == _T_15[9:0]) begin
        image_2_565 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_566 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h236 == _T_37[9:0]) begin
        image_2_566 <= io_pixelVal_in_2_7;
      end else if (10'h236 == _T_34[9:0]) begin
        image_2_566 <= io_pixelVal_in_2_6;
      end else if (10'h236 == _T_31[9:0]) begin
        image_2_566 <= io_pixelVal_in_2_5;
      end else if (10'h236 == _T_28[9:0]) begin
        image_2_566 <= io_pixelVal_in_2_4;
      end else if (10'h236 == _T_25[9:0]) begin
        image_2_566 <= io_pixelVal_in_2_3;
      end else if (10'h236 == _T_22[9:0]) begin
        image_2_566 <= io_pixelVal_in_2_2;
      end else if (10'h236 == _T_19[9:0]) begin
        image_2_566 <= io_pixelVal_in_2_1;
      end else if (10'h236 == _T_15[9:0]) begin
        image_2_566 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_567 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h237 == _T_37[9:0]) begin
        image_2_567 <= io_pixelVal_in_2_7;
      end else if (10'h237 == _T_34[9:0]) begin
        image_2_567 <= io_pixelVal_in_2_6;
      end else if (10'h237 == _T_31[9:0]) begin
        image_2_567 <= io_pixelVal_in_2_5;
      end else if (10'h237 == _T_28[9:0]) begin
        image_2_567 <= io_pixelVal_in_2_4;
      end else if (10'h237 == _T_25[9:0]) begin
        image_2_567 <= io_pixelVal_in_2_3;
      end else if (10'h237 == _T_22[9:0]) begin
        image_2_567 <= io_pixelVal_in_2_2;
      end else if (10'h237 == _T_19[9:0]) begin
        image_2_567 <= io_pixelVal_in_2_1;
      end else if (10'h237 == _T_15[9:0]) begin
        image_2_567 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_568 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h238 == _T_37[9:0]) begin
        image_2_568 <= io_pixelVal_in_2_7;
      end else if (10'h238 == _T_34[9:0]) begin
        image_2_568 <= io_pixelVal_in_2_6;
      end else if (10'h238 == _T_31[9:0]) begin
        image_2_568 <= io_pixelVal_in_2_5;
      end else if (10'h238 == _T_28[9:0]) begin
        image_2_568 <= io_pixelVal_in_2_4;
      end else if (10'h238 == _T_25[9:0]) begin
        image_2_568 <= io_pixelVal_in_2_3;
      end else if (10'h238 == _T_22[9:0]) begin
        image_2_568 <= io_pixelVal_in_2_2;
      end else if (10'h238 == _T_19[9:0]) begin
        image_2_568 <= io_pixelVal_in_2_1;
      end else if (10'h238 == _T_15[9:0]) begin
        image_2_568 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_569 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h239 == _T_37[9:0]) begin
        image_2_569 <= io_pixelVal_in_2_7;
      end else if (10'h239 == _T_34[9:0]) begin
        image_2_569 <= io_pixelVal_in_2_6;
      end else if (10'h239 == _T_31[9:0]) begin
        image_2_569 <= io_pixelVal_in_2_5;
      end else if (10'h239 == _T_28[9:0]) begin
        image_2_569 <= io_pixelVal_in_2_4;
      end else if (10'h239 == _T_25[9:0]) begin
        image_2_569 <= io_pixelVal_in_2_3;
      end else if (10'h239 == _T_22[9:0]) begin
        image_2_569 <= io_pixelVal_in_2_2;
      end else if (10'h239 == _T_19[9:0]) begin
        image_2_569 <= io_pixelVal_in_2_1;
      end else if (10'h239 == _T_15[9:0]) begin
        image_2_569 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_570 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h23a == _T_37[9:0]) begin
        image_2_570 <= io_pixelVal_in_2_7;
      end else if (10'h23a == _T_34[9:0]) begin
        image_2_570 <= io_pixelVal_in_2_6;
      end else if (10'h23a == _T_31[9:0]) begin
        image_2_570 <= io_pixelVal_in_2_5;
      end else if (10'h23a == _T_28[9:0]) begin
        image_2_570 <= io_pixelVal_in_2_4;
      end else if (10'h23a == _T_25[9:0]) begin
        image_2_570 <= io_pixelVal_in_2_3;
      end else if (10'h23a == _T_22[9:0]) begin
        image_2_570 <= io_pixelVal_in_2_2;
      end else if (10'h23a == _T_19[9:0]) begin
        image_2_570 <= io_pixelVal_in_2_1;
      end else if (10'h23a == _T_15[9:0]) begin
        image_2_570 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_571 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h23b == _T_37[9:0]) begin
        image_2_571 <= io_pixelVal_in_2_7;
      end else if (10'h23b == _T_34[9:0]) begin
        image_2_571 <= io_pixelVal_in_2_6;
      end else if (10'h23b == _T_31[9:0]) begin
        image_2_571 <= io_pixelVal_in_2_5;
      end else if (10'h23b == _T_28[9:0]) begin
        image_2_571 <= io_pixelVal_in_2_4;
      end else if (10'h23b == _T_25[9:0]) begin
        image_2_571 <= io_pixelVal_in_2_3;
      end else if (10'h23b == _T_22[9:0]) begin
        image_2_571 <= io_pixelVal_in_2_2;
      end else if (10'h23b == _T_19[9:0]) begin
        image_2_571 <= io_pixelVal_in_2_1;
      end else if (10'h23b == _T_15[9:0]) begin
        image_2_571 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_572 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h23c == _T_37[9:0]) begin
        image_2_572 <= io_pixelVal_in_2_7;
      end else if (10'h23c == _T_34[9:0]) begin
        image_2_572 <= io_pixelVal_in_2_6;
      end else if (10'h23c == _T_31[9:0]) begin
        image_2_572 <= io_pixelVal_in_2_5;
      end else if (10'h23c == _T_28[9:0]) begin
        image_2_572 <= io_pixelVal_in_2_4;
      end else if (10'h23c == _T_25[9:0]) begin
        image_2_572 <= io_pixelVal_in_2_3;
      end else if (10'h23c == _T_22[9:0]) begin
        image_2_572 <= io_pixelVal_in_2_2;
      end else if (10'h23c == _T_19[9:0]) begin
        image_2_572 <= io_pixelVal_in_2_1;
      end else if (10'h23c == _T_15[9:0]) begin
        image_2_572 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_573 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h23d == _T_37[9:0]) begin
        image_2_573 <= io_pixelVal_in_2_7;
      end else if (10'h23d == _T_34[9:0]) begin
        image_2_573 <= io_pixelVal_in_2_6;
      end else if (10'h23d == _T_31[9:0]) begin
        image_2_573 <= io_pixelVal_in_2_5;
      end else if (10'h23d == _T_28[9:0]) begin
        image_2_573 <= io_pixelVal_in_2_4;
      end else if (10'h23d == _T_25[9:0]) begin
        image_2_573 <= io_pixelVal_in_2_3;
      end else if (10'h23d == _T_22[9:0]) begin
        image_2_573 <= io_pixelVal_in_2_2;
      end else if (10'h23d == _T_19[9:0]) begin
        image_2_573 <= io_pixelVal_in_2_1;
      end else if (10'h23d == _T_15[9:0]) begin
        image_2_573 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_574 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h23e == _T_37[9:0]) begin
        image_2_574 <= io_pixelVal_in_2_7;
      end else if (10'h23e == _T_34[9:0]) begin
        image_2_574 <= io_pixelVal_in_2_6;
      end else if (10'h23e == _T_31[9:0]) begin
        image_2_574 <= io_pixelVal_in_2_5;
      end else if (10'h23e == _T_28[9:0]) begin
        image_2_574 <= io_pixelVal_in_2_4;
      end else if (10'h23e == _T_25[9:0]) begin
        image_2_574 <= io_pixelVal_in_2_3;
      end else if (10'h23e == _T_22[9:0]) begin
        image_2_574 <= io_pixelVal_in_2_2;
      end else if (10'h23e == _T_19[9:0]) begin
        image_2_574 <= io_pixelVal_in_2_1;
      end else if (10'h23e == _T_15[9:0]) begin
        image_2_574 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      image_2_575 <= 4'h0;
    end else if (io_valid_in) begin
      if (10'h23f == _T_37[9:0]) begin
        image_2_575 <= io_pixelVal_in_2_7;
      end else if (10'h23f == _T_34[9:0]) begin
        image_2_575 <= io_pixelVal_in_2_6;
      end else if (10'h23f == _T_31[9:0]) begin
        image_2_575 <= io_pixelVal_in_2_5;
      end else if (10'h23f == _T_28[9:0]) begin
        image_2_575 <= io_pixelVal_in_2_4;
      end else if (10'h23f == _T_25[9:0]) begin
        image_2_575 <= io_pixelVal_in_2_3;
      end else if (10'h23f == _T_22[9:0]) begin
        image_2_575 <= io_pixelVal_in_2_2;
      end else if (10'h23f == _T_19[9:0]) begin
        image_2_575 <= io_pixelVal_in_2_1;
      end else if (10'h23f == _T_15[9:0]) begin
        image_2_575 <= io_pixelVal_in_2_0;
      end
    end
    if (reset) begin
      pixelIndex <= 32'h0;
    end else if (io_valid_in) begin
      if (_T_90) begin
        pixelIndex <= 32'h0;
      end else begin
        pixelIndex <= _T_88;
      end
    end
  end
endmodule
module ImageProcessing(
  input         clock,
  input         reset,
  input  [5:0]  io_SPI_filterIndex,
  input         io_SPI_invert,
  input         io_SPI_distort,
  input  [10:0] io_rowIndex,
  input  [10:0] io_colIndex,
  output [3:0]  io_pixelVal_out_0,
  output [3:0]  io_pixelVal_out_1,
  output [3:0]  io_pixelVal_out_2
);
  wire  filter_clock; // @[ImageProcessing.scala 23:22]
  wire  filter_reset; // @[ImageProcessing.scala 23:22]
  wire [5:0] filter_io_SPI_filterIndex; // @[ImageProcessing.scala 23:22]
  wire  filter_io_SPI_invert; // @[ImageProcessing.scala 23:22]
  wire  filter_io_SPI_distort; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_0; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_1; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_2; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_3; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_4; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_5; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_6; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_0_7; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_0; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_1; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_2; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_3; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_4; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_5; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_6; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_1_7; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_0; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_1; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_2; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_3; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_4; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_5; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_6; // @[ImageProcessing.scala 23:22]
  wire [3:0] filter_io_pixelVal_out_2_7; // @[ImageProcessing.scala 23:22]
  wire  filter_io_valid_out; // @[ImageProcessing.scala 23:22]
  wire  videoBuffer_clock; // @[ImageProcessing.scala 24:27]
  wire  videoBuffer_reset; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_0; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_1; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_2; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_3; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_4; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_5; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_6; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_0_7; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_0; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_1; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_2; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_3; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_4; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_5; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_6; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_1_7; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_0; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_1; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_2; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_3; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_4; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_5; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_6; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_in_2_7; // @[ImageProcessing.scala 24:27]
  wire  videoBuffer_io_valid_in; // @[ImageProcessing.scala 24:27]
  wire [10:0] videoBuffer_io_rowIndex; // @[ImageProcessing.scala 24:27]
  wire [10:0] videoBuffer_io_colIndex; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_out_0; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_out_1; // @[ImageProcessing.scala 24:27]
  wire [3:0] videoBuffer_io_pixelVal_out_2; // @[ImageProcessing.scala 24:27]
  Filter filter ( // @[ImageProcessing.scala 23:22]
    .clock(filter_clock),
    .reset(filter_reset),
    .io_SPI_filterIndex(filter_io_SPI_filterIndex),
    .io_SPI_invert(filter_io_SPI_invert),
    .io_SPI_distort(filter_io_SPI_distort),
    .io_pixelVal_out_0_0(filter_io_pixelVal_out_0_0),
    .io_pixelVal_out_0_1(filter_io_pixelVal_out_0_1),
    .io_pixelVal_out_0_2(filter_io_pixelVal_out_0_2),
    .io_pixelVal_out_0_3(filter_io_pixelVal_out_0_3),
    .io_pixelVal_out_0_4(filter_io_pixelVal_out_0_4),
    .io_pixelVal_out_0_5(filter_io_pixelVal_out_0_5),
    .io_pixelVal_out_0_6(filter_io_pixelVal_out_0_6),
    .io_pixelVal_out_0_7(filter_io_pixelVal_out_0_7),
    .io_pixelVal_out_1_0(filter_io_pixelVal_out_1_0),
    .io_pixelVal_out_1_1(filter_io_pixelVal_out_1_1),
    .io_pixelVal_out_1_2(filter_io_pixelVal_out_1_2),
    .io_pixelVal_out_1_3(filter_io_pixelVal_out_1_3),
    .io_pixelVal_out_1_4(filter_io_pixelVal_out_1_4),
    .io_pixelVal_out_1_5(filter_io_pixelVal_out_1_5),
    .io_pixelVal_out_1_6(filter_io_pixelVal_out_1_6),
    .io_pixelVal_out_1_7(filter_io_pixelVal_out_1_7),
    .io_pixelVal_out_2_0(filter_io_pixelVal_out_2_0),
    .io_pixelVal_out_2_1(filter_io_pixelVal_out_2_1),
    .io_pixelVal_out_2_2(filter_io_pixelVal_out_2_2),
    .io_pixelVal_out_2_3(filter_io_pixelVal_out_2_3),
    .io_pixelVal_out_2_4(filter_io_pixelVal_out_2_4),
    .io_pixelVal_out_2_5(filter_io_pixelVal_out_2_5),
    .io_pixelVal_out_2_6(filter_io_pixelVal_out_2_6),
    .io_pixelVal_out_2_7(filter_io_pixelVal_out_2_7),
    .io_valid_out(filter_io_valid_out)
  );
  VideoBuffer videoBuffer ( // @[ImageProcessing.scala 24:27]
    .clock(videoBuffer_clock),
    .reset(videoBuffer_reset),
    .io_pixelVal_in_0_0(videoBuffer_io_pixelVal_in_0_0),
    .io_pixelVal_in_0_1(videoBuffer_io_pixelVal_in_0_1),
    .io_pixelVal_in_0_2(videoBuffer_io_pixelVal_in_0_2),
    .io_pixelVal_in_0_3(videoBuffer_io_pixelVal_in_0_3),
    .io_pixelVal_in_0_4(videoBuffer_io_pixelVal_in_0_4),
    .io_pixelVal_in_0_5(videoBuffer_io_pixelVal_in_0_5),
    .io_pixelVal_in_0_6(videoBuffer_io_pixelVal_in_0_6),
    .io_pixelVal_in_0_7(videoBuffer_io_pixelVal_in_0_7),
    .io_pixelVal_in_1_0(videoBuffer_io_pixelVal_in_1_0),
    .io_pixelVal_in_1_1(videoBuffer_io_pixelVal_in_1_1),
    .io_pixelVal_in_1_2(videoBuffer_io_pixelVal_in_1_2),
    .io_pixelVal_in_1_3(videoBuffer_io_pixelVal_in_1_3),
    .io_pixelVal_in_1_4(videoBuffer_io_pixelVal_in_1_4),
    .io_pixelVal_in_1_5(videoBuffer_io_pixelVal_in_1_5),
    .io_pixelVal_in_1_6(videoBuffer_io_pixelVal_in_1_6),
    .io_pixelVal_in_1_7(videoBuffer_io_pixelVal_in_1_7),
    .io_pixelVal_in_2_0(videoBuffer_io_pixelVal_in_2_0),
    .io_pixelVal_in_2_1(videoBuffer_io_pixelVal_in_2_1),
    .io_pixelVal_in_2_2(videoBuffer_io_pixelVal_in_2_2),
    .io_pixelVal_in_2_3(videoBuffer_io_pixelVal_in_2_3),
    .io_pixelVal_in_2_4(videoBuffer_io_pixelVal_in_2_4),
    .io_pixelVal_in_2_5(videoBuffer_io_pixelVal_in_2_5),
    .io_pixelVal_in_2_6(videoBuffer_io_pixelVal_in_2_6),
    .io_pixelVal_in_2_7(videoBuffer_io_pixelVal_in_2_7),
    .io_valid_in(videoBuffer_io_valid_in),
    .io_rowIndex(videoBuffer_io_rowIndex),
    .io_colIndex(videoBuffer_io_colIndex),
    .io_pixelVal_out_0(videoBuffer_io_pixelVal_out_0),
    .io_pixelVal_out_1(videoBuffer_io_pixelVal_out_1),
    .io_pixelVal_out_2(videoBuffer_io_pixelVal_out_2)
  );
  assign io_pixelVal_out_0 = videoBuffer_io_pixelVal_out_0; // @[ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25]
  assign io_pixelVal_out_1 = videoBuffer_io_pixelVal_out_1; // @[ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25]
  assign io_pixelVal_out_2 = videoBuffer_io_pixelVal_out_2; // @[ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25 ImageProcessing.scala 36:25]
  assign filter_clock = clock;
  assign filter_reset = reset;
  assign filter_io_SPI_filterIndex = io_SPI_filterIndex; // @[ImageProcessing.scala 29:29]
  assign filter_io_SPI_invert = io_SPI_invert; // @[ImageProcessing.scala 30:29]
  assign filter_io_SPI_distort = io_SPI_distort; // @[ImageProcessing.scala 31:29]
  assign videoBuffer_clock = clock;
  assign videoBuffer_reset = reset;
  assign videoBuffer_io_pixelVal_in_0_0 = filter_io_pixelVal_out_0_0; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_0_1 = filter_io_pixelVal_out_0_1; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_0_2 = filter_io_pixelVal_out_0_2; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_0_3 = filter_io_pixelVal_out_0_3; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_0_4 = filter_io_pixelVal_out_0_4; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_0_5 = filter_io_pixelVal_out_0_5; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_0_6 = filter_io_pixelVal_out_0_6; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_0_7 = filter_io_pixelVal_out_0_7; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_0 = filter_io_pixelVal_out_1_0; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_1 = filter_io_pixelVal_out_1_1; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_2 = filter_io_pixelVal_out_1_2; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_3 = filter_io_pixelVal_out_1_3; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_4 = filter_io_pixelVal_out_1_4; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_5 = filter_io_pixelVal_out_1_5; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_6 = filter_io_pixelVal_out_1_6; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_1_7 = filter_io_pixelVal_out_1_7; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_0 = filter_io_pixelVal_out_2_0; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_1 = filter_io_pixelVal_out_2_1; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_2 = filter_io_pixelVal_out_2_2; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_3 = filter_io_pixelVal_out_2_3; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_4 = filter_io_pixelVal_out_2_4; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_5 = filter_io_pixelVal_out_2_5; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_6 = filter_io_pixelVal_out_2_6; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_pixelVal_in_2_7 = filter_io_pixelVal_out_2_7; // @[ImageProcessing.scala 35:39]
  assign videoBuffer_io_valid_in = filter_io_valid_out; // @[ImageProcessing.scala 39:27]
  assign videoBuffer_io_rowIndex = io_rowIndex; // @[ImageProcessing.scala 26:27]
  assign videoBuffer_io_colIndex = io_colIndex; // @[ImageProcessing.scala 27:27]
endmodule
